// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AEuiH+Ynxc0Pp6zXZVMNFJ+l4dwhsALfPYFS8wtUPxzYddolsgtmtD+HXdPBCib7
z8in0+ovwOiVF3EVqzUHas58J1/FRpmQIXB+K0YhKlH1jMu1KXIsGkpUM2gjlhAV
+ORaO0f+7RSx+Iq+mDrhc6xTiTUUpRbirWfGKxCzqJA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2038688)
xn5c5yft1Myj4HQhp2O0nS2+c75l0qCDrfmNHxZGbgSpTfvH+bOJ2/R8S5SrWIeb
xkdUU7uo3G9o/SLIfgIZWsrk357A+wtdy+FYVyFi1T1gJz550Oawt8RoMVfm9hJp
Jjwg7pdRz9V9ncgiB0WcitNGuo9JJlF25+nmrReW7hR6eCEwtkI8kKzXL7O+nq7o
JmLOFqc8OpqM4aw2GzJ8vCilDIljq/TJualE+jm0u4scypzvE70CDz95aTTHrGDy
C143Flt1C3mUnBhDLe8tkRnPDp7jyNLiIH3Z03t+Kp3gamHK5eRANAg9jGEkfx8C
oIcnFqU9Txayi067PHGrzxLGya7lgJW7PoBW22CYo5sh62I1o/Hxs9nrRMEg51x5
UooV/6ruulpWFIwa0+sYByf0m0JsM91sX80W9xOkkzPkx9ZICiryK+DakOSxkDmT
UX2VLVDaUALu+SbsiLiFchqMsmvBaiOrOq/sAAyGVjo9M7iUWAg60vVGuJg9ZKx/
+dULE3mEXt2qPq8to8OsnHuKaQgLZG9+74qo57xc2vi4/cZ3YL2ZRf4vqE7uLWFu
i8KLSYjE98tToi/mE7MsW+VMRpk8gELr/M3Ee2os/AFtpOiRXPLj5oZ4f+cIN7Kg
fUkqls4a0OQI2UhMfxRlrA0N7OKNgyyyNevBAMNyagOdGJDDhHkRudptTiiAinNZ
z+kMhUp6zClE0OBkyldj8NgoY2zPadGncpreuFe39qxRO1eUCWDyIA+gZv3/6qQ8
GxoxzCEXQWs3a4l9ju8jVaCjDXldoGUo6texJT2FUeChTNkjPRScYXMUwJX6Zyhu
j58IhlWfQMky2n5ivXenQoeF3xbsYmP0Vdp7ul62KXcSNm3pZVbleFJ6zwSW5T22
yF2pfLM80Anvskh6tSHkwk9/y/K/LG8VhRvnw6+mq0LPhh+OcXeuKJKex8zdz26C
/4gs9KmpXouzpP0gs0LBlsRAQzlffrwZIZZhG0FyIxXDuMQfCyzUC6g5K4PLMiCg
RdDHRvShcElIUT6r51BVCJ6qjqv5oURrIoRuiaZ26YfNk3wl+RLFnDyP6AfGv/WN
YHu4M4n8SVjyVXLSOSVZZnPM+ErD+7Mwd57au83EItiPEKRG1ZxxFExIP+VOCYD2
F9UJv+iYPVF+sEr9QMOPK9dHZX/vrx+KDzt594WHgmS46LGxNyWnxtX6+PQoSONR
AQhxwmNHPBxrvAi1hstcwPLu9a1SLRg+HpR+dbXqsLbigfk8iwV4OosWW2NiGZXi
UUEDo5gEqvgu+M2oB1WuEfIpfogkyFsZqcBBlhND5X5vLxwwzN1uEeoH3laq3IY0
l3+N0x0Es7V4ku3gKcKWHn1hyezvxRdorsomjE8GuRBlFuKYBDNOp+vanX0Q8/kl
cUNLQPrUrGAs8CL9WOauXexQ7H6+L2B5n9kZ7Sh+QKeQGz+LD/Uo+wL1medUhB6E
OHopatdYgwTcpmVnTEeupIPydtU4lo+E+/27fNqzWwh+F/JnTyS0+dI+pl5yWqCf
FT0e4WaxyQOI/P0zdPYbMEk/Da9LxlW+aYsEEgnZRZbbxS1ITMLJ6Xc1F9aon4ec
ZKmIMS+ef2KgZtvAVxVv9Jhj7Iq6lKelh487zeYCPUqZVo1HUg1i3gdHp4vWjccf
tOY9ppZJGKCcNzHB5+kZoLiZWN4lCe5TxuqPjSTs67vUNaBSFRDFMfCKt9b7Uh7/
kTqFL2ctSBKViQ5Zcl/d6PLFxB/+N5aKus6M4iQN+lM1Z/QtPRy2qVF0uyDN+HIm
qoumUZxQmHNMwwxktOav0Q1WtkeW4qZQU4AtBunV1rACyRO3oYhmvdj/T8XpP67E
ArUuwBhBPjKrOYeDR+aASaHnAKxg4ce8/wo1vB1nGlHTBOjE5JgkJGzgBFsbb+/d
8teUASTt5vGLOBa32w6LDDEBesc3qw0YN/BOXJgkcsn3wg8MTzhyL+TywT9nkkWc
odKz8Ptx8qeR4/YZtluRDUlYnp44Wz1sh+/ePyATB5EK6X6BOgsU2nptZchFCLWW
kNh7CvVvjJpxuakFyYHt2A/Jzkiqm4lWZimj6Y086jZXvQ/8EZNEKv4hhQxG3jDY
eX8GiKD1BnqH4arKI+C0pbYNE4BIgHTHjm5JVa/vgGCiG6MuA7c2F6kM6YzTKZCh
dVguM2FVswiqPkFu2V8hYkvRJtTVhwLLiOmM5YMXnQnm/Rdf+sR3NMPrQJ1OyLu7
K3DdtuIs/zWSK1XxH1n/+GenoD3VMDuIcJULThEDeUzdBdBAzUX+GYf469tZJf80
gQ6K2sLDXdv/CeVxV15pJYIQcGIEYVHHaqgBDFzBgNUPEZR8jV6IPi/dCHxtxV/4
Bs1Hhu9WMeawZ8y2dBBMU8cRq8f1mjeykNmHj32l8Zge68U09MGoCfhlwr6Mh4YP
jlPLQuYfapZTIT8awjVhUojv4O81p8TOuC4dzwpe6T6A6dXJU3FcnkbVPvN6s6nB
WXqenPc8pgXVLnMK6WbBeud6ifhMOeqS0iJSuvLvV2xIzzVK2JkaoGlUXBPOJoFg
/1we1ejV8KPQ7VzGX9elov/uWt1jUOxSoYQBz3syo0dZQbz1YD4I5M9sx+4nmSNR
RAMYzzn/cicx9vCJR+y5qfQ8z9g/Jsl+ZMMLjoXlpRBLrIrR/2yQwvh3M/n8TBSD
M2twWXuBXHP4iHS89VCgatuCyExEF/5+K3lq1qzofeMEBsayJzX8Tl8e+fFXz0hb
FD7J9Ld9MV/xus8cbMSTPjcbYRfjUBHA/1+2OCLBh614AFw+llbZaxSxzxCbcA0r
hDvC9XE5auxOTKYgaJ6SbOfXGDQxoaZm8MMd857JUaJVKTe7KIb+iu1cImDKHE5J
l8QWudrRQN5I4ADKrxry/eEeZ1dRNDEP11iRpUH+j+E6/+zohur2mjYLryVSBkii
329fN9QXINe4LQH9AZsNCWYHe6PiKB3XbCGennawRtrZVf2ysxAdBSbLVURycBk3
LSWYIEJcHbcYkfa+vgi2JPZOUnkCnMcmf5J4nnvt5qDOUotr3dNXazynWy9o07dQ
KIVnCYimj/oVPPRTlTJ3DsnMHnw9rf3BJ7ao388+NmIwwRMxB3Dusg8vK6sIiIfZ
uEW5ZUazzgFYtB0n9+OQLqbTk/3CyhV7WNiMv6S7TVgSxkLeQ7ReYpT4/lkarkEa
l8nYnRZmw0geTtPE/CpbzzaACI5RdOMSEUyjRnd1QrB41+HoDW4Yv0lUiXbx6Zzn
jZyv6Oh4VROqK6U4tTP6SqKY7zVuPvhedSbqbZyhGrNNWSyomn1qGKEBOL345S56
BDhrO/ec0VOM/mHwcrJRFll4MuwwaO8N1cq7TvZEGtgwCkUc99+Fz4XEKJq/IIMm
sA2UeVDQeU9+xSTpqosoRlWvQb5qqWqJm9NtDtD3P5UizC6risbpRZA2eXbxL8d+
PXVk0kQShZRLs4Odf16ZRFyBYiLNSlm0Z0xWTj2zaTAMWFHvUlyBy0VlTVcas+o3
ZEk0s3XZfez4P6PgJQdB3JzD5hFi3lxrrdlAUaeEKxcfII/tj0UCAiaJBQAoZs60
m8ceLHhxCyCKcp1dkYSkA6Zf9vgTFGzUDptE+YD550Lelgl3poenTQ0QjRNmLGqa
iNeXuOK8GxwIpd3e0eIlkcXC+d5Ek7FbCB+q9iQfgT+KmmKEHnTj8wbtf8JPcKL1
1ZVSBreYwGJGHLwM+z3/fa1krFk/QeTkWs9c9ndXX3lkaYQBWxEZ0NVY63/2WRyy
R8BG6GdXJOfygDmo2idXap48Dj9W4A25EQ9IwpyTWloBMkEPhDJGJzLahu+QH5uR
WomrPk4JPr88tt8YeJSEGyhLPW4JpiaHcPsuNLqz1zETLYK18mNGbXE2AmHBUrJ5
n5A9AWHQ5HNAmSeQUZxLLCBSKvUcIf+wdUR9TTWMBcy/D9f3R4LYH7DjNnzIL77Q
xnXVJ01wNpEywJYWTYBmU8qJrMx7SqentIRzlk6v34EKAoB4Can68EkOOIy57VP7
9xHzz2zuN4XXexgqDcD9Q62FucRmaqXg2Wo+EJP+ZOCEAcpxPxIcePqRp+gRT+H9
11mYSDmohFSbffqzrFpD4Xy5DjKq6TMP6l9mOAzjaqyr3R0MajQWV4buHO8KV9uT
wXpuLQAsG9fxiC9XpvUYLJacYvTc+WymEzZ6l1dPMS9ih/W/I4VU91d6ruM9IUG/
/LD2jdO/JtGm0kWsLXKrNH92RhxHIwGx2ACeferTWNFEk2pBGJJ4CLKyaLNIoLJR
2s5LuISDDUaEiwUlZRtFLahUSnxJol9TGCkK7nP2Xk0jPcYtPOnc01L/jj4yj7nP
wrPdb+NSXiKDBKGiov5kD7Q3+hThv7raGj6JGRt/NKOQT5UZ+xdwn+TZa0q5245v
4n8Y/TvJPOn6K8QyGqzBeFTUeslTtYD0ru7tsL6S0o9x17Dk/z2yESgdDwu8pHtO
7G40x8INcF+wTXIcovLLrq3dOdsBJiH7RhOP91nRLPs1JXtFIWt1H+ueABX5t8XT
m2JFpQDguBxurxSL2AVoZlDu233gLy7tUBgQ7F/CoBiftDzL7Ha05a6tKq7vRD6c
s6348cx9TYhh6q65XG620CDhNHQaPlroJcw3/myOsV9RZaKKIWq0c8h0EibHuq8S
9Xu8PHuwfNG8oshL37UcjvoPNvgPy6ETfUH+19L5lRsjSDI0vjPsW1fvegc72yB0
EHJC/9gulcMVdjirhuXe9J8v3CvkjjvbrjtlSYp9/0ElnLSu+FnVqaQ21H23yIh/
1KJzzuh0B1gR4Iwe3xgB27TYib7TmqyXtK43ozUoGDyb/6lVbDiuNc3F8Q6M+4WM
JwiRRUqBLM0XeYIcQg9T/SpgXOrv2Le3GPzHKkQ5eDW+jOIKOeuFrq5lhrMSTKwJ
UcZ7h0E6Ru018nGPaIKz9GkYXY6sJVITu9GxvyYcYmPH5uNhlOXCCu16MBtQBBUT
O1/AP74vakRN7rSkGZ3QYRK5f6A792AeC6KaTRP082nlBhOMg5j5bmWRO+sPTJRc
zUJhkj0fEReceeJqZ2XpTbgUnjHOHmbn21ZLpycYXF9ZZeEVGRj87zIuQ8zS0S4j
BKzuBBjrJOqCctRT7LZszHI1bHaTP24BJQ4fYmH8OQNBKvCA8+YlR8uAzc/dzx8m
hJOMtw6X2EJtF2kzn8XyzhoffNATibDQPJ68f/+pMVMchkUl0ovk55rd88995v58
AYQe0766NYvmjGyeW8gyVWcyimQkg9U5rhvev7GdzRhXVvXQmAEw/zyqa0k6K1Nk
QQHNNTgkRv0VFVhbvBL7RS/42vmZlZdhfeYaFHbdLMTq+W9K9Dj24Jt1jKJwHxOj
bwpfsgkShZm4/YpSXCNiOO+ktx0+gWIRdiXgrijp94KjzgLtPRGcVx8YNT9eX8lP
nJ56BvS9SRwinPznJvDYNECnWe8a9Dnqob44wI7+7+C1n+jlEtjqUKnau9qQ6lAp
QthDFO8GqPAhkPh5kD27f+7TpXMZ4bEmCv8mzN4xbvfYxAGCpKs3WTYP9Zc4Ik4e
byYz+GQr1Dfs0TS+Ad6tT4YfFl4M65cLBaaxWrX7rEc32+6pED3talgCIYua+dUh
nTH/C2Xw7eKQdKKywNmjPeumey8RSL3kaKccmC0I5Sg9ErPibqy2ldSQ3QR2gD80
H9E/iXUgmQrQkiiSPFnOukd0G3ERinTB9G+MJ73T9W63vWyAnZVzzBbrnRrt0gta
1/YuUCl5DJQQioN+mS0PlrpIIdE5iG9DZ7Ui9qo3AMgSZim/hiRjX2Mi1s9dg49C
N3EVwQzKIc+4F62u2Wpgm83lNCTMIZ7tWq+oXvqxZOW2QwbuDOkJbTBVZlqKDa98
RoNrhWvDqxXwOZdru+YOaT0P8qKhGYBgiCQU2RLW8HxFlbilFwWyeUKRE7EzN37X
gj6hWIvrjyAyhUeGpqKysszEwXB4AEgakSlJbnH59dKBif1aVnrpwRCkivyN7TMf
SztwBHdUvE4kfzHaTqWs0g0RCcqjiToPCopWqpgmij3kJKFwU7I/19JagNynbTDV
yvWkBVjFsaLYD9VF5yQQ33SDbWojqHW3yvMflBKbkW10qQS8z32cAzys30Wbu2ca
DyXR7+EWDvWzuq/o9/gXSMR2IOrbK0pErBwcw3t9CXWpgDBE9IPI3UABkp+3Qig8
UrRAuLKI4MPy2Kxv4mUi8tjX+G6Y9GSG7G09VJfqw4vsM58FTYFHGI7tEeRjHB5T
JJ1rYYJPeZXDaOsYDUKNNepc4TXrQIzTpXPs4YXdxiT70qpj122ON/VMRFI1FoyS
15euqddWljOk+1MdJ7S0aqlKseHVC3eLoDCjc7xCpigE2XOYPmvMTrvGbQSl7hJg
LQrV2LIzy0JI3X1/i176AAWdyZfoFdQ6wKn7rMW7xo1Xmqf1V42QMN5jgObae4fe
wgEfurGkY1FCPHCJFcMIWHRyj935EPWczuWnUOpBLl6Jc7Crqh7d7cgtY/7r+FvC
LqFCiVSjq8sFz7sotRV28bykjj6utBKLu7YqXnumXfOtufPf4zpF4gsvMcguW/LR
s9tPhFjNfMTGxn4OjWArGG5U4TnshoMrYVEowfzevppP++mKAIfmduVBjshboE/G
IVHgNJEAy08Z3N44QeKvSIY33gSSgngQPJHF9UO5JHJ0pTn/FZj3nBfWYnyKbS8R
MjnJ6QvbSNQt29z4cm6Fq/O0+v0pwGNDPQviUDEQdeNaF3/w/xTgY8P809pd1z6L
M4mvF1MJxQZA5wDVvOT1Rj5aHG9wkdcwz6qRmON6ztU1jLY26FDpRZ0KtYdVgqAk
5nuQfjSH7at6e8GjX7vEGy/uVaMNrxa5hqVwQU/dScb+cqU5HVW4AKH0hjBArFhQ
vVX93fQ+dYG0fzkhdfDvcI/6mbVn2g3vLV+Q9/PVcAw6WUrnA5VfeztKZap54rjS
bxivLA6Sr2d+9BhZJZbqDzHd+TRsVhye7g2cgLCmbg0x500ts+6cr43XBu9OfdYG
ZQvR1kTvg1Jou25ml8jpO8pouAt4svqzzsS+PhjyGcs5ZJM5XsG/ir7W/WZjamS/
FewPN+HaZgTa/H5Gmvp+GFrvTH+0d3dm+PXa+XdYr8yL8XR9BmhSA9VW3v3xsF+g
2CRFWgrZPFvHIsB2GIpIarfqpnKlFzuKyt1LVgolqR49ru2Kj+9Eqv8/XwbkWjRL
t0+UPnjpfyTSC/cldTad+bTKBdfeTmG5NARa/3X5AnoED0GMk8SGTtv91k4Mv2ye
WyPBi/a4f//0n2S8wEbq+fGX9HYvFcvj9tYUGvS6hQyWHNaeH3MUqeFV2wrBloHg
Y/f9VWXOITyQRnQmP7KHaGg4TVdxWDA7flFp5rELNl3ZSHE4mylVpdi4M4MizPaa
R9hRmMECAo2UCipWQCF7xYGjmaC9HoaQeZV4Fg3Ug7VnfPNedC6/u7C1t42YcyLm
b7CPSsdfP32FShhbaPnrQKPcZWFYXo4hujWhOnBqDhgiT22ef9OFLxtyQKS/XVHV
RBSAQlFUnCngYlhrJ93VwKIM7clSLVFhtip/Kb2mnJBhqiNk+Wy1Psc1czEVfZ6f
2/yZ159Ts7X0RlRgsQLIV6U6N1SFprrsjw6G/ADUP/FdNEzo0OYR+5MYCjbzdH36
2a3TBm7IBaBrxniqOgQ55Poza4teua5ylXQH6l7KwMtlry7G0ua5jjIwDe/UCr1x
yt4YAzk4zJ9Ml0GbZ+oVI84BkBYCwque8pekMSK+HUJaF1j6FeWp/zExjwvdQAar
za3gyCjmAlBCAbDnkX7qriqXRlA7PR8aTJ8ITkUTYyiB3gT3aZLaRV0TTOT+NwFK
4Q0FTieT/KZC7yXGcVWOgCxHnLLWgoYeSuR7oICjW6wHalolcZ1UlY3iREf7BV9p
O453qo6qWfyicgjVdg1Nmr1D7JPi5k7IK3Q6+JRwE90OEZX2uanWjaGz2OcXdppg
j96N5Afmdi/7pjcRJLN8v7Qg9pTOksP3vcdTX/iWU1YpvH3ia3i8juWuYio7uojB
UKMhPq/hju0yP8y7WQtIIvyq2MrGRfTy8fmAvRiOdQsGTkG1w2Umr9FNDj6Z6vv9
rnSEPIA7x0KnpZxuJNic/9Lnjot6CLw6kiQIJZBM7KIT/SEYMrfndrK1spzIOHfl
j8m9NCRkrSkze7M9cyBs6dTdsbAmKig00KuEN9AA50RQRbyvzIKzhWmegEBUa05R
XnMIYPMRqZ3jFQxAWL1EGcHPDOuFq3OXbTunnqGJX+BlXUTylpbvLCZZ6SpPgPRY
JSMUADdoBkiOjQQmx6YzyEzJvqUDmkTEvoFGL54zl8qVqGZxCypU9m1kCnxK2tJO
DCutIGlV893cXM4Sbv5TN0+PvrvZSd2JYLeVxnUTZbiJFLd5yXJR/IChTfBtCmLl
3aFcjW6ro1UuJqY5elf/iBg1sxTJkVU/0lFm36khbBbs25JfmJVPUAlBOsWgpk0+
Hu+bswPFN490JckDR3zuoS15KH8FUlVttufTZmPYHXDCRkQazxXAsSoZm5dzfJbJ
cEtwsziIY4+Y3wyKsHy5SHssA07PYjypLDPnkokjKXOMEk3Chbs1KKKfcyymJpf2
L9RajMogKJm0tPpbmEn8FMZzatx7CUOJbZ5KzZewLflIt/z0zvhzFIi09JBDyOIH
37KdHgZIhSVcAohyO6/Lk6HwJagy1kCkEick8k/QocQJ+6Jlfyv8yGZqAROBV2MO
FAPyqrF56pnvthXUtJF7u2TLSfP6bFbZwEjtDOKLK35JJab4lrfTyOUyl8ERorZe
iM/hmCj1LzQwSdycZppr0hnUHtAdO4R6C+4UpY+wOwKJ6hQt1jnldg5BGHaBcTN4
gRWyq26YrAxWssOCcZfwWzTh6X/Ch5UgvFHJ/hSoitA/MnHSjuO+Sytk+WbY+z8C
HUtH8P+ceiiwIEKw5+I0aWib/eDTsqIY+x0oSdtxXWGY32c9GHVos6KmVY7s1Z0m
lbpY+9+d1soS1GzjW1g9l0YvRRThzlmvLyec0FVYJm51PWj0orMmTu36yVhBBVsQ
nAkNLs2HlyKnGjYfucDx3PCnhItDHpxYvjwMymlum35HHw0Y3zMazmh4YZbf+Exs
AdPnleXNKqoINtLFI9fqH2gw2pM05v0jpKMDVPgDHKr5fbmcBELW0xv+u6OFrEgq
3shqknCEMeleUTF514i8YO6DJ66uR2PGs8Hq1SsQRvILlnWv2ReFpfJ2xrOvKvoc
wOn/YONqze7+U4P/qjD/HhEXplIu3k+A+kk7jqhLLHRXS3WjwLpJHDlbLdGuBz2H
DchBjWth/8XTzawwiU7tXyCh0habs6VFagivCXcFgJLD0hZ+fq/kRf98+XSc8mhe
5Q/DvC0JXczntR8RprsFJsn/SAAMXUXTCHlENhsJa0awxrQ/sDJpVCDpUkSAOlRT
YN4vY9Wqv0y1OHitinTsoeWbPg5g0rcawChBs3FkhQj0XGVp7ZKA5piYked/2Mzp
tfJ6fxje93vEpKuBjBhFHGBibgL86KJuBWnKE2oqMSjKaPTv2JCJnVjlLvrGIhA3
zbPp1swyU94cUshtcSOBNiwDlsiV7sc7ObjSGmi4dOnaaBCy965YEqVvIhhA3nvf
5vvaWpyqS3RpIyuf0l+qHq7SqNjtrmO69wnGftTJ0j+hnqqewo2BtutcwqAwnnhA
tI1rhw4CVEAH2HfgI+lMEhgod5o7ZjHSXFmJZfHGlgEKFPVW1yYlvp9pBtbyI0go
G/AMAJeS01ADXBmxdy60zIigMPNS25akSX+zbrvxj0yUOJOLMCD8bP8kVUy5omgL
MXp7MNzYKcLkU/qyrBURtl6AgBf6RnYubJ/u7cEk2+H0/hC9BIT1V3GARU1yiTpV
5zeWyqQTQ02+LXsk4J0bPkecQSg6BYO/ZQ7NIX87GxqybN4zbVToDF1hEqCF8G2P
ywnMoEWMxv2DjkVdNGLW6aiq43nKt+GKaDjo5aRlkwlGRwtoF1RhGb1x11dKzLZa
yVYs6O8KXwzoe26zQUzom8wcn6U+STc8UdwOWxeCCmfl+DvWwiV02nqJ+WMaGIOL
5wlOfdfYZ9n7E2AtGyuhPSfo0L7/28MwfzCraiIEYNfno4L6ciaWkUPNy1hpDF57
4wm9l/5o0Z9EWWygVB90qMzjSjbt0mcOj4KdXWJoOwLV1SgiwJjchX9c67KSC3g/
sFjnr5DWvPFXrgVce0Z7DE6RPaOiJdWfC5wwg2zp6W55t6F/vUs5lvLZR8htuvp8
IcW444kPLVcAMUSwZJYltJk8sf+XUX2Oe/1Yp6WfwBttPN7zHV7xJCLcYEILhtX2
G2YZZdAWYFOBIw0ZZewXF+k6yInrFhaRMP+14RA/8f2dPmxzlfI/OetObqUi2hTa
/BA5/l8tcsQ/7zmhuIi53wlOjpg7R8Qb8fr7BDo0pzKTmiMjXreU0icKz2q97M0R
gaWRa9kkaxe+JT9e32kG0A2XRHBZAe3j9mBNuHi9abUpRQ5ESAH6f9NX66vZyKCF
hzG9ILkfI2Tr5LW2MsRFpigNcR9S3RuYgDNr/QwuhV/MrIS0oNo7mHOn/uc/YbbE
/QL6iG7NoChS51So39QygrhhtS4FYC+9w+5tEUdlqNV7JubIqdaG4AU6LM0jjeoQ
o1fZtnoyRESclZ8C1tCpoQ+4VmNavWQ5mJ1R86DwHZwD8ocKBnpspEAoUmqr54Zk
tD3zCHMdUcLgMzP3saXIgwirI2aBXyNJbtFwK7LJWTAl8pLkaUrjs72ZTLflWw2R
ygQmYTcsCCpPXR5TBY2h/0eZ7DShQbwQbUu/1LC8DWdmOmd403W8klfOeQ9bYflU
Qc7wBBYjQBUQSzKPX2QuwDKb1ryUjbBCgfmjpTflt4ZxTdr2mFmM2CyCHnyO8nqo
O8o4UcIIsczrZ7HtzrPAXAclGEUDH2wcXYYYNDSyKGEwQv6REn/qPO+rJMo7JrZS
/ueWddi57kkJ7T5b0JiUq706qnhad6NEBCy9p2Xu5SH6cQKDEasyAiQiSfct8ch8
44JxbtBYzYSZBuA/jSen9qD1FnWjhwmE98mKO936BB11TVWw9jRA+z5pbsHPCdUP
ShGYxtTjPxVbRALpKCdswcNCJiukN57qYDg8cbYg3X5jqFFUAAH6YxU3Zwhqw2Xk
KmC+ddNa/c9K/zYIkNS0CmzD4y+sHEuxIo2uUGPh7SDRq4kkQ+P9xfj8A47k4eyP
MaK9TN5xEMIBwVLXhHnWhkVvtDNCXhkXmgQpCN583nfmn1pNEDdwvkluH+SY5bdW
jEUdnEqOUvJyVnK9LsQh7rYlzkNV+XO17pDdUTLXrZTFwWBVuT+TZRQkGH0kp4QP
RxayMUqZk1lOr92tR/776VpEkSm862WHBhSUw/nT3EJHaYfMeoa0JdGXCloCVFcf
jomeXaDYeL2FoDg5fNxxcltVf3SVd9tXsp/4uGhT1PctRZvKFwaSfAshfE7eT6zK
A6jmzHIPg9rq397yi9dcvZzcPm+fWAmpfON7DOsOGQN/oA5PAwZZQ6VV4qjO5Vq4
gsN5jS4a96Zaja6jHw9iyi0xIVJfX0sywKdAgjp+14+Nt3XRSfvkozhGVCF2VcS9
8HX0+iUcJ1wo0dK0Yl6LneY4oGb4ehkdP7NP1lPeqeMFf2Y9gf1DqfJtkHtB2n/C
X1aRTqxfW2QiYWiZSHyxACPNDlTrj+7o4lflBS4q+7uI0YDFTbkza9AqV4LP5VsV
deEQF6WAyYBL7iB0ygslf5Xf2GgZ0BUjfrWsTUvycn6fZPCNCjpVeOPw50cgvS/K
ez+oTZQVLOvZOU15WO5ezt3oRYZGZ4T9jlT5Uor5hq02h6EpFOXY4hy0RPuYJ0Ji
hshcKcCsSv9dlZicRxlPEK+QtaZylMgkRPuxNxuCA6j7NQDpjJezyxoDNFF/p+tX
yrabKBsff8uDC7z/eCvZzADnfGEh0WG2MlBKUjwzctX64ckI1LM0W4/AcI+Njhgk
qN2do7gopVrNNyh64lXjTy5CeQaa2HI5bmbMeM+4oz3uCDEtrjqmqWYCPGTNwTR7
ZP7tcNctxQBLBPPmcmfHoRn/+LI1KRxZq2CZzBVuPZymb+RghqRNE346R5SdGeO1
RrLyf0UuWN+z7vR/x8xlPUxKe8hYnMaNVO9W8OCXIOgSiutu+4C1qa0VYQ4SLtTP
8KteyAAEsqNxuCweCZ7rfjMW21VmNe/Pe/izeJXZpdybUF3MO/b+0XDpGBpcMI+Q
7wDBytWOAwEHuuL9nYlo6DZ2GkAExW488wiPZZPn7vJdat3942WFu/T3Alz7Ue50
RVvZ4SFTHiuvVzH4Zkmvuc8r/4dhHRfyvUbyZljskxTNcd5cQTFA0324hFomQQfr
dd1OLiQrkL8Y9iYUXRShexwdbkszrHK8ONz5jFT7QAC/x72oArOwqstZuEnjqqb2
I/hFDHnRWxbXGYADLWLm9U4Us+dovq0cQAoB4zHVRjv53+83uwAGlto9SsItVdMd
KgeDmAmA6XKyT66EgiIsY0u9jKPo5OKoKc+b2fnmE+PMbzYbF5qt9qM8DNGyvb7a
KB68zI4UEviDtuz7Sephe/Oecvy0Y/z2s9/Ml4EkxRzVJO+Dj1Z53ejNrHri7nCX
ymydNbMcEixHGOqIi+84i9hdkKZB98IZv8chLxlRS5/eahLIfm/LNjslzEQNwu6T
DwCPIU2dAcqVrkaSQRzoIKgA0D53KyZhDfWnkbyKi+G1x04ngXz6gaZg2zZo/8OM
00C6cSgXhYfSkg1jOGUV1kHdDLy4PocS0MSw4UskU7fJfZEZjPbPiWJLLb+2DCRs
cfbzLAXtB8ZCPaITg9TMi5JvHu15zASHtnPyLyp50/xC39ZxwVPi655NjDN1GzFA
jETZBBUpnEwCax7hBZzsO104ev66uUOkWodIG2qOBPIS31G60RoJXMTq6Mm7Ri48
yV7wqgL2GN1cqGiky/JhxYpJ2NJ0z5TebtDd2zPMcmOm5F/+z+EWKz4gOIZf3alS
WjahfB/v62VrrKIHeAcSZCH2OeoScA6DxfJlOeEtXJA1amWsP2vKhZ5zCze5AhPy
jQmaauwtOuzJfkeR0wzNOMLrINOqb+/nPUSu/hnd+MlcLoH5yHdzQxGnANerH1Xm
U0loVWNgQBHStDzjso4i2eZhK3Rf9hUdSqIEWKI6q7XSXjfZai3t+ngdpdUDegkN
ACrRoyNZ7+i+nCMPeUhgxFqUFM6QGNQcrHQk2dP5TzJquqY961GlSVNJ2LSuDR87
CLc4qrCijk8hE3vFhqrGSihRch8bnBHVaUSMbNzenqbNTaN3HhClue5Wl3iQewQ4
qx7aTg9CkrjspEfkJOt9HaqjFl/CXSRAvPucew+7LTCBb0cPvKg+7kM7YSwQPj+G
HMI8gBFms7tuMR52wYRHgRx0AOS8xxrHNeFpxu+6SF8mBb8cyvhxeWBa05pW6cSP
V+2rV+3gYsN6O+9D9IpBKh74rwDR8d+qWd55ZXMOeZU0RNI1BdYforBc9SbOErVb
fnmEzi1gmALigrZKCpiGK2gVDM4Kq6t1bdIGNA9rsr3zrQ/4tMdepur0zRtcefDN
oBVQ5COoiL8Mk4+qXR7mrRJUn9y+4agtPlAU6keId9Novq4SiJk4NBlU28AtTrA5
FJG6rNjZBVM85viEybYWM85H52+fxLMlgLnBIAwtQdl8D4cZWkOXkCOPqg4b6TvP
S4BpziuOTmVGsc7TvXhKqCImENYWfKMTxS7Cozpa2BKLudky1XkYadtMMDUkM/Jl
uoIrlF6mC7412YSTYyvLVfKkEBPyhUJD+//GC0nvQ7tgU1up9PSUBQUOxmQtSG8N
5mtuXZcUHIj07pp8lu/pq/U+ZxLyDsEkFrdxiSVVN57OODRdzb6+BvGLyeLCmEek
rc5HNAQG3KZ/tgB1pAGmAQ5Strr949knugAbaJAzI8RhXRYQ/6+IftXiL98bSFo7
HCqRHTqUiwsHTlXQiYDjL6AEHYneIQZnmnsfUzQnntUGUZtUsT1FS18P5Qc8pj+G
0+YVrKeEsDiOWftNBKCsScI60bc/BUQ1/NyoS7iW4XC4wE+pEtZQ3ONNCjTbZYJz
+xgGlNuASgvyePbO1bKIXuDSNqEFf6PfSYkcMStuOvzeqIcnw68BR62XlHGLnDeA
Q7FfXqjaRJulGczHGDKD6ouqQZ5pJwJy1tzmTDUWdqCbXxeX1J7Q4hAt+3AQl7AH
kz7paUYDZQGFCq7MjCmuy5VDG3vHA5PiFt6hMAtwDCyEMoCveaNa0VTfz3P1jUkL
FipkNGVAuCgDFJoaOhV8g+TbCqBwSk8jJ7uw1z86Nycg28hRO04DHs4OOfEqmiT0
/LsGvqot6BKI8KVXSKUhiJ84u5OPsqmHmTR6IWEcfrmsh6u+0jxypyOgA/aKCyx9
juNBqv7n10Cs6p2oCG3jZpS+6h/9xFd/kgwUnCD5Unkk9phL1BpiJmlr983r3jVz
fraL+W7tFQ7lWFy1LOrMBU7i50r24mG22Mhk2nvWZPIvbGJYz+QNRZasuo4Vx6JG
libANCiH9NTYSX1cRFEV4UyAl6Y44ZQoq3sD0foGkqG5U06/Uf+huO6tU+J4BXpC
HVxThwWntGoxVYBkxC6oyeot6VJ8GSGv5DbL4Ww0+w1+MIyNDfBSyiPgyH8HoGRD
DZMzMochc6Q9qBFdztHdEmKoCrHuUPVZwezqyc323yhsUB66z7C7Syel+0bczg+y
Mwt8T5oXI6P8Dn6OW9pvph4Is3DNzMytcmRTfHShzbXWH5qaWyJ3dK/BK1s5DQrg
F4ell0OtlmdF2yYNSi27zKY6F1Ob3nWKcfH/v50KuLk1mUcVMqOFfAsXvbRqNPzg
PnZZVSQAzTeWHPvQPMjRLSuakI30vdiknhVlI980tAyQva8Tu/dRu/+Dd5xciy0W
sNigPI0Z+aA4xuPKogbnGCsm7cuiph081+gMaMsMJqNIhdlI7SSxTNVDrp7gaxCp
z+B7h/ZMzmIAA8yjJeZvl3ghMQjJlyUEYBQTlVHcWYoG+gUxcPZRoDC7u2G5353X
LtFtzqIneje9MApPu2w0IslMzuoRO1chWGR8rcInaxMYS2au3KDeBcZ+prjD6o+I
P9K7VVv0IoIxISzU7Az5x6akz59/P41lVpD29RmixwMghWY3YxhTEvDYcCk5mBA0
ZcUg7T6WIKEAujzXCW26tU1ZXSqNQbT5kSbV6/krVsZiPPwG6yGBnW31WUhRSqwH
EuvdBM4uMWA9owDVsr6kI0rzPa+LUNSvmtMnyl99Jm0Jen6I35ujFWI5XLSy553v
E9yXv0mO1itZf5npluHuSvwpYqS+LeJjHtC+mafnIFdHLotbgknZ15mm5zEVuF+o
eD7q3FJ5ulq7XWnjuURvo04HXYSMSEQkhTmaleeo8M9xu/lOodtavY0NQ9oBlYA8
r3RXNHbthGz1ncjVnIlyzxWjoEsIZzY28GSkXdpCQmwmRkxiiwz9Sy9NBhBw+P72
3N8OxozDcejnnKOD3ONzAFmzJqHVk8IP25Ge1kAAXB3j8lYylS6xPeu2UcYwN3bM
rG4rbOMWQ+AGm4VAttL0T8F2aPI4TbHReDUdlyw+8iHzzCH6Yb9tOCzSf6W2sO9s
JeetrGaXNFLebJjQ93ihvjmfiXIjLe+zzmva19/ZplezFsiLieZRx0AkTKShTSY0
hHTzDxHGtVq82QEmDSmgOUq8iNFhUcInlEcSAiVxrzE95BGGrVyBvDoZjXlcWmBq
FUXwrr7v8+8mUIkI8S4eoWvmI3wqHIfF4GTW5w6MvOYvVBMcllLk81N36r0FyIjx
jaujUC/iK4yqr1iiVTprorMYtduYICK6p6yq/IxSXFH5GLgNRubKxHBN//5VHqSZ
bRakcyN6KImaJc95AxaDOGJfCLhhsnLO7NQFWQoudb4nuHC7c3rD9ttrzOPUiYIm
qXLuszAH6AG0ALL1jjrONUo79TVYK6Z8DZLaEBkiTo5MubQUDBWW0rFOK6LNnt3a
nCfhmXMuHo3d5HfKpIwOhLjuxXURF45IH1gV/70c0baHQCd4dmoDAURG0oGF7AUL
vA9TD3DolaWjn+h8UXDO+DSbxo6AJCI0KaemmbuYnJ+XOCU+TAHcA7ApLx174Q1L
YKxoHEPL8yc/iiVIBYVztpr4VLacD4Y9BtI131vm6ZToL7T6LOr5WYfkTJY46ZDa
yqSorh69RLzCSc+J6hHVPF/kW7rF7G8rmmGBrTomegPMgwxHywR/Ypd+qyDGoP0w
Bi7BOTESCBOQlITZ6dvtQrD/VheClMEcmtct6zAMy5PQZ2v6GJ8ydZ0ga9N6s4Lz
dd/Wv9lMNNQywuwPWldwlPvMYDN6zWlZITKsiqEhJnBDQZAMDYTGtXQ4Y19U34Dt
lbOj9HOP0MDbzdgeYJQH+t8bJpG2ppPqJaKdYdhR2qHKpGSxHyCQ55yuYaMVu7zw
eDgLCv+zNDra5dDmhf1DjrNaf2QeZobSPgwfDlBBkQlfm/P8BqSLAy82jmfe2zPa
KSOl3PfQLoyLsBUoak/eEmSdXCfkCMoz2VLbwm+LiyCza0mip9DXxDqOJtj/LUsS
001p+mgvMF51/v0xnppsL7CwtLzKdTQS1CkOYkeGITQvawhBOQHc9RU27rlywmTY
PtMUb58+1bAPqfXKaMBSHa4ndX8F9SNkDgfHZy+il9oWnSSjenZD3G9tznncMZjF
PynM3hL+F5ubXwSkyy4ZVgslD98jMQKT5jv66ndnFnddbNvW854bXmR481nO8foL
d/3ah5CD2G82d33l4IaI3Gq0b+OIseEUsM03hazrJQu3TveADoshtV+iL3vF7Yup
J2TBaL/Nci5+BA5oAKsf/k1nCKd3dbsCdoSzSLbgjn5GyWrWZYA14czDivQy15h6
PKbSnKRvQgRCs9Gt16NDNpBIRDRHP5Vxy6YgU+r/XQc4S9BCuvGE9V1f6YLa0+ea
xf45c0Tvi5fSZslOswjgFCXTqlXe2wdeS2vCNqLTyxDOoYOxHuhPGYl2DCRgvcvy
oJLEsWOww+7gPa+CODmBF+ja8sPd887uFX2/k8G1xJJCARcSEJdjPe1dMgEqmpaD
IupybytOPrGI8UFWdmYeRs6D0e0J7rqRKAbd3Ml1QE/a68z2lp0JSM6yN81FsOzM
2EBpidJumH+KxtV0olOanhDVy+4TjDtw1FDkISJz9CmxPw08i8tq5aQUex97IGa0
jCzqR0GTWmeDauvbI5YuGLqkb4wSb5BMvG3N0GTMfA/eh+BPpjHlkDfcLbKx7nev
pbF3NNcWAAvLxR/w77SHmgnXs5ktmfcrONn+kg3xvgVrPbw77migD0m1gDuwpqzx
DBnIBQn5eb64/Z12plLg6sLCoIycSt8Jod+wZXnKfN1Re3Ogc9axg5Jq1XoZ87ez
KtnUkGVhjl2WzhJgZzU5Mrllxhctm3qVFG+KRjw1XZ0o9XdNQdI8W9qvl8s6+u3h
aQAyquoia6xGOUdJkErejiAYXrv186jE1B2k9O5bL7D30t8cWwKetG7RFtTU7vN9
Jmu+ulUXokaQ+Sx8fKFr2tX2/+dH+RegYgnQ6EdV81sLZ/JQjOetdCfaQNef2LfY
gDJAEBVGbnSdMRUa2nyXZEh4Hh0JaALpm+zBJU7HL1/uaiUddfsYA3WQhtdWhQhf
0ezm+jKSTfRl21GkUuChkyiTp1f46FlpsbB6ZDOvnKoLX22dOrmZZo30NvRM+gwp
MMSgdMn3U3YhlGbku0xmMyEGss7Um7IvXHzcZHd48Zpd4X5DsdClQe9ZM2j/p+19
AHJ/EcLHVHdQY7Za2pOTNiV1ys38l7NU413r+hP0+HcNIn6J2Qx66XRBPMQtTX5T
aCNQN9dZEWl2pfWmKzEXCvPPFgCnYhVXmtfTzz1+aIwZl6qvFh0UTYqiJtRLh/O1
ic25eVqJeARM8xv/9iGz0gEI+3UTlatPbkl70e7/s447Ivl8+RI/x/Yx1aemmYKq
NV2An0aHQduNdC3zI8n1DPPJtHmT+rdSGkBgh8dPj6cJZYRKm6PaRQJaExweM0k+
vkrNpbWnhzjr7Mm8PnDTnfbv+AnxtQtMD7pZyE0L2gnqTL+kgCogZAveWQUTFhiC
dQPolAWSM0D42emQDf+y/xDa2SoRsFV9XtdomFerrJZOXMSaAiCeTj4s8ZxiAWqb
B30lpThjsDvt9/6TolvO5phz5N0SymdlF5SH6mv7VFvVTW14R+zdK/vKXIzWMhY2
BRqA5oC16NAzUFWj3HstNct0C39NvvLrbyDl37SbkCcnpNbwtK9eybLo20q7+bR5
5HUyQvLZ93dZ/embIcOYcjwiED7Ul5+ScCqtWIJaqcla5jJrk3HVwaHSd8cln1Uy
c9R4txjlvKvgFZAbAngW1oGRjOSaFpG1hMjpeN47dz6nIsQHS45zHz1O8uLvTt44
oWcHCmxX8Z4JO4BJjXMitxqHV8k/nlMw/G8SSCE/DZcGZ/KLk25PVg95LAaOjL3r
LMJuoZ5rRF/02YGxaiIfGkwJMG8P1ScntJNqBDD+B9nmMrls69zd01oGNKRmVRdC
HKWVGwtq+64vmO3C7ZbdwrybPmPVsh7u+VlCz83bnzAg7y4aSre+K9ctHfj1HXIw
a8MHOKx1KgsgSgZDbnOWHhLiMgHa6SPueRxjVDo327/5o0TyWsMn+SvLZ3r7shiu
n6K5bsEl0zXVWTHw2ww8h9Ky4udusZUHH9pwZJwq7ocq+HxqXPRBXNYjZqSENUxX
C52XU3Wm584/qJhcneobg00i+mVJpbRgfGMC3JKJ2QWsw3oMT7YXxEhDjVYH6RXI
joWEKu66n0z09aH/gxsKWc0nUJlqzFvIC3sNbMzjQO5d/bAr1mglu+Veco+dyXny
qA+R2CL1znMGbLxA2SYNDnZwMQy+BHLjc6tDhKj9ffDDvhcS67BUMnmrwpnVE/ko
W7XTi0KU0f2e93yjfXSU5Xb8uGvHtxbJn7swtpnP+8kT5XuEkrPHOfX2PfwY2Kxh
zgjdfu0Z13cyWBBbW1r7WNIV9CwT/qO7sU0Jr+yow8GGN0mGrXnHATF/MVDc/9+d
mqie+th4sYQD2Hp+AawF7A1CKhRZl6Ga98Ed4vfBG6Pn66mY3JMw/96fe3M+29iV
NDI7/XtZEsj62xcrgyHitziugQn/I/DytLGpdu7PxuItCqn7NmRAZI9R+4Ki7Y3L
hU3jYiIm2aWhx4JOdy47S3N8KmsrijeqfTTjCJX0ZQ7Wy/MU30Gnw+U6JzILVexK
XfAB0m+Nh4xtWhRM8cboabpPtSqqW1hlJ5SBuAD+zjslZXSmCom9GvRkIQc2uQQF
Psu/ul+HJY4f/lSkxIzc+SDUY/cikBE3pyESZ8mDKO08DCYx7aHq2cz1LNN7jY34
DQXXPGIWBALRyMVCYFp17/MkSZCVwvwpLarnCVummYY1e1k3s/BVD8yslcNbLkWU
kfjNky66GuOn5KAXggOjZll2wsSAsTZONl5HCxLSemRCeaPuUnXFLgks5MC7y0P4
f/qqfgeElpbDSeCG5yEpnDXskaq+AJvNIQ3B9xXb8Xs74idOT0NtdY4p52HAPcR5
HFExnKJH297vFTn3HYjDidp60Aq80AASRZRUrgFbVxU+RCXNixZB7hVHVTHv2/Jc
eJZ/sB8RbqSk4p9iOq4oh88Neq3hFPw06TOKE6UP5kUslfUAr2nmx+o+8+/WaAyn
PcFDCJFGkHvlSAbiGVq4M7UOCmCEVTEzHMP8zzxgjVZkOR5wrBDQwuOHdSOKxdhB
TkzscsGA45Kx8T8NKto1/4suVnmFT0dHB3DYWxm7P1PoxjqM74KW4NpSHK6Byj7j
dDnX6prmp3D6f+Bl+sfjmWBPiAuP/+hwkHMbfsZH7DbTeOi2NfSjt/ql6fIcdYJD
VxS/c9ahkdg0rLHssJ2oSeZQUGqvg8hQZR+njaBLgz6QZVh+UxGoMX3zrXFXJ1Om
o/sgi2HJ3AHdcBn5GBv5frQan/216kICwxZDy9WREusYNNzXH4vSZEp8kgnuBIiS
q+iEz1f2Zm4kEtLB2WYezlqVqd2eIzp1uXTvoThLAQuD8Nyg++B05SGlqSGRLrZQ
n1bJluWYzsWnbHmXxjJ1TZsps5h0AWLilnZBYxSqFyoJkeC4tf3qI1cn7b+SNlw7
vNoL6/UYYcQXWv8vY6Oky2fcSA0IwMpHLtWk5PHRajR0reBPxEhoFvNDM3B/oNgA
jJhjRId3OazpCuxMtmNFb+XikKcDh5JFsyR8O+eh//T8tnUok3akinTO//YoEZLt
2ttM2tTWYJcE5Hi6+eLfTKZo7IJPdrRTkREyWQXgnqpWO7swATkNQRIu54cMvMfe
aQrWO6YVWE7tatzCsPbDEmGK7qsIl04eic8AUteojPfhjweakrnuvusW2E1xdREq
sGsO9w9hCgWq8xs36NgKH/5pmVrHs/ohlwI3DbKx51PMZ9x+IDM5wNFY8j7Mid5z
OVwkGDKXzbHcLnXrJ10XfIlgSnrfHCbCSCuv4EWjX0GgWhAU909/Nd67eK1i1TOi
DlJs3goOyjh/v6Kc4rGXKWG4YprsK/1+fu8ZSkEaUti1SdLGA8AxqE6hcJ4Fegfj
+ZEqTk0JVyCl1oQbjK2wOYr8bxha5ZQBlwvkx45BTubygKzMiwgUqQBM2vQo51iD
ivThaSRxhYuKkPKlRlnJkx5DmyQtGStrjYFY24bTaf19R+V/7HmtIE2gqcfHM74d
DcZnamGaEADckmnChzs5sP14oGEKw7cDklkJVS7UqaiGyE0OPHBX3ixVBJnUuUvE
eXI8yjoG2emrEYsFAgMqPd6xWe10PJaA/AIObBJu6M/NtMDB9mFqirY3gny337H7
LSt9VRyDU+rARHkHIQgIY8gmvklHaoiLvYiVhQF+KyM9GbVV87Y3EvMCXDCepB6S
YboOHKZatiVpvNJZP4wE68+D986ybIQifiJq7JfsDfw9Ok0wpv5WeLplOBd0KxSy
EZJxCUNmOBcQbQZ3qDzPdBvTo8map7Z6tr99e6yf2lbMPBk9HV2AfPT8Yy/gqHCR
Cu0i4SFOjnIG6BJfO7+lg/oHwzC+YEvdREUjMdfgoSYz9R8YxMxfJJZQ53AZObjx
+RBbhqqkfOsuWJ34rDJnlOVAC6NqMhozXc5o+MxJs7dJhHjXXPwEzjfKKprJk9mq
0EHM/MiiMvKP0+Wr6yZzPEA88qhp5AiXCFn9TuMiRUT/yBlsvRhoXkr2spHNJFwG
Qu6CTozcPgiiV+2o1rJRMppqF80dlMJsYVobGKZzJHO+0YJewKEAs/ByRR47KPG5
R/gb3AsXz+wJVUBju5qbL4lCRcgVoskAZEIXr9i0Cl3YqwQg4p49rX2fZv9uXerY
jJ6GzxTq6m/4IvkxqXIbYBIZNu5oF+COdMtLw61wk1ga5kUQb/QYuV9XQOj8W+kW
xnZpMZJRNXzWwisjJ59Lf2KU24eiKVP7aeryK4wrdjB1fNW4/iyC7ToaDuOS1eMt
av7g8bDV+nzMu3pznTi3pdq2XFqR+ojWU5b/MSYtNj6HSMAhUua/CyW/um3WVDQ1
wGfKh6GPoJseqvDk3AsCch39Q2m/1o35GWV9Vpxey0y7Kct79Dme/zw3DoO7JZmA
1eMA4E9zpJZk7YKor5htM177zH9vD+IcMCxhV8uNJXDGh+62sDBflXqLG5caDmZ0
ynC2KOF1xaE9a0ORw0/cMtq3pPNnnHbqkbN6aBfyyLzZigFREjj7DhITB7bDHXGR
S8SgtsPtICbWJGZNUiVTQzn6POydmVRuaYCvrt2Yq/bzsy4XbfnQ1dTwnd2pAWzt
9RuXNsRoXj3GJq8a91qcIQLd0U6sopDIuhsHlLH5x22iey7XOGTBTDxnRD/yEW5P
3dxbcIuewHmQbsm2mVXTIKntXfyJZBMd+4uoo3oKFZJdr57a0cLIeSdsnedGJ60v
0O5AohsEQUmDYZhHj4BB6LauHQIVhwjRm8I1ieUfiR0uFN5VIWSwXoORyGZ8K5m4
ZUwi9FLtVphnLumCfwwZ1o8K2IhiYHwPHD+BxtzdWzs/KWsutel50AVIqyKMu9KK
6qZ4wldyA0/WrOFFwRlrVJYK5W0qmLCMpUuAXwkEL3NG4XtClnUE1bP5In5UE0/C
cVIBkL/NowCVsSpP+mATP+84em9dC0wuoINx7RJrt9zr03IvpzBTim+THkjFsx5e
ERjLEhT9okDcQm7yGiIJ8gPSrJMGWlc1H26vmcbmn3H+W+JII5LoJuKq1/+Ujucv
c0NUYwf+tcKOKpYHIcnSKKmpF8IxGC01htPkFVaUiqfNimda1dIf/0bu/vVBH8cT
DxnjmANZW4g5w/XeAsDcoBk09pBnXcnBSUshRRV9Paz+beT4tAGoV9Ot0XwmH4JA
8y6LV2nA7q5PaG6OSTRrrAJk3RGetsapGK9WaOtKWK+y22tvUfS3WZEM+hMEI3aM
Q3pK6VI+ITRkdOmTyOTvtPxYSPVgdIZtuVb0fCjiVijq7CN8+aDBe+Uy3yB2Rxdc
xEzfxBMcetxEKfvWqQM+J/ELNN/hoDkmaR/vGS2goy0ebKzgv9UPzKAcJrO3pgAC
yd81Id/bbxvStkyHnJ5fqgzL1o0e+TI2JLCHXSbG62UzHohrgubFtHrJTyyT9tuj
ki5HXuCFpFH81QUbZP2faJvRyZNeL9S1QK/PUsN2H/0lALdyDgHNA8tGozuf/yMh
O9RPHNPPJfVbjN53F2674qI/ae/ngLboC0pinq/nQUy7iAXMrMzY+3jQPkVHYLjC
xEzdP3tNqQsItU/09QO+lTDuFKe5u3wUUMsYYlj3WecErL3vyDPan37EufAMDzRN
EWO2zdYIUFC16L8uzT+qeCUjL1taz3JN2+jDX8K4MZkzS5PuQ93qOgkXBvtbabof
bFc7qM6cpBNPHKmiAidt+VHwRTaa5HtdgFERowefhvYyOck2DHeN8edNJerFpvFc
/QBo/oCkYutxCVVH8usJ1Z0M4w9DuJ+mO+IzoJjq4pwiFdiSIL+qTB5m6czpoKIR
tioZMJJMM9xYy5BPWx02P7W8Ros1d/mmY2CNW2bJLdcD15afXazwRYw9HRC+35DT
S8qV8qY6ZF1OwpNAS7XzLDfisncKlplXCt9E61PJLinIOvRBmwqSEHrNNRKB9aBW
z41pRXTnOHh9Heq7qVF0T8XUHSwbwlVqtBqA5NQvybilp3eRIHx35dk4xOV5a43t
l6ih5gTOkEhkv4aXYGLI/jDL93gTu6SzHTx6C7DAKt00LEXk5VdfGdsBulK8einl
4FZxoVTfGiwlvFULxdfmWNPbb8qBueSHm0SYMp3WmL6TQR47Ksph29jrssvdOs3I
5T3TlmmiYo0kIAFvdyFMa80N4if8zRdSPZNhaCQLwZXhREd7z8ZvyM6NQD4q7TN+
fGFlzHthEqKV/16AYD1TwW7rLmIP4fbc7sHw4tIXKjoT7hJKThYJQvoWVYC77ESf
sltSzfEL6qQM4y1Nlx34/OEoimSUkZ1WjjE8/iyB6nFMUCk2DnElVuSFpl0MufF9
HyybOSXDf7O9nInfjqP6ZVk3FFECk7ioN0ZNbyK6K/oETbF4yPYG7/+IcpcdU7xU
ybJ1q5gWk6CoZc4r9ktkGHeXTX9Rpa6whLatNYM/pijjD48ySKufkkDBShGsF6Ay
9M0EOr+Jupe0EnC+uhpwzmW37u4v0Jgzfw1WlKaap+79PVxAcEDep0AxAoqX30YZ
sWEn4j6cutBKhHRtFEqDILayYpM6qGsXmPgD0PXs9mWpWTtms9jKiA5mtOxe20wA
KBgngRB44UWhg8FPjWrumBDlYZnOhE0Gw6uG/4hX0taQBPmABqCTg3pDIavk61ho
Boea4VYYIQ0N5bWR+ReB8/34QBGw1zVd9KzL6/ex6W10/yMFaEi8sd8twp+wVaCd
zcw0jLgQUNKR/FEcqYHQq1XPLsBLJOjAx34fuBIYoexd2kUfoFC4RNOyoq6DElvb
S1XXIUWgqKZEBjTIEQjh5IaXIlzQdTQpNMqSvq3PJ2z93SirZxaMDpI1dvLzcvll
PBvtEHrRf88sqHEt0DLm/Idik38j0IzRdE9pbSo4D4rTpWqsf+T40KVzQaNMCPbe
9qXOE9WClVy3boQqrNwS+VKRY7uYwNLI3dv7RvpU/fCOcKCvYE4jyy5EdV2CHBKk
z94fyPit8DzHDRGaJ6hNVHpjuMvA8lK6ReM0ddPwqAx9quTaXf1yuJjIWtBa2V1G
/GzcnrX/NilSi8Q+ZF7fV/tICOHcX7zeBq30llNuj4XPYfmN2bPXguSqAA6S4oIN
oNZrv0harEEXSG/weKskyXBnq4N6ATsSFx4TawG5RiNk8ynKLJTCFVY/Xra+XDWt
daixK8NAkFviFrQPmtFF/Ye+Bu482ffct0mjgB0Za5AA2BMmUzurkNNPR8W/RdGL
jXamrSrrz2FUPC22m3f3GTaHibD77J+0i58saMwN3eYA7TO67QZBFL0lpVgcllvX
4x2bGmPnv1U45Gmm4ILiSRGNYYzKmzxqzPM2vDRxWbtMe09iw3N29HYB0wzK6se+
gFzdlWIRw9G/wKc99XhPs5DBs5aI7ob4GNKMfcQk5d2OuiPjxMxNNjNFMCgeP+hb
4bXI0shtU22raAQgK7KwdQlEPqeoyuvDEvm+cJbN95lJnj7lV/uQ5N8GvxuVcRen
GgRILp5sB+5IyT/eYCDiSvm5BD3ht2tPkfOa2VjNH1NyqYLPP9pfhC2jNF3ex5KM
7/vY6/n+8o81L8MEq9bsw5YI7iCCdhhihq4p8Z69l3bdRIbBWQM+6v/1f8/148aO
pnbj9+9XCg3OP7Wdj1thusogC1+M8QzMcqzciQ35IZpjNI9qO6T4O0p/enGrnyUG
yrT2jh49bgqFxNYUn6CjeDRGgkDN5tTzLUoeue7sifSvNZddtiIk6EMRUaXAozzI
KDP+Zh0B6yBVPBJ/G8Z3Hmq865MZBOduLTDh1IHoL4FOvZRj7jQhLIACyNBDKvuB
6gnbmju/t/nfTA5PEDROwIzHeoKolaxFkE8ChwEPrDQicA/EN4vEvVd70ZQaOlXp
+R0u3dwYkPpQpUwUXG8l8Bh6dG7H8xqgcjyRwiyquxTNkC2f5JcLpJKfAxAihQkF
Pps8C2rRb2+jyenn6INS4E89WDItOG8sB4WS7JGqazwRtFdlU35MWV6LaxeW17Fa
KEh18GjK7Mw58FJKgah1mlrAQnJ5DVD/2Lf6YN5KMkSgTdNJ0KAyg/CD1fK9Tk+n
lqStj2nFcO6fZIxXZvbZbjkRbJ9/Xi/7zH7vI0RV4DWfqdvRuieWqXWTgRYN5CXU
z/8747yELNe1aeEhj5Bf/FkDxt4rwiucPd5iay9pB4RAj3m/0aRYdnjG5pA9Jdzk
0G5/9AvUjri3E53O2ZOX2QnNNmN2xgbYu4J4SCNzisD5ZPjvkTTqRhATXIdoe4sr
dzikk1AdD2KPoHWgi00T8w+/KBUdXBMPxVZNnHWiN64YQ3scn7frlnShYpKnmqt+
fP9Et4WHuGTw/dofA8McoxNNjPGdQmACANUkxxbTObU6MuLOc0ueluGnSgLWs3k2
K+rPNsyp5ro7XY4rPT1kvuSCiod0Ht6czOSO69hJdOyvRcSDqWwPyqQwfgwMB+5M
GWiUQQjrFQ0uN7cq6547zG3loMT3PjSgxo9Wv0DSJza2f2j4C5N4X8UbWQq+Z7Th
ZJmqL0UHo/qSepBKx9Hal9ZHJ9tcTA2P0FBy3CM/mqVOUm0Uhv5m/d7mO/7Bn/eU
USkm/USMktP4gfYCx7vHpbJSsUBikR5BhwExUGe2hyaA6Za/oXYkF+GAhZ2gZziA
wNPc4v55R/7EjCCm+u7w3xp4TX08aOhNNtAuBJybUGR02MO5uQ1VeRzYwYmQ0CLS
36aXUEu9DGt/MqCdRlWT0Dcf1JMg5phElmLILKvk4Ke8I3KguOtb/Pm5pPNroetP
rC8Qi2EU2Sk320w2HrBkB2rChqvemulUYGMpWN91E5yvZGMLMM15UmeM4+9VxGwO
Dm8N3h1sV62Xj3HmXZtBcrEHpX3Uq2RTQt/RxPIJunh6FQWPrd135bT0kre/zIUZ
2+Dk0/bUI+CbWdHMVJ3LeUBqgtbjLqgel5rs1zYdKELcZMK+mMy6UVok8mjyANQ0
LYf4j6WIFUZH+ic7Kw4iZMKgqyVfVV/fSPtUxlPkrF3CYsN4AgPUPibXnwk06KoY
4eQ+if2m0F30zXmuu0wQxSUZCr9/uCBu29uGDz3CBQJ3XM40JHZLUJojCdSgxo1L
cvM+Aqy8CRdgKV0NM6dLD7sp9Tq8b1PuJad7XOng61SYjMg9tSPm/RLgV4ZEHlQJ
10CM55Ai7Wq9w1IaxzXqOHN2hGnUtPd2n2QgATKfUNaCcA2udp865+1K61cq13I9
MlkIytfMk4j1ToUyyfDeXsvjHFm7t7tPzSNbwt8gpkJcLMy/guhcIhBFlF40KbLK
ffXn1Yxx2wJPf+4h39myxkMgonomPXwEZHdKZHt3UB9B6Q+63MA0LIRJjI4x/vxW
2PZEANqyePtcSw+PShiACoyaAoGu2/jpu3YVSRAarxQB8PGSb6Tc2hBsyR1kfRIh
S1/GmzW0/LC9m8iqG/4ONDNBWr+yO2QP1QUgezVZQM30pHHO5R3wQ+wEPOXm35OD
nfnk17Ttz2LkQvo4y5SWKZu7xU9bIeulxzB5KPWrHXooP4SXwpS1Bo6h94D6b8J0
0T+8v4QeOiDBgEdADUyR25gr0K8/6Szig+D9B3mIIVXFc46fnz7VNgu7Z2ChxI9a
/uRMRZKaw/S9FEcgfSYPurJcplafG/4yQcX8S1mrWcQzyLHMtMTtjlGYJ6qCLI+4
r0qYKnOdK074YWEmoos1d/A9X7Luq3s9RlJ61vkl2gPXCoRBsFDs2PQaV4ZkrBNt
Bl1D8iFoNCcPIENA+75glO74eXQwo9y1ZLrLZjlJQMoLoRPZgcFQm7acOtVjbOU6
0LV0Put2Yp9yC+EhunfdcKoX2RzJ2tvZxfa/yjEdlUCIm93Q9roOkPd++NnAxDNR
fTRCmnH7mbkXjirwB7t70+V+P0SUeMuHAtO3JQxuAo7K+InP0jDuaIna9SIZMjyC
iP9QKW8sYiz2yGZ9kEQz/2b1yEwMxODCLteasSPxn094SBc5YXlc6T1T7qztvstb
vkWNeOW2Y249Epa/VGQnGiNs6qUrMT4BChI8gRQbksKzAMH+Ge0WER/FoshKLVDp
fKI+3zlkplyHLx23gJQNx5Af+SWRI/PaiVS3vd5HozjbDURwYcPHet+gqWpjxGNf
2/0qjJosdBzLOsdR4ttGggYCLFecgXzByAfWUVlwFhmxGzm4GwitgSc74UM4+5SR
pDOiNkh6POeVd4+0WxDuFVg3E9XjCMXi3txqb3G/UwKORZ6w8wW6tvk+Fk4KhQTw
C1bLF7MuFP2gnmx6gU790uWQKBLRasH+TFy8hNGq6xUO7etelRFK8ALFa9DHy3JC
p6UwyMoin7z+XQRwRu6H7LifAihtmqxqibOBkucv8PZKY2Hzv069QBkNTZSBT4iM
EB0eZDP7w/idvYUvOdKQ9QUDHJfc5Fd5VbqRzpHNkxrAKKSVt1K8SbUzTGBlDWTf
Jmvv27h1RJKruJy3jPlEeip8g9ZlTv13JhkXUAX4tsopvvz0QCeH/7m3xrQipKZ+
HITyHS/DDu0LUKYga/r6heqbjFU+Uinr2efETwKiwikN2+dpXzPHv5lCfIg/uwyM
ElB82ITp6elb+N9kAw2XSCdoq5QfG7xyRoNIq1qo9pkq7mW7oUXLISC/5g0uAKi1
b/xd6yypUo5YZ1P+VdM8wsT9+x216mHUVENluAAeLlvfS9xV1lw70dBI138Uvo7P
Nlq1F8nIarBMXr5S+Fnx3wZGNE6cCQkKSWdAKmd2B/nev58TCT7vOglfG1mzOF4X
cSi+AcXOfHICs/nGzOGerzIZwgk+0U7Lg81tnw1Wcna+yIMRf7oVsVO/h4gJAm9e
yEY64ZMHzalxqFkICiZWlV8QeKNRQBfr6quaviJ79r27VMKwpYeoG9bcLJzr3VS2
v+uavZEk5m5P1x7LEXUiCZ595g3zlKlBoc63tI7nu5c7dQfjYlc5qHmRBEQX9YkZ
YmCqMXkSUa42yi00osvuVUvZxdVXZhQLWh3wd5gxWhMn9wgmKSO47vlFTyxFmcc+
WbQRSX/rUQT1HP0L9Ko1P226vShyMfKh8/n5xOs+BjGFp0W1KnCKzh5J3d6GzeiH
D4xoqaw+rsK97JTDJwN5kHPJAxCvexQMv8l8+pCr8LPRRrjvIhz76v6yPXjoc4D0
4Raj76J1KkGq8+r8DWV1LIkPi4Kn7VjdDmw/4GZDw1sBpIbtxfTj/vfSF02Qv9eT
IbxX0tViuv4CtCcqInL3QfZdTFeWcJYBoZQsFGLNFpRYO5oXkIOgwCMTIifAMfUR
vMzT5+KhQp7UCqjkh+4oYl9fIXIhVSbAkPO9T6xXoCB4buKInvDU2fiYjv3Qvw6s
A5BGhJFB3dq+82ONFEazvPeChgI7nm56GRnfbLwHggC61828liRqnPyimh6AUQCI
Hah3mvWJOavBN6nG5yRkA96nRyB3DjPmlY2wrAvIQhE8PB8Y3POZnxZR6TjhXJ9O
2SXvLWwn6KfLOlUvOtMgFBHx7TiE9wrdy9n8irGUt2SuJEM5L693NMWptS8Ckdsg
Wkz00H/P0vr7s+Cq+bkXBWCs9BfRaPxlMfS85AFsmmU6NFPbhYgrCxvAx/Fb7waK
qi7aRZPEImdak6kZcrMcmSKwH2CFnmtTCSahZGeeOYzkrIbdi6NDTrpP2Zz/JwqL
9yoYRDaeHLfWBcw/J7FylcXMV57CrrrrakJpOwC9vcvxG22D5a5E6OMe5P2CYLug
SD0NB5x1Cd/5I1wEvlAF8d7vwGeFx/wjtWBQ9aFeqOP9WN9GAFQ6+JShkD4NxKkQ
tQn9VwskEEawoEuHqK4Hiffh0ts+U0Ec9QQBYwWVNF4/3bpf/eDpenSQgEi47jer
o37BWWU8TyuBzvstUo0/AFcnx4fKDzODJsbjNSHDZuY5ldXKQJXd+HC+xupUDJ8b
IIAqwJATIzxUNQs5GeFZLNo2i1u1cUdL6rG6802qsiCDb9ZHM5GpYqHHQVYW5R3M
JwEquw41eRu8B78aI63U+9kyCpQCpjikClGWFarlD48eAeHVF4LFoZ8EwpPAxO4H
lHfSZu86mOzmt/zewKCN9LGTvd1vaSL7uz6jxpQtcmVbkTeBdNoxDKlNLQUExrth
bI3hneY9EmwWdbywC8fQEgctKKDOSGvdSNeXmEiJlALjDNj+zn3qqTYopcyXEj97
k3BdEkkEmoqfWnK0TRpPFYNH2wNhh8PMVUULYKJPOwHUkIO/gkck05SICNCNCIo7
dMlFpgG8lnvapZkAKo9SfTJYVEGugEiz+GuBMgym7uriV5jzCQ60Eos4JQ8FfRbe
caJC7gXvQ5OfhSokg0O1k4LSLhPjT1hh1VJ5oNg+pQv6Oc48V8oJp/cLLWGI5QpO
CtuvmW70zRPDfb5wwMVYeY5Zn5brdzAfRrZGvf1n8wzYuMgF60ILkg3+hY//qvXx
vkSBf38UYlSTN1lKYHLOcLrpEaAaLJVdcfzxI6GmeRQ573N5c3DoQKFay4kfT04d
7nLJSLKvqMhcuvuEOEHOi9+wruDWoI9Y8aORxQk3pq7tF3mh6RFPGX8E/6nsnJC4
W89yhUygW3HxeHu2VDzYKE2MR94B8aYBvD1OipGu51VNxa519JiNj2TY94HL5dPV
ntZfYsYZM/RrjWnD9T9T5SCvFCBETQj2A9rYtdlV4ezCldb3wmaLtxS+I1Aot71z
PNwIDe8Wr8QkhzN0w2UXCG3uwZnbLKMEcj6dciu0XWlnQ1/VFcnYw1RKkEsZ1hz6
Z9n0+/4Rcjh27kv9ZrdpYqWC7R/rmezds6f5tl1XahxAplvTkiR4ro4Tq5qrHTpI
QaumcRcNFkiMcOKKzwKaj73GA/J6j+pWRYSe8gdzKnUpMjL4AgwJdnMlZt/f/77M
3P0u3sSUsXwARY/ImPRWOxDhiOVvHhuyH5n3ffm1YogMwVa9am/6cKC6h+dpGGa3
6l5MQ03TZbI3DWbNC8ONin61mhiVV5IcJF6YLg18ufK/YpSOTFw0yLXOYM7AxdS3
5ZvV1nwi/1VktexuAAmNRDM/4qNCIxtplDBqo54LQ5weULWHbK0X+e/KWzPh/sgi
djTtTEzZlrePzDguQOsGZIEVfQ2PEP73ynYDGb/7KVXn99n7u9IPzvVeShvGuBk3
elYvQU94/3m9e+6hN65OJkHcxrSqGGVUgBpfNtcoSrMsffG3ZWMP8Fpl4h/o4qHz
4GWyMuatBFi84nFOaJr8qTmXBJRDl9H+cRbqntmaBgI+xFDzvXUGJsknaTRQlLmO
JhCPj/G/3InVXStU7TwgaiFPaWyIKhJOrGbVtHbpKuUqpysDA6HjHBHHesshNEWK
logzN+qVUeYaUhgyOQSZKgzKW22c48uC6L8l/g4oXlVWvMpQwWXvQsemTHRIp0Jx
ZlL+XN+CEzDoIMo5coTS8Wzd8qtAaXkXsJtTkYqpquD77PjHOeSBrz39UB3pYoM4
Pmf6tyWLSo7lDE+1dHLn0i9njKGxZ5y4J1YEgiTzV4KOn8NgidbjOrY/ePiuXMWF
rObhz2CoNjo2S5Zn98pfV60F3JsPb1f0mRTyHQyWq2IJu4VkkjQHH3lEbEP4Hj2o
9xqqYiiVZuU8fliEEZNhlIalYvq3VwEoS7vmJ+MenUOOLEdCHIl8xCBPMVW3Tucy
z7xNUFxRczvHkOcd5RLJ8twVqhXt0L5r/lgTAbhTI5DNlkFKLq4tusiKpcZetXVm
K4CvTNrqoy3S8/aMB7/7R1r5F6hrlk4lttm/Bzl6RlbnSk4hukUGDjOGzLUEnpDt
JuxJU7ToNS/DU7qmt+qfBZzlyweyupKNHlxgoLhuVoLUO7K1Th4P8c26GdR3x69C
CBvtNIQTYEsTRMFGxGsVDYTrBYDD5ZYRGckdKcCeTlSBIuLE558yjZEJ9TiKWuLM
Ih5QwAldaPc9Gkax6ldPRrACo7Q/UDCTMimXHz14tj20u5RGWYPRYwCTa4H2ZAUi
qWHqDrgYdOz1x3zMFkCe1nOXPByT1MWXxf2mOUccPmYC2DGGzW6pn//X9HbQn+1R
us3vly0w6SThXwyqMCygB1uKUeGaBc7d/lTQataOMAwZJf3b/y5r6oe0u8N1ujz6
ri1fmEcZzHQ3MPH59uTyFfF9C53LucXzhz7Z0qHo7d2T2CtKh5+RzAIMRYsqZ5WF
BqxqgpfBzwZcvwJTdAiA8OsIgwIzrWa4v96Hc0ZYM7jJYpehqezkZQ7nUWMUAgCH
/x+G/OcSRszNFGIaxLjuQr4dqGW0Osp9DHKj7lLlj32saogeEaxGr0pjXVceB38U
oXGiEM3IZJGN/R69SzBIA2FNqxW7VAI14Le1UqWrSsNQqpw1FEbRZ33GWV3NH+0u
94liUeRgN12bZgkf/lNePWAEf0kWo0x0sk8KTegKfTeKI6rEmBLKMhNzDLErX0S0
mUgy1QFvZTvfuWVzyHLmc38f0Q9MTppUiM3ky5EtRlQYz4mPAL4BdrlEQm8M9+w8
UUhBDmifxHWHkX5S/XAGx9OqkFFThjW+IMiyq7oHdDVYXWK0pjxyv3xstcQiAjVh
3VboNE6842vBYjU/NfxP8j1tqbHxefm3xb4gV+FXdT16RT7/J9D+kWGFFMnVaSLO
L7CHiwHDyVvWF53fbEwB7hIQyEWKPsHYVY9eIC+sYtp8vLaKDVrukL8CX3eqfzRa
K8e9lnkSMwCgtdGkCn/vAh7C3RgIDEPPfOucX3HefALMBOkr2aUPYd+AaNGRv0un
CwiTYjwVZz/mAfx0mWtleV1w6JbSmIEe2L4/kwdC3YmD4bItVj6ri0CNlAquN+6f
RVdACQhVgqH7nQmdJrnWSIUnomERB1TLiEiZrZ2F+rtsJF6Ag7NQGl6+YeDCL6Zy
wkgbIrFS8Lo3AVI17O+6pr//7UJX/bDHHCe2q/DUvDpPZyVhEMSJizz4JrpTBmzJ
E23O5C+pBOvk0oj5g7jebqHGA2GST6xshqY6c+CknAMOm5EAa3uPUPuicFpUajik
EY1U+iCFvDqhJXZWSpWrWUbJBLzbYmDzA2X44YyBqRneu0DOhL5tKmmJHoWNkBqS
Et89NZVWyhK1uIWQEHxu7tuDi2wwhDcI2jH1tQqNh8MVecFTZlp81HR0VdIGNK65
jllEQ+PNtq0JBn0j02SAhAO+8DA67nM5D600ZC+56J1aM6QBIUGLw8IYb15QS7Lk
dqbr83BX9gU6ER4zrqjXKvjHRd0gpSoCfgXSg0OR9Cq24LRRSvkehMJ/sd2zDOu+
j9lRpokOoiRfjI/MGgq6QwySba1f4yNCbZEZ+vcx7X8YKxdrOqoXTfqz9f5UQGLC
VSvwgML9A3HMQdfLzXjxwS6uo0ERSlH5oibYboEM9lmsRiiDIEX6WIjNO64Fjgze
EgiawGQLJoG1THFwgKSopTT/fsvfzlqC8iMHUx7Tf2IKxARyq8HtwIruRt5wkIw2
bkreaa2D5Nm3Gawrchle9wKLhk8hwoIsR56kZwqHh1wNtW0aR0lOdc/O9cOKNi4R
A85FXu9ZMymW4MhX9NauePtyaulckbDfsSHUrYa9K3u3FXvFm0tZBLtk71WkqOYh
4yFq6yH73RcfR41+6y8NmY3XHIi0ti2g7rLZ0E2eVxbclXp5u9oUy8t3462OqUl1
dc4LMw4cGRYaUlF+Pz30WDyU/HdsGdDbnH/LtXTLSDcSGDjt1bb5GGCy24s8hjYk
wVM9z85YsG69Tdyrl6m3q98+9VTpOMGniazKRVWj0OF0e/tM8e6em94oVu9wHx0L
7mIgE/zJsQOLxYzRG3ErLnfxossKqkg+8RCpEKOIU5e0tSAjJAZoCz+KpPZhtvCn
iw/xTHYN5CZKMRMTFuSSoJLt+fT0QqD7JNwvZfSVcNV6ONeihU0c4tl3rsc5L9jJ
XcqXzqiWavShNqgtFjNtfKuuAox4ytQWG63UPfGs91tvEq1TxIJsmkQ4OEZx1sAS
g45jvHliNcjaiQ98ZnDwrJ/qFtB9L2/AWfPl/qq5n5kCTgMUWpxcaMwG2WiTEWpB
XwicxsZanyXP2z2JWWhj98fXlFkCGUViXfx/wK7vGYNwtOKcqVWsW7/f3jPI2Woo
YYvukJ+PPa6QbdvGMsALuVtNcKZG2wcb1EQa8zIjWOUP564/ikRZKp3ymeSxVRgh
d7IPA6ifBlettxRCourkAu6Hqiu/YgNY9VkHHb+iTLFfYwmTJkCLZk/b2LRhFByt
xckNeHJ4tOo7CJcH2+A4MY6+Wr3pRGlxaEAajzOJ9W8MVe3vlp9FAW36gAIrPDf/
ZRW50DN1xgCWVRUk+ppf0/bzjYC0ECxuHvh2iDtKO+f5+E2zApTHu7cetVqnKfqV
Mm6UK+x0wAYNxClV0iMt9ZlEYFD+a85UPTLb1N8k7kBH47Mx9iKekdZUkZ/0qCgu
2tXPW/79RpgQXFk/88gEbgLHfTbfXaUzkHtQeUT+YlFxayjXhVS/RHgu5+MuW2I1
xm7BkfQ2Nh3E5GY/tvJPr2PTfwrSrh3G60RaXpIYIssnNU76da6IENGfxxCANu4P
Yd9TX4mDGm6Shcxcok10xXHJL3VoLltbCWAN+++gVAEb3ft0m0hpIcNZ1yXKhbeJ
viTqbFNnQHCRADtGWB0/Zz5GhuUlK3CB6AKSe7oEHvppyfVe/S1Y0W2AIX6IbDND
LCk9CpcaHda/CHfdlOjvA9+KdFGfj6y6h8E6ie6HYT4ViHTm3cPw+EK+tmG2yBjE
QXj6YmVZzez66S3F+SPS7QlANc7/KuzmUdX8C0yFCs4AR5rxCL6h81wumkTc2Lf4
zOPYITB/YRki636ZP42gqMNq/VCKECNtpJXU/2cu8yquvUet4ZX+dWKGtnh21q+B
3Mp2RqvlZLH2N/G9C+NNhc7xgmviFoWlrsD1TNNoI4C9a1UOpoR8d7SRqupd5GPd
pd0MazBePKiRKsNwy2IEKju5yzKpGiAx4l/OabMjyfi4nQiQiYDihspm70sRl4WD
a35rh1NsLy5wi4CpQL4Lalmu7o/eX2OCAhC880A17yxeGkZMDXenVnHZTeh44kgG
hiJI17RH6KwQhqe6Avn5CcPpCe4c4bl7t7/gw2DOkSkC0nI+bCgdQBDbmHiKJoZp
RfVYsHDYAD/bfxlMWOT8StGnZ/KmWMn5fnSGo6pR3j7848YWud9kxQQMH75slHrV
+wo1N3rul53UOzisiFCfKJWyxxp/U9CXakSODuNhT1tBZL9d71/qagceXeOxXRpJ
7zD+1ZGxodON5N+9YPeMe5LSq9ymzbB/RKBxM2nTYtmOCouIR5KhG/Vy03Y2ZeGj
wOrP16N9LW4c//FBw/DnJyM+7bOwl3zM9HfOPouUhJZRcSvF2nrc7ou7B000+cda
So4rLH1rJ5ysN6ZLSDv4XH9BT6AQ2M70BBmWFt3/tA3YUBReQMs9hWQ4zSgCBEzZ
O5INvIf9cxuRQA3fTfIhiOm4tuIJLeFdonL08p5zx7yolvcYMkjOUNDwhLW+uFQb
BUFFehwstc5gcjFqQIjsit0NxI02rv+y6jymu8frtul9IRwUfr8k9RmGvCmKBWRw
ZhWdgUIInYn0t7FnAga/3RAF5WzbcglAZiiQWRp8CboLf5yc0iAhBvSiiR8dOd5X
cSdrpJZMAy/CbE1AcN9GI3x16YMdhxq3ZiDlr6OibLCxoM0k3FG64GLjJduK0VHQ
36NY8AwblhaUoyUTN9s583jHSqFFrf85SMDDjSZ41t5Fhrvtrr525FrflucuYMJW
/CBTcSzxeq8DKF2aqbR2uQyOAUIrS7iSeF/lqTdKT89d6vSDUzdRQAI/OQ+4CNym
mU6swoXYuGB3DL0cV3r/B2bnK9x8NRu9+M2rRI7cXMD7ZvJnp0or0mdRsHIOokR6
APZKiyN13YjqiHiwb5QaJc3JodxGIq87ZPBL/87rvwXwODC4hiXrRy3H0Xtoov0a
cdp9ZdZK9NzN7GWyZqhswSou7kWOMXEggjNKImGEF8qPJ/tvr7mMbM1RNgZtwOtt
qxy5a7WDW97o+32aR/Xz2Pe8ULAeuW0by1yUYG3CPTDSrXbxu7Ad8fQAv5kBaMZY
4+PS5bBkImSGMaqsntKuWUGNbulROCsEjJ75221l3WiOSCZfU/QCBFZz9/wjdkhA
1eEnyvnjmJoYYOwzRRrH2NUVjvJweRyygmeinG5p6Gps6CTc7+LialcEMHZJ1RBG
EmUUrSZ2bz6Sx/9YMRHPDAVW5/bfCpl5LWRtNe1NlG69XPPsk/VW/4H1VRp1zo1Y
glbUpUCdewlWOuDGdP6isc5liHwCNPDcsqArr209embK/XaViHINj2Mxm246EEyP
jupy07vHOvz/kIZQo7GHgqH6EnfdN58U795rSC9TZvWm87yHgQXrPlpR1DZhk42/
V2Coofttnxpdy0nDnax0W9t1ZDTerfm3FlfSy6MboutDl2HF6lQOGFXhRQmlgDZF
7H5tMHu6JWlwqIGUs3Xe5Ms5doIyxiZQ53Ag1UxckzR7mqgwAGNykN4XCKBQMhv4
0qO3OIe3I0Fwt2/mRVNYJjf5+rE0/jBq6XgrhemWFsZu5NFA/YsYT/S4eQK1bkQE
qY/ccozgvySeC7fM66RRmVJmWeH6ZNJRJoHcx594u/JXju95u1cqet2Ynjn2mdQ6
+Gfmn3Or15UHtZQGrx9Xi4x07PRyI1N+sg9bZCGY3CNYnXBDmBUpqvy0wo1740HL
dLpP2REi49LfMx1v4e8/Pva8A7Nu2EuBBI928L5NqNbGZHI5jM2b9d8uI4XKOszj
dtifAKDlffugIbxkDF1EeyjwKE5xS3D3XDH60LrPPKwi/TfOjK9WQD4sqnr5Fhfj
WAUuIHP6V66p/2B3xRn2FvrRtjrjXxfrIwKUaFzjH00WtiFTJr1y7tx1lZ2UQWQP
qOrb+6unJTaf9FsfoesEtaPcvx4dGi3TJpZ29vKUqL45QiHGR+Qj2N8pAdYSkRPR
g5yj8987W5yhNbJGwgTjkkd9+4LAg3gDg8ccZBATg067GY7IPtvS8H39KdKhFc3h
0YWqoaoQH2/t8EHupoaxf/XGbUlC/LMUXmYMetC1aQ82Ji5FeDfl6ditb9+p1FCb
Ewq8rAZIwucHw/0eCEk4C++O8fAWFOi+rL8tUfsUmfw1/VFqGt8feknX7zmH8GOA
bmyDeaJAf5Lph1dwRaiScyxsPxEXe5IaAU/Y7vBmlUdCOKf7o2Ago5H+e7xPce6U
xBS8N+Wos30ikaMyA/lpxNHcOMl80usmfHY45d9HJZilk3vP1P0JHX1jmdGXHcrU
EBmyBdhWjeJox0Anf0e9L7KknBClvyROTZMeIy2KzIxmGKeBlONgHglJoK1ziAMB
6l23so10Nec1FaLdFDB4TZ26mXZCFGPnska5MSCBoVpGNx41qSpp7UQrFkJaYBCw
i5O/S2HsshDjEGr3KOUklze8eeP/Grri4HbYW66DLzY7KK3iFk/6SHdc50uOETlw
MoVHb9lX4UbWgfBaxMB3BlZNFhhyXq7VSGu0W+pSXHSwwOoFb0VxZlQjppN8g3LQ
SqugQLGgD5g8HsPVbKMPR5B970lREfHZe01b0oPMD8H0FsKJhsCJNHa1UDoia3ye
ZwSaQn8nZsgziGWGomr+Kjo/wcL3KMBXU3DKOoy5AajYa3/tZ/PhwX+/OUvZ2jLv
R6zLNIU9UROIREncCsFJV/TB6EVlAptZqTjcXSR9CDkb0rWWDG2WlTKl7KugSTix
V9u+iRC1Mb7XYOb02yWcNkPjg2S7z1vXyXDSmWl7LhSXeyhohB4MO8rFK/kSK5Gp
z56fkpsoyh4zZfEeKqAMLlYZ2DA+/6udeM1bYKc8sVZ62Zn7Y1/PKUnZqCr2XY0K
3c7FMeacSPsfELhk4eOlK8dSzgDU9QUzoThIvtKCG44L8Gd6s/QMUQQIJh3IidQC
WHNnPXIJqnM5IYcDDdtU0CDOyuY8jM7cSKhRHWaNnw/EDouoLdCLF8k0D9nOZ0vb
pxkUxCOc6AdVQXzJ61CpS4eqBb7Hoyywdb+1TQKGR/W3HsvNQwlhuO+UT4tQG3A/
7KfiSKGzcU/hLrimhbtIoduRVdQoA7ecvI5Dk4EIp1Ame2a/6Xo6Vsx4HSl0AOSi
Gx65URhv+kvpxBqjN0HD/vaoLMA8YVrBnfbC5EAZfRTymqJkRLRDA6CpSZnJwNYb
ju0pPWg5Dq/yE19++2da0ceMNRn+Bs8Sg5LvRgixCwQdOJqaedMK49sumpr5VLuo
6FOWxAwMDWskxquwJyIeMgf+XIci0bKFZLDPE/NdTnTv05p+CTFquOtWnEy31eSw
fSdf4gfWhw4THMYFTFcDwfdw/pafOM2JcLdC2IRiA/3Aih7EexGHw1sxWLKfueto
GB4W2N2VNGu8mgFXApoo8mEluS85IXA5v4ocj9mlcapbizgxd24J/xwAPeU1MKS8
KpZKU9BGVUO2NpTPPKoBf6MmRBd8MsQ71iwTHeyIONRRwP6i9I9qfMyyqBEDY0kJ
zj4YUkXo+WLKjRT03cMeO7oSNd2D4T3o0SJK89C0JQilCOQFMyWNJ9NWzaAE0Qea
ZJqFYeWER76pm2hn9XgSqyP11DXoX6Zap4tChfVJ9ALR/aTU9Aql25N//UUheGgD
4RUohcuwOcDqDw4Atp0Je2ENuhzHwDI5ZRaw2lDZMMZ5B2x23kEtyGtYF2PUve/n
nAVW+/8xVzQcRlkJCUHi0hyt/dx89ZTqUa6cEv1AJxEvS9eAsLR4vBl0MX+Aft/Z
2ACiZS3o4UTLAw/mBJ1wwkZ0L0HdOjvCcvH7poL3R1xNQ68D8KKIwIrUz+2pkMMG
YExm3gsUxn66YUnZUFtrheqc1tFWsYy84KUW2Dn5g4jF2B93AK3dBdHO4zYaJC/Z
yM43FLNxzsEh+yKogbGEGBf4metFMEnMnR1HOaPcuqYrqL+2pDUw8tXkiUjT4eOq
Kd+vvMHc9Ui/WQyx5f0UuzJW16eB+HN+5vB829vxw4d8RRYn/opFWvHGr0WA8wfl
nzOFnFmHR8E+GIzH33gPlX7TDIP13dmfC9UZtrJIB99WW+emGLJQI5yHkWgkgwA3
vQ9e/DnfnGuVmRnrPF3OXQGafTgDJHw1Mq9q9EQYXN77u1sXwL0pzSjOpBP2IMoD
gehDpAuN8dzdNw/bredqJAE3+zLFdSkfCkOaqtfDKkqjyw/g2oAb9CU+lnABxQsr
fmA16ZP/pmox3rbqXMoXgmliTlFklR3uI7uvie00/3jZ8N0x5/K+75U6TfQfcZpd
yVJdvODFiT1itIXQkbRk1q/N7eBoVizOGpkPwQMztn+MDPrJkKi7JiEsXoGT6bug
AfWMND/RKcTfKmVkbrVyZMrajCdN+dVqNfdx+820Vyx1p4VN4sBfLmsOnJ54YKbK
Cojrr+2pw5UxVh8W4rk0dSa6nHiuqgpXAcm2Eqnw8GemlOH3q/AyGryEmtfqb9d1
y2hXO8S3heQosgC46Gu7FSnP7JQqI2nW1iFh774kZpfZHHPoaz9+2Wq8gyFYzORL
z6qAY1nrlIbJgTcVXKKg9S+fAGT2Z5+LOPs+8TBYwswaxmnAxaw+G2cc15CmP579
mATqWJ0BYc8er2l/aHHeCYedfWCMzc3DZH2fphzgc4aIaX0dnowa8r+dfRC0BRKf
/mpTqyf+4KnRSmXANpocab2fWWAcCsyGi+bqZ/5e1sbb/PDYcdNUMgHpaSQUX6mp
1RhWEbWQf8Om62lKr6cM6SIOaTy35mhgAUG6Ciu9l3rVCT26YlDoWzLHo85GgQjC
H/TOwvg3unLgFUoLUvogPOBtXO5+esK2N78dESsCtXhrkwolnefocIdpRufs4Pj9
jKO6ACYa82yqVoaMG3+2bTP5NJPn2dD3tcHClOLo3QNFNMNgwjAPB7GwRomVdJ1q
z3nhp888ueL3pkv/ZWIzqF+8zAcSXdlzmJuVcOKLh95gXyfUktKXMg9qeCNCm0ZJ
v0Inhxi8+CEaaElc7TTszPTDUN96HdAutJQzubZ07+cWXpeul4/lNq3whQwvscZr
/FbcAQg1144kOYO8eGMhbuINyQHvLE3UEr2V4wLVqCHmHqRHENefG7eV3d2RnvdB
zE5JkJ3ODGVwbY4U/HFt9OV5bQhvBHtJGpnwYFhvNG3sSoGtyvPBBPo/OKR9q/YU
Dppz3Qad7QuHOm1ak6bXDr8mC9sYuKPRCqTv5ENvohMI1fh7bNytlxZhdG2Nq/dC
kKwoUSe7ocqu9U65gY9CqW6bfNBn+exWJeZwoFqvx3FOAq22TlRE6C9nHNFaWmtP
t2xbHXg7Kw2im4nxekgzqrqwamBd2A5CWCRb8zBd6iSxWH0hjRS8IwWFjCuF2awc
GDT4Y9VM9pT/lqq48Rdelsr/ynijRjx0KcWZvu5UrfPz9ZvOUdLnhqsSfYG0pLHh
DcKrAZ4H9q+t3drFFbrNj99PRi2a6Xcf6kkLRhREbmlN2nTvRkhX5RFBFYg2eMJg
BbZfnnMt/iwYDMHS4nG5el/GzOJtlNquqzwxYj3MRwBJbDz+SH/XNF+srCK813AR
5qQbcbz6ovjF50QKeJvo8VmUyFZCS1SMDsMH2C81TxHoEZ6aM9isZ/0hEowZQDj+
ZYEamDpmtogC4xg5uLFD1I3FFeQawQrvc+hpQad6oMWlgz+poYoRB5yJK6bQa7Qo
ZLb7ib22yS/3z43/kbi/KO5WcIKg7iRJy+gyGRTfJoRWwCYIbk/Y+5KOpJ7WY0OP
/yR8I0OmIojWzCBF3SQhdgnVb11ccUKQbtUhjbQmh7tmZkZooc+/WzNLbhVnHcDd
yDKUKt9L1vzTCNqWBbosOkob0DWb55J0EpcGJR/FLUAv7a6UJBGOh3whLBatiMPR
Gnbdl6dZZAqV8XLjLNNZrIhnmHEMVO/uv+qGFRDGauhOmsDCbgLnJIhe3tZ1oVR1
tNYqFtSzAyg6kdigqKwFXygafFH868lJEihk773fWXU6asU94TFpAWraRu8Q6l5e
Ivj6sClIf3MJAXFO0yeOHTbxzuTmZjG+uqsKOqoMqcxNKp11ZX6D7r4ZNdFVPNTS
q28I5dAtv4faR+syne23VaPxgx2I4CHKzDdTuIno4w6VSVkK0NknGa6VU2a4rBMp
BIHI0cWMmd4gH/ce1oRsg6fLMjFshzmT1HuJN+Mro2EVSgT9Og+ffr71XnBVna+Z
IhE+WlCBgvMBNiiPbdSd7/WhDZpuXl1CUVi4ffXEqmnOnbQ/MWN4jqdPtir66TNM
IHBNr3Nnc6A1bdTwTuTmisBAQQZLK6NBYNzj1QTsOCIZrbUCMpqwssmArOj8k4Ru
FcLDrbLHP5fSIheiz5GwPR18pbjNdeGpks9DCKpAel8s5osAGw1W0eDi3pQ/EYgw
9Ee5kma/ZONlv5QzSGfMMyTlpOKMr8Wplx2uKpq3/Wq6Xo/X5SLd25whSdj1duq2
L9O4t9v8G4Wwatq6DyUDTjApEhNT7RoXNtVPu22Zg/XFvlVaYSoV2vxOXwdjwYDE
/xh0Zj2qgI0WDu/5tpuwDWcu/CJxZ4GrO8jfjGZEs2D2UASJeqy+RNct1mKogjHm
emrP9StjRnx6QsGToHP1WMKN4d1nbg+eM9rIg04PqGv390P8XwjpS3ZtvyPkBPlS
kGNz03CxtlZwvQCLnwjoOkqp/AxXLnvvRnTLG7NrFX4zebrBSq8/lehpvvBnrssn
XvcXMpBPD1Y+T7m+1ovxcFzpHJJSz3lA0qc9ZfbcThweR3H2PnUDd1QovMxYLiUh
FubhKfRddJ/212kJjOyuPcQCt9NYC0QnAoVhvp/VPDY94C6ZUN2zoaE1NIaUDJ/f
jl8c7IOOwUOc/C+y6vgal4sLDpHmdgdQVfIweqbeazaQIpxbksyQPZT+LGZclRWW
VUakjOMntC2SpKKx3YjeYFJffthtVxRtCAZiAjHGGf0qKMF3qr8hMKR4abBjJRZb
FkdnvvxLGPMTEcqXnQJDRERVM6OHGsuuF8mxdQhqBRMPNkz9ZKmWNtXV4BUQJkgB
f7dKER398WuQ4isTX8SE/XdAJYDpdCJd1PmXh1guEmDfNnHss7Gg/guzB5Z0S16P
j3MulUpgcBsD3aM1gq7zyrzkK5Yzt9tpDGVILe5634Wrn4sGaX4g81qkU1AyprKT
5tNu3tZ8l9dzijFVXS7L+VvmdL9mcY5b9bLFNFwVmIGnBVVkSrvbSPWLKEESXLRy
teL45bdGfMG9HsIoxaIGwEcLKRIXNKFaJmmKNCxZlLayFN/UM2egpQGQk/ENfbKC
sa64swAcPvE5su4UIAaqnahQ0+5H361qQxbPRyNAsa7xP0Em/AVvwfRpPQ+lgXJq
BoeEAhWvOqNfGfvezRq4530h7DvMeINg5rAqZKnALeI41gboLQfV5Uvthgxh2wDw
b1oyD4YPed6JUfQ3SZh4f+M1WzimQI3/tVM8CdmW56X/o3StmOlW8oTsYy/QrRyC
msKIFhcCOdB0JIEfttXSORbUAlN744oN76p9O0mMGzRPVrLXpUDQ/6pb1onIgjTM
LzxExq9efMfs9Ye+y+a1Qv6/aBYZSuGKxRb2gxYwvczJJFbE3NW/wmgqkpne4bli
T0Q/03dRKLAdr8unyf+pjX5EfJEePjOQ/PVCNPQcnzx8tb1BpDZiG27F6h3T+9m8
Cz7elmW2PCUsIF8wvr2pBRmP+6jLW/px6tdVXDGm9IskbyuVFw+Hl/Oa7km1ZK9D
fXVLmzlfGMlgLJehMC0z64MXaRKVpkmzkD7YGXdaBYDRKyLk2jUubr5n+wlmQxlE
GnCf1rmcsVEjgR2szaTgf7j2MxQ6XMl/h5SdYyZo1/S3VO9E4HWcsk2JM+Egy4yj
g6+W3AKcp86c0p0r6KaSkm5J2pZ7Ojy45zYzXcpQtvVEMEeQnCdCsCm0DSjeFIsf
VMrcKsTLr0K3Y608oB5Gx+ffKz+WbGTCCTmbQvpOK2vUkBtdSLfdqPJpcfN+ZBuz
ew1Bgeb6cF7aikeRcO+H1GmoEsKDva9Ek3jbS4QvFBJy84Y6Fr5Jq4EAUD7/qEjT
MTtmGyRH0RqsCuR6T8GhxtRiw4/sy3F2f4xdiaGjCtTbGhzTVudzC98EuVA+jlrn
CSsEuOwL4FSP4PsJCjGwIxTc30XiYbCXPZyNePT9FGugRaYOC4ARF9owXM2jh5MP
hMzqSqCBypVB4clYwL4TDAkpC3BYwg+9+mI+FnCympz7YQPM27Ju/FnsO/nK1uZm
Ng4f9XaQqiDIN/8fOMUyB81yOmvG6wIQXZ8dQ5g1zKAAGy6kL08nD+YuX7CodGbL
53JF99sv8SZhH+ddRiq/+hI1g5KfZTuB2W5GwFmRVKxWA3aMwprzZpeOGMMeLXr1
+bFkEqTJancV44/LWlRCuJXVgmMhg4RUgYFxshKBeKLkqIgo5OGSe1lf9zkVmBrR
vSzaeFj3ov2jTW5BwRGJQ89W+yESOubkpHh1Y7sR4N9IQwIMVBJvXc81Pi+wJLTO
fs2PLTtlHCjm8JChZQf/l7avv8sgBig6R3XwydVTO5Mv/ixOdSqoQC4KBlmf/JzE
/xT8ZMMDZo1ezOxvjMJxXPtmqKxrAk9DVbMJPx+c8mnbvjpbi3oQMLRkW80HM7or
K9v/9RSLtxL2yDd5OtmldKQHesohfRLfu/ZOkoPu4hx5851QGdw6ACqQQZ+q1/OS
/ZwuJ2G62jVOjB7nTBidScHtirHbwPwe/dclqgJiLCS3Nt1NYQkqtt5j8YIjqYB3
a6II9KFS8sH8FiOtw0e0Q3wV+n7AzzVYdjemGYAdOv5fbJ6y/bONysEJPvZc1afp
qT+vVfe/PhFJBvt8OxW26ALrcD/55DD4zTIn6P+qtP6JfnIpQf1vtg0Sz/9hRoYc
S/BMDV84ZpegTJm/iPTETwjvM6nj35p3PUNbxrJ9JEJ77S8OirLPP3ucVlKcC/zL
SMFReH+bJlb69V6jf7w0oJ+U+DdJBcaFZJXCBcDypExZ1iULL/2fswe0EDdcnYM3
tdSSYSFBGJktoKBRa75IJx1ld3Gqps0gI8EPOKWcUwip8ki3ZR/FYO8wOO0/J1hw
O29dQND8eZRbs1kYMJs14hB4RqDT7s6F6DEJ/iqyzUkjxkgA62LrEmSDaNgn5Urf
hzc/3qhfSqcGV3Sag86y/CVVTJmEjqJcsFN/resG+iMtWEHUAkXvMzj0KLHC7VES
gnVj7bQfQE+On3cRmlSZqdCc0sftzWOeehMiJ+kb/EuhejE149KLZJwjjZVrtgTr
srHbo1UTvDezA7sEtlSSXyJ+jcIeNIbUknnWbqSz5SgiCC7fDRYDqghVsJiQuEnN
Lk12tZjKlt54AisRC+or9YQL/hf2E7mGNtWe9OlvIapIikencPDsnQ2xu6TQJqwe
5Fk4xhQ+X04JCZzkgEAsjHX4NWg94ZIDikmggaKknJ6+N3VaHntXnEHpoONSY+UT
GpQyeDX1ianYJSW1wmDljtlQa8FtxNU9JxcE3NLc0KreGxI4dGEhg4+j2UJMmbal
Km7vgts/wgw5yJ8FgN+1s+X9J8n31iO/LI1jRZshSrWfkySD+zBncghi6PlYS0RI
GXCg1iEbRxVVxoOoKzFW1QAE+80C3sK17m7wJ/9mkp/KP7zDAOsakoQ3JDD5pr6k
cHwAxjktSbpIutPfpZIF2nKISGxUmU+CqlpVS457cQaJ0UkbyLoJjuNaEDbbOM+O
lpsvOVXvmob3OjogNSdR8FGY4dUIHQ8+Y9rZyYHn4GwEDEOA/s9ASdnGTFLuQyqA
82eG7Oahlo/n6DdHwGpP/Tpj/jO4tmBGgNjk0eqfIyG5AI/PYjb38PjUASOUKKV5
M2Gfp7JkJsFfZAgMq2LDQm8CprIl3rTCf5VyXed/S3p3Rg4t/cjjfuUvkGuSFtRF
P6eADSJU51L9iNlMSdtW5sGUkWjOBmaiPy7iseIT6Pq+qqvlN5m/Q9YL/B0+ABS7
L3K/t5JuVA5gC+kJIofDTPiy+RziPZnrNS0391SEGcDgsH6+3FUFAnQPU9rlM+o6
iuHxiKSwi0ta6SUdo3sF0B/KKuun+uiTh9yeVmUIz/MwMl65SznOovNC6Kzo/ZY3
+fJD0GClDbrXeTJ1WlIxfyuIBpEp8lFxJ8wTWVp4h8orh54C+IWdf9zA/1VoIk0A
yuVXfu72n0LUFU5SgkCcTFtlt+DbVi/bcnJ1AWrCHBi1GeEVPVYungdQjOzOl7qe
xee1n+2AJyOWzVSNTuIypd0HT3QoeTpctf5hmmxdrA0SWiTF25SKxVdg+CeCW7ze
e2JgBD13ohDZd2xHj7j1XrV6dqSPXiML7iTHOXG6d3tQXqHyXv7uzsuVxG65+QJQ
vBjMeLbfgYXRhMTutOeKEZZAOQieUftdiPFKNq+TRl9l/I3sDGmSue1KmlvG9brl
25kOsdZOBQ7rOGdQ2ENDOQ2w5/jc80uLKC488bqvcVWtAgf/f9ztjt4kDvjGqH8k
H84Ui+5JdMIexS1eZ8xwdKzNFRZmdjB7ST1PET9cDNXTEIkjaluKlsvqiztoh4hP
+fDClGmhSuyZlW7eATwuNpNiQaKoJMssgMpb2erHeS68lDb3+PMnMWGsIboH0kWR
3mCl93IvN/9lSYLL6F/V+V+tclr8zMYahIBPrx5Ifz89KDkmFlZbabbuaAvTdWqB
vEbKvUFL3w0y5RSFRw6H6/d/Tj8qaIKD+mmYcBMu+fM6wSK6MVSs9PmNIjwTCVNN
+MtXADjUlIxIQGRB1VAUVZlTtsT0yTP8xqxBxjv9pROAtoaj251PjwEWyY4ifCs+
7zUIyr/6+y8Yr0WcxffNWG+D5QE4HMvxmm+iRMgp8ew6n5CfIc9NUdFpJSpC1kIk
oOkdN4SKRNwcnfCec+pcrD4L90c710cLsbQeIxDlT5zXdvsZY7DRV5GV3yrzUcEn
awIaQDs1w/trg27ghqi2onMrEfFITeafB5a/HErb8IE6ppM5HVjAIFNbhZ0ik/5V
AMwMvB/wYBrO85t8sN72n1XWjnlqlKqLwkfI/ryrUzigcGnwYB5f2lxyJjjs0Q/5
o7SYh10myHnPIckPC8A7cORoebcenxJkU6yRX5snj7KrGfWEqwW9qsfXtm9R5SQL
RML8s04ClctFHEZ+wAUgfzr7UQnr3trRpYR56ZBJ5QECt6x4xfn8MLiXWuz9xlnr
v3Yrjvsozu3gyYEzout7UiqFzVAk/NbqL7oSuLbT8eU/kwaSghP0JXtWJw3qHFQl
+k/LXZ1U+VFTFbeDgor1IjVb277vfmKpV8L2Dxj4Ej1o3ybDYWk5Wuj985GYkMFL
uDOrZ+ua4aVbhJUy4TgwRG1sNiMYrq4z96xcuRn/sAKY6FzSW9Zie5gm6ZtSOkaY
frXVIuKl7dICP9yyLRTOeRzfXSTBnDk8Vu/E3hiJyi0IaYHeeMc/rdT4DktSHR0Z
8eo1Gg1ebioTVLE+O9ctM5hYEnqmbqWtmm2gq/nQkZvFrLvw3neXNroLrXdGbXTJ
vxMY+xPxQqR/uUQW7vlHE3UaesasDH6TUMfVf5xvyGSVJJPenn69cElVrbRo3WEf
HBHfxfcQe3PDUxVpX+o8nhTJUqRIR+eYv2K1feRZY6GfWrVaIZr/JMBaxYGUaLaw
W3yNojIwp6GxrHIgCclC2X/NR/JSd7L4718b5qs6l3I5rSy84p9SQpQoJTixpbb3
D95qVMIT9l3QAVBAFo+5qucb09i81aI9zVUT7i0Y5CWuvElWrUcu6edpdRLB9lFW
UbCE85EoY//9BpYWMH06+acMJjaIwByAOcQd86vLvAyZsMdY0QNnlBclsJQiTnPp
O0B8IzkE3PiqBXWbj8SCVbrUsQjNyaZeUk5CBtWllAcuSmg9zcmayqZgXMU2ZujV
wENbjoiixq8Peanv/Cx9w4bleS5Z4ARbwV8HrLci/FYVXhbrDpHExtes3zNo85lC
ByNKaFKKuKCjsCDYQR5mcZ5uwnNG4Uj9jcWw9C40iO1nfwF5VwvnpZLxVTaXc7W1
sBdV+5nqhgbrcSj40jTP03cGID0k4uaQV7PYYrhkO4MMUOeo/NL6i8pU0m6MAWJQ
LlP+6YUPnAoaFAjWvoBNVeMehZ44xEBhtE4kyggbiIwMNXwSk7iOz9KR2SerQl/z
7DhfjnOPL+5FtB4F95KqgP8RNEwoNuuRQYKJaNykOp1x8RPgtGXoPkzm7t9jiwCc
g7VR+GqQy1HJDfeId7qpkyrljQPQNAxAFI4/gnnIMF4mMfmZ+9FkUqQ3+UYlP2FR
qmPknSvKyGg65GISMi+rGHBiUgW4N+6CcSFjwNxZ4CPfFnzqrqD2MD3yrywBVxMt
CHIBNJb9ej6r37+JvPoKQD3K4s+dQ9OxDeCQJeSUYHx5bu5GrDR7GNDoQmwawxbS
R3cr0XIC5rGc+ZvKC+VE+gVKzQhUwU1LXZHlsjZOXX4n2HpbOAaDyM18dCFLuN2s
M1C2b55Axc214QL0YH2U9/NLbonI22elRYPQAb9HjbmrhCHaHXtkEYzPzZGBXCuq
d9Ig2C2fLriCr1AfFc1nTjQFSr0Bv0vJ9yVXGxAOg1KWsO0ThxtLK8Z2PcqQ2kfo
wd21LFbisEYk6QlM6pPWFae9jKxfnX6r0TuMU9f3OL/VYhHsbWG/9EfhTRIrL80t
Bw39pE8lBDx7FDuV9fZC1q4l91gdhxoU2NEuxhYCoXbKp3/BjtbOG28iGeEcbMPC
EMcDLqhkHB1Qa6ifaLkrPQBbNIBSyhKa1oxu33itXHZvNwokU1lHMMDlogNaNTqq
dYAUld4tyBjXmiI53o7SzjH7cISRGlTb/3BMVNoMkraGyVw/vxI0rqxeRPpOF2yp
KJmfQLTuCj8QqhV6B1myT6d/IcnrgEno1/1dcp4fb1HKT1lYh9l7FZQ7nB8VbgRy
sOuFYjwhGDLkbbyFq01OAARYg7CYDcjIra6mvjxBk+M3l6kxdO09oPQLwek7vFQN
kXVdxmMmwyyCIm+JJv8xgdVEndK9gc54cNp2J0ElWd053js+PudDwwy1fA/D2FQW
VSmtZaK95YZm/qtobzTZT7R8EEgNeAlKJ+PwfWZTErQYDJOEYUtJiZ65AH2ZX8jn
XGMMlz79EeLBwl5LdsQUlQ6rxghtoBHxk30vLda40qxYNo//bSuFs79aFKC5aU05
G2EzRz1ixVlLTWtoZ5g+hmolGJhvo1f7XZPrjkZBsUD9Ut+4MbTTccvdYhZaN6+8
QvQgS6W9NpCDYxis+Y0q32pkYzkhoDEtZeNj11Pgvn7xJ5h0wMiTNJ+DzNEQXKCO
vWq+sIS6DM1Eyofg/Ge//XEdPnPTWZxIeAthMWEjGxykopQkRQLu6xaN8ZhQ7ZAp
fKzSHU7ngFOJR2Xj02Rm0sx5qNWjXZSnRwYMhPqLzvUfdnWHYG9DMsTZg11Wp6QW
cCjIb5S26dzFbhfEDCTm+E35RrFeml/X/FlF6oTGOW6mNvUTTuPwSevKmn904Fhi
FpulgLDtwCrZs8c1uMK/Kpsq+4lbCajXz6WzE+rr3hGhUX/pP9HS2rRYiifc96V3
E3pqpIMpmdZjm5eVgHw5zKMcp7DIK2ZsxOFWIQCsTqzIl+skHi7jOCFtRyo0n0oU
e0hTZrJEB4lPPaILPr5SO1kkVTzcnNzmNhgXZw+kMdV4t/wnX+HqVJa269bcRblA
jzPWWvpxCho3uEuxtPYzjn4DIthHpEx0HR+ZdkY/6P3qjJMcUuEWOEihRlbRFTU+
4hdx4bNKxUQoGDeiiQXiLHIsmzcWzGYngrnAmf/kPtdoHUky+Iy4W5LuRZOwU2i2
oea2+B8wdSdu/Olhtf5d9sCG7QWCayAhGvUqjTo6zV2QTMVZQoJaAzvDrCzzpv1I
3nrqxdqqc+eZKOvnoXwR/CpsVvz4kbgWYPW+hQL2hQCE1dphA/m7eVN577Do7k7x
mLC9RQYHQyTyWy7RSKHENqA/zvheqglnPfI+mKAfTCTH7+f243QOka07XXvhu/IV
T80epsvCb65jmPEw2iww5iyo5s1i10TN1LSxjtND6nOIfnhRZnS8+0P5MvjwAXl5
GE4v/qUeOvK/7pVlhrXPjHyouIbrFEYbiWcuK3YPLXplLmapf3Fi2P+2mA8kaa0Z
PdaaMVRJfqyit3xobAWrkgVdv5/OM7OwLbgKuiL05w909V9oiDcTQbSW0myuuqsr
GdbINvXNAPyES+qJf/Qe3OOFbqNIMeF8Mbunh3PI96hQyV0oAmsSwu41DWLnqHxL
Dpel0wBiPxphl1Nlu0A3z1VkGKmYKUupqgVCgJPJm3sUctWp3mBBTARPAzAqURQA
E/MB0f20caKPTqcm0hotxQyhSx0F6kgUMx8EXfpafPOenTKyImodqSgfrrV4/vqr
bZyLN8Em7n9W0DHNFt97Qy08pnT6PsN4bXI8oGnHepxalT+ZesP041j4fI67r5Bc
7pmw7YbpSZkQa0FCMVAWY5qa//DY4/wVU4h/7rGDSCsdeYBFInZ7+2kQb7Dp8QCj
d3oaomiyDKJIKn8pEEeK24WJ4IIEn+i5ypq14qO03axQkaIm7VIBamrtuR3CUQDF
9sRZUev2JvBaHUslIZUyY9hv+ltk9CNNC5NsJcEEtERqE6Zt0k3WMCh2ilewETeC
+uO9PVXjEudytLRQHQVTztadYV7HZ7ulio5Kceu0ApV2rbw22Q+3t93xypJDha8b
09JPJOwoIIM9fR8ga+hRL834H4NZuWWJ5zqDzZb42KvDbNC+xTrSqPU/r4Ouvdup
OlsFzXOtYTjr8AWyoInYV7ux4BY6nTcRYy5b0l3lMFH7hO4F4OBp/tShy0i4aN0R
dbW14xSvxjkvX4mooTFwORZ1l2385XLL15B0WFkP6suWDc2I1JS65eY5zYlS5R5g
gIt5e4gcpQCNatK0GWF2wbAhKslfOE5FUba3pnPjN+wHhx8u2326WbBZvlDFjc6j
T4xPiEJ8pW1bA0wQGJuVLkLunFQTSTMnMgQfFnVfXAsv6XuNhxOtQZWzH27iJAog
eB71GXGJ9fvarZMhm377P+slpfau/lGe+RMvSkGKHh/qf8ZzQOfIMBORi5mxuiG2
DMJjpETc8uBMC1LgWIat1Fw/Xe+/uL9fKAVvPi5cQKP4NSWXXdwMPzFOyj5sw8FH
hOTZuwOO+4CHJTHr0C/FXcDOyPVvRW6AEB+p0VdR8yXENhVp0AqahRztGOij/ICO
OcF4Fso/4tBxSZaZR1xs7kep9JIzOv+AFZ57i9hbY4rscQJHXjUmF5f52uoi+61Z
v+dELKkoyF4MKVrwgsVyYLc02pfWNc/FSSrTU3l/PPGRvGmfClNxffEeSoqv9Y5F
PVXqBB5gShm8Jrf0mH9+naXMUbR38L5FjIH/1YLN0jEPk0bkeRN0FBb+yG545/Th
PI9PFZEW9KfDe1Bjt/8jYKS7OwV/fmnhA8RqKzzLJribr3um4ELZun9A4etal+Rf
wNvZgbxDLYtUwosgaVCjFT53nxgHCOQFWWcxKOtAFrpYxjZoGE6/g2D3C0H6FXo6
U8q6I+9HbAQlzhnGYmrPZyTuwuVS0fUbXHwK8Rv1y79cirDpcQXhbeQ/fktxlLLD
0hjeY4KEW7nEO8Xgz0607Q2IU21yJisBk0lzmB2/6+gskwbcsitt3Vam4tLzH36V
o/ZiyUdpxGO5ouuMD/oRvUx1D2aXfn9HEIc/4cznndplUZaYvNZ/dVPi/B5YjwN8
t/ZQD4xInqUMhMQonDW11g9/BqkRFzhASzQFw40V0nCHrxOxwuC7rrBvC/whJfLk
dMolIPxzsJ4C6Smvvs2ILOtQbchwyqSj7DLJTnJTFv0vlNZ3pqvTrr/kORcZqffm
GoI5XzCbh/zIvbodJ1UcxCBIcTao7UZI99NYB2mw0h6C1IkrVq/1QRlyg09JP7o3
0w5GeLSFKgoKu0qe3V2xldl8mGkx8xgWGyBel61StV0yb/EpuyG7VoP0VaWaAhhT
6sNBudj9726lMda5X4+DkqGTuRd++D8uQZ9T0S0FUgeYKd3WgBRQP2pNYKDLFQEu
A7BvmDAWSNjslf1yviIIqxpDFQpBP0gA26sxKYPWyLtyRnRIlM5kHz09CJYhALUM
66HKNpxenZ9CiYjJuC8vq5h7lZwIdOt8WytLv8NgwEqHTT3gGmaKYcp0FH8cI6tc
/k57OvZOEwkbsm0URxP93bkOvGPOBJaY1884cnwXnGv61BoZ6i+Shhv5+aVUw1FA
Sb3n/UwgLCCa2DFyhqZOw5GPrxoG4w1P3HF9A2Bdnzm2isvINYIv6ZahtVZFkomE
jcXkMwnpxhTY2mhslkTzn3GTdGfVNQs7/8jDF45oR2Vj/0RmGke+LiadgdiizQxN
LLZcfnVf6KmFIBo4qr1d9JvkkZmbc0F4dpEL6/AoNXXlwKXvGf18xS1s0w3U0WZN
32m+AC7W9mR5N08XD6jWZLWU01P9eQg8ZIk2ffcl0LjbEiazM8kUILGCe7TxLRF6
naXdjI9Q7wGY1BkGA7m5eWXZfM63a3l9tN9T4VRjrcAewSJhkUmKQLidSxPo99Du
Gef6S31ptbM8rW5UOAfiWI0mAcGKOI36PYV/PPj+QKKLrk3k27INlaiuJeDGSOnO
MiS/hsFW00+AHfqqYdH2MU+hIR4fS18lq4i46T2EYYAea7R5DFMOhmv5jr1G1AHH
yKeYYcmo8Xvb5Il1HQ6QlDkLVSckAwUgLUDFKL4Eh0Y3J9OvAN4M9tTDm+pwNIY0
9KUhR+NrM5mJhXzQLLGOZOr8A73UPpXRLFXv8Av9W75abds1q4ZZWD7TdDKu7nwZ
TYWF2s7dKHm+6EBT+m2gsMci5dPXrDPhamD37k9u5NrFTSNgV1w7is9eJfpccs1H
9RB7phMQQ2wXTWlgJLpkAH1MBWBx5WX/5bXgtCqJwXtXwwyj+/NmsCEQrYtlQbFT
1Z3cjquAoabjzCD2KJD9DgaPynVL/Y25Z4su+ChJQ51H4cZVFaxeEFnoLS3RGxaY
cjkoHmHWedVTLyMl8RAwh9RFwKxm11bVG4acB1UcJsIsZBr9x13u41HxYzGPRUq9
wvjqoKjFN2c6wG23u5iSDpWDcSOAfuJUy0mIfacv/vavkCCu536aSm8oEHvdfGPx
kw84K4zuwEpytzLfeA149S4Ks5xOhVKfEZQEdz6zst/xxNh+6NzNikWjsktfmhiq
Od1xLIaT1WZRgqB80jEtzGy+8bGgb7LyFbSrMJ0ERqimnMiq/lDayulLbB/jNNYw
Ph8Arkq3TdBZEw5s5VEkndZp+smfwPuVIbMCHVEfcmxZYeZPiyWsDcKiFcGHBQwK
WdyuN74xB5+dGC0BUhz7LSkX3OeU8fSpTZxCY6pO6kGzb0uQyJFcPcpKRbOwJRPb
qEZjxFTF3fU2qArFVxrA3ULSPSl5pXejyzFwPZe+R/yo7KqHM/aNqyxy3dupgWd6
T+LlfGvI/ny8m52bmc/x+rNlB9AWCp7Jsy1hYnO+F6kx73VRZN9gS1RwFfdquwDV
/dJUfv7F3KfHuGGscbIGBP/9mmsjvhUJ7jCJ5l/xkbjWQCHDFO54/BrK5uHJAL6d
07U9yp5nQtwmWV9KjvQyLwhjSS/9vf/6Rd2TB7RtsxsnOw1QGoTD//2cHiHJMpZ9
J0rdRatsmv24rJCwAv63NsCqIj24Vd5pbwomQtAJYR/ByGncZ5WFRqI30SthWlee
/tCRMQ3OZ9i85KtC4Rl5RwZ/pdBOENxSvieIcQHJ5FwJJW/sMeFJoSuiRsyvPXRp
giRDw5WQGfEYSQ3geILpofjaWk9Nbo42p/0FRJvuH8YLOZo7eJoC83CX447la0Gs
q839+12KV/hGZtFGXnw8SYfPWPNpRpBlFVNWDoSPG4qxyJqOdycbdoaz5mIFMuOR
ud3mZxteXENcqMwH1NgXHuaPWb81oZa1PKNAfOw6uWKIS2SaauLTzqAhtUJEPGcD
ihNAGlvnpUDci2WB2nnR6hMT4XpX3onhzpS8rIZ9/D8CSsf8KMSmIClr3gvSLK5E
TZYfov3/mzReCE9TUfUDkOEpOfPkXvAUyH3YLKS3NukXmbnt8bz3y9fDJD6ELMlf
K1eXvhb1SxD3u7yBYikQI2P0wZJ1L3sn/ptUqTj0NimU3c9mRDDwwbJ+M08auTiL
JPGc6L0JUqjZ8g5sgFldVkBJpil5g0jkFXBqOXdM7q1xu9l4PlexqgTOHjyBosMz
54tgBjq8my5BXv9c7j2/u/WjlEOLNdxDXRbjOHhh7FkF5sPzPxJ7AoEgDvAjo/2d
/Es7/tYxFovKgGesHtUI/XVCd5K3K7p5HGer9PDRsvg3VqAIwfR80sCw7raSpmEx
N+CfNiD3VGBlueqIR72jeDgEGSehwB1lZpBvSq47qpUTq8rXmQB4AzTkY2LVSEI7
okKN+cj+jW2+mh/fSN9lIpsuFOhDG8J/v9lELfyq+AGNdb3WlkJ3cAEtb4iyz3Ob
4z7S9bE/jVTNe0y2qKHjnKbwiVYkJCpiu2UEcti39KoTGhsYTc9bZWx19cgMCTF3
dgRe62sBwe4DQF+EBJRwE841+Pj5URO9fUTi7DN0tRvDTKxdybBs+4TobW/3VEbr
3jJ07ir3ls6cHA9hcZrDTm8dt5BgAgdGGwYp+uh0u1Ld7C4hUvcKGlMcfG8hduXD
ErWGARmjzrwvZHmtlamQOCFRxk1A5oT83nEOHdS5x+LORAlAyKtVRCfeTztUuJGZ
4CBwOUtsSwa36qWM+W9g2NPIeNnMxUcGRVwJa6rhhau428AEJKBQKh3zcvELV5az
Vc4mTIjwfIJan6yKG3DJDphxeXX+fir+eEZ/jY1fgJL8ivGh3AMgCGEHWuCOjSIQ
stoxFEcLwhcPz4LoTOBz6r/Zc04nUWJRMvjKPkEXgtCvyOB+zrpzfnJurio3REGv
pLxquRvyxRukKoQg2UnoH15NF6LOvBheRRAdYw+YsKqJ5ebYS9uedL6ZRnUXrS79
yTYnL4JLyCmg+FULk+dcPiGjC2gchtMMNcyBhNvj30Iq2Lho7f/ezO028SwTNS4A
/raFCORlwyAkZq0Vnc0frwnxsLkp8I/OO6LahCmb82lRbWCe0uAwmguNyu+KwCGh
0HCRuJqiSxIGCV3fMw9ma+Wrn9wHM8A90KzvlVthOfZnTIlWMjMldikWN0RZSXAe
SXVdp3zLi7y/fBR4g4pWGF8M7nG5mJY8y5zkSN4TM//AWm2T9EbeyrOofH1Yz4F8
nTYz6oy7ijpTtfORAgCBIdduGDq3JgSUnbP1aUXXfwHQRh3j0MUNAI5E4J+FlGWS
ZXQJVog4M9aohL1Pp8TJY3S3E0CCdBR2f3imm3Ipb21LgxYDwe6PszKiXMnHw0IU
85JieRw54azf4IvPEzzddiV4rcc/pCmW8dUt2UV/YhAJd4uy30c4XjitHEj6ep7N
3b5HBdNv5zHrrnzaPv0ZYCZ2WEjxII5YD0H36Plbkd/5xcUqjmopspLevFK8MVrL
bBL+9B6H8tYdKan3cBf9VQGoRwqzE4VYS5hmWpzxpatQqtKxNhJBk4jZ8bJdTwbj
K4eYus3ZfePauPxFUluMcbgsWTu2sDKNJw6T7KFSnXpxjaSl/fQmqLYie7JyZXAT
ALuHS91fXAA5Ij8205uYgrk2PAxiZ/spyA3XepbBjUj0leNIMsBMUniuLPKQrKnw
Ap+/mJK9gEZXswd1/6+iy77JBRD5ZZrpoV9qCZmXzb0CE+H8wOMm5BAT66ztQ73W
0TcwaqZyE2xeoVOp8jMeW/t8/WLD0wDLQd5SsaZJq6696UugQDjsHh96anwmwlqH
zgF9Kqo0qQ9Yo7YZofBRQqGWMeL2x5H9AmfUD3NRsmi5F9847l3QyPLjMcncwX8a
2ugVucAcAukSoYnbGLGVd0NbMdfIKuteO7oq0F8DZJ8vi9xGRk4mBHHD7X8rfK4w
IixNZ3ff+gjfHiPqhZNgMcyZRZc1OhM9xxNjvBfwzYKcPM7sqx5sydOQs8zqVJR4
SjqYP/j+XkCFBqM4UJ2IP9eEkE5UanazM+cKpvoMlY+Vc4HPBbaNzKKmss1yMDD0
7NMYa5GdrWn6tnzeimTGYbdNQGaDIhkr0lyfWYqfsMHcW4w7bYzo5o9aYvMsoaTQ
nwrPN7sOi0c37usuGbMBHGyHJMm/XyE4hTP8cymwlq7pZJjKxjSOciU7mIOxSEnY
unOJNOV/MHFW1vj6hNHo7eEST2QNeaphQYJc24pRbktVfZq7/P4pjdd8a1nsRXW6
Z7CFgwz0M+fdPGnklrl+Ct8OOlctumG+e36iE/5I+PihhIT14DLUolh+ZIb+xHfK
iTVp8cmP+sMvrzcEIi6sLcyBUv7QAU1FxTKZeNV0JeXLSeB14KLvjUpAjEJzE0v+
WCxiGxTN+qUsOGn7iCWAVEqtYwpywyOIZtdHqutYbuUEbOPD5CYtuJLPw+Co1StW
UINSAr//fbf6dfFSAtYc6656jDqFyZ1ewQUflFQs1ZRwnbwxCRP2yjZGs939SX7x
Sp4SksBJuVWDiv0K8KjuGg/fPCGw5HRxKvf4ie2YQK8AMOJOBP4gXeAoIVFf9z+5
lBLPv4gLrRKb+ODsOGXLb8mlgUIFakMNWyqaGZxorswZG/OjIimV0UeCU1+7VTxS
0C6sa9Gab/CVD0VvSFu4sgsNiQ0nV5m4oVhnhFfJmVzB1wmuvPJzwhPisPBxC6Ym
DnHCu6ErbSaJW8UU8/xbiTOuF0AtKv/pnL6MdOiF8dtnOsd2VJckXrMgPQafxwEF
ktZaw5LoxdlBO4AcuopddLqxWkpvb6jjShsSGZPinB6NZZr006EdhrX+tQTYXW57
44uEMm4+owciR0vjZtWL+knIR+zy3LvosKkjuXXBhGbzuROt7mcwUe9XJE7pvJDP
vCylgC8IU1cfUhPWI2PTXz+E5YaO744KzsPWKjh/b0j7K77yYtMIL6TkbSHDEjRi
VGxnWsPhoIqavv0C1M/qY6aHOXt8VWXNDiBQ4nDN4qIbD5/d4GxACvSeBL2cIlrl
ixASHWDSlJkpvYpGvf9XyJFo7M/5BMWILYUjlROiGnmwLYAlOH86QGW+gqy+jSmf
xHto56KeupsEL1Nl83AJliePYNXgKlzhqvak/0sUjcDlMz4cetJtR1sB2W0ETZDD
A6lZKY3THlTR8fY/yMClkeb1eiN4gjNgqn83ZkR+vAY0Y2UBpPMormPvKqB0F5XI
KDfIkirjdW3a2qxUu4IQ5LXj6zIULf8igVQmATTF0/gQ21jFNMGlgR5SbbmcK2I+
dtVYpnb5adP9YCwHg6/nmL0I43ZgqvvRsfTjwqH7/uPJgOojpC3aeBagufpK/JH9
T35NqZ0Gf73UK1+9B3s/zG7e4cJ5hPse86ydkL5UjaEuNmjb9ZzDrD6Yg0rsIc7y
5Ku7CaZUowt57lg4qFnlA0Ym4sqkXsja1t2VJjPjZkKTlNu4XW1XBdW7t8HuN96X
JY0SW0fPnF80M0hLLJ0AvnbpbdDalPV5G0r9lWgMdRVqBwcmzkpfK4PS61/jTH/N
qOIh6a4aCm9LRZHLHqKNOc3KQyX+EplEBjXf1h4CwxsBRvm3BuyezBULiM/Qde6l
bR3znO6q9JpVeB5YKHep8sNTtvuex29vq21c7bMtZwxOI0v73NUrkD/ANN82BswK
fFH+gKv+OY4Sl0BxZvQL09r/8q8Wh0jfcGyheJG3UtejTuhe9MK935QOJbKgsKJc
HJBPaSYiC9stpp/fWmyUYOZ2DOTyrgodlmM7geDuvmuzVoX4lpQjhIU51lLKM9Bp
LsPdx6x7szbfPdJAO4gq0DCIBDsurp39co/WcWpKt5K0D3yl6FKrnKobZok0SJGp
N5hiksGO3p5SRzNCnTqCCcVzXr47XhbNY/nuPEqPXdXWF+4kJ7EvKCFlLa0z+dil
P7IPjWsse5WqCM63c4h5HKjp5e3dUfBONg34Y1M64ylMxGngKbbTspTD4lMlBzYT
CK8yF8+7yMWSe7XqzRol//pJSYb6b7yJSCCleyNPvktiT/ibP/l4Xtd1jsCeBEa2
gCfhkoZfG2rZGBL0jNkW0QzYIxaELAHT5CdKx+uRKkm/qCTMf4iTHYN4BFQCLg96
04pZVC+PlySIS+4BDuD5brOtJuSCuVv1OQ0gU8iekeiUPfJUT4oIUgTtlt26RcPV
STb2bC0at9S4Io6z9vwhESrc1WMF0sZYDbbyHk0kgIauiUDoPvCtXQUmKNPJJUrN
Ueh24vQNz6aQHQ7+VEOh/dk0cZr9lwQ5s1pb/ybbC5sfeNo+bNkWIPgp2pQ3+2CS
Bi9yLcpdfQcGRIZG5MSP+DORVgFi1Jfx7WdZ1CvW1gjmzao26wre7PHHiCtjZbRR
+o4iwtS8IioxgTh316f8OEnL/X5kKMpttep3kOI68X3MAhhloJAEwjnrHtak1p3A
MBcAok+aq0N7AJpeEnBqsa4R4JBnMdd0lSkV97ds4yKCjc7c0OmD4TqPVplksZOX
dYVUfJK5xE4UA3XuDYpN61pgV93iBGDwovaWCnWD4noAKpqqxXAWRr6Cxzql1m+g
DSF/nAOodSkv15fBf/6SBa/JezChXVjjHYT9buOWu9gAMDY1ewqi8oe+MjR6zZpx
uW5f38otd4KtOzsu0Gsew8MdxLzMUWj2yBx4mYxutT68gNPFhcjU2aSpgP60RLgh
CcyUuM7+ibZeL0gbEEmBioAdv7LoHdmDKYYKmXo0rgm1e9KdQwdUT/l7MyzunwRp
Fn+mJ0YZpxT0aJn5gQ9k8pfnARUd+2saXYK8svkd1uymRKJpSrkzlMNURPL0ckZa
FMnToHsU7QxzfLrTWFDCoWKNa1lvec/F8Ym025kYcf1XAXw5bJUhRNPOg78s4GPJ
tUgybEeBB7SYsU9dzkoEN+n4OEB08I3It5/a52lVerZYwh8YuUWlcVVe1kpXo/wz
B3e2uRdZpBxr4aGkSki1v4bo0zEMrCmOxemHySa4/S4/4FmXEWicdf7lZaAcz80a
MpSYBKrXOLCqV4mGNeVEvi5ecTBaaf4P+F7gvZTcCK1zl2TPKBgHrDbkhYXKamci
JiK4tYTvwztmraMXutprzYH9AG4ZuzKRD7l0IOLbkRZMa1mE5GwnGKsgaFBCWGmV
qweaSLaCQv/S/k82J3HMmwRxMGoUS8LA++DnkQebfyO9DQejt2gK8ZLKL9tH5Tng
CJqK0sYW6dVP27XJkjRVZocKyFCfEOhKSZ48xaIC4PvnPl7gukNCrWXMQOLzKpEb
5INW4ZXCUnhWwMBjTBMhsUwTIJGc7IYHk7cXoU2Ch/jTv4fUkY5o33FkYNuAOWs5
qvAAy9Ae3gqMouEK7H7243HosLXOmznUzZFAZjIzeCdliT8LS9GofOiTGk/3ASNH
7F321BhF84hH/EFqtdEyNIGRXek5VDRVjPRt1UAHWLWsN9AxJS0MqXHo9yb9nTxa
+9QtyYi/ch9v9RhWZkZhf69oZrAHSW9AtVM0uxNoH4L5aAiM5kO+uHqhagKEtrML
UuWXGYhNp4blJadsF+cjBapXkjogj+sp7uB4kNu93dQT/xD+tt1Poydndl4xvJOt
IYkfspkEV5oFZqn/TsDyqvhs4OScgg0BncqPIem+okGhSq4LRGKSzFlfY2UjEhgo
jxNciz43ha1k44tlBibjkxrbnySX+2ictbqErUsVSQ5uxl/UKU7vYRmVhMUbGVQh
SKuYa06ImXdspktmcMCe3TBhrMVnCeejpd8Kw852zBceQcaC+GrPKQrD+RVzEfip
s+JptmObQFBR5tiKtclV/qUe7YllXi6cvMqVKeg53P2a2MO+DbOIXs/Zd2CJkNh2
0dpZ+DEX995vH6XYusXA07jl0XmPEplW0yV26U3+wVa1GqyFTzF1PxtPm1WgA/j5
9wimZKL9mot0jk37+fSYUMuhXVtahI8hPdZ0KLiL4zjl8E33iswfpiZwEsynErle
63OuL3Pf5DOduFbh/yDiu3YhziSN3NbEpm+tU1dm4QPxUd+yp3v1NKjLBDw4HmJr
yY6V40VYwZnh5N7GZyasylfYJodjX1ffz+SJMbVR9ett3zD7QbX2D60+2uJP7/KK
+cAugOnZCayNom5iqKnL4ztA0xchTbhkMbM6xlziR00UpZPjnkHsYhjuxuWZ/ox0
Utjs1V8b4tJUYcM7TOUjVSmATvpIGIN9UT7TKLXAdxW5iVdNFTYZro2SigzcJUgB
U9Ma9iCkArSgEkRhFdptbtH/FMBKEnaCwvIa4Y9ejEZcGdrZSO3Kiy5wrT5ISDwF
ahYmVc+UtWuNS17frPzxYwzgs8eqXAGDhN5D/sbsp/r4E3QyoBaLisMlixzo/64K
J3iJYOSrip64wqFfWUedGqJvNC8e6vlf5ghOAr+FDI6hcuGCg4nY1U/5YWYYOKbi
gfRZ/UvxX7YUJnokqFvpN/unRohCOaJpFmqHN3OuIM3lQmfONjfEG3RQUkmtwZly
vRmxnHg4l0D5Ki7QnpkwnsS4gxtYSuhtT8V4pBZhTmHekqvZ27tdyw9nva4HZRpK
8y35Oq4n6y80X6Syf9EWR/FRgkmvrdt1TCvL2/caSL/Qce/8ForBvJ6N89cOnHOl
mIe+Uodhi+kk3IgBiDb4ttaOZULSzjjw51/B04m3h7O6v5ZGCmxJneFXZ4sG2rKD
w6xLdymADxdXDuKW6IUYkrGpciMXZ9mfPYGkws6I916ekD+ukPi7ACVxhBAhkuMb
SzL/eHBOXH+ahTvAOfA7osiMG/uMuAsD6dR/g8Qqgm5uUNZlelX4nbJMP/QYOI1H
xi4PHjl1i5xa23JHHtnycJuB4FNLDzaIwqlFGawnZjdOnyL26cZMIV9lv3VT1gsx
t0LU4YREyHl4rXdVE7k4a53S1Vchf9sYCAhDeB8/4L0uz9KIm0TvI7/JHngvBLRB
tVQsPBfGhhp7cgr2mgLiL7T1yn0226UQ0noy+F2jpNSJ+JQYdCHd/XJWRNKQdlwF
p4955LqzlcwCMdmHuizslffe2pT9iXH6DrAwAiHo2qVD9IFh/ddAjgZUptbyBjOX
elMMslq7pneeLQSO3J+/EjMBhSUNq3LNjIbNp6UwCJEenuml4T+GvhZWECbQ2SLT
1d1YGe54ihTp0FJvoT/4uOXjaKSXH/4z8QTeANVd9NvdYpnpaUgBRl6j+vGC8MVM
vgsLcVDXILBFUhGIDYz9MUFNbsqFLqMDfsWZK4fE9aaxk9iHX9Rk+MIHuQD+GeG7
Pdtf8Jujrda9JszQKfH4GprBM0KcmqGvaSNsw2MY8WnpHbI3cFyXwhzQYpC5keSo
OX270WXtlzkIINlEcUrTQmHpA8iVPw3HIy9PfDVQYNgyvkyzD4I8JCgOV0F12mZP
Pg4k/GzINwV+XL1eHqa4r2VknzB0gZC6okxRpKsX862sx7In9E0M6bX9yxUdTGig
0PlEjVDzdkwz1OgO+Z3emY3Vytr3ITvu5A7fusUBRJ8ZBQovR4Md2nEPyLuOyp9l
AN/Yaw2Chh/NBzpY+R1AwwEJrcd4iNEdOIcGnhSGO/oK+dbgPZp+dT6RJY81GxdS
p5ZtXutdpV/hQb+i1uyY598ZuwuIzNtDPiGZ9tXhMM15gS/WUM+xADNrLt8JWKWD
TwgnTwteK/9qRiIkDwDJMMSFT3DUDt7yXloRbzUUkndORQAn7/uiq++cQv1GDaH0
/o1jTbwkYl1TDFtGCIPlZP6cS+qzXPjjetbUMc8m5DPRQyTTYVW96D7TvYc7jGwS
mK9JliDowTB6dgiRvh1+J8IXxwNEVnjIhoMyfH5kx8/cXOF9TyICtYu79qKkl2Ej
Skk5jXB4XdbKfnmxMXqy3xpRu6BpA00BB06pkI2w7WyveJKqzIL7f2Wu5XkxMTuU
gNzjwRDfH4KigtV6/+VS55JYjoXsZ5nEpyMuDOayPC7a514Adk40aySLXuFRvU5D
9Y3Ut4/P4lzRBydjdJ44KvLn0mdwpJOs2Qkt2TVbafan/QsheEQwsrWU3dABxjuH
AxvrdonyKERt2zaf5UX6K1ro8rN3jRt+9qLekSbH7MbMVXwv457iOKGX+UQz9UJN
ufL00OCTYKX/ScjPC6ElRpn1Jy/eQBvJ1qmqxhm60VnaWFkK7w8sTjNPQqb+XdXB
Q4kuIvzP4itWRAQ4mYJPh5S+Sy2c5LRGC/OAKlCoww9rxYVQg9ugblPoOMAKQFv6
ILvdbSosPy9iAf8GLMp6bLlQ7nIYsqSmLT4Y0RFajgi9LXH5SpAwfNEV9brKSTKi
cuB97yFR1XNyZVvZCBVDLo5PCRVXCSxkvmut+TAciCXG2vfcm4fJPktiWoTRSRaY
WHu8lXZPFpJ4mGdfLhvlWW5ngNMuEKFvgUUYR+Ajd8KHA3efRCdQPE3aCWJ5jyg3
4wCBVn8sBBNMpOBScD+TWQcPUzVujnMdu17pE0dlpdAxRTDjMOWdK+NEJ2zLJgi8
Boj9BhdVMvbgSndzp603M0c7/AkP3oCtRPzgSKkaFsHtqyU7qDajkxUeWuscri/T
TSnf2b37fnWtK2agx+TKcBBFUx+U5RHH1i+p+SvDYHk2OtoLAI5VKSchS2Hlb6kC
x1/eQvTKaeP9mmbt2QzD+11V7xOrEPKT4cZH2387pMYDGqTE73m15tnDyScwhtFk
LXykuqHCYSNA3ktWLlAbzeQ2a8TXf9FsJbCOAyUukQXg6x/rKF40U4GWFd/FMbo+
8PAAeHNwNlzthG/MHJTuBZWJbIiTztrXSUWbTnhljkhgBAEMrDASxDHTbryfvwj8
SdqPxTcjA+LuCUjnhFnoGWVV6qHR2gH4Y1rKUHcsBcRWdj+aEBtZTYR6hWikKeYm
KMa3LPMPxU9vb/4y3udm0BykDaKyjE/uRtmrxrl3AJfNXvrrj4kXY+eNesO4ZPPg
ZjOQn7EKXLvETIgAKsNtpoNaWB7lZCiRz9+wfdCCFr1GdVbMG7DANoT/btWeKq2X
GC0K4zICPhRbNOLxW6nGgjoktYFuWHyExYDkFEuA3IiE0tQEpfzlcCstR1pRP9Jg
6dV1w6+7AcqPDwkXLM90dS+aK8DF4T68LmhEhoxhe7P+QUHeJjyxr5sext2MHwwW
4U/DU/u93jZDEaIAJqEzJnOxhfOzvChRb4OfvR931lJuuQTSQGRXnhX5M8TbTFkv
PKAYFJ8TJXd5mKZluxXJyhZy1LzbDqaijTEMRE43ldSBrNg903+iCu9V7VSuXkxN
aCDFEMOXjANxeUn+BYWrpZl/F3fAYd1mo1cVeLgBTLEUYfn0+MxtjBUwfuV2IEE5
jXYxDLh2hogXFXIkQwaRYkUlb0YQz5kGN/oBrPdqBDXZ6rb0oyXc85mpr/38xIJS
OgkX/BDRsIz2KrJsoQarw9e9VuXJEP7bwFGpiHD9Ip4/FgC1ClV+XrGCnJnFN/Kt
ebuYOFYGaEm5xGUKK1sIBghBE6U+Z5XmaWWHRT3IDaCGZ74mcPMfJ5R9/iZjrAto
MBx1wAKiH8Cztz5RNXn+UCYycdO7saekvwl6Z4y/ZeWx0gwmoeoGzotKTLoHduI/
CJN8ZDLOaMk5mRRaTE8rmJGqdpvHnqhE/AqQasyhpjCWrbC+dRhJ+CF1lEa/4FQE
a5qiHjVtgMHCMnhlZ3Ayub5dlV5ZrdsPBEM+gZri25g5lvICSm8+T+QfPRle/Mym
/ddyQ7hs+bWzXZk4FicxVPsmfrY9rr9E89IS/EQaccGlweQHUcEkAuRYKfrGnHSM
Uut18PvXkloCb8cu9o7XojHLsy1Qp65ZujFATH9iRfUmKEXBicky+0wbtCEmrE7V
6gNz4XUvimcrIG3XdQ7AnbgRZHSmOsvCgHHWV48ZO1Cc/Xy/O4nGhbaELq89ys09
OT/z9XqH5hlj50piG+tnhhojojrPsi1p+HORLeVWIKZ4bk5OO19uYD1zRmU6OEAO
ST+AJzE8IYtHx/Amkl9dCxznF4QAPnyAIQ6j+i/wJB1tNIOv6Wi/kNC8CCbLfI+7
sYHlfbPAmA4IqPIujROko3NtadnN6CgmE6iGzVYdK2P0MV8T/ZozfNK2BfU4E8mX
69dcV6u4hHzb6Q0yW4NqHqO0j/u7Md1YvBXsHH08mCFkAgBnxbInCCuwNZhwv8kM
PEBI5FUxl9VmkUaK1SlZfwvHa7gngLyARWJuTfxRD8cELgUylVg3EXfWgH9cU0Xb
XdVNnZ5R0nMnWzG160OEPUoI1vgOhHccNYnITm/EG+TcUsUGtere3xXflOtK2Q9a
lXOeF/3MqmhXrMgazKSbaYM4gcmJubrtX+04BhLRZV/lG2xe3e78OW+MieiCgv0V
Ojh5LL2BbRtHpbkba5rYvaqAQf6/zScLJOtU+uPkC5e7ACBLcwVblDvU3aR2izfA
ZPEfeowADUFoy55K6/kGvDTF0ncsmfp7qVZIew6Tfe51SYuWsnjar4yXeFsMdVtw
QrdigxXBlJoyHfsLRolBinddJoxQ9R/F6avUCCEU+NoCAuyJtAoy724FnUjLpF9R
t1fLK0syRIcbq5+4C8IFLYWsoyHkMeQvbGYNNpGOtt9PwB4l2ypwKJRZpnp61gmm
+kvi1aXpZxbrzP66V/q8RPDocvhDW/aIcOu85wiEr7h6ieHt8yufevmYs4sts9jk
7b1PMkN1yJbUwOXRUvxgjIvxg2kKIl1WI1DsEcN7WBCzLaLlnCa/CxZ8+9H+WTBE
bTX2zCvf7n0m1/Ym39WTTn/ZdJCA+PEPFTS5zmvR+/4Yxc5rWC52Wri6lH20J8Qi
98R4q6QS4JFOdb5DGcIKiVHY/G++p2eLM6BGE+3+5Pudc/35FbPtw8dHitt8SIUc
x/CD5UmGxNqipiUK9aofj+ZPCT9m0F2Dx7PMC6ZY40TsRfabwdZsYsz2ZmN6lQxm
dWAY5nJ7rq1l7gFZ+tbfxFsn0wLNX5VHQwQlwceg0kU2lrDUfe+g+Ef12AM/9rHs
kWA5CCMnxwoQhd8L2lLsOyrNqvdFDpQLGb0b3s7a948N2FHYuupwdDkmfq7FGX8e
nz9KGByepq3nKF9t0O1GhunLkvl52GZxdqwpL63rSL6yLfS88fQkV8ML6EdcEkZv
kRZrmr/1XvIMBisEkph6gUKVV23dyZZ1KfEsbGY2rKUHSLCUoms7Clq/iU8n57ih
bbeJ7uDuPy/1Dnm/ZZ9fajMBUygDzGmDQZbLKmp1ufhHaBY57pJnPch9Fkm4j3bY
tEIX+kSQyR+pmMOqlIu7u5KJaCR2qxsLKXMr78wH3OSMhq8vxtJoZ70PH2cc3KC4
bB2B2Wx9zXi6eJYsmgL9CPmK79vtMkrYLN+tebnNzBjl7Qss4N3E3pc4oVCnbHQz
4fEbPUTFJtKdI2cwsojlFOMaCFqyDrET0C4KM5wO75wkb0/ljQzW2sNcupHnzk8B
QkuiVamIEvNhCO+klnrGvigZrWjCo4cwlyCs8fI9k5d927werXz2vH91frd94DFK
qyianRWtuUD74Lh7TuwacF+Nmece3ufU4IMPFQHamXkgt4DRGk2XzqcWljFov8Mt
YSx0ZMIT+dyxtEBNWR+f+vVL+FfQSkwYCIBqsqR2ZWk3I0KCsLHAn+YFdn+HBqZ5
8tysdSmcx+n1kvwKtSpKGW9lHMCiNr8OvHAGmMamyXDkP/OsXOKAOE3ichbe1Q02
HtSH3Ydp67dpzWoicCM3BcWO7cU2NXKI2fyktmS94/+SiOGMBDi9NKj3T9NpDBeB
TdSn487o1UBLPwnR/konAcMQe7ZEdc/NA1rDEYqboIqT9TwJ1mpNo5CIHGJWqf8T
H3WKRcjnzPu6qwJrP660o1+E72O8HDNM5gO9DnSEoz66G67jW/eOSXEyVXBIXsnw
/5gU5Ppbx0B4f7hsbOps9iZXxqc+/YHWBQXiQWCgLOyz+nhmrURoKxuL5573HCoV
2g3qit58D2CCm7n9DbOh/GzPY0rkJSssYNeZmt//qcD4kLHf9myoVSZPQMy7XdQG
dkp+9an/pVmddUfzfEMO6PkfUBbt6HONxxJbLgn+LSi8RPedMv4xaHPyI07YFutO
mFWSnz/xzQx37Y1JJW5YVm9ZXY1dh05ozeGR2A6h5Wg4DXxdj7AArIldbjOQIdcR
PTMwi+/4JNWMNg0XsoA2NFiBQkCpHjhQx/wm8urzGfhkn93GtYS1ANSHDPbtlyoU
kPeD2vdVujVIyV+N9PIsLOFROKRcK49HU7VIDRWGbEd+EDbW54W9xQlW7z9GNxbo
xzgt9euxoRZ5bXDCNRV0C4H/rimR1vD6fxcDRQSG3Bo4owRq9eI+0s9t1Cdtw4hv
eryjNZnOu/1eeKVC1XRtrWp8bx6FRNFY5CFyfbpZcyKPoYl+IwbvCR7gGmb70KTS
TfbquhOdCXEleobidfzjY0B1sCYMijW888b8JWb1cfjHabCqoRpgRpu7S3x4ylfv
c6bGxeMBxFnKyKA1fw9xKqT+HeFWxMS9RzJjyKeG90kVpZ4PwZKRIOqqCrGC5OOE
wo+w8MCUC6Q9s5s6VOmcCI+/AXJ2FpmI5zQj0v8uXqhjftuYCigZBBqT27RBIg+O
nB++tTIq2A7axKFvv0rjqpOGijb5t8K9w2Uq4t+kiKVC/Mdramvgbbt7t92Od+K3
eO6x62iqEN2EnNSwR7s9kTC5CLE3RL37l1AFcLdSm1zQRTQN9c1UGyp7RKOcvtT7
PBUyE0EXC6/R3/ie7kng0jNMxKZpmmD8R/9mUQnaCeNuNSgqN6mfefFP79Z0fdLs
/S41Vr9rG9Xwdo4KYrfDXhiBREpbzOIjic3Mzug5vPNdPZ5AYq+WynFjGLCevG9l
BQPEX489MxiIe+ppKFuqwl67K5hJFjkkUN5Th3j2R6yhSt7jsgKaBG0Tjg/Z+/jm
ZtClktAGMywkkPZaoP9Z8men5Z9woLnaMoU/WyFitKEli3Po1GlXO+aDGHlT6Gth
rc2VUVlsTdP27NpdptHNo9KvNdqZBQgUOBXpo4bI9GyDAQATIGZ5ImWbsc+0WBhV
5vlEIHONeG7gnOZ7SrIbFYsZswOh1iCp2G10v55h8zen+TwXWntNOscSHm8fSsRa
1qRMfzYf81oQRC2BJ+NQtbeU+gNLFdSC8s7CL57RITEme4kLzbTKkyPAmyeJ2eW1
tkRjkDwBZz0PiK+jQFz2iH6S1jiZ9DYzfWI8KUYzrj/Dj37L+Sw9qI0foz8FY5EV
ZPHAu9+nHVLHxY53zis/o3RlKd1zi8JGA1d34HRd2DoXrQK/72s/o09Y0NgFWAyf
dVDdIxf3XaDb8ronTiVl8WKjA4tm46ErBMPJprhNlK10xTitXe+LP/kIvNhNDsok
dxaSv8LOBAlovYVITIOtqhfXCFV+FNhCPHJSPxyGmZgVAccr92fEK5tuukfqP6rN
6SHDLf/28e8Cx+xMgNStfn9FPKMrDK4iT8uJc6WGJ8XzG0FHdnj9PdAsRhsTllGu
Of8iqZTpg0DYyN2wRRzSKJNMsb6Qhm+RLFD2edCYe0IGxhiO23alEPjQ1VggVqaP
+Qq64yP3hV8Q/HnIYg2WHE07QtgKPzKzh67Epmont4pk/wpHLv5ymFGs4Y6m9x2x
JTlZqMRr1Qy+HB3WghiWMy8nF/TpG5eA+hyEZQWc+5+IsiEy8aKb22HtzVT/EgR5
HppM9BY5X8xiTVU39Sh87uuVLzjNvF8tbINK/hO0u67wSWkOPeRn5T5tlu7aVKP6
FHxKE2JQeTQcQq5KT59axP6VVI4RPQw/yCsXd3XSwiztovO8v24fj1fENGQg5zEz
kluH2FURPVv5KzH4pW9cPwiaGJe8OdwahxOkwS5EAXNPUJpS7yY9It02l419W03/
k77pNfCo/+VsJ6Lg6Ms3IJ5swAru0dHGeUqX7G8gro1Y2agx9HLUaJB1XUj1xYyK
HL9X3Bk7wJoDoagzYUagqZEGMUwsy/oH7aIkb4zTcAIpRj4n3Xukxva7ZfIntz23
/np82IQqjH0G8sbrS8eqI7cufae+BTyOP9wkVuHl7++fbg4UEsemYjuFie1U/tKj
WCJki1k3eLKU7+VUPd33qsewEZqXOjgRuxgCOQjEGRXt+CTEMt9q8NjJ5vITCllR
MfayhMUQCZLgxl+KBlCEEtRxvWFBUFbpDY5xQkVWV1URS4krG0f5Iuhqt5lCFJ+D
yAVkXdZmZnx9nnWLpDxpMONqjLZea/lY8if2wxNiiLpUGZ183B1gA0Tetr5HZoE7
TeQ0sHhyK41D3TIyKrTSnSs3xdIwJjliW1PX2uIjpAE0ux34UL4tvoq0bLOptuuK
NHrv4jXCKvccvPgfrRHGCypMEOUSiieSLle+InRVsVLBSkJoNTs8AaDiI9/IzqfO
X+5dFxYnWPwVvb6AzdOEDZM3nqIoG361jB0Rf0UjtHEpivp2zj64KJp6ORWNsN/r
umagg3/Gjmvy2eYm7Yultdk/EdPuo0sVVe5q8v0fiZNs3G6e5NqbTA6ntXbKmVE0
zOE4V7zubScmZem0nSfuL2Bk2a5ytoVbCZqCdWS7Zh4o0gdRhO1+wyMAqVpojk9I
pLbkGaoI75cQCrTVphykKKM58hZ/Cy6ZU6o1m9+IdWWJ2Gc0lM3ll3q4UYO8R6HV
fLEP9CddHwUPZmpvesv40ub1R2bjQbPxXltJWr5nPupiDvRhfydBeJ97PxSPa9rx
eZRWz3zvB2tBGEy2VeG0K84jUv+sO5nTEWt+YD+6asy236k/jH2Tc/DGYpJT//vO
chcCyEKF5P9XBKvPvNC+iEfJujGF8YQXSW3KM2zSJuiK4/LG2kVrKo3RqrcErTwf
x7rt+h/nBj1ZjogXsfCtm8L/ZK0JeFVhjtKxoKTm+vORRL/Z+5l0NCKJ9z789kB2
NywaTJj9uLCaEl4ZCTG7/+vefiJzZsCndgIoOmBbIOro434EjFVmHYODEqMYLtEM
RS6p2coslIn6rGB7MaFv7ct/bAxwjeX9NAQqTSm0E3RKk+WyRLVa/F4ziUkl7G9b
QRrcuYksVBunHsQyXG9i99BW9zvxt2VRvW/tECCb4uXmqEjBRMw9Dg4IOk7CIkHf
ZPcViGbhDD9qPEuoBWtCb0k+un9hFJW7vtUBdXaoGV1XBHc9+CJtx6Zgqcb+BWfg
7gob8V/GlmR7WXxL4YWR5yS36sal7nfphSCDsnS6hgN14lPbpRyuxYaTRCMtsFhH
Mns+0X87/4r2ATDo8ftw+vFZZlXdDu89ZarU70MbT19wuuDORsABvwhO+RimWEPQ
gUsIX6NiaadFZoDOu/sJbeg6Gl2RKG8JB7N9Ymmal37dp56Fj3UFq7xM7YQ1o5sV
9bKnZG13x/VZJSXkltVTHg/jgizMaThEIxpilX+AVaa9j6+qG5Mpo4lUKrNuQpdy
2IBuwg3E5r9O5Hof9He/+h1ZZnO4/VEeWvJutgUVjTUwsq1ukE46+ShbDmxpg4zt
gELzJg/d8WUWTE99/4N6cOa8+71lVviXaVGYEL6YfqfeZqOc5K0eSE7w9tIm1kzp
jjEv8WS0WZSvjJPj1XFGZCX/RNZspRJQFw7n+K1vycOMG+0EW+luSaVhMtGF3Qpl
+cOyRebJKhIcu7EVQC+H/XkwadmoCkAMNzj8Grd5Z3Fm+vAeqmEhwXthptNX6GrC
9uT0zbxY0Kqvvp7iFM5Cy4ViG3957HZvkfvQQF+ktt+OUab/8XU4AQ7PA/ZbdwEG
C4QavvdaCsPcLAkjzojQk/qhysZQ6gZswyQ9NBKJOtyQ9H5ZxnHJeZvtJT/UXQKt
3C8jvrgYfCsy1KDcpvkdj2BMsap1tB5kaskKpsWkOuSJN5Z20zRQOyFOBIUbhV0h
WHrKf+5aWeEX9kQrSL2F9b7N6d3FRsp455sk3P943E+AXwfRKuwqvWh3csdG6R3I
OV+zbWCMaRYuzF1CBKZyA2BVTbkAW8w4y0TqXp8dk7FWrr5UefSGTIE84ji41wmx
zsFKDPte2BEmt6c5AFOCt0Qf6KCn8jTP3GbAmqo60OQQw9zqhB7E7eaY9a/41s46
hny0XNlSLmdhqZ3g+4Y/rIliDV5jLxcuzyD/dCB1MOaE/81dQeGbIuSrBXEtLPqw
bf/QKtb/6M2wM1Iin6tNbWOSpOLsw4C6He27OwojnIYBXfPuMYkOTBF1+wQkZs/t
Nh/QYFhOnkxBKHXZ4DXi//yH9yBcB8RiSpnXtHUwt/6rwpsWpX2WmApy7lbCVcJr
AJJ0Hh7BJYcm9trOCqZPy+S+fPxij5b/gsixFluOhrki/hVwitX9X63h8HYG2g4B
M5W/nxY1XZvr9l7z5v/ytuHANb+2TDJe0K6EfSeXilEJojcdwsLGO1WLpvWygETm
ZdNmCwgjWP+52syMqGMJ/L/2sM8tjmPDN3VFcu+c1Lt9liIobxdFmWTsmemirOl2
wOE1gNh2mGitkTqRYAhd2ViSrVZOHgc8XaP3bcCFKbV0z/rqS7mSV4l4S6xAvxj5
zDz0NAoLtL2C93TgUTnAvlXzT1EWKOH1EstJrOKPjFgS0mHEb2OEh71opUv2k1y9
CFmvXFuIdZyFZj+jvinNr9ESGt1DIeFFPwPg56UoDype8CiZMTbyCKK6Ax7nVM1W
K3QqA9ZuKWWc5hmk9ceZ4o3NkEtXp16kva9WjZfcTtCmiVRgg862KIkKDyI8tEaq
54kRIzD4GRn25s0SAvVDJkL+Du6Oa5hjPqDEzgRwkpkt36+H02JCOUCg+ZS2SAIj
VLsaaOhPsZqvue2+hZt4l/f34Yyx2dQDw9AoS43pwjPL4Xy1Uu4FHbtef8U3/XGF
DRVSRnFAqLTTJgS+ovEZfT0ZVcxdXWuBST2r8Dx8kRDbaactB58PRI4seUKHSnPJ
F6jT8xbxGPmaJb+Egh2tIsoab6ZSbvDuSb0ollvBdAagzbVrjnY4fxEefs39Ru0o
97eCPWEG9ZeTKcQyoltyYp1wU+CkDPyRE33Lb3KSCuzv9PA7utv7tWrLmQeaRnT6
PvUZuBh/M/LP737z/iatfBkB/Zqgj6BrRxgg4jHFyWirjx6vVY5WIF20zo/i1Zh8
HphXTZi1aYQeCPoq7z4T91oDUTviz+AfgCFfOOaXpVkIbZBZs/zyaHogVCJInu1P
MAH2NqJEdU3mBeZbW6VYoUX85NGyQM4sPK4kDG+Sl+fvlZdFXRDl6tCDlWt57lKj
HYnyr+B0mrL7dwwmxTeL8tvANEqHSS49L7Edw2p0gYfRuaQ7PK0WUNU81t9NZMI1
Cg7kUzLS0c/9zWhKQPohG4+KT8FEI/RYk3eKl7+RNI6iyb8/2C0oZK/CcwnczyHo
qjM1yM9e0FZIRwN9nhkhxerMi13KkssR1h2vbCfx8n3kk329NS032lKXIjc6b39V
MhHgE0uaCRh8HyvNVgf0HWAGCP7URKXAHt1US7+59LGJN+1ppbk47zlppewWCzCU
hd2+ZVSbS1KxXKaXyqCkBlxNbEPwa/UwCwC0XNvdTtsYFc5Kn86s8dmBLkhl2ZD4
ArYGeQEsx2ZUwf29yLamYyfz0m+NIsUb7wBdWqpBAs3sjy+FxGaAhWh/RWFwJqtN
VIINqTJJTOuU1u7b/iNopAIXXp/5d1XmfV0AYdOdnjy6wc7hOt2n0tAZSMxrkRrK
Gyl6ONOkTocw3wmKR9LjTdDEPMfsIm4GwDCuLU0W1c4q5IHVFuQMj8GVwDRa+3dF
GkvOHq6dooN/wM5juAsz+9tWDx31VyUNnehhIr3fxrdWEDiybKnpZSQkLcPXeT73
ViRiV2K34NYcFIPxQZ2qh6oYpC8eTeu9LaxpCCNQhZHon0DHzJ1xPJfpkMm3CFNj
K4UX5y37s+xWFlaHWZ3sLQ1F4jL8cA1NGM2bok4EPLJQJcdszMryg9csOpZv6PdE
jine7ZWx1qdNLfhLR+nrLShSVZVSGqQcURSZEXmZFhsaKpmRo2YlqzJr5oDBXtXC
srN5b4jOy8F4AblFbZ8DsDr6QZxn4/YJ0Ur6IGCOVsUHH+PTUJ6VZ1cvT73A7CtJ
OZJJ3ufwQiI4ePv91fXbULUA5UJPedqswO4lRoQbWoIBLtvsRUPgXpl0B9L9pQ6x
x3Y8+f/CDM6YGhB6xYC4/hz17oSURnglC5JgnwP4muLS8U2CJt3NJYs8DB2H3DQh
far7l8t4pvrAN3SWwxF7TlcCV3P2OPnx86Y7vtxIANAvIu9rHqgiI5NvJ8jLSDXN
icxIATEcx2Phj+SwctlvcKHAiqpBxjWlTQn3qhFDSgt5HqZpCyO4BT6wZ7yvtN1K
j9qBzmhfbMfoid4wMNhhUZh8ksxdbQ0Tz68/sLjkogOGPD1WKZWjoFoYuaqGLh8L
Y+NY5SFFGdwN7jQ/d56fSDCrB7bSa7f3hE6ZqfQhySqidLEVwgm2WdM35Ya74LVQ
FsrV7CJXPxozZwHzTire/d9UmiIcvkWMGYwK/38eThvEgh8wYb/7pCcL5mvGWH7F
u/l6cxUTCCVrYuaOwa1kaRZKtyhizPhby0u+ys6JhjiXbNtwGe73QGHcWIY18L7e
aR2fEoAudoZsFrDxXFrcMmrwD+CRu01wmiwWm8hYn3k2xJBkvtGCmp985yGlG0Iu
7na6ShiQIvWDpATcG58kga7z3HNMu40FxU5HEF6sDDv8m0zBj4DCkBs7DdXN5Iho
hQGfqSpAUjaQvyCbQiQVIvgbDz6oVImiQZysG+XmCQ24WoU50Elk3GlrbTq3JhRL
GUxvJm7Qi033Eq8EZm8QSeliNEGiV7yXCo1WAve/KZD8aUb00OvBn4MMyEokWOmB
QcH3tLHgr8IRLpdwrFaStVpxq1AVPFFUwEOXE0aJu/7Ct5qFrfIAuESnYKPpPmhs
xI9p+tRJ6XLVLyJDQOnixrxiKfjpX1JISQDgcAFhpqi7HR/wRNPzhaByc5CZ1GHx
NdZysDSOa0wcTL34UkBPGMaKC9T2ky/m1I1BAsT41JNajrHgH0GW9LTKBFASot/T
uv+bb5RABHncHzXJd0FzKOIzw6yEdOzimzCw9NBQUbRsgD20CqmmxpUOfRQreGbL
xKAONHLo62odMuls/FNv6htPa8iJmMoIX+ODCidYiyfJNeceh/YibT8zqUknx1dk
WkT+GgQ3fm4+EY89voEI7SzDmo9tDY4/ddPnnJe2V1ryYjlVjAir6YIZn8CiqKbh
kfVmksb4aeKc1wwooOX8uirAKxzKofZj8kJe2vQiHFbtSQIBqE8MfayctHJG1e//
gTDwbnqRJbkXBYEQp+09eoojGskSbyeYm9niOT+8YGZGKePazpuJEiU2bbfxvA8u
oZsL9mcfYiaar44no18X713esOundg28QNvKJfvWHC5rXXrI4gEu0eWLoa8GUBI/
qvv8dJ+EKhjswlLgT9++DBRz16bYbygPc7X68vMBxQQgY+00vK2GSUy2VggIwGYq
20Jjhxcb6v744KC8X66k7St5qwcp09F5FQvk0QOwBB+OrYJfIj4QgsSf+XDCbM3+
OxntfFP3Ic2FZWdl8jWMzKgYxGmfMZVDtGGOQmuuVtMLOxl9TUMh86EcCG26bqsp
IM8q3CtjDMUQ0MOQPi4y8pfS1wkVCga7H5cL/jvAghLvVEp2jstG+ansMplOK4KK
0KsXcBZchuRNh33PY7bAFWQmFVYKDoX+IvcZ67O8d/XklF4jpm0MsBflza6wy9GB
ZuWl4fNOaJUrzEl+nlYz39iiagmCrN82XARf6oqYGG2213ihnU065jQl/o+TQeZ+
3yoe+W5AyGtoPUxTS21z49Pj607H25KOZbPrzzXoD5FP2pNQPXAWwXF/cr5cE3ob
a7Fmdl6q2qUkK0oViFxCUZE192RtousqZGdI/nndLBrV6bjNdsE5XQ6kqbyh5b+v
yjDIgYWHim0ylUTUKy1pgNlpCNZ/JlAKYnci49i7rV2O5rovsID5nXqjAWfdCmoo
g7R7TsIXNcGQbxf73ir0HfD6MXFZ9BFXq/rrl/Qn6eZjMgYUiZYfy+ED6bNeyYfP
n7P6zlAbQYyZt/aGgOvFXqsmL47eFAckHzFy0kytN/PjzHpb60ZPeuf+GJ22Ajck
OS77ATl0F3s7xjNttXdXXALMufTGOR2Rn7VFJL7qUWJITw3xYLb8WOS39IIm1KI7
xosUV6oU3GPoFGoKFf2zUbF51TkngKhr1D8pkv7QtrZQ3O2aZGNsecZlq7csiqmU
BEHjN4GyunkaJ8GEr3cxfaiy7MtZo/DSSCmUHjOkIxFQ9FX7Gc/o0Na1dJNz2pRP
kuwcEp8TC9PMzBYZqB/bNMYePk6M/ti64CFWfW0tAlfkEPNhreb8H6+Udw3oNC3x
ab1FjY+q+oV4RDP+U/0IzdreNh3XCmQTDl+MPinqIyhkcfrJB7Vzr1bAC96sslfF
HWWz83t0bXwevXx3cNLDNclc4moNPOLF+tZtzjo1Xo19u8K/1m11hxob+wDq0XPq
lWtV0lSAyeSZUMbafpSR9y4C2Y079aHI+7495LNXKV7AvHA106QzoNc6hrjOjIw5
b9KjsNHhTogp0rNd3vRpOPHQPdf/EZ+D/7o3FwVQ5uZL2xGhVF7m0lgeVkPezlZ5
KIQYuvCjS0nMKu1+v5kBpQtGIna1EI159ugylKEKcW9TjP+sQm7naNlaxqvuvr9g
Q+g3hiAGYZZEDa/NFopEooMCRoCc37TVSVVsjmF3Yz2C/7OU6w83HlEW/82Dsz47
DSboXhiPtqzTwCdsAnjFNdLvnaLdxpTkTh62ApFlt94Gs/JOlj0W7+yHMIrCR7qS
F5lMiWLKLuPYSyAMc224Bp2t4sQ4pKMfVUFvoAw/2C/nj3th7nXFcWDF2LaCuW+z
V8GWjcRvXTQUtAklvfOA8rTdhkNj4r4hYwYCSxfQ6FLlyWQqJL1aEuZ9eLO7F7Tl
LI2UjoTMu5iB7xOpP0M1lhgNcniQpeZZQNXqwBeeQQlwB22wuYeGWBje9Z1dc7H4
PJ7MEoCu555SYm6+/3P4gFkGkR6CuFIM8xVPJ+fGW/3HgA0qPCDy+MgOfDOZRhg9
AP5V7b28MXelB+mQkF0nbe5VRaIKOrbcOol5NZ6saPtzvU9YgksrWRQFaT/2Tv0G
TAQN/JsMMHrPYqbEYoID8v8s22EU7FgPRr8KPkglElWGMebvdZB+zvlV5VF9aVkG
TGQXqbxBGNUJnqG9XmoXl5Cby20JHxjfoyM9C6pPC9POhcWy0YtHm6wwezwl30/m
5zIgwXMN7cUzBeOTK2cN2wgqlHLMIsCP4Vgl1xy2ZmQRJayjV7/VgQZ74NhVFPN8
7h76+js7ci6jomxuncQDoqoACrB/shs6+JTLYmE9Nq2Fwlj9T6DLtUhls3GibEXP
wxQNT/Y3hF40x6qdTWb7T25v4+KLTWS7/7QqumNsWqeTg8qrw5YA5xO9v4Jx1rZN
8kNp8a6yVqgWU1rqUwiTLKjQ2lMpaWbsSyShBa6/4ccNJjl0oKtSveWLmNZcaoDA
+HZEY/q8U91v2GiMj0Uh9GAuRsOJN0BFYmb3Jd0IzQbSKXojQDdTdFW4oawMjDKp
lNWDjVPUpEPDQqDo4JUDfBEV7Me96nmY9BTl0sNF1fU0h+O5WuluXTJU6VvIo89z
dEHybLN6b8qZ7fCEYSrDWOs2+Pc4CdQNSOX6KF3NjqQ5hgCgUIoA45zt4/3X6If9
6jAOz8rD8nxvt3Z8bsrLPCW0+xdFls4Fm/9WSZUfkm0vFX2ITJ84KGGIWYcMSwtl
WoBd5T5ZDFraDX+QDpBs48GovBHLhfdkNigFt2Ik6C3j06YSguqYx8uv3Xnf0Xhz
1PunYsSiHTbkANF3/uAQXyTM75bon5Trm25PNzq3hTmc2RLkRd4CKRCKQzqK3eu+
19tsd5BmhOfBtz7hs2dphDiqT5uS1Io0fj+JCNbzXT2frrvoHM5fuaIdH+4Y273F
wWfIhGvn0tu4GNoub9jZiPUF+SA6NdUIoWYtfDtnlAWnN/g2SdR59x0gP5kvD333
VOvSWb+T0vOVKbMmkVqD+7kvnvP/FGwlD2jKrsp7yqmtsB1qyk/jfJH29JvzhYUx
dyb4fY4s6PtyqVkm+vpeNBsE2mEYQQPqRcrKRfV4tGLCnRZiHuKuNQ0wEBSUKGr1
mc/cJ4A0e082KCwduHP/UMnYupmgoY0NOj7K7Xs3FB1xdgNpU72pZcczZfEoSz40
fnulPKA/oWNbSlz//0miEjwChdSSRHSo5cM/7ojItKjxagsXJ0W+d2hRZ2X3LuQv
ETIsJNNkVtJIlywrAfnXfeWrOOG5TBaUtZAIngidfzZZ7LmwUyY1+mcPiN8AnO2K
UI4lAhhqVAxBFvIDRXZfm3q40kw9fccyUuOsCFKV+FaVFUIpRQQ6LBIorSDbo0pJ
kmr+VDd7YSLuY780EhAa7aXNacHxiET/EKcomz9IMiPOjTn3pIElx6Uvkbi0m7pt
KNrAK0XDhXQccm4lz5vJJKCwk2g7jTGrRCiN1JK/PH/QvLhvMdmOzFL5z8x70Zi8
NpS9Qc+KHPQBegxHfa5hnqTLDX2sFK0yUKTcL7utrUF4o7iJtl/STS8pBAx/O3Mh
gJWzjL/rhPZ69Yr4d6mEIPBqM71Cpw8jH/5bRwun8Q2LJzuCPbEvaiKejDT83n+O
crHYRJtURMLVCE3a6V4yjhH8CNJ4wUledo2a1lUUpvlAzcd1pFqV6BjlVGjQ5Swj
9/8/8ymG3r/wnaVgQ+mXsVqSILSsVYuyacSzr3UM+h7iRT9TXMoCIvDlerUCaszp
QUrCI2Q7APvBhdF29gHMh3SH1ar1IAaatYZh78c9a+8CKjwtHij8Vv+XvXAsKhqm
YK809tovqOPTRbsJq8uI8YI15Fxieo0/AZ/mswHHC+XPn/Gln6eIbAD11RgteF1V
VYcX8Q426c3rvBGXUqYswfckthcImmPJFXvWCkQgffDKT5a06PTMOTikoMwUSyMQ
aT5utBYhD0TsIGmCmbOVlmr8embtV1YrFek46AIyyCeTMwa2T6cctISNge/lCh7f
xQXPRIxpXtFNdttG3HDjbJ30wAKtq6+u3OPZziZa0/Btd4ZmdBA85iJUkJxduecS
eXwv54/DIOZLKlIPqIc2iyfIZP7qZZVksYpGv0ehhNHOpyYWF2RuP9+nSgRFXOcL
yAzDwF/sIm/EcEWrb7T3UOi4xFMli1Gx6sm50gYEREFStd6NOAidKkqWHuyu0CM1
ItkrLNSzHiqw6HE85I1haZoBCsMIawg2wtaDmBeAPgE2m2MGqyxhRm0CuHVynIa9
enZweQBsnW0rMbEU/lI1lmUQZKnXPuoEfY3t+ycHPHxKbZ5c1XYvMCa5RIFyzaAj
J5XP0A11SAXPqnyKoGmMqqLQ9ZunKkCLQNXm02XGEQN3wdLN6P/BPjJNTxIxWj47
kCEC0Sa8azKjQbg6RieabG2EnKy9FIx5NAhyyjkz9LTv3ekPAvLpP/ym9VJfy2vo
KE7ew2pvKT4kwmB2hCFqLL9zI9e0ntOhukwfF/qAWFRfQEwIu3WrBVf556nr6Ghl
21wM/ScJNKm6g5tm1iHGLEpm12EI98Mptel8+U+ci4UVsPU4L8D1yHKjFQvfrYdc
Yy4CgUwdouBBePDApCOcp74OOnBOyEXtfxQy2ZxfXyFDMGpu29jglZnwspCDORmF
9dj7KZNgP1sY05O8Uk0jcBE9GExPJLx8BXLp1oONINeRUU7x40yilBnrc5o6hi12
cOn8IClqu50LthteNxITZ9NniJzqa+4lkn5Z5uZ0CONn/n3AoGxkkaQW3nWZosLs
LMpSr5QIux4seZ6b+lOS33onvENc2MHaaE9Z0Ll0W+8Q7XDebnDkKn2Lp30J3c29
BgVnzMCVoUy5vxKS2maTV7XdgYUhy43VoM4O/qlhpL5sNYQ4TwIAJjthQ1VAKKN1
jYpoSpkMW0xrmtYjU4x9NIaeMAOTQN+0wNh1IL2mg3kvX2OxSU5OfCzZ41HIJDDF
sSJZ9s62uZewWIXcLtooCOfFkKkJm4CnlU7cWVZEBak6YgRjKNs7ANm2HqXUjbkr
9YO8q/t6+Gdz33wzt50kZEI3qLv4zMSV2+tEgpT9jUdYcTze7CiA2mwDW+3p7qTc
Ehg+iVjWdxX59lmNQ1DZhgU6fGGuGfyhEBqW/2/5Pf3dKah25eyxfn/ML8sxzuhk
9Bu4hKrB4YRbi7jiGZtVnVQXiZt0z+zvLuzYnq+97VHWSCvuySB7tc62ZnrNlnpO
OHcTTDW1LI4lQhzH7X8pYZopuEAe8QsCBhvgeSAaM+aQ0CHgP9kd1MVZSjSyhC2n
CP/fmJggPLpX5j7SvI0CGDWTm6az9fGIXXAbZQ3vOpTDVYTUe5g2ASRxU+i/EFNO
fh2TSkpM65v2F7z9Bem/KA8RIvRQNdeXGq8TVDZt/RpXNdeLNoec4Xvdx1ROiZpB
yx8C2Ga9ketjvJKpyKRi1A9Nh6V3MRk1iB/AGnhRdG8zYknJM4qdtJygEZfV/yKB
T+0SexeZUB8TZ8KwaUbldZouZSWYobBkdaWtiRgAQLlK6RY9PJX7uJkNQIXvEFJp
P92xno6Z4AcjaklghKUz+39LtZOhTnv5B+SGAker8O2FIh4peIUxyly8kLcrufGv
iDXRl8k33xk3/YtdX/ql8FeCsaeQ03zhjp5wA2U0eqVnd+hBK/CwU9c2uwTK8ULM
ERQEXBhIXjvRrF+AwfnBXfFqfIVCmtvjmHvckZKujG9Gmn9wY8SxxrpOK0iTGSsv
6p7OFnuL6FfR63swUMm4hYTXoE1JrUnCYcA48+sMpFljORtVgBxH6t7BOwSYyabQ
ESDpZdXMJ6BRYdck8d2H7cCG1NWVbBuNgaHf5aQu+duM8MSORGiTpPa+zXhLc3OP
2KGNqWh6UxrXeOSgcHlK/bTGd9FEl2SqIgYl2o7zpf3U57z9Hpdf0EhMobCCx89p
5xQcLFSBxY9WgmJmOFhux/dC8HOTkbcMpuiTGX2r+F661i/JSwAJmMUYrXQ0J6Mb
bxPoHm3yJdf2MoUVTK2RT5oBTuwLKgFqbrJMrIOcjvp0hHDwQSyiyTuIesK3T/AL
KjGC3En1hXBxaIgybjbAVFPxIW6tW6MANVz/TFkWIFdBy5Ecapy2qwLxxzbbZ+Oh
3uzvJxsWDv85b7TgSD75k3GzePCdLsX6LoMTKffi0Dhg8XRmq5IOxsZrI5oLUyCn
rVeGK5Ow1Hy8ZLV2RxLnhLY5+4Y+TK6yNS6R8cjYScuu8CdO0RSbtQ9MiCKl/9Ax
iPWxwtHZDg9nrb5k/DqJ8UOIvd21rBrY520SsQYLUgY0qHFkSfIBJipBdg6Ij3Pt
WTynnwGNFmLEXIEvWTEraqhNSY/a23JMYZ/JBEsNSNj0lkb4gdSHSvsvXQT6w+3g
fH5g6Tw7nujMNOVFNhh9NONm47aPgb1wFKqr7DMvvQ9nYNWsCe+tpuiM51H4ej08
Sr5OUHPq3PFcJj6RU6tgPMnNKal7hQr+qeEYBeB5AkmmjmKZE0n/MH/0n0+qjf8H
xf/mv9qL+ZMBC+N6MgqlhjN7qN01Q3u4Im+vM72oh7QjLktshmI+RDtRv0Mjm9Bx
JZaS3jlautqVHldCNa2WM2fGTQPxrgRYpUMf6fNSGfIUNILtktScGQwnvCjcNruM
btnM2MqI7EuVBvVMubY0Gg2eRcvUJoK7xDqZokx+DDHodIYnsHRhWXf0VnJR4vvd
iCBZ2j5VKFqQXfXD215XNsw/YWcs8k8TbgcQOkLJwIRdlguVQzAyiAg8lq0ua0Fu
y6Jnf8Xy9jIEpXXB90OuX24E6gIG6jd3bQYc280l7ODsYFdRW6EUEOzGuR2ldnue
QAi0w2g9+2DH2IdGboBpZDl5Eyn0HuXzrIwywv0B/IptCWtowAkMFuPMZx2roWAh
JNhGvWnEEt2GwIchtzRgVbRLS2tJyjZIstmujX9vqt+fCf9loWcpl65F5Cyi2EeQ
LAvmmqmGCVQSFDG4CXsQPDbFfJdrK3te8GaYKH/vY/8QNOOX/SXcLYHtUpXkw2sp
uxhKXai1imne4WcPWZR8cZAx+x4Aroy09bOZHwBt+KQ6c/AyOQgxOaU8oy1klLVL
rjqfQfKB6uQRnofu5SbdzPcXiwALg4UW1LODtjsUIx4Y+rKU9g82WBssOXtsjnDp
uSSxg974g5i1tmAmbwAU86lWWZEz1yOQgms9wBfNTaQy1qGpFuLYtR4Znm2p2oYA
Rk/AwXu2xh/5p7SHxVC2lTgFPixoegjD8vUO0PCkE/GS8dPZlhy6oddEkEV9JJUc
I9vOT7nCUSx3NCHZ3578Q5yP3UuMAZDCaRCBPELTvuLCgeMfefVYg2pZedTPnVbs
3HhHzT34JqTV+0I0DoNAOkbEplSt8CkfewkkaIuuElY8MoQAyEbY3HCwWabTsKCK
xdFH2FYZqVvE8pBdEtPBSJXUNo/yHWsL1OL7n2YuJl+o2e/eYJHgzD8ti9cNTd1W
vY3U0lkqi1g+l86Fa5FvoUm3IZuweJxP9QrRGVLYNsjMDD38P/grhF0YsKARgf3n
5kEkbYZqc3tN9e7ji/yTcRWoYrwUrLEOK2hvPOThnFTDDJbw/unhE59f2SBaDjKb
5dNSYu1825xSPwNk4wtT7BbtjfuQuKeF/62+0PL6EaXVOEIEWGsOuPqivOt/zZ+9
SD8JiosQ8YQHvNxZ4ghhpaMejK33zpdqbJ7NynMSvyd12RhHPdvYnuvMevZUBotf
G9cxTECJeLdp++F1m0AjgxMh2c68YiXTkX0QrFvSpYNA5eGcgq2Jrnt5g8ru4ObY
i2m+N5pF+FeAd3ej5Hc7ARqVfFDf8T4oeVX3k+9wdr/ygugYsIigwRYDOvV7lJyW
duRVaxxHI+gZhZsOAVBIHH5EFFaROpjXdgN7ktWgDQlylbcve5ju0axSrrrUF1BQ
Uikl6OobBF1WbRNwKMcT8/Kb7QYROahX4SNH2IAGfNIVIE0P46aAztx4OO7QqYGy
tdYmt4rwEKVDbbdewgfU/99SZp3LkDxQ9OFfZ1xQlYpvjh/DsCJJPeVaY61Nsutg
WViJq2I3jCXqg/RQVOu9RZUR/eyPQT6y66CDQP2TWZj4+quYWnOfUFjsqU4QTbq1
52xil+0xH9HOC3IiDWjI8KiaIOa51mdOH02V85Kq6oQXsSQKQUeIx9cJi3znb/Wi
xyLi+tILoEaZHLOXipEIYUz8ZiGWovn8DoklZBFZijenrsBqHwUVXpJxX2O+wVgE
oaNsBU0tWCEFvOWPBi/2vogm6nn8mn61uUmcrmLb0uUHSstwp8Xpchd+nG+wJB1t
/fmvmZ36FQJNjmaPV0AViSvt0L9YUl9iqZp8YayIzkRmTRz9b+j2x6GBtppNMvCw
SEMX9MrV0xY00S/q944peytV7NSFJaD7LEcgIysO/KbakZMlzbec1YYWnRBMIHGl
ojKrO27jZvXgsNlk00IJdRQ2FcJma6x3D2/WsCCHo6s2FYPNUunGE2DlRfP3DzwH
VN9mAHeSNXjmMlNvF4d6v8DhB8GTgnnl2EkQfoP5HL8zvA9lxATMbFdYDg6oGo4P
2ZI4sqigx5XMQbm9S3U4aF+3oFwo2C32qVFE9e+WyWYL8b1kL2hijA/gyBEwxjfh
+B/WHz8mG2z5uD4Zl1xzF6kRoEfviABvE7GycSkALvjbgt2pweYhRbDGmHBpE1tG
1gAy63jhS+jsYGKUtUJMnRCz+A/uhe5xEfjDR+2onK13A4pbFPebYvQnwv3ZwRmN
nRaSmP5O9cIFsx5CdmE4VsIjUZuTtDT+48dOcKw1ShPBb/Iav458GZ8uCnOdWts5
wMOa2XlM/6Hu8qlvueqqCP+12hU2TZA9iArSfYo8FB+YD4ifTKfmAj7iTk3zUZPT
nYk6UzoBXX5hBGMikDuVOiKPLMHXMrADLh9PpEdliDeZsqP+eq6aZ6eSSRdFV/CU
8vCbxPov6riXyS9fhzD/o58LC+sB0pUUusidPaWPCCd7JIqQTr+5Tou5uOWtYUpF
WrhWDQZPFv3M4VetHH3HJ0MJLiquF+EZy/zIMysKA2YfHjHPDM8zl5c9D4gV72Jc
/KuKkQDsFEy5wjpDfkhy2Y+kekcPKX+TIplOcZxEoGxlmnyNP9UUTcHeMyATgkFj
pZR2v8/7b0DQw8oZXAiTYj5d/+9JRepmgXV3lpn4rct8vgAOuuHh/TAClaFtX74Q
pCbTA2rKyqYMNKWLfwc8h/TSgMgf/lHcerb8zCNjwUCGxeBfqIw4HJ0vJTJvoS7Y
0qTs0gwsU9HgFOOO0tFIboKuR9nAmQ1GN01rVoHqoJIdmS2vJI5lz21Nf3FZV+2m
/hxWbe+0T0umPonfaW5SfQPc/lZbdLHlGLr+RdlmKYqd6BhJRIJ7BiGNkziVXNCY
UpvjnQtNOXMfHuXdyzan42zwyoq9MvDPqQesc9h0S4AGItOQWR2ELSKPvsYjdPWT
aoP+W9W+T47orsVJJdZRL1U5eCBpegeDI6ragSH19qBgHQKkvW5Q9Ap2Sxd8210E
cENzoAw0YM1m/M2APNwLahtq+MxWBOgfatid767BS678hXzKLNMHL2CASWsScQrt
fG97loo2ZSD0mpEAwNOX8Y9B4UVL+o73VVOhIdiPF+Tx4TZ6b3sbAZs3YJca3sjK
W4i8gqEMQ3vwmSrUY+BRKpYHPCS6jf5ADb9pCX1JfEnsJXrQVJ6IyxsHrmq+YvPY
HUgcpWFqDB82NIP0CBjAt+R9yuq/PLO9oY8h9L3HxWrcx5bHxj5LrZsCd7h0YKjo
TKeivVtfs7n5z/E8UHQGuPhbZiTa2iiJa5TPxIYdkAJIWyrT2gttd97Mu1Lw3+/Y
LQQXSU0d1mmgQlIWEZFGt8jPQaJH7WWIS9NDo3LCdtuGMl9v/cc9PUAVqqDTyHe+
Qb86annupVqkNKCrMhFdubZfkmj3gQ+wwf4ZrY61EjpqEeHaedyYjuUIp7iE1a2e
9a/gE1H7Dy89GUVvo16kP7FBDjmA5vScFziuhAaJrWeeAvkgC6EOuLtaGHBEYX2q
xGoPJX8c7yySE/dHDdDtQMFhS8EOcsnOJ7rGV4wpbDmEyjUQmKJuvi/C35yLtHqz
j+KsUneeENtewVpLkwpErH2saTZw4dRvUn3RsGrpjTCMaqvVYWX71ZhCSxI1FhYv
jNSsUTtjFCvnygwdU3oRiUZPwaagVPBCQYYXqqR5TRNUS95QuZVXP3+vkhuoa1v0
jGssVr414LW7XSPzH1Mof7NO/mCy52K4a7i1siuIytv+dyb6tMPFZxxiex5NuIh7
xZnlRRmLQxukJQrVcvXY9NjDhHng9R5fwmiTx0qnIDkm0nncJcyWrnDTuQ3KP5z/
nJeUOPfXcoWyjNE5tRo97hFVzbpsybvW6jL9Qr4FDFEfWCbfALdGBW9Ig0usdwpU
PkF2OFKsXGOTU3wiNRIU96BGTlxS/lKn91XiuHX2bGqRmYLAKyJTahKEycuR2Ro4
BjhIC13/0KYRE99ACLtvD6A2iLi9yM8lX+QpIsH5QeKaj1JeyGZ2gTaZBySpE+g+
usWb2jiq+i/7mcPDkbjg+1/BGuvFq/TDqoZ4lJxyjsWsvvuXj07BcMeyb4DVI+gZ
uLSvB0PaeMJyRx7q9p38xsB1uiUSBTtr+4vbbXiusqQyw+P6eX2SJai+nMDT10Yj
gDaRSYz6NM2DzHUUlP66mKhEVwlCx0d5zInIJFq6Egaz/D1z8/7TxZubey34x3sn
J9aJn70CsRU+GLlJOgggrcNsHOZOHzEmgxq//PO3PZlmtz0/CRixVsvVDR4AIg3x
IwYMIHtBLsBNITLiq7c9f82ri6sDBkWWhIb1ofOfVXES5m5rGe563UAU0hiOac+6
SDC4R6lKx2WolwkQyKyPuW5TNHkQ7A/aRHDR50ylp5HYfax7cAjiG4YSl6Gv0Nq4
5dyPAjFdGicjpyLHxqBd0Wz0zcXoh6S7wsS7HFvc89CVZXHl3CVpNVytBV57+iFa
jpn3UzhDzNF+Fpq7dmOTzSWEfCd3V+8dNEZTmvGEmPXw+DYHB0Glpf0SPZ937192
bJtaUBVGjzq5nhf3t4fTFKXPYB4d1H6/0APXf8UpZsIBxFDtZwiBfMj92jw873QM
SSV4BvNR4Z0cHCwvo/EV4SH5ZDLDitsPyn9auLREIXhHmNvpjeIuzzzpJmhSAOqk
+kzoI4TTYAjsigVBtCWJVM9TAKrq3xUxnWbulxx5Uk8b7oYNoLiPnvAJrz2dFDOo
e2UOlzif2rh+HrOlZFyAOyMJ808NifQg1z9m6ggoXgPDzxZcZ7owCBuChiGxvS1z
MBZuv8cPsUwskKp2U1PuS/71/wAqjPSItDlGPcybS7lAf1eaosfkxhgTPc4zMJ+f
EoiL8mxOHL6JBVtqy1iCrq2vn07835A1Jmd+rpbI+G0mFfUXrVjtIdtQTOHa+VEl
/nA6F/VCRnqnwmWc3DCpjCAMZJnP5nCDzGLPBvilhOVE0T8jGAMfhyD2OXIXz3bp
y4amiTEC5si5EN6vL9Xr91M1s4fi67QS7jsyQYO+ylNzGM2vfS9U+/vsDxvUR3tU
/Px93owblyeiPnjOfmBpDku8TMBdCIh7KxYlf7e2dU2w/J0Me0a3VBl1JoymRkJR
2Vj5wK36ZQU24MvqjkL441u+sefBGUaZm9674QZruUyyNuJkdf1wItXwpXIuaDLA
Ors7LInEXhMLSQDlPlGXnIdHSJtFEInvAzAw9+99XEZLOew2tmG2l2xyMax5LMSl
/7/8fa/ZbJHIe/GTs7+UKWed3ccq0a5gpzjBjKx/4KuVxYvbvG2UNstF/cA0NSv4
X1RPWAXsVopXnOctkOm9aiTVNpgWfVN1k1ppL03zvqWCIHo/r2oBqddxaEv5YU0k
3Gxu83TJFvEKnjM2T33PfX3SJjyEv0BNbITotF3T7EX1eLJDrSDtDw3+HTOSKNSB
yQRP2fN6E76ZzlLWiIq31DVONh5lNDiAn+5z/Arb5S7Cs78iNYfQj1ypGhoBy4gq
g7gu7MwQjPWKcAqZMS9Py+1XaM0Zuea8iTsidSPfHqtOclnsSzky0QJx6YHSJiuy
ZZwXKAVc6WNa5X7vlUGmXHbSxsbtZa13aVauuqc+Y4vrlNy8xU3itt+dkwfrqH/u
B32mtLe7COCIkZABzjgDvker6uBWs9w+UkCXedz6ZfsnrckKzwHqrKFdUAJemy0q
LKuHpuuKjKrkdf+WuwyIkQkUfxq6ftJTX/puAo8gYqWd8LnINjSQKJjY+XHS4/9Y
Pa/dlGB38npnFQNwnEIZjeVy+o2FVBjsdszkouyASkiNvKmcUqIi/TIFczm2fCv8
Rx5B6FYTDMVTNvGl0S1lbFnJe0zXT4ZGUILnukSM4wXOuWqm6C1UevGbrNK8fb83
iuN4sEg4eHcxIA/BLn5QHYOXJQbHAn1LxJtjqbgnxpR08KhJ+62FIblWl+R5BTNK
Fl7UbvTNjpZnX4vRC2U0c4J25tE5or5t+7n80rMlHHlteU6TbBgNrkKjzech6om0
P0BPKXsZHF1MiONL59ppfiVF4C4YSkZOPcgkinl1ZkH1SiReu0utgTdJjSZQnXH9
u/VgnjiU6BZQIl/LY8D4jvI/XEG7we2Ve+lfgn25ff5zrg7p2tP4IcHqw8sXM7X+
X56PPJiRW6OCUTgbbOb13rNzOmirrkKqHYK2vFvPL24eRq6L99lZroG6smfu1iIi
NU6Qw8LxpIQs3wTWBURM0pWYKUnazo95/EyaScvHuyQ5CJp4ztaO699eQhbPbzN1
5ZTSlWcK+oo84xVWkbu3ILrZO/3LyY6yD4pIgu2HgmOr8D5S2TIJNTn5HgY1qnUl
AE+SCU9xOA5ly568iSE+W2AQEqkMUk7nsltN2OJEMIgpeoNwUsTG1J17EtDXWFSW
P9CecDLHZ4HPO3sGoDIuX+2rNieRyQjmgUMj1KHc8Kp3LZHtkXtxcxWE7wSvzztU
1TBt3jmgTzRWE5LdhmWEy7RWCGNkhUuJhivB8YISvbfm2/Rpjpzjxfzn/fDS+Ap6
NncISPmWb2Vl/c6p/96KaY9U7Fe8rr0dVNmAwhnQ7CLK88hOTopWmMoeb0aaPcfA
zemAgmQ+ComSSSRPUpcbQP6/94xQimxhNC25KTU9g7eWmEvHktU9kTQhRs0QM2SP
/HBYEwcQ1xFcFsduswZfWFJUCsMJkGueARGo7LZkgYVE1/+vnetXCMbLQgQCeS32
9CagO8YcjeJK3LWqpiVeo4B0p5R82HQ1Ke3L2XzJ/0z0C2rDSvjiBD3+ue5QZF3Y
oYAEsoQetwHbTeUkBBqTkUE0xmORhtHvswwPCEMJmrlLrE2ItLkQfa72HkoZZxzP
VNEdQbrGOlhonwfcn/Q8P1hMeby7QBOvz0pLdemquEgyzSPgUhq1d2zRYlrcc///
VXu9gYOkI+e3EAAmTQRiUbfjENqANCPZ+nMe/3Wl8PTRA2JpYBjsMiqSLfi+QGHt
IGlMnuCKIXOfkoCPzD8lT25fuM+pVTQDzwT9Klswydjrj10NGzPX9CGJijKzw2bN
O+k/ENNVh7Xebi3/vAtk4XWILrzKSe2MXPuJ2XMg7Di9Biq6xtWeGBjFw68zq7Dk
v2ZJlGNHd4GWricV4Uxhd9NymyQU2Az5Sv+dYCDThw2E9edbDWtOu18wEX//tncb
0nd9mlegB2abgVkraA0BfkpjmEG/p+OnNgsNw5NgXDPYbeoH1f7pgYow5wmZev54
jN9nZv8d+d9C6H72/K7msE5w8xnSf3gbU+y7lc6xKfdyBAoCtsvbqhTWcmBFsafK
cunO5w9tYQK9s6VgwWNK76upRRiGJgf8KBpnlGUhR0lhQJhAzPlPQQRowRyV7xys
BgDef/x3jhASaQ7uc9QjXAGgpdmKoVZ4455izZ5OvXZf3209pDu21dQz/uaf4X25
n3IdBuv//QeYhufroDwTWL5aNsD4OR/c+ivH8iWOILSZshnu0rOLVitig1PJtR6K
sSefSKD5ZG7UbzovWErbeU/kIbmZp3X4NZVWYoiJ03xjngT7e1q+GPAnhtqnEE+e
ACyCHBmT0O79IDDmuhRku7rDV7o4v0GXeuP2nGYbmWRzxbKDCSq8n243LjUPrLvn
D//rqVmSl+0AiXmgWkeGKqPc5RzY1wbA2djnYVGlmEw9maQHSIKl3XYZYhqU/219
abSyhNPVchgueLEZ1LE3Wzf8u6qDDMHNh7qcbrEDw03ldq7T7ZsCjY/TKPdrMuD3
CtzmVEcpEV5Xrgm1WNSkbLbNrbWXP9A0F2ESGTM3oNVG81JeO5OQA9FmPnwpzBLV
j6HpM+Tjb6M7+BpEofE74hrCZo9jvaGgMuWarrKtzLB81q+jHg7snF4UsTppYIac
e0SfexrQK4GgiSHxq9fmWkHT3x/Z3WP/O5R3FtaeoyXkUBesokNmNQVvZKtrjzY7
zKWwJjohZGl4aoAhKPvt1P6MViRb5oY6i7+5DnTMeJ9Zi8ZX2xl0czsR0Fk1mn3y
Q7Fm/82D/nG1uz3xoRWhowSkcq82uM6WJkeEIeclBG7Fbke80SEJKiK6eOgOs5cN
wcGyADQd+qMF61MRoYdGsGMgpnpO2QJc4+OtyK5j4C3aH5zySvWGaIKH6OXtdHFv
jCSwEyzRV1/FqR2ABSrhtH8jDfeBOrl/LgaiXC8z2RMWFQNJHMjOwwAc9QYf2Wzf
wIBmouPnWPF9Z0VCi7jvoPyF9nA+Xh6qdWyunaNnenS4ssVQQW8rkmHGlauZ00pV
LCauH4ei1DkhwF22YwHFEE9iNb23xOjZlI7CvIH1tCz+OqXWbwiOjoFiIFU31t+8
lbsBMryHO7G1G8QopAj91fmPXUlrgIFqEneJgwLOxi8ehiw+KyTCXiaxDOziPzlP
H+BTeKP/C27ydcwgFV2n6nfSbJso0L13bt49KGHYLWnr2Nat02YQjnuqYEJM2R94
QlrBC7BMhTufZ+o/OY1RShUXFenAGlNgmC4CPb0e6+DtWAzwDJRZhWwX64Z2PzvS
em4CiQIRul9b6rejouQBUCbTfsRt+A9dqwrPuWwSpVNluFMiPdwHdLIeipfAPvMk
WwQwXf3rE88brzQMUcloq9bXeTPPsRq5JcRF9bjWFnyoUllSOF4ipcgrblrPecWI
Nj50d4gDVSEBAMlqM92s8e3VcBeLSh/c3lt66KCCUcNzS4XoiEXZgh/sEhCUrkwY
2Eu/u8NSDfrggl6N5Ru0yrLHWkvAyXJgR8gE2nLkVPyCr9UyI4HeiUM5nJMrHgMb
DruzD9qKJrMd365s63G281NcK50bHFcCM5BPi9rltVxDx7KxROJ0IFi2E9TTbM29
I6XJD5qLAZXUQSw3gs8LvWzwXUGwPQdjDub0ejayYRKr+XJToMRgSAq+UA7siVAB
J8UpQMlaWGiog0+sAIsvB33m29Mzky9y0CVJHAuLXm34U8Lssyeaplqs09KY40dg
YNpr1KTEIk+tMEVGWdGTZa1Qxi3SovwMxiCGi3j6YJ94g2mzQSEnL0Nm6hDMb5+/
Dg0SHOqZxV8kcNwyklQXwahiOhgLAAOVGi2R632pDpco8lohvgjae221Y3hooHu+
QtUOP4UhhHnOhc2klNE4eyq1mw+CdTPGME4+BpX0W8D6ccCV4Xgo+vZaFuScSLdd
wmp9Kf91+YjM0JP3u64Q154kBXmI5mb7oqFZU6oxha/BCholznYGKyynmxqyah2B
sYZRrwZSEo0JMmTEDdfrC6EhnvVzwzucvhZG5nncy9FRqCpHEFOoYT3E8TYo9ZnS
Wn62qDsaT1ooAw/KvCmsBbvPavQcYCJpiRwpTpFg3CKXEfzS97hkEDOFzDzC7VW6
GOIGo8G91U/gWrq7/GZcW2Iul/HTk/6S/oNvFE1mBmYG/SRsjH6IvnSAgsYc/8bE
eWSmWvUpTVoL6GzGP4Ko37W8kzyxKZDpJb8fNezbAYt7UXxYYMM5h1JuiwiVYPFQ
TZgAo6Hdq48NsyeF1wDQGKiWaZyGKuwrWhlgR2G6T+OCkxyt2RruhLzFTvZWGy8F
KUJDRhyRaigAAoFZLrQYtQFn9O5olfDw8H2NRfFjW0uewREuELb06O7QoudAYvxW
qnpjhOPH5ORnWglAYst94W8sWqBZ7oMYWBmK0NYXVygmcEQWEH6WwLpNL3lWsklW
uc1Th2Su2S56NpbcIo+2yF8bR6pVjygTAPIf8he3TnZFVjMUZdrkqfeRqi8pFvv8
3cJsqR7HlZDyPAJH25R2Atu4BjekHvLbW49ERSKkVNUTxUJ9dCZikdX3gMw6I2Z5
xAj3+OhA9QxPMs2Zd2vRWQbIAedrHh8VbeFqp9AYSVw9XF919mVTFwYnM5cnJbbT
vBAav0xenAoo3IGMzwMDsrHNRKO2qQgBOMPrpLC8nXY8djUZcsJ6tvBtNbBYxBme
VpERu8trRpTCP5s0slalKHY8oYNkCesoegOFeZPFuks+Uiv0hN6ZX3WvUhjgHA0/
deak1uCeoGCKhrNC3MXUxr1FLyN5yhJDpYLqFs6fSiIhIH4ri9CaLyegdkGINKE2
AGam5n8XzULYnjjMQXHtMFs6L37yfjdPyMyYRIpm7a/J5IsW/ex/LqEm8SO8P2B8
XiaBsTCo/Mtiu4va7zje9IY3X+CnF9PxpC8yfbFWqqOgvtPnEMGZu3VUBotspxNa
XKbbuP5ixAZ9dcJkrGuCn3JfPbigpoMJ1QOF6wlV3mmErsAq2aJCuD3xm3K2qs8G
BxXEfP1hD6dH6tss8vRExZxQuVUROsjQ0j0sn3LqSmiJF5H7vjWJEEdsAf8oPutT
x5BDrsIxhy22JVXURH1iCRTXgjetoFKxrZuoGvTnQ2piMP1iJXNxMDg49UxbWklj
rpojvQghqeRheJpe14/r6twL63EJSYKqmowM3qRTBq20P6L0haFHBwKpE+Zf3ONO
Ol3gsRcuQNyL9/zDfttT/mQ8YwBbeKRtH5N6TDkgU96lAhcdACZT8g4IalRzIcCq
vX9eloo4jR5FVb783iPRQw1f7+iGVlqfGIQP09o8zS6r3tQeNExyLZCmr03ZkDRn
PO9d9atzLj9XO7izXq56u3nBWVqggsRu8qV/iIqWZvLWeNPVOwOs8mqIzlDcrQLk
C0ABWgD2wbLP+BD267tLUx3xIxfWUg/b4OMRrKkE1ORSUGJ4ZoY9tyV9nPb3AhRR
BHK9pH/Oicj746CIp/PdigIRqipwYr3US40GGkGixwjoiy4KHsDkT1WW4b/duqFM
j10/QIFqPtVevvH5P55zuGa3spX28mmzgmLw0uqt/yUKnKz9ZmjOnW8SvYVag5Bu
KWi80cDt5yJrcBp/kUXgD53a0cQGjEwcbjAD27+flvhb3B8PKgcNLtJYMv8RQD1n
Ty1Jo3EpagVZfUznbkqj53D0lnlPRxjI4984vWjfy+jqqJWxBSC2CmVQ+J2wItQl
o3/U6f+5Gcw4q5R4kJV90N/WeRPWKlgIQY6+DqStPiQDSjd7bnkjPVEoATdzASwz
owaNMk27CnqHIFpK2S1KzqNM2KmP3P6DzbnbrA0a3x2Ybq2YG3Y7D2hemMxQL/Ga
uj0dmIaNeg4mseLg0I8+UuygrkF9JIvFLKtSiczddJIWvi8R9nHDL+SV+caIkP82
M6erUcxIVSow/i0dQi6ITfCRDxHHTSnwicGtRH53Qf+Nck9sxMNv2maHYjt1H1RN
xn3VE+Ugc7QCNBeyypKw38LcMZHbtYT7bhlBbtXBEDU5W6WujhZ6vH/5Hoi7V9uu
9eg3qvtWNJa2RJj5j2Tg+CcbI0CsASFn2vVlYtbfZReFqzxWs4Or34/Mlw3nRsII
G1P6bugKlzM7FojrLgsrxaCNk9I6SXLb8U2yJQZS6502SrTvBVNCTuDWSGPLI2rt
fh3gXakgkGCTLq99sg5KE5qR8G7V0OJy5+aJDCsvXrOBc+C7rdqpTYVs6DOWShoG
w+yTNI3hVgf6QXYj2C2rFerKYMln3MpncD1gi7soPcIJtluxGveutw7xZ7cG5o1G
f/pbdBVn22HXFX4dDAZeTJ9LyjtoSx/DS3k/e6YaTbC9fVCacaqXyu/ekxw4xsoM
aEb2Mdnt++0A0NER0rirsYN5lOar4oq4fGqmrBN8uQJWlua+PnC55pD1Q8UGclWS
Fa0jSRggVJB7c7C//iNvIormG2UrtdCKgfGi7lIMMMHDh53petpW7rO9MBDQ69RC
Ogg2i2LeJtcEfygpTAZA9NrehrjEh8bYOHM/GK/zU5ZWCPV6LEv6UTJRzNRcXdWi
ZneptZKRqFReStfcnMTH9F0CIJ/6KR8yFJHsEVV95F0EVoFzMcJ2969Frv/WQiy9
Vkw2HNUCYpsQNWZ0ZEAnVeeE2NYa19VfF89TFuCtwyKwsFSCUFMOAaens4elSmLT
NFnFplKyou3Kdj297wPzC8Yw17OTiZRCS1UGfHTxFsia9lbnRIgA1J+xE2jShbtP
dWlQw5FADHx0qv/WuDUB75luq5G4Q6bwTQ2Dc9ctJ1ZT6/bWJ6sVCmbsIEJAGETM
rgmn1C2ogjXeO0yd1bOlZBtJ1P2pFglgKEXAZiaJHTk71RdEpfRh+0dNQd43DUhU
/C3Nx9B8oc/PxS31GI9m+eaoWNXTKJ9DCxLNqR+Ed8ebFIHdrCNz3ln2T0G1AZr1
etXBNl1FW53pma15FepGHJx+cq83PsRRkUVvOGoK5P8kPJoooq8nUnKYAXUw0OgU
QfiAMOp8AMFJzXIaHSS6l2whJC54rK2Fk6GYXeuwQCvzRFyiIluXFoyJt4pfdWhQ
H0fzbam1FR03sW+uz9chR7T7K5BXp5m9HOO4jsABk/vvjoPTCTvkCug2bhzfka9k
LWTYjWtgTdmT6YJg2yGrpE1J+Z25jiJtXZ2wxyujdydg7Wg/mdgtRADS1OigEYlG
WfL8xSrardj1w5F4IPjNJd+4YbylG6RpghehXYbV7AS7bOI+3zARbw+x/FWJYXvE
AP4Tqg855qwprRvuk3fNIevJmB+6eGWsr9WuVxKCUGrkSRoG7TkbYIgoriDSt+6R
OA/pkvwivPXd+Cmn+NMx3dFPmfXnFfoJvmeh2tJZt17qXVX8d426PTf3U5KDN2rq
ZvAvERHX0Q35LTE9HSVijofqEEZyQBd+GfmRQ+Ic23dtTVd/glWWskiMe5xwgUxC
Mejt4ABiOdKM0WKaJ3dKgleFHXvKS8ObBy0y/skx7Pkehk21/v//sUA2T6Z7gx9x
bOsGePtXEYATBXQeCbrYqEXHkaLiXbYNxHBBQrvm6FYUyt/i/cYyJ7AH9z9fAQLL
Vh1883Rjqz2i9UwnN1ygf9269tnVcFVS9Adlto07GDarC+PzkfboQumVAiL2Mc67
/eq+NN9Q/Wmkts5JD+r6cVm0ROxxOxaB6goRY/Xhj1prq2GOd2CkWrkegTkTmXFM
C9Z7REppIw7O4qnWJCzLXWG1ufZ4vETN5arjuE+N4PHg80EKgeaGbQK8gOg7fQ62
c5dsOoJkw/FMEtFYN4NhKHP09TmIvVvi/bf+QcNrV6F0GJq8nSDc7/vls814tHYL
cLxGy4BBK98fSZMWwLAloLgmRERoIVoy4K3Pxeuawlh0ru++1rUyjNy0a7h0QitL
qyeFEoUkek/ahQI+Dr52html96QrIpiuqBM9T4BRWfPaSjOmZcCCz5UAPGXw2fFa
NsuUp7gFaQ2LkuoHMJqvV4C/Pb6kvpr/0RNRmpaBB3EzqVhFUpvyG7B6+/+ZtP49
wl/1Lt5rTvDSzXkgM1/Z+hF2kyiDMs48sJc7iHn95bXeYBwHqN+3+/yH/WeWcKz6
MxlTezoWffAGajBI1Npyp8rjWz7Flm6qrJ5iJDOJjrQxwksJXiTfhmkk/8nIWvpf
NtH2pQ7DGR02IDktzaT8uAqkAlqZgM/0qV4vT+PWQBjzXpIIPQnNc9Iil5sXcJSZ
38Wm7DyAzI/c89ZDhDVZvgNfM1JvuUQvFVbvlFXO+3F0GsJJTRUakGQZRtzwot2k
yzGl+RmQN3P1oxozCFVfr0MVXoOJCQnylePSRT+2Q7j5v1+HDSfrmlw58bEiTYsK
kV2TvYxmnIbCC9x+fcDG+rJ1N+lz5yVcCLKCmXyiqCCP2HgyswywhaIIiHjNs4jE
RFqy8WNyqMV1z1xncCZtqCZ1KFGsutpkReXt4+5D4UmrukOggfWdLPGjxuGglXZE
CXlmEnwSDhLebMWt8gzCy78SkkFY0Ij6peff7iqLzrHB7fsSi77Q2XCEJOEZDaYo
vG1QWOml+icqoqMSD6uWvy1CC3IWRBBqssP4Axxig6TxsBleTD6aqCHIgqnVnjfX
Foa/QW6/raTTWg3KHvkVobnzFRe956rM4rSMUdDmLhGVgfqNjtRNbSWdP0XHRRkx
32g3ep/B0qNKy17qXqlnJDMfjA4ZQaF53dv1lutgCIG8wd6fifoc+sYEGJaYIlJp
L5lqHyUPq01jP8O0jAToWJcBV6RHA1t/DEXeynl+TXnrrox6R4WcPxcnZNRGTDb4
Bbd3HETAGy9qK62WOjXZKSFjxR1HJv4ChjMvYT1U/ouaog/ZvhckHXd6Vc3hK1RO
KZmxziLPEFoR7Dew6KrsIXgOEKlT8gRcW3r4sP61Gqg4F4NpQvx9VeHnzm8JCwQN
jR7cly7WMv/Loxpf6iPItAU6xwbhLFO3GsUzm3qjif+oST9jg69W5J34qpOvhMJZ
rFZi44gKQPSQVBOBqGt3YFigk1iKAcRBQBPxaVH5eWaxTTAEhMpcoNvnIs6Ecjh6
pY3VUK8jFbfRfQiMvdycQZXs013tXrLFSgLSbpfR+OwmOKc7dEG6iL3Hc5Yy/mbE
6vAbQo1eUrmfVO5FRciU+kmRsYjJ5D96McI8Vrwngqx9Kem0DC1N5gKuKEPTfbrV
08/znZUeDoCH7S4f6M6QKDCYaQyHDWSDMeISIMyMwuA7W+0BO9tftf4z20DbuD8d
UrHKXrhAsFA/WZtmOkuPK6O3SvJvmWpS3I1DfkIFcpHCpeVeFk3NtM2bEWmiieF7
MJXjHQK8tlGdB7tVVR2t20hpaSRH8Lhh2TfAJ3LJvh5/4gJipGp/Hb6wJ391b5Vo
dy075QlVYzJ/q9okZgixGzYn2tpJQunhVZYQM8M58NZhBEcMlCme/rc9Ssq11Ujk
FY8VxOFROGfOPMQwt8Lefqqk3QDk6PS6oSp8mO8TtMnTUpMc6jMc6Hnyv7lhi+ou
xHhCG3oPamUvSD4aROe3Sc8/IrPvgMumRI+d0zSAky947aendUlc80QpJZZuD9OG
ZtTyFgXYHR2PzKZH7PLsjV5X/GO537g9G4AdCfTLAyg9rt8RcS27pvpveu9g93Ib
wG1s9005Ax6uVg0e51HGDu9gp3M3HLcuHnL2gDqmuUGC1pHQGJXXgbaweLWoWtMc
Dyv85mlL2NzsV/ME/r66CKdGTJhjlArsZ5h1jzhfgRclWWe1JLQPxHGLnSO690+W
+kqmPufBMNYLCvAyWbMopqBSrDFGS6X6XfGgteIDKPyI2ze3huiccWnR9noysnke
/Y8IXxDKKmIM7I40CgdU4POULmawowm1FldGvzoChM8GhG1ssHsNxiA36sd/aTfZ
gelM+T2L2o+9qGsF+aZVhAZFpN1BXIPeK5ib0unluJHxEzhXvls0DE+UrktB1UaC
EEuc4+5ctGLLtHiFWimIzBnGII3t7uSYoHcfaly+/lbPpJmBDN+1uWodR2Nz6691
qJbBM3m0w4lKbOHNtFTh5z0ospNeKNChslgwzDGNtnLV/RRYxqtRvj08Q2j1cPzl
Cn/U3G92UUT8ZFPfgeUIU1pt4WN6o2SEGsVmWrW26TpDgCzltq2Tbc/JaZKs8AnZ
8jaeU8hSJ+WHF/4yMWv5a9RTxEmEJHd29Iv6zLZ7494FMDuCvCjQNiuMt3GmbECU
GkX0N1qgwQLUfEbtUmKVHVnnC2fTXeT9bNw+Np1YNU5Bp2QOEShnEUxnusbHY2r8
+UnyKSFc10R6mz4cU3ZtQXFp/waH8H40J/gMhZFVUlK3UoyiA2lQ9tDrlDCrfoch
6wXhQma8Wz2tA+2bNs5j9vVGyAi+bjRBY/Ju7cS49sySu7EVmppadG2eBPkL5cn9
QnmALGtJAN4TkfCkBslouZmz4G19CyQDG/IZsNVukJOabliKPiF3h6UHOf0OwAp9
x0eLJJ91znjGa6fll/H2FzxQivxkRwHturrTe96zWAP0MiW2eGZxvfGVKS33cat8
av+MySazjoaed5HZeeC2bPC2kai2K0kCvoSVpob5waACp+Z210ZOXS0cpJYazPMh
Qwdwed0vxOXKnqZsLM6I7UranoWw5bsgqYtsXJwZ1EOx5ZvBHErJrCku0txvb/MP
rw2ARv0HI/JqFF3/X9n+auWbi4m2vgTBc7J84qSCdoST+lidMvtvbI37ULcrsmW5
9pNeMkjE2bimrN+/apZjFHhfpXKUOgnb5ZiLOm3ehSOLVgkXzzSBnhRCSUmHpwO6
XGNBg7s6XBDlIzknVwAavQAmYiWbM2iJ6e1dv9X5F7Lzp2v9nQ3fLtwvSets7dan
nf6Fh+884hYKc2RIzRCk7eQ8TVbG9Pwmr7n8FVmtFzHcmrqkAcE0vrlJlov6lMml
tvjtNo2/kK/LR2dJpGpwq2blxZnmJ/h4XLZI9PReOsrLNNI9CXlE8V39oQEYIXtA
lhuEiCCN1yjpo5zmsFeYzB6yT1dXBjguMxOM4tGsp2mgNarYpZk5mvHmerLI7gKN
lfRH+Mz0rQ5UtFAaWqGtKZ/0eVWQbmhCxxH45laBICY7tojNE0wCdtprP6bH0T/p
VQBU+aKOhCm/zOd6EDeObguiJ5TXyD5du5qvAY8aI5pYmCfSTi+Ex623JKEpofY2
a8PiDDOvt2cKBetvGiMzTPuJrnc0ss5so+QErW5seMXbFJMvB08lfDLIzJ8NVopf
xa8aH6TBhObWzCiULGsD1x9MBhmEwGM9ysvqUrPwRH/engI4DyTFM390YIJJpg25
deoYFUZvqwDbHxLIrY0B6QUNUWWr2KoM0+fDJEwd8hJqmAUJJ2BmZaWIfwb+yJRM
Ckd3gh4jI8SCrdY9rd6dBwtPsxkNs0vA1EwCNl144WaYFSpZEZGLcA8ULhA0yl7d
Jyh6/+oADKCqlAhO4eBy379nHrDcyjdSldjah6Tv2+uRfCrmxxoZ0Ck2nePS3nwP
kLUq357oWNMGggXLcs9vudiYt+iypxxPNqZKHikBFkblFvv+89la9rkeOgw9D/YX
yDxh2yvWZCD1n5UTSLR/Nkg7oUlE0YGLpb+9+vYuSEp/lC9no8OIt1K6y0MOWusX
fAixNxX7GxS7PF7QYTcXbqECvmS0qVkWW2pJau1zMgUnDuPShmFaDuWSbVvvU9Kl
SQixpgWO8AAYn9hPI8KqMLo/rBC06DkM1UpCy8wGwvmli5DYfp+B70P4Gw1X6rqP
AVOI9OYV0GNPjz9iKxK2GtP5tlzHuCCVGtmi0CpVSUhDkekLzyBLIZ1lfmRkE1zg
B9tMq819DR3JifSiWvZ8B2vYozHf6RusVU5kB1lCo0E6ZTWKqomJAIdR4yDiHRxM
mkxJZuXCw/qjsdVRXdaLxdxYne4UHidnzIePiCYnWvHuOGY15gc4MKx3G1U4cO02
N8TZfv0AX8gn+nRd0UGfnzl8r9lP/UESep7brjCyDfqfBoRBs4G3o8e/WO4Bg78A
GuMdILxrGiA/Zkh262n0xGryAab9xfZ8AsiDiuhHIZVvs7rLOQgI8NLPyTnJGz6d
ypnul9XyC0vd2UkX9zMXu0I0TsDuJO1HzEZTKtaBzvNvuWwC4O2jfrOQSqQXWmVh
QvVhoGWFlG46+EBm+IqRL1q9uwP4v41do3Xi/DPQmlUmD8xFBsA6exPcNFNpRTew
Y0A2RFPSrt3Aq3/dn41TbQW6trefs4dMmMP4KeOG6jci1oNTw9HJ36s8dLxYlNrr
Axgzo9hijhipUvSsHlKHiwz11NWLIfakNenEEkkjt6pk3aA9AZ52Gl1bnLg5edkZ
mHTLPCrefnepgo0mWR+V69DqLpO1PnedztSViQw4SLMoMMZduuz+adJwR10GlLya
b0CO+3iLe5O3NWw9okf/4Srqc1b4m8ShaM0RH23ZcZWbyPy2CkAOag2/o5HEwbi8
udDLMgZXlN1R6qN84s3NN1TkewJQoUKFj1C469x148ki1FQ1tAHboqgcg371Dgwj
jViL9fkaDni8yJgwe++SX8a8i4+q7uelAXpCVcocgNDn6zM0DsxU3jtwVl6kDBQ0
KbdAzA3Xkuh4VJlOrjaP5EdbebjW4bL3etWY+Q3tsIxetUDYYT0nQgX6Sn+YOQJY
bLK+mjiZUxvnTonYDCqe432zkcs3IqOuUHJrb2FFeeTC5V1KddgTbT6WcgUxMNeR
FlxLJqF31y15kVWGGo8b6Jhj2s8WxBs4GCs/JDuVawKeYUOG6XEKiK9pPDydEzh7
HmbqKt8/Pss9vWwD0D3KaABp9KhQceQ3K63I6vlsHRtCOiv16cNezwyBDkSFiClB
7+cTIDodd71D8PXOsA9wdHyCh5pcf6b+R9D8TDqvzmFLE1gLGnu+pZMoH5dXaIsv
/1yDhjenbwG1nHzKgn+fdYmILyHW4HzK0rv6x8UoNGP1SxxhkCAqyKzHqktp0dw7
ylW37uIz+aB9HSeAu6/Lypj7fb/aFkRDDvwLXSIx+qG07trid7KgXQGfQEgmgh8Q
KwaTe7PfnytM5tO5X1kQN0krbWWMRFd2Jt4gv3bam8fCA5xSdpCd7IBoqG99tt05
XaTVj1ylGCNnOvWJKcAtUWO8Zk9yPowZbWUiZpcRU5TTndwEH/pC127NbnmApxue
C6R/FSu+zyfkB27qrZcu8lyXIphjcPRzK8ORQjInRTFgYJEmPEAhb/oZ2+iR54Gd
ylH9CvbO/HpLOfbmt6le/jdbzldNyDUwxYTkEZxgMZ9hSTszYSVC9ZDeX+/nw08p
xghfdCr5vhEjqHI7h9IsJLWNNh5UpDqBkqytU4OlnIPJ5BJrtWuGxnvqKWbf75Hc
kFOqFgmtgA6lBzzHSO+l0aCR0TtyTb0odsg48NjvoUqDPcaOnzqooCUv+hk5FqZF
gGKhRQTvmF+ptUjQnXi//az3IeNPQ2mhfNWCltSb7Gn9k6W4x3iqRse3uAh9usCM
hq/nn1TRu77NHAZ/a8GBOPyQ5Iy6/41VvGwyk2CY3G+DvPjUmJVidfcx46eecEXf
NIXsPjBNwGnWm5jhZTNtG+7GsiwlluaiDdj2XrzFfHtnTeltsJ7avyNPt3zeDhzy
GeSyokt4dluQ9JWPf+oygYxrPadeITUjQQD73cQj32XYPhNHsM4GAFgrhE23ViKj
cqOM7n43VxyEFcS34Zr/YtX0X92BGAZID5yG29V5q/W4x8u/BcnePT+XTPWV5+FF
PpO9YfST4qgGLPoZYL5DWi7uuaTmUdhFpxhV2nEvDbi69meYjFPhf6sq1eQs5Lsv
O4Q7Eo5o0pZw3TBpC5+JbzZV7YQt753lOExq5D22dW/q4OI+aENVN/0nXIqcF42j
E6iKkvXfFHXdVnCjbH9YHWlpYaPaJMJk0psselFnujam09Hx1mRwZ5IZefB02zHw
wO6GDHcXA2+zzzy081yaKGuyZqqEMMB2Cy4oCot8ksEWd7+aGX8K59YMuIjlYZOk
np61vVr0anOmrB9HHjzljBMtwiEuFiAK24TPYBQqj5bUGovmdApXiMs+NmaLGWLz
DJb3qOeQ1mBpNX1KuS1/4cd5ssfKFbXNnVBskE+7wCWcN6bO5FJv2lPEaAQjT2+k
GH2LdgtWdX9wl4srBXGqOGY6M6CXzdMOaQdSn5wLy8EhWnJ6WxwFN/Z4WwqD2s6P
sDtqJc0pB+fj12p4VBezuCBppSVGzSgrg0Cuf4x6g7GhTvDc5UvDW01zabfxgZQj
CNJrWucCcJ2OIxEfCAnTGqq9TkQXA6RkoDdNP6QZOuCV9JQdmuishbt8j4XAAcDc
/e0E9HBPBkM4JjnimkiuwRw2c3LmRY1sj6lEtPJET/EKrsq6USmt6zCFeEidk/Jz
PTsNGvBCmglWpX3mH37tfO6gykidSonr1mAsV7bwxC8bxR/I7LeFFAJ6gDrGaczb
XhmpetWiHCQ1R9fpm97a8EIYTveDNX39nLwClttQJyROVEh3Wt/qX0Xq4zC1pugp
BekMlvZooLsje4OSdgIbziKOyg/3v9bC2O8P3JyF7K9ShVmrNwyCWcwdSxx124OT
ZxX3ld0dQzGH08ZwTRE50TyTBTeJ4Gm5RqqtCDxASBjh3lJPCCr8T2gBKOQ7PNAj
0nFhmBNNiV3u2/LMJFuQK+I22ZEgCtVyFlpXcdOD4tMtncjnkmuT7DBkuUG3hhkm
LVGKgeDS1b2Oc232lSYWNq87kU3qK86Czwnt/O6yBonJdbL38thQ7e06WDBZW4eU
0Ej3HYnX6Ld3lFGcrTbXP38f5gwKWAiOMMPs/Gu/XyJDGDGWAxdfX1VV+lqbvEqJ
qp+PN1xPIwNq1hjqh4iO+VEz/ASWQOQf3OF6DvC4JyCRNl9CxDdk4pWmnhBncUEV
1dHyQvoRWkexAn6+Bh67ZgevNrQL2BeKgZGTCC52XwJRg9hpQJLUZhO5fhGJ3Wgo
fEbB4/oJyBUnVLdxuMS/XypyIn62nqGIU8ynuANKRSNghme+HjqMEZuwQPE6Ts0G
LLPSyIgVHzxDZlmqAorUV6XJh0IolqHM9jOoljG8t3MwCfHN3s7lU8u5szBHisC5
GSikZBEkpDl8hiLc48y+jX77LN5lBeOp1MR3bqz3aqu18rthaUgOB8rOh6lARCfH
v/MEpV/5duMVHWQ3n/lN8Fn5+VFfV8CuAf6Bi0jc8sBXX1ETZJ7ZNanI73ylZbzG
3JVVOfWFHaR1mU7v2qvsvJ+8PQ+b2Wq7ccd/LNxMOxRdUHM1Cecu2rq3j8cl7IE9
BuNgN65kzszAp7gdR/oC1YpGwugwVoqplItgZDPvnb0jwifliIF/rnpzQRpnAw+E
BlzGobCnIxBSDjOL/LM9agBgcVIhSfDVR+bF+DqwrKBQndtV0ViM5fjdVMS/+9qX
QpYNJw3DTWgVI4TkrXArj+nSnc44C4Hy4gDD/jv8r+NwTNjKP0ZSmQyCBYKoRA5J
8XUW0UkF8mKu0nvg/pwAXIqMIWVy7EnJKPTsNqKsbmnwfOZ6Bn8AXQ/TnAvvxunk
TReOD35byeI+KIaOqB+55FSMeCvfnKy89GXIQf1qIrc+z84SqaSjD/th4S7koH1+
K3dj+6h5Hw/8i/vzbnF0bs8Unjxh1l6eksD2d04cvIfnQ0zLb5PkutvfC8ca9lSQ
2dKfUP6GjsO0/XutiWph38IiErni+S7ua9HCiFNeZ6HPt1O7dwpriKv9phMQZlP4
M/MOyJ4VNcNK/PcxfpJmF5n0+QOPd6V/6EK0Uh/au65Xtp8JJNP3Iq5PhzGRt4JV
qTP4zsCA3tq37GiRcGu3xb19j3HVrADb5XN2qGznJxYX4CkKvA/C7BIwmFK/UhmI
XSpvXGMw3uch/KDmL1mnLs4UfkrwdYGDbIbTnYF0V1yPmYeHDyzoB34MVSTNrf/G
jDE7I31PXPdrMx5xp0WUpHDQbVqkTJaf1VCQIpOXI/qM4NcJiHGzLZEQOaXwUe1F
oLhQYvjeucdmkz9O4Zce4RxHD4squ27X3CJjwBp3GJlF8RFXasiQFvQynvULBPqv
Qptq6VQVPJ5oEvcBNOSJdyZyOzDL8lSDBzuM824PWpAmEFVkR8u+GRCjatc21Jqr
uQUi19ivkUUisTpSevgqfyQpun42owQRsKohvJ2uMhAUy8LA7xwrhZW/dl0Wx/G0
oogP2uHGBZrNR/aBZd0Dg14DHg63QxyOSeLY0Ohs6YJGujpVnUP2brRJzDmRkyqu
f1HDZumVh0W69sx/h3Zacr7h3u1ZnwlG3ekwVfIEgmSPGucXrZ+f3e0+lsgySdxQ
emu1Q9GfEHGR1vJKOk84it37STr4jwrzbcLswOo+i/MCmKAHKx5GTq945QEG9u4k
0ofZPwv9ay/ysA6FAc+xbG4E3cQJolVcRnDLP9DQj3ctf4+TGxHdTspRZwEvonjk
jdXTPHHkRtTGYu2LUpRbp7cgkKIg5QmGkr1tarVbrB18ebVxsmtWViCwfEat4Kyq
pT0pz801x2kVFEu68hAUlczpuTDpgvRZErcaPaDJDqftfBQaqwo5o0GwrwJYqjfm
HrbXA6F5BfTDi6wWLvJk8Sb1EN7RkbXhjFv/F3Bt6dQYu4q0Pm1mtAYOtCtLAWRG
e11FJsKmBH2h0PowKxQrigQjlPrBDm1i42aIfP59zJCJo5NbMdLe3mJ3a3Wmr+lO
UgRZ//Axa+tWhXY51YUklLBQX+sKAqBB4KmII+5G7EB1suhdvoJE8P2/Q3OQvUOd
OSYe5klqn5qcC0Y6pFaGK8hsrog8ZZ1iRIfrDhTpRpVsXzgf9LjeDExy5sVGfaDp
rTSGzcP/kkgCzYUHkbnuvbQxckAwE19B8NrVxSjqKDkDbD+MoQEOhwKSZGLkzc/k
ea1/oqK6MFx3QDNOT+85yXK41bwPWd+CIkNXhlMedep1UKeyTbTxnis/YiUNwMjE
fZjoI33BB9YvPxiBKLrq4w/0MRMxDxYU/05K0preE8fPrSKHVuMd1QeaobHAApnB
kL4tvlhR+qilqzxSRK+v14wI/aJdCzfCT2wQpyqMFQfb9wRp5siTqQ4ttd5lTi4L
oMkoPWBV/YGgsw3LoVPLh2W9SXcWDErtAjY+X6IbO98+KUJYeG1z3FHzgACbZZbH
FF/sPEw2AJlJiOiWOwM2pX1OMNFGBa6uR9mq0ocp1sYrJJM7YXoc10hH5+W3v37x
PqkXxJnn7S65Vuobzs9qGFHbVc5TpOzHVX3WnP1oMVH+j59J3cmmYUA8h4B+vEiw
eaW28W0V/D91IJLYy/AyD2zLKlvMSLKVr03AeYTBISN4+5yDjjwnVDUBRnMmrif6
42gWKZJUwwouzO/vzHN9kLsQBovR5zCLhQpr6hSBVJlKJDBA0ETw5tpU6rhfYJbT
r7GwZLi6bac7AXkw/UVYESKsYRbUQuIgx6yCCgeN1a0+RnhJhvtqOttuwrsbmAEI
oAI0KvXQm8hy+z63dpMLP+ybgA0W/GfGpnk1pjPfVOuLeZ8OJ778ChLl26r5ywkn
6DglA3lB1Q8m84feLV223cXhl9uXH8/4Su0iJaZVMzVZxlYiojonj+Dw8pNlpasc
rnu96leUcizWpMAf0LZ7hsRWlkvXJ3tZMgbmzYnq/DmB2h2bk415g+9MHeXYZqqL
GE3vMfhAIZYhFJgBmdyWWE+MzwBYYNHRJUvjfq/MdpfsEqBIIW5RMT65mXSr3E3e
ZtnXamBOzAxM+rNrRvBYPLv6+TG4wJ+WwkPQJXOs5BaXju8V5m+ozKnphNhQMe6E
Fu2zkqbrJy6zT+YWl6v3yw/AbtvVCXO6xNHSVGOL+/Fkbo6UiJ9uxrMR/0BrzKVP
zJVPymxlOp7YaPx/eT2VccAoSO2dTiTlUijtWnnRyGjHMrpt5Um40319dUjnrbsf
VwVpsJom1uLGJN2c2SbvNHmWxFP6FYYTAXPFE38vIXYLI5fFA964XvNRA/z446xl
ZAmHGt83WrAkCiXHthmkX85yBdJMvoUryS+jgSdkg6VJcaANBIQxhfOuVQH7qO9F
nHhRrmnpcMdtwu4VWh6teFBppU4A3CPp3eZIr0nhSgCiCv9iMa65zAtP3x6tIpP+
YNaK+9yXqPhDJbzK09TwT+xGRZHYKsIwp9BEw2bNR/Lp4fCwYy+0xjm/2Myfn34x
ZOLaK5uja8jhzz5XHhAFeaumca0PFTrtrw2x61mbrXGo3A+d6rZI9/PIqEiERbp8
xrf7/ue1Exod2L+sr/zaKRuq1KZzFa/y3HBapCttZEaM7yqVgG3MxjsU5xJqIrkl
M4J3qcjljKxoHbJWeKo16mtohL/uHrL8bknS2iasPvyku7KwvRNNPecBUNk908JY
cQeSgBvKpjTuSL20YIaqoHTemr78vMiEGMWRnKPJwUwmBH1DOBxd++M02PzFOS4/
P5AsRkpESEhqantHzYIRtfkhfn0qreuakFSaOTUlKlIiTxOcI392f9WW3NYqYUOD
XT9mZ41EIxaFd4eJ7WZXN4jGlT+rZSwCtlIQgh5ZQD7TQ4nOu/WDMSOC0QATlVYi
2PFO1bT6rZIVH8supxhSy5jbumJ1zKFp+H09h7oarHMHNxKMufrYZD4/NL1gSDKr
aCvh9cCiU4g5YmWbewlCG5h2qltGNBpevSTSXr0CA/NkxVLkclN77nsrVgdQhXAv
zM8EwZUYaqKE8gUz4fgMvpJnlSJUH9QVK6rU8I3XrMNxPYOfVLesSEJgJPNK5N5H
d4dMa+oym4P1PMIEe8Gv80WlVWuqJO6oRfOLYgaISEndlLjOt/Yfkijh45L0v2aR
j1UbDrQ/INcyGrLbuf3yQd8LW3sgQuJz9mZ6OrPSG+UGDBI0fFVU7j/jSgGwxFrD
hxxgqn+z3qNErHgcHHxatM1aKF16OA87E9sC1H+YhrHgXEuhSCPxsbq9nxaSJ6Ao
YdFnvN+obQsDosR7r+NHuDBcbHQnwa3Y/AwyGaS9ubfSJ59x9B+mUXac+iex9igS
ghT7bKGKY6zCPH4L47DmtOJ5yCCHXIJLX66CYHH7PAYssRKZVJyx4RYB5dv+UwvT
if10/drT5/1KAkstIGU86bFT9wNOrKkbABy0jcj6u9YaQ92h7BJn/aPMNNYV/IC+
qAWrk3DKznxAVwvLRnfvUIL3BsTejCF+3ze8G7/pwoSKqU5GVGGwR5inqOOHzqLT
sRlouIRQhGoj5OUYXgC3NNhsi8PBQ3fn6tN68qg+QkTMkb6mtOFZLJ96VsL0gASJ
C/TMr7PS6mEc0DMqOaDAk/6/v2qPtInc9ACDas1COGB65BXUnO2E++1A4KWogjy5
rlXzx6QaB6ryswMKif8EeKG8VIQP+/4rAb+IexlJ+FVN18EzlSu1YwBkunIfFNid
HFxTaEAkHjZhInHCo2IIeIJz3aLD9cagfIeh7yIEx+8K+A1p9avagHjRzTWl52JM
vRReOK94KYQMuGUj4Pf0sV04y8atTaS2IBaY2/AIWc3VXpvK5Qt4uZmIpT1HmCSW
Y2ElP5bkmEAB9dpg0t6c4zLW3OMyONE+kijtDd1JRWwjmZO4CbKbTTrstxHgd6+G
ZIbIFtUF2weVRLgCJO1r329r5zFWYfqDIu8pPE7m1OtWKES89lFOjCMxmbPOyVkI
qszVrVSVtY/4Edq5a2fY2cGEkJ/tUDnQc6v7+jfGMDLcrYaAOScKQKYizmAldnwN
9aleiVQQmmVOrCt1IZweuDVQGWAFUTyK0dI26SyzsERiRT/aQ/nPC+0qhyQmw7r0
g1T6tKYhqdzX99ukzfNWpr5TEIYcZP811fWfq3nAutHn5c0Q5hGbnQyanjEgKB8a
RwHIhWAnx1R7fR8vxbtCYQ7T2+v7Pej+oqK6tRyxTk1NfhsdB0AkOjTmwt0PGY5X
IMH5qehhL1glbTw8SjKASS+46H5qfjRbbNz/KWwKBGiXDb/5hsCvdcCALtEQ5o/S
/PQIxaHqqHlxKO1ZaTla0X24bWBx3PTJy1A61OmreHKa3JmiOcF6BST3m85DcXzB
Y4oTWNM2AKUqxQF40OPPxehpYEsU0CNdARarrsrUZQoHQBJGzcJ94ln7spLnaXgA
uT1EyV9WjG/4mD7tAP+LEDFDPNMtt2Kns7Ks9ntnbsPzmYs17P/cvQPRG96PR6CX
pS3bm+OVEtoypwSAzxgxGeHBeEdDH1vlifXzGYheYwTY9q+MGflyzry3cg0H59im
q/zvfYONDkh36A0F4zBYDXE1vn0rkPEsW1GWSikpsPfOy1+Y+9QoyAMoGsSeBTcZ
twUvfS+DXEpq6MhSv9gr0SbKqbD68zjM7u/o5qyUnaiNu0nhzp34KiFHpdniV1Mk
Kg2TSgqWuKviNDUDefVw1msVLYyWlGj2d+iaDoi+TBcvAsFI5RFmhhcoWAQ3Se+O
YIGb8VwiUdM3ztB6xUZwSd0d24bLMR1d1q95wREnfLkApvVApHhEmkvGi+k20Spb
9CWO8/fVery3EFv4CqFdw9sSQng/XWB28qwaZrfxAdXNHjTDqkeCUWUC3DGG89hW
cavLTdfu4pkNh+k/B111S9GePQKqZvp3CcJsdXYKWx27GbYPFaWGGFmn2JjpOyAN
I+HUtqT8/gBxDJ56KedlApoqZiTbawBn7sBB3ZMarHMUUf1rh6spp3K/k2pYsGbr
RFPigLgxIs43nrCAuC5F5vFXQRFnk2DMyrYd+t7avqCa6nvS2EAUHxxVSWPNoH6n
ITrD55fRcedJa6FsbvkbHMw4Svr5rDlWTZ2ffVZL3yt2XrKIVYApECcbeCj50i1W
iOmO469LxwNG84cRg9XN2EGUZaf3dZEvpSyfpO9WJL+30ks6bECg6EG/ng+wuOOd
180LwOtv4tiznMOtSL3Fum6Notp7H7h6EsHC2UXJr89dX59Eir7c8FaQs5K5fPjB
SOw7gbOzk/y78OPtiTV+O82b4+fZX354KdtvfJBpq0rPlCHMyYgsxLvX8/kbgiwj
xoOcH+7EIlNonYwAA7zgxxQGGtZriwAG33jrE/4SKFiDnhiwwey+8oLblrLiSFWA
8JY/d6wN//cY3LfNqnuuwpZrgMKsv3F1/SXnduQyxLUY42b7K9XD6XihbUJh68/P
VzDW9U0ylJBZxnJovHoNDsORY2QoXa0MhsuMlwhFt6XBfH9UoitKKsu2y18/P5eD
AYneMOepwRZVs6CaP8KkV7xLVLb3XhoM2B2gOhOHooLggE82Z7ywhtWn6oGB+zD6
J5AiyIYxbg8CHGU4CYGvFUvYnsRQT3U0p6ORbmlQfh0pev3GacCQNnOmkgM22mYd
luxWq+OLY6me54dFaqDAtjMrCZe7dcTrEeAshVY6Jsq/QjmvXVPsKaQNqhVs7j2E
9A6Z+ZI7Eh2m7VbMcN1acV98pLzjewCzLmUkiCJa7lWNfa728AMcM9G1YlwRlnnh
1TdVN6Ce9uQtUWd7NFhMwe2fnkBES/yYf+VA1Rkg+ooFSO2Tlkc4AGE2tiVBt3+4
rqLgQ0DTjkrd66v/QHXzStY5wXJCyq8fMYQ+kp3Zbe2VlDrWuV5v4q39c5GihOP+
EbO50pwYSAqfo1FZy/Rg/4jjFuKleKaJ9o86Z/uEmEhppzTurxFN3vpzTgpYGWRO
toUT2THmtBPf4tmTnZ91L/QejvdoecFqlh9+sKKxzHOXkMfl0cT04tN0oTyzneq6
U//yH8AqCMIs7ovDY4qYpQkrW8utzgsNUukHysyekQGhXhtsn6Ajk9guMrVXYZk9
cqephyjI+3OKgcIperNYZRwlgQFGX6UQIMzsln+4l8ioRxN9ZY37ZyPgBjrvX6pJ
F12vmoPPugpUF3wXqKfpqjCs9Qe8YxFP5krKmcswuDRPAyaJviwMyxFqnYcxFvUQ
xm2pnk8rxUXFKfx4vjftHFC+TQx89qdj9PyqGsS3/gwgLGqbwR4RWoUdYsNCgH72
54KdnKIi+36uJWicJ0x21ybN7QvBOAyvTRbCRD9KxmfVlA8hqU/GxItMWhna1Yal
3bwZ5Y1EFF1ml5B/wG3x7VbFJOjhxhfGNTJIX8Z4xG78ziIKqUu9phuygPg95S+B
ZTA+TWRH4mujO3KeAWiOoMrdhZMb8zft98b7yjHY5ovL4/VTbUf9yYg0n4lBjJFN
x1BaSzaNepX9Xegp/CcBtTrMRJ4+LdgDi1amX4ymdCWhViOPbwiIdfV91WbT0V7c
MpxbfiwsX/20LXQCayjaXiViPMzN4/+YbjjsDHOfeGnGd4FntsYpA3qHvV13+IHf
Or3ll0rCdehr43WlRHjVCjJBtpDosnEV6DFS2yY0S151J6ROBB//MELNyOYmXG8w
psZ11mra2Vi7wFqhZobEd2Wxjjs7bhjvyLQ7zCrF1JfFvH84cQ6TVwC9IKAAdvan
KMpheK1CYUcWDGByMTRiTJ+K7s9IMKBAlJQzEWnSsSUqWd9bXL8tO1W4ax/ELNnf
xR6Wz+aK6bRt6HGHzinajDP4NZmVxlV3kQimqGwYoh6KRTLIP2Fp8w2Cq/sLJ4Za
IrxIi90X2kTU5peJqF0GNpFqImAsITZLlzfXjQt/ONczvTrpG2zMO/kOAn2r5kyf
5J+uWqktRVDg7iv9Gl/Vqd9XYqNTV188HprLSMBEokhAlTJ+tCmcxC2hb+Bf8tIa
ZNrBecJZyXCzyaeouHStc27S3XWc03atRjsfqLoZzxs1SaKLPwCTV//ZblvY7YqC
lM+KJOYNc+fsMJc9zZakAi0BnLfa9jEMTK+4I29ptBxYVAXLiRuGk+iY2wSEraNk
mozx584HFvETanNXJzLHrmc1vO+1Ksv4zUcBMpyOTI9hM/hBLV7nilD330LqMu4u
yxawU0UNRjkV0JkPHjq2aD5WXWYTOIe7EU4+bgaVTVtFOTLOh6ecbdFCCl10dLsc
8pDqqVV4+XGrePlPcIKd+2CI6TCdJcfEpl15S6UmLMeQV0NAlnyNjPG/cnCztv2B
xZeTlEBlIL92k6Qo1tmFH3O1biHeSz54emAP9VDKFgbCGU4EbEoe1wZLE0hjSg1J
iCaMD/kSZjVbuKM9GW+D8POt1HsqkFOdghp2CBHhWpvLY5AWwsvM0xfwM+z8lOzM
Q2GihGYe/CRWJEA8FgpZiPOmgZ/DhEnt0sSWgUAUwkUanAEVtqvJKeUjMF4iFWsR
ARyrKq2paWX/70kMrWlbW6ecp6vSgKGkG7Kv4PhfkJuTzt+ArYzCKkuI/rjwhg8C
G41fSMnGIMKnxiGXD4pIj/5gUmYbYLc6nRha7fv0OK7JjtTWL1TjnOOfYVfCa3Rd
/A4K19kn2b4KsQyVEPqsH//lxoZs+diymdPKEMxbB2VYd6T6ZtaBudkWg3pBx2sw
J3TzlvtvmVaglU1JEq1TMSXuPiQj1L0q3g/UB77Ku/7HPjAYYGuzdusrhKSQw+3g
U2fiTkzgpKFu/YyaNRoORYLhG/lAKsRffdNkuUoNVJDlsiAHtHwtx1LQbyBwPLbj
qWWQ1Cgu8R+amQSVZ6fvWM/nP6jHbHaOMSyD7xZTNV5crwazD3vD2rBsFfEMivvU
3v8pT2rfWR+k2SDch68/vJB8Uah7yB7tSiKViPpk1OfCG806cXx5Q+hgs0N9q8bO
dZxFvyKLNpMdPEulCtmq9zL78uobuTas2mZjGM86IvH128rqp/davLO7lv5cNBNU
Pk2pqbkRahgMTp6DS4+f/mImQeRYVA6b5GA2rxaDHN2OfU84nUHdq5mGmOd3Jzzq
48GudQ4kGrUYM4f5riGOEwy5GRezRNtcB3d7zlhWDN62O0w5rFTSQaAwKKbzKGC/
vbZ5Mkg0QjIEkeo1OhIVsB+EaHNNt47ZK+ymThB7V2zHzQ2nr+qwj7cTzFwB6Yss
g3zBRGMy/rlk8q5EKK2r5SVQ6F3HNzqAfyf+eyWE+DKotvC4cFMk6+YCo6bqycPC
yQdSyWgy2hrAsS4B5+igxjIIPYmrrVbzt9BQRtAaiWACGu4EKTRYmq9WkmVKsccl
J+jGjiDTvCQO+rNB7DKGEiMIVho4QjxbD9U5HdV1NubrUSYSsBA1O/hgH2M25M+g
y8JEK6gUwCCFKW/S4aQ8hlablViSQ5VBsaZX4aSB12vx8EO8ckGrGDY06sxR0tJP
4C8AEzjsc+lyEo3PVFA2WoWGxTeK7rVbwDpgHljLxS0waw5OFJG2cTg8uhiDZZrM
FxY5cpUKbyEtGznaFiq2z3zNRimKGZX6PIRVa+V2aVgg8NXbxdmy52IWo5dCWird
K7xjwAtR7peN5G540+P9pzwWDTe3HYPh7yXO5OXpVHgz0Hl8rAlci1KIS2JGmwqb
jo1RcZ/UD5ggdvLUizvrvvfl5zgGjO6OtqLudEVJauaCXhrnuR64z44reyB86FQ0
v0a+E3IBl/0y4VzJg7MdpUEl45dn2T2kcly98QsW6qtnW1k4rnLNP/I0CEMLFPb9
sN/K30hs6xA9HtfzXpGJnE/hI6KjJ+CclDfJYyohpEsbxq1qN5RP7l/9TIVbqyDY
LtcSn7oXaegVxdEYVgsjEs/+WOwJWTSoZbPthWOI6lMpi1c0MDNIcaoVuN1+sodM
MtDfU4jCEK/FkyydI/z64wB8F8ZbuBI77I1tTGpKJxXlNY32Kr58ZVGQgUQ5c3Bx
ddpa8QgNKCKMHb6yQ1Krj014welSjLtJ0Al1oNAmpc2aprvSopFUjAbY8PEavQ2O
EEYEP0VLw79SWeNEY35EnEcs0g8husQmfbgcSjkeJM9vPnYMm1VNLOkTyVLyLxxa
Fpm5HEbJ8ouRSISaPicMsZkWTerUlxLv965UnFx2oT5+2bjW36W6SxHSDaMoYbuh
XrLkHu9nEi0Qi1J9f7mc+HlrMP61snDraM40sbFGRyDp1ZGf4Y+JPFSivr5UDhX5
o1O/tV81xfkfbMgzDq1L7byxC2icApeLBKKB3CGvFbQ6TXQK80FCqy0ixemlsgn9
+MGPCJzvzQCvC4oj4yLKcHjtRPn64yNgT43qgpGj7VdKG3HfFZdbPKaxQcaXDoZj
Rv3ctqwZblT+07LS59GYRK8zUCKFAdw/DDd4780sG5AUrh5KgdWq9RmfSzMa2whP
R8SUQiFF2KS82K6KJf1z2CsfKkr3/hzH4o1oy/001hZit/4wVW1nC6N8mYk75fwU
dfpGKfgPRLWZZ7f7uDMpTfz8A0sEvwGFFOex12ugUg7Ax4KkbniMXm4dMEUi9jXQ
pRJaUcYCzSJiFNOm4Ln+WOSM9Z3+EEMU4xkfQXWEQG/HAzYSRPxWSv20yh4a7t9s
ZZJ3IadfvnR4okkDtypC2AFyufbtB0VoOSL8kTKxjzTOzq8EY2gaCcsBDVc1j0Xi
iKxGexWgZ+eRIkBux8jvDXej/m+j+yGYne6EUQUMStXYAIoAuJHG3B6HA5FitnvG
76Lp0YftYFzQ70ySa+1Qxbj80mFTXj/PtIvLVEcYAw0teySr8g2GJvTrEw892GuT
S7ORWLCwBnK/dLf1SNRm3V83MkllQ2P4I5dNUuqguOzBulTwmjJKn/GBv3XDRZF7
2w7v7q6rwb4x+P6GsFW4euW6/w/tyxrZBllElhGXHxKvlYVSS6WuDkHN2UJhiA3w
OBv0g436TeoehsyIvRlbdoAeDQUbIksvefKCkMEeyF8SmnoKGoLcNgKeYuxkIfO3
ZB65X4sDaS724Z7RUF7b9Q8elxWkr/iNBC59rygVzVQIp5MaRNjo/k4JQYgQWsy/
NeRNV2CeKqjxK5vDdYyX+6A5jHtldNRYau2v6glZNcrxLVG94/qjY7HCE1Gn+oFR
CX7/E6K35p3CUGdAdxTAA858RJHzS1TXm2c1ulLvn6o3sLwPWG9Yq2UR/i9GyBJ6
BzOof9r8zuKAZYGGnNPKhM7nS/TUaSw/90EPFUsY/mhy580Qx06Az45Ga3GHYbnL
BgKS+u7RArUkIm/wAvdlmlnaH8UOW/kfAMstWwO6GEhqfWVcxDLz3dQfgCP1D5b4
RdD/AUMI8OIytt28ATAw+V5bxd8g/9Xvz1WE58tlDqznjyHKsobS3MMIoQR3C73m
KSNEHGUMkZATfH/g6F6bOZTW8XOuNLuvGL4pAJqr17l2Xc31EmatdlxUiOBLOhLR
Jbzj0W6vqwgolLpcM9PNXv+1xgBHetrifaRic6fm87OMK8NuqK4JIrBAfRjnXxsO
Shz/thv8i91TsDwAJN/ZpqkodSS9+y7JLxNAgx48nQhavhNRPqO7MGfnuQBwVjMU
x+FHlHw/8Gaq+trEhAot+Ie96k5xG08JV0vCqzIniGkrv/kvKBR2yOfL31XJVEcm
FisYNdhVcv2zZZADYZSmLvgSWJC36e9jgCgZRkpRI0nONZd5WfBKc1dVKl1X0LF4
uTL+WCbZ3MUlnEIqcO/D7L7Vtymko9O2W/IObUGx19mw6swGJDneNr5O5gqX6Syq
MhlW2QvZS+MDxkg1DV67d9Bt1uNEHeDI68njqQXIi4JQ2aIFFomDdLWAZjbqQKO7
mCg7jQgjU79nOihCwPRTvON6oOptCwrSWDYoGZ3ZUMEqy1mf3s9gOWy+F715RzuU
Y4l7+o+shktd5ERwlmmqaLkcwMCMYW4KY7oaaNYPA07Y+vnPs9sjpBl47c6y79HD
6DEJD9pZQCjoChzdqv1xMI7ZA2c83X1mOLN4VeD+4XyD2oagzKOg3beQYMf55EdS
Eckbi2p3zuehcqrjmEzI2YUvOpAZYCsfNI8166zwCGiJkxn3SL1Bk8U8G/wVCHW8
2gDtP3nnG/K0Uu3ynQJcd4Qtd63itD5CtMVkXOL7TlAqRF+njtIN6sMPVGtnO0wK
p08g4QPJNcZwGL6EX5y0CL7GnWjQlE8U/ZrEeYEggXuaZPebLalnk2QKnTKj77gj
QZlTLbj+WNKUdau+MGKY9oZ1A0WYOyN6WPGPS+YasSVoRQNMGJmklJLDJPkE06Wm
w49X4SU9MiIo5kURlmS9TFQW4x0Zjl95dHlElFcWRzHawq0z6RVgdq+BCryNd+GU
k/eLHASkB7RBnK5rgozh32YPFl1+T01YIQjEW+SwSBMxELxsgMs/Dfh764e416zC
U6rKP9gxmUauNE2j3YuRc2VGH6BUW9VW3VHbbanF9uUwKZBobLWX92aS4JRD2fem
J3wVNQSx4UrJluYYA88msKFl5Vuut3pSCYzefzFeET2b4833iiW7JJ5oNLk28KmF
S4bcy3SXV8f16K+RDE1Maq9/IsWQ/MP07Sr9LxMZ6rbsv/r4zZFyN21Twf6GRlUg
vp0+6nDr50dpJAwjo7EsonaM6Rdic6LOQGbWjVxWAjnST9LVvXss22FSvLeR0mMh
UEe+CptAkdrU97YJGShjaJA17cG1ptZzYGPJx9AiIpCLoMWSczofI+W4pT5/mXQt
nUoKnYL78k5rFkBYP+EubH9x4jyW1YoPrkJRQfmPCFx4LC33qT4Mma9xHZp0Iwsm
8+ZCN32LYSltCsCyP1TYQsVWZoqX55QpHJ7+K/IG7HF30ustwxNYFZrpQFSVOM/k
39Wt6E6qiCjs/HogAKNQoKBILi5dZR8YUNcaJmA4tN5savQCod5Q7337X8VqP1xL
i2rP1VFT5TRAw9aTMSCl4btbrA8loI+HgPqMav+Lq+eb93XtIMceFtLLqqnKP4tb
rD0eJT+m34CAv3VdR83eLuMvNe0ynAXuYytIhPjETwWwWLTD5h3TrnkUUW34/pfS
QExGV8S8lTUDhJ1UdZTIFSp9yqosoQGhajFMMkzYw9pewBMEGvyTyTZvqGg1AFE+
AQMIRGZIxke2q5Nmt1vT7D0dUToNzZMhstkzw1fpQdq4r0NLeG/FLNtAJEx+BEHu
HippvMK1RyD2B5zfkQWR0/aOIcunQUMZ1O211tWJ2HDX4EkOPihwjNw/gD4gxgF3
Qozzf7XvhLQ0hLC6r+DIDChvPgIZc3uwcMm02D1kKzGRvAAdxUm37bsKHE+2imS5
P9PzG19LbVTIpXJFx233xn+JESox08jmO/DwXxcbJ1JEVukxfwIcvdrXlVC4X6u8
XeoteYAf7GtwxHoXoFWsNC2lkTiVQekU4V9s7s87ooc/PYUE7hxqt70w2i3pNxDX
iQoy5WosLc1N1ZBegHeEkndLW/WbZRquotN82qJFCPGo7WxJXyxveEf/TMeXr4b7
0TgztA3PkBZUIIax1e0crGvjtGWsWVrbK8oullmyV20v4xrqQVTf/EF9IczxQz14
uEaphkWIYZnlw13zHnnmn2xcMAIBZhTr6u+jenWape96LnHoKSG6Q73J18ogl+pd
+kKq0UHDNBYn+SWJyQYpGISvXium6NRO2PhQ4EX5Rb6j1FjGTe1yJy9Qn8IX6dw7
8ZNGBr/bC0nnCIK5BoaJt7BrFtTU0lJNrLXu7295HJBIICCZoSdmwblIvvg4yBfx
1UxtmqzP+/m9nkPvQqGa7mS7NQpXnCRMkezP+8y+yU74OvZADwTM0NYRf+lvXQ2c
yovjSc0kqVFD+dTr379+/jLmYp++qrefYgxSQ+MxopOn6PaoTWvKOZsfr7gkUeMP
jdgjHICcbCw4tGG56DBDT3g1kV13h1t1yJXiKcTrrMyO5AdM3wDs7gyKG1zaJuDV
5fZbdBQrxgQ2gbD1c2rSfjVVr+sDruy+6dg2ri8kKfZZ8ybeLBlox2hOotOtB+7H
/ZNUrxqvg6aD3r7f+hqm9fqLDLyYbgoyYUnBKCnKqrrIrOVpbXKEdSAV8t+FU+Uz
nIsYvWV4BxE4G2TAHdbE+M0p7CaxgUHOvGcQqv7pYcnFZtupDxO/z90VGb8dn9wd
nH9HZQH34Dis/ZaRusDkMd8uAFgtL20g+6KEnFRpsMRhdZwuGScnu7LDsjUIiZN3
TGBuceAjdNI6/r1zSlM6P+5mymDnX3ZxUXBXJQMg4GU5OCRi49PHBm7zXBe+DKUi
Z5UyD+hzhDpO62DJHSK9k70qS9+ToFrsYGrqurov7Iel1VsGdWBCqGFtRj/Lg1Rg
GBvg7jYfxrlfQzspWYeawur8vrEz4WW1XwWW3x7bRwJ/nyKbSgfS5e1lM4/AXikD
aJad1wnR75ZOGn66wAGrH6+UD8iOQPVZgKctdqBNtqOme01RuC2Wn/w9twHMQs3Z
l+fVqwLSvvL7t9Bv2ZzrPIVy/jvcIWxDO0aU9PSFYER+TL9ahaHLgQKaSuJnKruL
tZg/TC0j9d1cd4688E1tD9Pakgq6uksb4awHI2tIOb1I0AB9Sz05PzjhO9Y5wDri
ixTkcc5CgQ3EY6bRNrcc6w0tKcA0nKDeZSewGsDqLHxboHkEqKe5dwJanYDzj2lt
Obw5dYCho2YJ3lFHvahoyCGShP/m3eu6xAlX5MUw4DdfmUtH5aM8XpGUWL0u+jQe
SBMDqL/7xfRL/EPpFVQIEXuqqkZjNTDEYfFR0+SUgxl74hjaTAynjh00F4F0g4cQ
wIwGYgTUNWhoGqbTy4hnAGJAI4DyQDhj3uiMsb5AA0M8ovXQ2b8JnwTmAz0YLUmn
5ss2eTqfMGkYc74FqQoaV4Iusm1qhfqmGC+OxwM7vdYiyBvq5NeHX+WVHg4D9fYe
k1cqPk/dt1IGfhXV0w4awNzhGSUDqJebyP0xJwXDLhLYUBjY4HLVNYj/3MUkP+l9
OJUl1UcYjjE1daXZIuRSIzHUU0pv9Kwz4MmN7oPMwtqitWbT9JLZ27d1Vq8AEIUX
w/GBxEW5UvTh+84fleTC68rTsuW51BmafRHQMiQvwsycqzZYb0DC7ZNZVW0Jk2Tj
cCPGLPxDj7Ntr/5aoClkYkFx+j3tXhVCWkUakYKIIhvK5nQlHvJkvhWKjQJ8dh0E
fcoH73YjhElg88FcIhQ6e0+uTz3qCrk8U6J4FAh/wU4IgHoRce8CW8bfmoOnTFdD
ibIJasi9LaUJwEK4pX4tCoyIo/osSWL/bu47aHY9s8/nVBUh351JzZRuXaN7uHQi
eFRFxfEvaAUghZslnTZI14ItoTmwUytRIy3y/qk7+2o3HSHemE1nBHMdn3XanuPH
+p2mazQPbBzj3S32aniLf/bREtOiDBc60rKeFnetDU8eV6ijRbCxYl4bXq6HWO9/
aDiKj0VWXAaCrDA5mxIVg1xGNWv/l1nx5WJ2/DWinauQvvkGIEM/uaeC5/8SC6yx
BdQIB35IpMIO3YQr7V3SXCuidWmiDLAV8Nx7speqEiFs/xzh2tguTXy0qax2FHKq
pjHwZgUIyrqAfAJAyBzjudmdC1bvLICdUhhn1lSCS40L4R15bcz4aXmwJHM+8g92
AeKYpUS4rDoAMC73noGT+3jwSNAlOntRj9oEhQ0orr42DhUyFYbZF8ML45u/5A1j
69QtTxZkoNPCdAVuUKIo0ngo7FN61Imw5prjJO+XY6lywKkuIw4n5aCgWHLD+Sc3
1SJ3mdJAUTeTZICZECxcZlW4ycyOyvh4geFKAts4Ds1Q0J1ePuM9WHzH6VAHH9GJ
7taDuEhowPYZWuR/RPqbzAESVv1izfbhFT2qLaIbdQYZ/U92vcBfAACnNhV3Kqll
/QPG8P6HXpJ6+HIqvtzPh3JmNx/0JAQFb0PuLKQTefntfahSiTMA0fs6ARy8D/Ze
Vaa9RlMKWKatapFxHa6DHrD2yqbn5DqD2CTuLYYZszM/Eiugvi+Kd4LRvXXocydB
c3TJ+6s3yG2IjGg3zyngRld2V5J1Q/ST3lbjW8QcxIKG3RI/JGczND1e34cRscjG
OZFJ+rqvcagfTcFTmUeLduRg6Wz5YyvLRiWWFM6KT3AfswE+WjLO7+civ0s+Mj3/
AlRv4oxKF1tJSeMzg0j4mqUg7/6yxMbge0nd9KS3Gr4smzI+HMdEvX4o3PqHUeBG
ciH7w/P+KutN+Zdkmol93LIxtDmYewreTPb1uJ/bd0Dvo0Nz7BPMdmA/e9CFV6s4
Qqqy+qwIxQZ6ubVWpGXSuhnzuvVIHs4OIjcq90ZubnM08WYlCpo3IWcSVyNqz7bP
SD9ECXcRGbhYGkcf8xrIZo1pxCmv4wjM2jr3ORfi91/nt/9Y72oL4PDRTcOG5m9W
CaiXNRo0kIEZm8rha08Qlu05lWOuYxcOWhsPwmR6786mw+Mu6oxK9WVEGg3mqli4
yZBcLlDAKOo9WikqC/038cLfD4FgBzdz3BJBu7LUUd89Y1U9ZJtQPHGq6mgBhTsm
X2gAFTtMwKphTdU4JBShkrYBElqc5cKBVKvHBZaTEPlnUFrJLnCzTL/atgqji8aw
oiVvvKJXhlpvNNl2oZZmxTHPappGOrmsWLFDS8aE9aM3UNYNe1w30Pqy6u2R9v/s
0qjqgEsqhfklqkxFkkzQaunjytAQ45KI7jutlZXzU6amWPemjglcGUdisXKWWVQw
6bH8OyB/MBwaFJ/I10K70HTYN6n1hhI8xXwpCZeLmXqoOzUXCWX5BOIVMWGGLUq4
mVS/6UauOgQellqkO3jBxSHkSgz9etXOrdcN0UKlV8IKrFqbgLeaUKdeDNVo9zOD
LSl8l9aQzco1FUfWsYDavl/tjVrlRWz84zNUypAJ6VnxfSW5BFgZheLsFTFw+Ra/
FFADp44LXZyUTfqT5wussuAkDkvERuNrfEp4hEx30vYqIoRxQZBSO7KlTI3dukqA
65+kVBDkmJiSJKK8D2dt5DxwheDaGULtmJy4QWJ3o4bpd/i+lJ08/lUuDnsc5q6s
avIhmWpOe381dkW4Wlf1xBd7zwuMr8PbOW3EJUkkmZMrmTr+qwanLdIvU52dkWs/
tUtkRd27MJpzOOz5MmJSG8ybpt6xo67TY9TJAzNSMe8+AlsCL3EvsxVd7jSxrmvs
5QYYOrU/x3xOsPPMFYef2vNTJzEnpwHGq2JMH1ZqNPLHfEH7Ll6/Mdd5GlKVgkxM
62Iw5malA9vRoKRCyT67Wr3l6fzPEN/bBnTTK6eF4c60xiTiGRnPRoWl+J+o7tan
LmrxKVtdQ4neQ04/dnXM7wjz2Z/Q08MxruVEk2CVe6eJMRPozEJkXfcoaj3uAc8p
czKBLNMLrABSWLi2ZXr9cD9uC/d3M2g7VS+5k8NoiOKATXPcJde8g8ddiVgP5fih
qe3uRo/W4q4FjPfc/7v3izJDms6dVCbvOjP8CLiT45lQsFSYLApgNmBb9BxOHEZH
N0+G8d4E4wNeLMnBNqhto563X2/0BSU8Cw4UPhfIF9ol+3HKKSNUOCqi3JLOi0ce
6yoPoInSsUY7lAQi2F6WUWpwvUqHNpWMjeiGlZES9x5Gy2Au8U8n8OcnOBnuLfaA
ewuQxbQTN38Jvwhtf0V2nk7u0cvF4MnaHY9le0NVAlxsvPNfFfuDDEdQ5SYj4wJX
xDcv0d0MbeWKaWar/Tgfvc7eiSnQodmdHeonY2wvi09uSVg585727jsfjMrNrrZX
RlNf9PZE6OlKWGsTYm+COrpDHNA0wLXu1yrFrgzPwnW0nfeD50aXOOIXquJmVXno
G7cemxz/DVSaLqhCRCnDnXXOF0RAqTmOpjzU02K830J5DDFVks/u8wnsXV4OCFIO
oQIjvUEGgGNr3hBduDrlyUE6RNnY4PqvLUFK98HItPAifNzYyWrnY93zXbTpcLod
MgOy4YfyJgmtSEwye9UW0y0wKG7kPUTuIrBN5NKnWnb36/1faSnLTc6tVMvNnbv3
25q86oFZcgC9GnAtozj5XhxdwEWrMVwS2+ZRl0fRcOBEzkSJFKdJpqIMn9N73Rlb
0OQUImmCtvTmVJ0G4X/tK6YV873WqGr+k2hMdPD6Ub3qOlE1vuDF17hIWNBemcM3
FIQ+z7WTWF4WblbST/EufHMaxmaJ7IfCz4Ed09X3xUgcwXskJHKw5A99Q+8Ww91/
PZKlYCY+Qq2bjpHLaLQgvlWIs1AVwhm8mP/w2PNMqkPr2Wxkh3+kyX+46yvXSdRb
RAS895m1usp/E5kqNvorqMsFU8bCscM0ujB9OtpPgvVwIDB3ggobe7Ba84MhDMrm
tZuCFZzOiuhhJVSCxNJ5MTOthQpLAnUjfoa8R+rC1y7xDNcfp9wjS5ObgqywUxlS
CpN0/snvRMLFAv9VP8V0UxA85MxV0rymepnWnQuXuM1IeECA7Zf98qBuzGMNo4rK
I1yleNHv6vINnNGT9NqKjxpAmWekIeRirh+29S3PcgsYzCvb6iDF7hma+31nUo8U
+Veg1YPQ/Hak9KpjDnOyw30WUdb78O0YZRhS8M2QxQxZ4Om76ES9FxwjmJYm+eGh
HGWlg7lQEWsBcoYBMxNkDHMX4rWNjlP18aK4VJ15gsAAQrpROSzHajk+wrhhwO7d
/aQKMS9Wla7k3BtSTbSWHlQt1S013w2yYAqAwU2NO5Fkvz7xpV1m99GQP5mKT2fZ
l95FQs4mffgiqRrb+6FP78FSohZQhaewXZm02Jv02yargt3C52iGzEkpfI4FwJTN
yRtKrwFK+rJuUyfcO8w16MEhjC8HMCFRUB1KwRQjj3qDH/VualIxV28TFiHEsJZ8
mwGfaq7ag4g6YTvrfOE4fKA1pmg+vHDblCYhhiMHsuc1EnHI4CcvrMvwGFMQ+7o/
8DZHdv+MN3+jLUvN+7Uvccw3IuwuOgxOi15AU9zkf5Y0Wm7arL2hZWEkrxKPT1T1
ySd4i7XCZKMNrh1k8K4C9vqXveQvsc1qXUKjog7kbxtLi3aoEPr8WiaJKW5YAZLy
DK7B1b6dRn3ZjSseOb9fAZCGmIzYogVdIUsZsPBSkMosen05eaJVOGmG0zxFpFo3
ToW1+YBcPQPzB56z7DoOLQ3fEMaVRwrYg3M/zmCil3pTYnOWTKCSiKZ38pADEZaj
jOyBpTaYG8YvWR8Yd3IhM5Pha/3Ryc4B+UxACctAq7hfoGgD4CJSSz4aavwQDDuI
HfJOHimlT5rgE45DVqZNIfHUETm1CTCc7TQwi0IuPZ1XkehgqexLNY8E+uWxYz8G
uwE24goAFA1P7Gd0BT2Xy09FMfPQs4NC5B897rFzaeOW+T+Rxxsz+U16sCph5dXj
UJFpxpbkf+gGvFz3/EV3pJ5jqM9aSNAlRo/rFPhg+oohTLjy+b/lerK2FG67sCCK
CyhGbk0v4Mgg3Jc/s0InpE1CmwmjVx6au3F5/fUaxRmEzTL1G8fh6HCfz3cSTGF1
AeFKQFyffDGextvPI92carIzeNocvWVsmb9TJjtcxtRH1khlJKxpZ7s/G2IMppBH
UY1e6uNawE5lijT694+1VnqUERfp8IH5jx2GcSck6mSMYWmYZOEg8sSVaysBBCL6
Pgm1cyVImS+VCiyOKxy92DIgEC0U7njLT385FrQVCzPXayRc+Ct+UWV096ysl7sh
6nt4eTrd2XViaGQW60av43WCJfxINrCUqFooAy32RqJdTHOXP/YOl6uxYFdnWgkR
FjrumlGnyft6Jj+h8ho7s4tVq73mv/Gzyu/gsYPj6evH52AoPXlTLIIsaTvuZKW3
JZqtqJRZWtZvs760X6CVkiB7VDnQjXTMdfhEX3WkwLKPuv7B8JLkmtiMnDLtdNWO
4NdL5Z+A1vNdist+1cc1rSdBmFaJ2HvNzlu1+VVwaurldR6/AkyH42tXKXiXrknf
DjkfDYXuGzZYzX0Ekvxba8B04pAHlAD0/jyl0NvZnqOag/iFDSPiae01TPvmwAFD
jsCjR5Vs2yiWBUb9CqcvWf5o5dpUUVbjs0o596Cx8h1CgdUpLwQ9OJoSbjYD9O7b
5aD7VgBcsrClXM6big4UdGYF/3ukuxKpx0yQ/n43dGpxkeyR+ixPIBh27hW284mK
03/0SHw74cm/A6Ywt36iv6FnoS+E91YWhchwItfIl4WLs8f8eRfxGeddSGdKGCsM
19f5OGMaJqPNcFj2zWVUcTyxkOFO7JFIg0bnQXQPWpVGg6RFuMF9dvYdyBWcTWdb
7BGwf54ZVmJipWS9SvxuWXh2+8h1tBqb3VlL5WqwQpWuqoVObIAWgT1FZeQ7iY3U
/Dgejr9ifJrMEx0goSSNEh6RiZF/I9CPimUzP75jl4D7Opv1CpBCzLMyLCG95DlA
plkKAuvh5Sug/kWmBi6MT97ToWxNd+XCQLKsLCzLBi3mbrPIaZllf+99sGENvASP
lyZazJR6H8ha6hRJ0As28zKMI1ILFkScBVo+ZhiXjHa/zjaaeQdjasIEV6UK+xZL
n5rnSmTgwwjN0BKmPYWR91Yhe2EnEmumao0UFbroW6lyRMVFaJxAZvhiX/waen/P
urjTz9nRFGFTHL/d/A5s6OWLMkLyYzjLEf1xKkzppDhbW2r7gADIrX5bUSHS0rjz
tkB3HurEKLwDHL9xNEVo+ciyuoqq/LDQhl8BahenmKFu20t3qxywTfiONKKX6Bs5
n44VNNehgq20c7uD3T/H68nDNzie+Falj+AuqDWT8d+z+B/To124M5+mZwXeo3K8
sVNg/XLHw+GVx/5wZRyBzlFDrgdh70feiUZuAG4+7kREj3zHlu58qWQYNCBVArZ3
67KfxD75KsTD91q3094K9lf6SS/wVOd/9vcMiKyTi1v+inE0AIqKA0AQTqLjz3+Z
osF9zsLCzn5sETMSgdSTTkU9OeQuK3Tm4+H8LdzvWjKMMMit0CcKEnxzN+O1TFH9
rT9GEE+fXVdJ4HX4yEEK7ME/dv9lhN+U2rlpW0hbeOyV/L7wvbBTDzm2094niSk/
O/BputAEVOZm7iCiHX1XmaiTyy7nyMXV3LPqtk984v5qo0iCzuN9tYKpES8lWFUa
ICwAVNWS6KHAfta9u8QZt3muSNyrwv6Y63rdpFtZA/EsvaNLk2yO7Weo0H7Nk5pE
ygAt9SlYevLQeFchCSsitJWSAElB5CApG43Mu6B3KpPQVObLNn04vEubCnc9xBgV
vgwMdW8LduE2lSWros6wydX0bf7pgKVeTsY8CiPZMam9mFKI/f+uuqp+w2j9y0ZM
hI7mhFjdJwPJwkZXpmpobJ8TFHIDcHErUZIoEIbJeFarZ79pNnqchC7N5ApxQFqW
sdd1dXwpTPKQP8aeeurX923Jnb7NBWFPXGfZAGFP04yTL1OITcCZb/w/3pH3sxw7
Qx1AnSqr5nvleAVRQnp2Qq6aCmf02b8eyOVaERgf1KmZc1VaS7EFFUucHJ66ramN
uU+rIIY99u09217gbgKjvlvD7/ZO/SrglJ4sBJfCEml46I3nquXLei95cW+/tmro
jrmzHvLq9zZG/JiIB0m9XAAK83S9KasWgirlC4eekvLTIVkURWgjf9qiWnye4Xsx
tha2HgGmwPaqLoNLqS6MrXgTaimEPziKq8ADiDdfk2Y1+O0jo2usM9omW5+fz/Q8
UOMyDmt9nzXDpMZl+EacAQWp4bQAuoF6pRcu49qutsy2J6VnplDHylBsupw5Zj9b
kAiQ/vAClLONtWUMkMWPB7etnyezpAcnrf8YEQyf20/jBf/N3Af0xyji+hxNbDen
Pgg57zrtNIe8WvZz3C05Y0gHE2Y1EK29Xi1WTm3WARo0ytgFEKAP686CBwrOS5gq
rYHmedRPskhGC8rzavbVMmy8PdExcwmMFY1AGhH1RjPeFEaoBL4QQW0EZgww703+
NSKz8sT9n0cy3hCjFtq+ybleAB5ue7v3aH6dSnCs3ez/FNmYJFnqjxwBx6jrl/mL
DbPH7F5zOpSAe31MmfBo3sw4oTYsnLDXgMFXwKCKZauD5IXFNLaum04/Q2ZoI2Ao
Brg20iDvMkS/0nFD1Nu3BXFl6TCGOU0CG/gLC1w4wYzM/Tbuqb25ElRjVBoFFX0L
Z4eMhjcp9ZM9mnfutshnH0mu5Wm6mu7telcXIpct0M1QfAoCjuiZDJC5ddpjKIIT
8wBY152rG3MKX7h+EDdJkVAjhdW1eTtGgDNi7fvtjGaYMzHyvhJqwOiTRvoKG5S9
tiunCGWOTQ0ouiZDwlP8KH+tEP3qP/GKj6ANE4Enq1PMLKadP5IEL73fgpYYbMIZ
dyBF5VbOwoYU7XH5oZgfQlvk49BMqpJccATQzGlgwD+TBz6tXUDKJcoykgm7ux3U
YilnNcY8dCMWga8K1djCpzLJOCSJOTQWtvtEjaRIOBO6gQLhCAo/Sbux/5qMKugx
1llnk5+B5vz53eaU/gHvSVMRMyydSH0Sw7cLg3u7ErH0iagHHjRsSH1+3BioqwFa
k291J4Z1kHIZe60HUkJ6eQBnYakvVheM6kd7Hq/0STKUQpmfRehGqGpmyLNIsWTc
UMzDGFXkdZShrbtzo29iaY+p62lx+YZ00d91IDyCjXX4qCKNcvu2ZwXLwjkhBxcH
6LVOw9ndcO9dcl+vMTOvm6kTxujn8zjmkVFzgYC8KD7+MkdE+OF/eoK/wKBI3GWe
R5leCByrBjBHAyn4YhHuCK7BGLDOM02xoKHbEAoR6I3rvfEdMyRrrRm6fPLSCMyr
rtJi4ORuX7eZ2r2u8pHNhb1jAIjqFIT0B2vTZ0WyKCKzkN0epqnYqgDK273Z3pnp
9gfksQ9S9EPz3GEs2oRFwGT+5XHT5I6y278bIsqoBySwPt0NrcukJFMk72gPNcxL
5IXfs52U0X+X61ILBgyK7KvCvSKsSSSx57O4J2WoJU0zMzLBmxcsQcuW7cNTUraR
o9lQKcre0yybbMewgX+lZxtxynCx2ihI5Fap71TS9U5JgTBUceT4SxRpSNG7aZ1V
HnxjAxmRtKD9oLWvyqJPcjB7Vxsib6jxLVrn/ig6oxAyMaevV03u80+kMiUzgiua
x8nq7juhCP1SkYxURDERzUjFpxunZqjnD0qLVn4xw5SRBFXKlVOjjVTj/fxmHRRp
KvqS8Uu2DuJZJliBmpLk9LwjSS5xCH3YXORyKdXpo+BtpA4u6pe14NsaoFNU4VEA
isvYJRIL3m9Rnyl3PEDJO7i+W+N3ZsNLt6Jfu1UdRLDZWtLhBkJHjIpt48ivdpqi
710oMzNWhgVMkm/PdAFVVbCHCb3lMx9CpJ7KTBXMJzcp6t3PrGDH0MqfjZbUaTBM
Bxyv9Nd8fWopo/gvol71e3imi995KdT+BzoAsh9NpjUBCZXix+DZOStMzpgsG0lb
SjDCll203zg7/1Ffr1nltOfH6lu8PinSW5D4L8f5Kuj5u+E+pvKM/OEZ3sunKGy9
2WdXqM/U8LglOshL2Inuk5Eros33ePlGe65OQzVmWRCXRgwdD+6zBEclXYJFeO5n
ndoFW171f6Ki43GdGjAtJNZs2VBYtKaWAJEeV7mzT3J26Pj5AarI7pvd/7wNb2Ch
dSibWQsUjDUtb/NRLeHSG370ED16BxRA3xEdo4WqDwz5dgDq09PkoQtY/vcZg6o+
RzfB0Zg7FaLeWChR5oPt4VCs4S9/JjXjXBCSdHTnzE8pwHdVI2EDL8QEKuW+655x
wTmdDRIQUnp4lApEz6J6BRxBQQy3ff6ig43avz+ZpdPmcN/qlMpKalQ/ID2icWLl
oRGhsef1S1swyT+9weEh7x0pF+waS2exoYf4xghmPy3gmVEMXswa0tOV0aIAIQuu
ruIbCYWQGizIZ0LWeIMuh4AojAovFmXC1NU0fS3Ae7UGL06nuxuMKozypay3GQjg
Fb+FMpuoVx2B+AAM4lKyOrf3Nga8nCDD6TCuoae0eWMpOsvRhgPrZKsp9WCFviwd
MhMF1alKJDBznmVZQtAnDifrJsj4COvAcvFFLcrw46Jbau9PBarcZhr8G8UyAl0f
yZQX8OTogaCP0dK9jxMwYSW4TDAmFzFs3UrjwEoePFpblUtoiWpvvoaN7zQYS3m7
g2BP3KX63LKHEqSBsV1S5QgvjaHJ/Qd4I6XaHR/d9bLXJ1ELIeRpYm4iFU2qxXwK
q4WxvE5lL9YMOJZAHkFYyXTslmx30wOjmI5ogpwmhrMOfaNM2bvIxcFY62v/zDmX
NB1aFIvmwkxUv+U05RvD9ortNk+fh4hMoBn9STIkXeteqbF5mEbkxEAEnnAD652/
Byvlvmh2WyPtd4rkV2A9gvxYqOsz1n9C16ItQJnlD9BBwaKAzPCJQaFsmqt7/0mC
wdRL1DSo6HxNCxvIoggzgr4Xnpb+PzA/i0xx2HuNRsK3KsbL1r3LmypvpWmf7wHT
b7lC+UfiufJRhoo4JPkfTc3Hsf4OYBgqN/4Y7o7FRqyrlV0I9VWzWoakZ0h8abzZ
uZ6UFX4en1aABIehTJuVIM8Lcuq9rLtuPjWuQYbmmxZBpHpWjkpXskwmZcuMHpM2
IaPhhVJTcDwVVMxKyNq5h+lycUA66VqOTUaoGgW8LGNQbHc16tA/vguHE4tr6C2/
ZvB2hfUOrfNd7afQQikJwnPCaj9moqDcv5QoU1lXHqnPOAbc11eBaLaqVyaZer0O
M2A1lpBcVXJLtiL2+uPrfa2osffQ3IIaqgmdRJIRFuDjHsIAv3zSo4XqLsW5r/VQ
gl3U3ElDPVq19Vk9L1vAqA5Cmj1/BX+dpZFFgCsXmqrsJSTHUh+RXDiMcAYFfh4J
MeurMaFOsdxCPq544vPFU0yKRJ+uImUKMfiWPzMdO/W6zwGIZTSZ4C1eMDLiHm49
jr1n/kIyk7Gaz/myxef8qWPspxh0wM663BDwBl5F2rLrumiUFDJyPnG8zsybEXOf
LqFJzKzCUEmFKnQKLaLqoh6kpiX92SSY2gQ8vpiIaS+hnGG8nkxCeCq7He4vFcmF
gYcWqbE5IHBJg3Jnw+5EuiMi0dbdbMf5r2uTTw08aC/TKqREO/OWvVo4WRl3fgS9
ZLXL5u33QEN4Ndojul4yLsPuPR+eJuDXUE+Tn2ByCjjO12dBH+5LGcmhX9KDxFYM
W6fNKBNeMc/CD+d7FeYTmVKA022pK6cMlgc/SX919AvaLp7MjtwopKUkdVWPCzaK
o7HYuCnR6R2v2gLC5hnjCooVbejUqAzbPfztZelwrL+y2rd4gkjP4/2GxdRNEOkE
s1pB7K29tEbS4fkQO8p/Y5r8FmsKEAckGvJ8gEkq7EovOCdLfgUgO4ut9eufR1Mb
z5zTipuY0LjHQ5NiyvKTaysbAmOuk67vgbhdtWPyFDKU4YauB2kK6RqbFgEyALjd
0EhpViReuFwR0t55i4VxQlWUyNBkMreq/QJoNsEuXkI6Inbl5fihDhpWmcwY6Xft
S4+NjZpzL5D7pl3sfSicdNVv4aETLI9dxjxzd18RePkXxHKdMIBDyqeEK1Q/iRXQ
8+Ak1GHwJcvMmubeQiB0lwyybB5PVwOeD4UqPIuuuNEztON9nlE8QHJdqMxEpzRJ
4pwEzgiTNNbk+Qoq5Skmc+cMF6WTRCBu37c1CYGUa8+hU5VS+hYk3wP+12r0cyfp
OHniHVuJq/AfDTOoetHwsLKl8820A8E9KAJrg2o9PuU7qm9m0roqjS9SR166oKhM
WNR3szIE14QAgFhsHqHgOgX9pv0IjXtdKLQ2LASCTYsRKT9slkKxJnMkOn4/9CFx
R3/Xw1SjNgDC+GgGpWHHuRlTgFiWNT4IIpaLb3NccEUY2JJpYjTujSxloqPCWTLb
uqU6tWGfYAuRFq0AGzO6qhw+WPEAkdy+01BRCZAU/oWOpNwf6svTVNlcgnAKbTYh
r//rmoiYfYOfEPzYVfCp/m36NEvu3ZqjOAM80BhzjOVcgCPRcDqyPfsWt/UQUHFF
Nosvmft9efopB4LLKhf8jkGCH0WsyHuruRo9KrO2VaTmwZ2bJxzBRO08iy/jti9Z
DgNb3MNrCxjCTQ8h4zorNRxSQGLLMXYRYlDVq1EpwwfnadLRaeZdwoBczIBpiRn8
kDJRQ/Y6ETwkNwclW08+aD4Rl8plco7usFIsFkqdR69899VcGNF9CQXWxdz+koW6
sHMl5qM0V9LCjR0q3RIw84qt9D3h7Bpr2sZC412GtSgGMI7fhhGjaa/U4WQ1FNKp
hy6yCR0zBwaC4/e6sizeHfK7xfkGm5KnOWg7pFDSSWkRSSkUhOd6DsjjeOJps8bp
616VSQCImrZI+sPXW0uOHTyjZW6/uz0IEj1X9+eAmROEk2Fprw6cy0pCf39BDhkm
uaep76opxLqOAUyzNRiQBFGFkDr19FE4FGffpwbGK8pOzc+hVFMdSR8n5Fk9vf4h
D4lmneMt53TZhb2vGv9gKIYsn2/xA3wAWZRyj9dJ/TyJAJZGxXX2lG6nM4D1jVqo
d6mGo0PVy2HPu7ZR6ZR/uAwbjifhiDO3bKYg0rjWDKhiTnVRmn4AkK1bvHvyv6IQ
Y22kzjrwcctecZLfpEfbM+C8R4gWHknoYbxS0V2UNi5PcmUG66dNGWFEGbvmEgCB
f1qL+yWrkzNTwQ8d0xwi7kdOpvwRKtRsv4k4wGO0Lm7LVH40+kyUI1kUkr6WujAQ
JcH+8yuB2Zpnc8z645rR+VC+NdmnXBR52a/h4kZ5rC0ViEor0/G2GkjoPKvI/Wi4
szWaPsmu5TRp93YBXaMDoWcKw8rD3/JG0zaFtcrQVTqJSAjfYBDy1uw0+G/YK0h8
7Z9LEBhae6rC1dNVshnf88oXhUsmKu+v15dIQs5XBeJEV31JPQppH2sOL2Qsz4ZJ
db+hnW/fr9ssydzf/DQgV+PQkDvqQFkL8vEWv/ch8EdQY3Zj11sl9FBJN1rBW6px
pnQ7GAwJMb9I9EiKgsYLHaU8Fr6zumalqfGp6getaOBOk9fE3Pml+dfBVD4vho9h
eZEB7eZNPRiGbHXNVYP3BiMXeT1mYG61u9/nu0qoSDnqVVD46jnc2LbVqR+Jj2O+
FLl+GWmNN5K3vDT3OOmCOYJvXQiQK9RNKhhLpZbvgeJ1Eu9neHYX3J1ihuSYcLHM
3CZEZx2siwNLbY8aJ5P+GuThClcqCBglULOAdUBFs0dufb5b3IpjWqspU3ylq7BC
qAsfx9wil0D3jpXFf2IIptUF3NPKvYCUBtf8roIk36LLQU/uGUmN7j9wLF951wwT
Mei9SpNjlcVoERrbhDFNwUVfAJYEcuoDJ3DVplBgTlBQFnl9Kwd3RcpiaqeYevTj
qDcT4WwNYiAkgtTt1ZTh9rIWWoGIw7n/C01vLh7cxoYKhdG9860twPuF+2QzulcY
TDCxPKnm6HVTjkv5VUHeGbyPUoFSwHK1z6sa4MuL54z+9bCADjt978cQPYRLe9eU
srJvS4N7QsD/wsxC6Kkt7KrjHm5hwtQ+IqXWKKQBStviK/HMlIw+8feafuC1QxfL
LIauCQE+J+mfTeABslsY/CCeZKUSaDS2Hqrshm2GcBUlXsqq7wPz99rtblSk9dAc
ArRm4aT3lJYQbR2SuODzxYK90ZZo4D32tHztuiD1Nis0V8mh2jVo8FzK5FMdRnL5
1hXRwYvXIrg0pLhPACgmOHDYbfH4TOf/hxqpqzcFvWaGG8p5BZj6sNttOlYricVj
1e+NCgDDntCFYwD4tsmtBs0QqttAzQgvq5hDEk0dnsTLQoE8R9u4VF5/WuADRna4
JLaG66GLMdSAUilxk5hicssPolT0dJ+3xiluMS8LVca6cCEDc/qjMUWrlv358dk0
VJuu3vuN9KcU11Nvs9amHnPbcCGHL+N3UNc/jdA+WwYr71Yg6kMP7gyfo8MEJfnc
ARogIiEXPlLK4R03ALHUC8bIH9QYpDn3FQW01NoqgdmSgvaVwCpJhnNkW3jttg25
s/0mXm1qSdLnO+lUcRf3Ublt8LoOCM/sk4eUcHBBOAhLUQTV+fqCzvWQxRcMZudx
lPiT2kp8dM24OhtHvgmWnDJAg9sAe0Uj14IwqmiwyJGrx/0w3MzSnMKpUGDCW1df
Kv34ZVsS876pkEZvn1UG7qX1NUUVKYYx82UT41TPmH3oQtju7OIgkgkKMtBx/0AC
V6t3XiAuXbQwJCBDHhg0yRHeFAN/TMPtK09Z9mG5Gk2k6ijcUkp5OdA+8E3rrcDo
0Q/QOCpAr6ThOautTchl/RyFy7dwQ86hrkq/ospXttExPeKcyixdCtqf6TtsxXUg
gBFMJ/Seo/Ew/O6Ld8chqQP1T6ggi1IR29SVk75eMnUOyitJ2Z7g02ihod8+/wCC
cTSB6VMuz5iLI+JJgk+xFlf9WRLIDyD1zFPCx9a2ARs82GIVcfhwkNjv3oZbqDfh
yTgr7n46cSJcSO+FwDxhoxTdXpeNPxqnAV13Zp02vgWzWZpDOhgshP8mgvPJOTpv
CoMSzs2IX1yu8XZ29yAzhJaqXi681XzfPk3sitCZSITE2NxN//umbF0PgPntisPx
jSUPF7/YKISkN6HQjbLDxyq0slJ6C1o5hDRTuUzuA8ryB8MW5Hty3NAvda1x+XZe
8eJ2rKu7TNzMRDzrtjbQbd1bFIEpk49hVe1JKXaMI0P5UfraTaJkOFfuMv0PLWW2
UdQM4TU4nrtVMoIwpi+yCpM29dNMKrIK+KlypB8BBeYcVcCZa+0Ey/zcmrLW6WW0
N2VkzgIoWgcl0I4tZ/EbZSu0BWjdjs2VeTpdS0GoEeXos3dLgLU7Z4O+bUItShTF
nZgiXF2MZ3Tsx0O1HCzJsxHbwHMjpKxmkC6ZhL+GB7hp8e3zgmffOCCDSxsDHeIo
OOSp+iSdL/DYL9usBUfcBKAlZIqCVr0twrnLs1JenJbK81um7rxGGajiMFQOuoSL
bQ3q8lDnx8genyyomMKhL31vcGvqBJ6kiyjCg9T4aYiMcqMzAvjn7Aj/fkKCxN/6
7gbuN3yDDeJWKKYT6VrVH3tafdIzgzUtgWC2Z/3FoOQh7MGc8/iEAvXVjcYvrSSa
m0KWJa7LftZZWXr7dGV/UQGRD7zZPIfNNV0OpQjkUPMPEATNkuioolWIVgzJ3Q3J
C0wahYOpIDZi7acutNlubQ2io+zcDraifKoWMOAjvv0Lj6dAef2/gG0fOzN07N7/
Hl3uYiEb6uXO3XG1xb2cWyV/LAlWebMykXMDTooZWfzkTyNm7yxhcDRY9mbtDVIO
YDof+93B0jtiVb7imA0s9uJZLrgA9RE2Y7smzbdi2iQgFUbIGXaM6iULgrc96vpK
2b7eRfXSJkhnn5/GvrPNWsyGCD+YZmyF/H3uqPRueX+3Bd8n0vSOZOrzOYIvmFKz
vIt7w06JITg1UOY/bhWQAkpNRfrP+T2E+ixeLqpzqymlM7jkupIJWnKCj+u/rKHd
IGHncJge+whAWOE19hJzOztt6ZelmqD9DlOhZRnHnz6TKRllzK7zKxl9YyP9g0Zf
YOaNKM+cBmDiN5/6q2Ra1geRbdlunA1dIGSx5zUplN44o2QZ0YozlTbkM26RhAjO
HjXmjhgNzUmpAsjbQrQC/Uz4GkoSEDRiNUF39DaZq3aVXdp9VeBn5bO0IaORbzGF
PqJhcXkNtktZs0eOuMWI4C+AbVsr9bRmdLuLBq80mvBSpbV6LBpY9k6wGudYcS8U
3/mPewWW/2xvZY0ejBosftum+h5DkXVqYdgyfn+Fv1PIiHYMHGU0JCeWQf6WikI9
RargJ3oZlbvuB/EmSAwL962USYshM6MiFt2ioTyJsw7931zDjnn2cvC9GQXEJr6A
fHJaA5q2RCYMTlOh4AXg3vWp8Yg83OcT8ytOTixkep80mqaak7l1Zba2VugyfOic
2E2lM3FOWUl3YH75GzFoNaUKwb3xJJCHAsInQol5QBmf0MbyCc+f4Qs/mdDcoeQA
PryTJVgIKQ7alUvbQFGu0VX3mGEnt1agjpEpXcEeoI+ANFHp/ELterFfRQrxZ82e
yhBO2OBejRVopHtxOhiQSebUMLme+wfOWSsGRXNsq3eRZl8tb3C8YCbkgiYsoDnw
/lUPHk/DQhwTzZY2YrAIUtG9F5MnrsxHW3NZYxL6cIF5IdDceoxSrP0AaOeC4LUk
5EPPZkoZCDQGAZHLdaPU7L9pHJ2dpvSsGSDvr4FoMYx+4uZ8xAJ+P6GABxdoqaq8
2udrhNP7dLa2fBTPaXWVlNBNdqjF5kfff6Hwac7geJwDqT+XkFsg/5N79iNpBQ3I
B907rH0/Dixcsd18bUxtgozMXOU+mhIZ30HdHIqBqN70hlwWsFeMPhfl96IiJOFF
22WUVsKqrY+GRXxr5pa3FEfByyhy2UWfYKBMU2XHwWFQqvXHgpoO7DPYC1MAhm+i
ogVt7EWgwJYJXN+11oHTPM+diumvH5Hsjlp23+nfaMDa0zJat6jI73qQD0eokUly
iEPNzgWceG/8b1dMfmNlbvGLwcRQ3h+zUcUVKmftR4cZuPjmyH90hOqGvpT3cRHQ
Am6tcAuqhntdIBT6L4jm4vENafAdFyQcZnLj8fxQgt9cyQX/Oljm6WycyhtTf+jt
NSooucFo3sMGxA4if1Wl26msfAHlME19RdfYDxH+dvSRuEq9KSTlSJ6OQc+bBsi0
PEUd7MkCf7MI658kbBTgRXJnJYD3OYG8BlzRdDT9wtnj1aQbq4DK4ySSkaMKOr5E
ildgqO4pAI3me7Wva4Jgd8EAg9uRh9doJy70lY1d9YZaf25+bW3f+20gEfha1oUg
QYo5pudTOjqU3op8HpHSzjn5duALS2IyIo1h6DXFzCrOhMYdQXX52E+QowZDUJVw
5yl993yCBF0Qn1BqD4YL8IgYNjrN+Fh3il83VlVanJaPPWMTOssrfGcNBo5+FiUq
f2mPD5vWfHSHM9KVo0DZGMVJqihkfueAvW7eaSOLNE0Oh3Qe0gMBSbhMMPlaOPeA
1C0kHQHJsE6HsOplquex1u2unnCGnKi49beEN1LGE8+k06wdACd+ZOQQ3W89vgRo
G+Z5OKcmYVSNYhmTWVygXjK509V9YG/TzXSU+egIsIOwxzsh7oyqcWpA65EEtccC
oVcavic93WaJ1dvMWQF/9oq/vXPu1iDp4seBRqMQ3tqsQmFg6pHJPEc+82sT2WNe
NPEBzK2WBjHTAfMEvTmqjotriC03rshELiC3bci6WS7ABmbvOB2suzYwo6XM3X0k
J+asJ1UcrYHIumfYmmye7udhoKytJW5muyHE2pyS5mR5HvRSi1TzAXXR2j8QTDHE
oaVVB+ITUogAXZ67w3FSsiLi+JepNrXw/bCzUjIYbGW7HY0s+Rooz3Ft2taw3KOp
P6o6DBoNhBucTxLs47CFd4euPYG+IqOX0pA6eLv6xH1WNVviICmKnfCiGMKFk2RG
PnWqa1rmOX9D2mdRGV9vQf8A2eEAZuVKd459tC2m6L8ema3RITfPXvgcQvN9hoIQ
sbIW7kjpllQPQkBz6T7H2RkCBUBHDbs040H8TopOJo6dir6WIuzyvm34kE6KuFzK
92Q813gS+LD/Yw//h3mNMA+3E461byj7ubiV9lF3JxAi51Ib99s0nMhl/fRrY6DU
48kdbrsMKIDioIyHX6YPof2/5dsr6aOdsnBe0nzg9zMBg5SsC1v4kOynNCFR7BRq
O6rjxom+kTRKRttU9dk1jnZk/8HY4aXAH4mh8SNKbLiAgIJOiD/PuM+BMAQRqNTF
WumRh8/zQWJFDkLJQZm7HtW9jq1c464X8stz2BdbKhUmYnAD8/rScpeR9/yaGYzc
cOvDhJsk47PjI/muryV316hw2dj4flwWs1er4rxcrOgzr/g30ZEU7HOjFuwG9rkm
0xrm5oTeAmKAsx7XYgkr2PWHB3qyMPSnIVrRLK9qAbFevBRUB7W0p9u6HHOZulck
k2XZMr/Bdfj1CIdtZ9gg/yxxNyw0aFCIPA0e8euGR+OkC/TQenvzH7bDgqzqmJK0
aNAg9WeOIZqHNaUp3gEGmyVqix86T5x8NDTbLFWmgCGV9HNf0QBVsFOuOPn75s40
/M/6HqUMrSF224XzJQaCqx6Jh7/QCKUS7VPvQHG6IP7iBp14sBzR2JwBeKsrtoDS
X+B/7CXSJaOAXzpz5EBaTxWYetZ/vX2azKLh37s0NScRlmv5jRn/4uF1ZxNwZWOZ
ABMlVSXI/kyh1JoJDnjILV700Jx0tgSblV21IpR/grcy9J+4FyQi08VyOTHRUunr
/pc3zY9r1bU6Tu2VAa/aekgfCmebMCiIIOxk6hUhCKDKuSkn5gYjh49gDHfTL/JJ
scxyjR2wzKuiDkkcbiBSYyLHUaXTpRKxlOWNVAGZMT3i3x/ndHys6Ddw1hJdHkq7
h/Iawv4lI94HXk8wAtLIwHgBCag8V5Ux8du3E/BI05/kLL/Qx1mSNbWljfBKvn/6
mwmv5uA8KFEAO3U9uNuatOHnw9zMIjpEkO82pLRsKYjUxvWmb+KPJ5zDMe1y4IfU
wVgUPB3Pn7uYs5pPXBDrcilBnhwwSHmzbqKx5UQ/ZuHwyEN4HCsS3YknxEMkNKGW
CQFw5BWUwGKrcgeiD6yL/1VA1T3rokAkwHEWotjS86kIriFlr16EGw8mKjdtYyCN
IT6K+5iIheua+r1UE+2xTovHPyClmsFX7WDn6QGtEBp3On2y/ubDaOYdhZUcKlNl
8JHT2F7pbWC1x3+gA17VEXW39851LF1FdJPvEKCS23EuTU3XL1JyiCQVkUBPzpab
n+NYGwS+TGIkVld3eRq4h77tEzK9eYclC63/zZ6/rge8FV0zbkvixfJtt59d3hkS
qg9kuBZW/GBZhWyu4g9yNz9Hf6RszQ3PJdO7rcjcRs3PF8lZbz5Eac2IY0GVjjHE
eHXuFAV44lulCvz3UefRe8t+5IyoLoOvxkNFX7mGv6AU5nBZyeBCcntbXYwygxnt
/INgvLTfoDrsFkAiJus6uM3iqVNPXEL76iVxWKEs9QOAH4/wZ4jEHrbdt+JaVYaZ
f6E/XsRHhuRxOqmI1G+MD3YgPdH2B1a5dN14zQdM3Klgm4dQtn0IXCwmYGTRjie/
c4tW4aSYZaBrWAyaUUx95vfRA1m2Wxx/1TUcuWb2SCbKdAwivV1KQmB2XczKtrvw
DQRPgXKpciUxt1RQMsDVQLsu2yw6s8DfC/k3wsnCMoZ/79uwtxdaLjBGeOemmvux
qGkOIwykNJKhrQfikRVmPm96D0bq8hEWtxWbvr8U77jGeS/s5jRbjotIe2XMooSd
KN+L1QHm5V/kE0u6AMOwp3D9VgIVg4ZyegG1aT8xdg2lfc+oQpQqbphipG64cHhb
97UY3XWn71NKvh/RKzLOQuql+8WwPPu8fCXJvy0d+/oh8W9Y6A+xFq3UUuPY8/92
4ct1953G+Pdpfgg5RRJTF4v36q0AO7qyGaEvcc1RcODf3wRCjQBL/OErDll+UjmJ
Uk+lLcrKFxgmFyNMTQaeG1n6VfbyQSefrZ27bBlfPTe1T8doY3KLfXUMv94TQvNZ
RuRCpBm/LhtHDEG31Nq2gBmak4pLq/Ccpske3KTl66VYVO9eY4CCBDPKQPn26+lE
QwvlenhksRCdgwZ+Wjg+wInlaGRu0Wywi2aS6whfRz5mrtl/Lekv36EirxTqhqKH
EsSLpCJIaTYAu2EEks/jOZJOFTlMP90outyJOUVBih1OBQOS/NoJyAOf157x5QdE
PNUpcFYcwOIOw9LSlAYX0YKCEzOxsr04pzwuZTyVioSnfloFxoX4kKTkFbtnK8QP
bU3QH7p9oABZ4Yj8NdxsYJQvL1H39oq/kGWGrzLUzI7y4SqiKvvNshE+wpPErEY9
4FjAEnLVOGF5gZEL1ZM64DhOqb/cOjHwH8tQOCWHN94MA9tUP/DlnungWI55KM3p
ZvWvLwbfKxn/CZi+DwhlwWzNNgOuBRq/wxHthcOD/J8iEQi14XKKPwP8shCFDd9r
Fuy9NKhUVnxflf9kZV8nrmu3KokdlWLmIWL2r/a8JlBM3Dw4j3l01ryQkCwczvaA
2RyRqEFi74ftjRL30HhByuiqMGzVzdysgD4iOCH94jUklwYqhLK+2b2YFDbTubxp
K9M3j/cyjyCode9gNER9/fRKJC/o79leVRCnuZ/dID05pculNcraHOQX8XVqoIwj
gumGr1ued0/W/RFSagvR7txODiR31Z0lnTjFBji878LIhqw1ydwxfxZ7izxN0H0I
/JLrkmxqmqHBAw6oRDlwDoMYqmHita8fl8fwjXKXoh60Xtdv8zytFSAJCNgZDQ2B
h4oAM2c+O7Si02nrTQt/oSJqyD1m85KD2RgANW+OllR0i/W+DWoj0wjyXa6NVt6d
FQ6lhQjZoou5Tn3XZFWyXjfNZl1o3QpXNyBbrUvGjM41rKG78OeykFkLCePqnYHe
G65/tSJAMpqY1CDD33pvW9IyRPwArswFsIgnQ3TpSPm9+0j1rn0/CKeW4Wn2BShm
iJnk3M5lBPVqUpydmK6diXuUz7jI4Aj4G5BXh53TOpZXYvLfcBAm/AQb3sm7feJC
fMCcnoALSC9qx8CCNW1OP68jGboNGV8ALd8ZdOSqMGVRRFMxoaboJks52EKDuPmV
Bs4g64gd7JGiVrXkiWCbE8YDWAzYPMxmDXZdUt0iZToltPho6Aag9I5Nav+No7Di
lpkuYcbq4gQYadH9+VaHRKAsici8JLCbuYT7jwZh7pcQK7H/jLheugE6tvw4M02w
bt6ammlSzJOmTl68L16DzWb43DMw8YXbK+eBXddME02LDpRbg1Qw8x8NNexx3IMv
o0FcRUnxKR+i+mxXws03RXDlAErgx32jbGmfvO71iySJLeynLKOScdizgs55QPux
/PYR1AIVK0JD5wEiosYQfifwyDTTha9jR9GTwbMp1HNAaV4G5W1qUMw9l/Lmni/H
BC/8yyqDdLyKo8BpDKNKXxPEw/TJlnDTK5EctkabMnL7aoEJ1k8kGjSIRecF6N6l
FluLD4B2sqb5EVuNS5uWsaWStxo9IRk9b8qB5boh7Q/oNTngGYjXi8SamJd/x8u/
C8bRDuewYdPLnuHMeRFC1FgrnoktIR7lfbKUvfl6pjegvr0M6SQiGAE1WfeDy36G
3rT4JJcHuoQu2e1+qQielIB7vSeAhI8FPe1cEzXNUzRtxjmBmZZxKcbRIysvst7B
diyc0OZpmFt0UyWWioo0ugeSaVY4/JeW+yj2M+0XDqtjW37sNsq3BX38MbbJkRCw
UDBNrwmXmVrAKqGo7Mpc4on16Lb3uMbr3L62WLEfPEmQSGKJ5cP44IFyOctCd+Wn
ecYxAkHqoCAX1jGtBHOcD27wy/m5IknCp4/9u9E7+SWreahTEXSe+kg73Hz30DNp
edO142lx+D42XdzBmuu6OeTl45lmljQdNHf5Yn4mVmzYkzXqo5vUQsLeSBbb2uhC
jSwR2SmPcWordjZ/J5hQ3qlwgTpdULsCgWJ5OBzPqwA4Wcx+0RCW3NFBRiPKV81D
RMvFYl20bSDfr8QDMvrBMmtu7AtdaXfX1JHrWoQ5l9z38mxtQskhUKDvbTmpEBaa
y2SmF23MRv3Wm6TEVFo3PY7OZYFbJi38+OmO4IfWm0ha834355PerZabq0bGuVet
gHka/WpSWargrzzlz9d9rJ3l35HG++VpOI2FL/CLORHOk/RAXzRizlW/sbmS2gm/
hYjzIU7FFT78LQWEQutXn+LF3F0Ls/5kx4IejvHxmp3fzJj78Vyji8yRuhooJ/NW
1WMc1tr8KVaUoh9eCN13xMUrFguKaCUTFkffb0bdwsq/+I30Z4WSgYebvmIZZTch
6pzkdtV8zEuXWCS/iG2jcj+/OxS4ystFRFXfBH/wBtlT9zLWB1e2uMABmTIgVnm6
KBmTKfB1o8PBY6fpc+UlVGihkCzditl41anKvoSLWEwT6LL2bDeCgwaFU6CRV9QX
o/81+5UstJbCZHHvlgZOhmIGXOM2ft3bhlPKYREsgy4jD1v8wYGY/S9eUNBiRQIL
ji3oUgInxVFpViL8SlvLdAiDY0mErp5T7YI2yTw9TnvYTcB9cKmPcsWO0dtz/l0J
J0IV2d5WZt/Ua6WIAwnFz3inGO5VYjoEgjW1h1C72KzlliDAasl3qjK9XRFp0ncc
kNPZMxMd+WVFpPGE4xntEtoex4mBxzp49QDNUsxPGfJ/criyxQ/Bi33gy8+dNIdy
rkIlns4jgzGDdZFabJ+PPmCL2JIsA5mxnTWuMXELaImigFyukkCjYvg5NMDMMCme
uUJkAQNwIscZXPBEo6yBrmIEu0KsDL83ikz0zC2ST7KwvcBSwSMusX0Fz0loFNzo
ADSodZM2ARHqO9vZaKKW9yLsqFO+/gxkiPu1p0Q0OOa0lov+kAW/eaMc4FdqB1Dw
uVPQhQdatokB2l4qqg/8HLUTtM33OagDByAHTcQZxFUzHd/cI9JI9TcBG0e4owS/
s07Er++1h/X0b/viENYaCzd0+c92VWCUwl5uvVzVfpISRvvgNJLwT4RqBgGY7F7I
e6pou2ZaeRAf7LKoigKFgkbSSYUN4VLrY9KuaCkn4ZaEmiVnMYIj3ALHdCOkWX8S
TG3QXl8OYjjM96L0jQR/TzCPi6DaU7oeFyuXAT36aS++cjx0eNH9Z/DogPPndxH5
3D/URHv7mOg97sJkAIo5WFFEBiebsD+boqWzgqHwqpCQIeF+pimvP+TjaF4+sXQS
BwXeJEif3OhI9u9OnYazG2uedGVZf53KrAZV5UG3gAfkfMmUjSNvYsCelQNV6X9z
i+7xIqxSveQIsAuX75hXRjfL0e+RfLD2e2N90RiUb5VV17PPzO8UJgtYBe3mJTR7
TYuE6LFzQKcLOh2HoIePjbXLXyAT0ENsepD4CpIr3NtGGdJ6qmwiP40Ek4LLV5FK
X42bzNceN65AK79wbYVc+zNaf8T3PFrMOzhlGebxdvlXJ5gpJ4pyim7tysPXgZOi
qsZm78Ar9aOZxitJrrJ1xh3bp3P8HPZpYZZR6t0qWlWC3fsRk6f8/5TTwub05SoS
x8whaBWq+KXHyE6YOjGbglWj5nfAW+8FGgM2Jx1aQctM1tLx5hl17TK/xPxDeDVI
L0c7FP8v2I1wO0yhsKCJzRmu5DovVuQPjyVFS3zRqXjRFDHp8o2bJIZi4+qQOLHx
VSMvFZkURc/NqcaqL5cbIPR5jzmKYZXd6ovCTHnsY/HOUC8snjjOVbSaionqp2bc
IwMVHEcxXdqHTpS/Jc+isAajfUFUpebiCCIwssVAP/Vap14hdKZCLi4E86roIa5w
XB508UnpKmJw72MN56dpNUhBtGuG9P/n0sboJ6WNru4IyOSA/YVMTZubX88af3bv
Ra4Yrnu0TyimUs3qXMMQRvh95zzh2UwjReGLW7BBXm6/loXbsi+JeuBrCVdUcGIf
I8nMQnsyQfKEeeSigAbhm2oxoxBoJX1fdpni0J/zD7szRW3zdLyRV3oXoCeDfUFU
yRgtmbcZYefvhzhpJhqHVPiSbS0+U/KcODUwQY4feB4TofGbSXHlQusTBDJ+QH7c
6A6xg8RNmoInelXPRFtamz82zGBLcGtruSIVPcn0EBaCAm2uaV3IpD9scg/Pk782
Kv6/nCA/iXbLTieGF2U19n91XhqXApxYmiX0J+tRRQdaETeuxWcfkl3rZJNbyk6u
dH+/oMadhl+xD1c0O8vlaI9hzv7xbjCwQbOkd/ylXjB2Wl4iQB7UjPf5CXsU138v
ag+NbgNk8jeGce3qOdvh9xW+DYEviHSleZGPwS+FdB7z5Dy+oKHrFupCnPFWnN9m
Z3bv7J7dbGJNxhztz2j7XeNjPbzhYpeieYXFHqD5gZ3nZjtAKV60+gAwUy6/b9oK
H1IxTEGjwqiF2QnHo56Nvo5KiRmle6pFJ9051CCkWpzvniWbp/R5fIPRr1E+N621
BPzhEPIquYVSmQfBHy4nojMj+JwLJMkDLmH+9KMcbb3Wfb/HjUrSvY2i4pNRXL2C
ETAsHuaJqynXjzznqZjBTq+hGQiPGDirR+c3ejFybTOq6xE3owFCoQdGR52MSEiu
N5+Aq0bprXc106XtnoeMRK7YkHNStmmMYWd6zm2QhuiCiwW/tbzV88N5CdLcrWDU
ewmG8ShrcT/GGiiXftrzf4KCsNAQ+b+1EZvpcHH9uR0DQ0LsMms1S8VHPlOXbpM7
/j1dUHaeUEvibbfmtRRfHglZxT+g3ZYHN35qYcLlufAQlRrAAyA/drirvqxWOWxs
VoZ44TfePf+pkKH5j2Hr/3L3VQid0AYrCQk1YKgScxHpf2uhYMrSh2gQgMJskRNJ
blbkCKRYpqPxcD3sG5WD417aCkN+CL+ySdCE9SouSjCXpBQpl9KOW47bbEjOuxzH
+0jo/hpj8ULK5Shfp5I8RG4AElfoRuIkkIL88oJbPOltcCGt9zVoX9UZwZB5g59w
A0duoYjoWcSYxAaO4lNm8MT2lU8xiTVB0IvZoGqotViZLQQfiVcOxcIXjjIbQNSg
zFYfDBsi2nSJrlIyIUHPONtcO8zeGq5+dcFJ9jmzy7C27yGd4N8ecmUmEoHUKg99
Ftv25gggMy9sfHYl+7+1Tigs4q7RWw8vJj2lm8i56T+VBLxQRPFXSVOFfPVLEt3P
rgDWsEA9tuuj5yz2P5v0Ti91NzVSfBOqsf5KJpgMQeHew/sznx6EzkcvseAx9NiX
GjGr1nTRFSafL+pEZ+PH1Gb7hABMqpTf8IwaoGVr2iq+WiLowFuz41aPMr1YRs+0
mxzQaQvEIx7p7Xe3RbgINWeyj4n/CPyApcPwEMDek/wG9pXALdp95F2QDsdPQbXz
9cbAQv/6jz6aKESD9KbBPLYusmq693K1Qd0z1h1g6zxGReqpr6wzlTka5SXpvbh0
ZMsdSbk73epypwFJ3CFQ56zhUaTY9ZhskAYP5v/4Q7HFXC0tsH6q93U9Sv1Zqa8W
q+3QMCcBw9LUvsymDNOeESAaYVmeYVZ5FNohmIy5G+sk8AkKTz9zls6fS4Ywdov3
/ddDhDA+NWgVG17C5ka0GBBoyvaVvw7lYhb9XjsUfe/v67FHIF/3CTLPcxX3hXn7
vsFUo+NF8huA7IUoVvct0X1LztZX0AzJ/ogGKTg6W6Ievx0AQwqQO6/SAYrocW+0
f2nxkTO+QckEww+9o/lSXMTKgTh3WkXUoKzmR7fznx+PpsWXw7A0WCcd9fA+JX68
X73tgz3P0OXNW24nNVEKpVqL6OFDIFKmBFk/5GimRuhAz6feSNKt2zTyObKQcxVi
fkEVbrGGZvsp3EBJuT68iwPHO/RJtMLz7bfGQwc3WoqcIwBtkoNf1cqHhpfByE/W
cX7qZmCFr1FtTA6ml1NItKmHjhBF9xK35EZDFH+Zskbf1dU6rwXbzNEqk4ZM45Pc
j/e9Zbgh5wOfoN89VX+2fZ1Fc3tevQnFiUpK6D4Pi9K+e3t1zXr5GOefXkqWUBW2
djgwzkA4/tQwz2OkWUQBlUZv3uktiQM7J2J/bOJ9NHid5lCmlP6t823YkiPKufvU
Ou57MBwPq0VcryzfefY5xyBo+zKHA4QMjgofJTGfVxTzYiV2Nuf6nS5mSzfdRm7x
xmud5UvONaRGPCKQfIX9TM0D2R5hiP8gFvqO0jGfIqMDChHNRi3dSRZzf3SRIbvr
qPaXTuk82nM7qJSkxI/WmMy6X4ml6JugUZE7EmMdLAd0hsmDNc3juWIzqU70TZ/d
h037Zz4Pq3zhavbYij0Fj39X5gO791VHSgv5L6pmDDokz5yTSx0WDgZpt3VOZli+
Vj6of6YLWPAkUktQQV9hDoIQ8d6Yw/FOxUIMwr1jdv1ZkMVaCCOOssutrBbegkLy
jr2AKRTExgs2Xb9gl3z5xv3EGpE5QIGbNljutpmoPQh+HcAk5yehzUDD1KN3rrUK
y4Q5hR7MFSS+1EM3+oeGsdXVNAVR2ZMzoPvfO+Vyw7pJtLwM8ispef5jZDLK9p5Y
/XfeLUzU/7qoEaHRcQLwO68/GZwTqAFecLHfgAGAXI8erEbFevBGrJguI0CBw7Ao
n+/H5sveho5UV+IP7XDkeQoeXd3Pg8m0ShfDlqzpyt5YjWLMK2RlPlVKBDaVyyRq
dV1N/BVw7X3CYlXp4BXHZHDCl5Du1VUoepe/D74jKT6V/55Y4ZKhPEq4HmC19Dzl
+6fM5upJW+4XTvjBshupQ7oxAf0IdUi890uHpcFCqpwdnaLTcX81K/PRiEH6Fbw1
L0+nXDKUZh8UlYkTsimwdqi/KEFIsiKryybmtkT2V5ORarJd5oVl3MTE4jFla7ki
zdmC6Os+lMVC2HAnM0D6dcox19EBwXz3WZYTfa0DDo/s/ryXFaVjOQaAETm1KP6K
TFxgVDWarbmi/Rz6AbSyI+Y4Sc4+O8sEnVoYwkau3ob/7Gi1zdTqgWqNA36lPvpy
CFH3ly3IG6hzz7G8zwIzORju85wNLu2szZYcrzV0PKKVLWwpp3MHbPGNLyzRZK79
DNeR9oVecAWbuHGU7McyJEj7X1CgQZ47z40kC8amKbLLBvbyJIPL2enjvCgnocdT
Gh2e8QFGpOfYPSA5zI+8SwX+ILK2Pdo7rXyLeK7e1TwaEkJeIa64xOfBCkak0dZp
bWdluoDchakPUCE7AMs4H3zVu5KIjsiIDIjoFHWIvG1Ef7P75a+X6Higer05XSaF
xF/eADTXs4WA0UqfpjUbhEsvXy/vGuB6JOFZJCf2cB/hJG68DI+9Yjb+sgGU5bbd
EGisb+Fq21rMQ70Y70Vk+GKxZ0/ivS4zWdZPlGwUo2lMMs8ib0Xj3CSe5WhjP0jK
i9GmEz7M3pBvkZQjp107Esh8Kejxmqr1GIGV2niZ2dK3s5xRPfgFylCpi9VgfgwO
U1BKiu75IAwfUYBkyo8uTiZnsWA8TIpIaxvfLYhLu16qCU0Cyt1EzE7/XZZ1nKZc
xuN1RuNPHwfT0SiXy5Y4XSHLQx6nRfJH77vRWO3aebCypxmeghWVe023LqsY7CnZ
gqJAmtdRNX/1wwSi9wQK935B0lphip9b3rvI0KCdUEVtBCEMj+aDCxaYBLxogTVW
USooytFHf3bok6Vb3DNUV483k4+XJat3gX6jcHpX+PJjXf4RqFbP04RaPhEzAiUg
SNVNUeg++4+OagBr+Y0ou56XcvPFDkHeTs56pqPREu6vcFNLyvqyMTLo/Gv2Vdfh
U+879+yVArmj0nfOsbFQ+R/giGFaEl6xO+/f9eKNCLyc2Cu/pfcQzBOMc3NqzDVZ
Gt8xOkBOBW4W+AWNTGcrCj66eyEHwlV0Z06dk2ZIaGFyC2zI/4GMNQjNlC0JZG2S
cFaK8mH8M36U5CUordww6xzl9u36U6Q14iIHb+LLVcDWCWaVHfSXsF2DRR2HUX5p
U8gwteKq+16RbqRvPj7fE09QRpzvD6cUgPajmM2R3TI/X7OC42ac8PTAzNsuDTAe
fu3kSzxXQuefF04w/Etn9sHI7yumptTc/E0CMF4xQPFEvh9zFehyCnMhtsuoyeZL
57UItIajOzfeODkMu46MKedcQVdpCjV4cX61KCkBgHv0ciGS0MeDlprHFiL286mR
5QdwDyxPyvAvV9QOzB1wmNkvSkMXLNKp2fctftHkOVnErfrhW9qYenptUObmF6EF
MdCMZ3aw7OwHxAUCL7Vwsn2C+UnbeECNU5u9J5qTCHwN3usSV0pSpQE+LpPuSMA9
iKBQjAr/KIWpwCSVSzh9dYqejIjcWpTH0S96mZQFlfbK7cUmYmbJRfmyygsPKKgv
K10Y7kJQHyWMSuvVGr1LZQiW6AfeA6ZFCLYzqDXSYUTSI83+IllrWhiCphLm2S3q
LATvEmyfFwWrm9EKpY1H8O+ApyNPHF5W4TYUvil4+UFHI7NLPmpkBIjfA3k2f7Aj
eX8hl34kOLicA+59diihV7wcTajywcb/bL0onx7nQPLGbxMLEmOWABB1oIMDmtN9
VXE6FvAAqtJLR0CUzKRFkhDwtkGv1e4/JzgMQVUpGsg9QlWFBuSXeAi/1XPZynLc
cTkDr09Sa3my8Nd3ztowKw9svtb0hWn9p4VdkQLQoesaSoS2PT7u4CqkMHmozQ52
gRRA0qtwr+gbNvYjI0U3Ai1+x1RMwtBf8dvV4cOay5Ckgd5y3FX2tktnYJybxbYq
MjC0kVilBRpnhtmcA2RcX85t7WbokdnwrCzb1QClw+gnxfEn2fLLmSZV4bieKGz+
zxfQobKkJCGAw2fRbwVHbnFnMNjlJ3dwO68pXCKY5wJTkpmoXo7NYO2lZVyHan6v
11ewimXEDHZ3wBDfuxcAhL+8aEAxff3tvX+NFZ1fYR27xv29uPMDvPrOpLTLIfqX
Oyx+oiDxXIAlZM8d9QfkKvKiSUIPWDwr+9YFGhZXRFDwKZHH6knYiTAxt8xrgy3z
4Yy1a77sMOH2gcXz8c0FV21L0hefFLAt6GRNMEzvdiz7Uw+JkjAnpBYkRgkFAZTi
0GIXF7xeaaLbGVrcXXNu909QAHazGSEhbduOV4Qkf56k9/Cnj/QFo6xIS8ueMRox
um5zbMI6jF1LI2EwrBsJ4m6YOfnfx+PXgqaK/m9JaUo2A4nJO7wwgBWEzI0tFGwT
48tw9VfSzAgKXL9sH8x+1VLUWQGAi3eYTYrGN1He+rObbJ5C7K2d+DIgzSDSBjJt
xMlPOLLbr/QOVE3wlboBaPdu1wbrpm2nPV5tu5Vu2d4kMsMtyFEyCzwoeKYFTEJ9
9NF81vWCGycNWTKPMHUAR1+tuRFPYoU4Wn0hqTPr1MHieppnC0MOJhKhjHrp72Og
kba8YR9l+wMYEPyO0IJcIVaWzrdSymscYINaryCsghLwc+lcNcSSCuDXTgR8Szvu
9SuOgc14RNyQrNnzaScARzdRXfwDeZga/YqmuRFGsqYy3zwnzKnTl8ARbWYG2fME
qqyjtojfF+a1gy0zNRBIP7R8WcFSzRUq0Q9Mk99YvciHv4eyWQTcLFUUkKRcc2ad
K1EDbz8TX/d+/IKe0aBda1up+vilzBgWCUhpZcOMGemJRVc2di0CdWf7//7OHUAw
sZpkE3e5Yz5i40EqABX3ispFQBi5Tss+/HKar5Eh49/MwfSKPiCKBGPQF2LZyBhC
LRSZYqkmU3uhpIMZq+10jxKw+QNwUNJJ51NUZNKKvxFLnUszAzEPnaBEvKtIGGOR
JwDsmEkk6VD36l2xQiPhf6Q8XMgYXqCx8BghE2BWI3jSBWx7SY/N2fVbKerBisA2
fbt4BpX2cXJO08wvYTvSgOVpvX+Zy17RDCBVpohMwgkmWS9y+zjbLCk1d0fEL49D
eL725TbnVzG4Bulv5ltUWt+4lkUE28swxSPHcz1neSuCMAei39qFqCaR/9n9GpCq
KmOdaAGAwcU8XjxTyuvO+dhTHoVwGfcqg4gheXUxIy1PBLFk3yOZ/MNZLaC7ge8P
Bfji8y404RJE6aUvYjpoPSbfpi/ztqQ9TKH4tC9bMDlu19n5pHRVQi3qAuWGb2zx
e5zcw0Xg4rPzUi6okD42ywYJ8Ivc5SQlSa3TjVHiq6QV+Ri6Qd++LANIDvIQV3C8
lT4HDBrbY+RycIWD3MYUwfuqjYLiF5aCspdSBMJfTiJ4O4jtGSN/ufHoelUI8eOp
DBNzN6NaDjTFqrtdg9IEMXpnrDfcwZ8XIHl73h/o/xgjzZMfn5QxubprOVf6Q6we
MYTrtepEbIsPGctdcJEmvpxii9Sht2yAVMxH2OsvgTo4KKP6r7GQVGfcLS7zIvmo
B1tepik3/9fXet+c9bWjQkFPNe5x88QNQ/uAf1kV2szlatCmuto5KI0Rdl3Qn6QS
eUJiVI+e0WeOAvgPRV2sH94nXb5B+0Uv41tGV2xCvV64/4QoiFV4rtgguKrO9tqL
qYGoAMxN8gl1mFD/F+9M9JCLEL1nyAsvfoJoJJwKS9ckzbSbWiSRyUadg9sca7cT
Ks9q9O2xYKws9tsQrkWLk7h2xWvEJFDVYaDpl3lAhnxN0nLBA5LH8nSn54ZKAcL1
8QiYa85wUpSKPPBy6MtQBci9gR45UvoK0eoEvmctC00aUlTceQ/A1O9kUf6BAxkM
UuiH52OWk8cbRCN35Yqs30dwcC2PSe9oOF8oWUlJCf7Mrp8LIebDz6WQnAPU+bTw
BwIqlWJLDCHRAaO+frg3gMDSWhBgqklo/rQpJ1Hk2a66jY4Rg9NxA2q4vOcmLxLV
LmN1G7Ba8+0zaDUmSxWiIe2Y8kGxmXglt9cM0Yhs0cfOUc6QrU5b5wMKQ776hMiT
Tjdfetxywv+MRinwrxTgZ0XwMHeC46Qbt1BS4TR/aU66vyZOoG2hPsPRgsSVp0en
aWLEKAncaPp/btxYsXQGLvX1Su4J5gVDLVhONqkwFRXTALZDzhH9iaNOgTZOOpB1
4cNcom5p0NN6mYLc7vqIrYkrO8iZtWX7/gZZBVzem19MBvDzZSMazJtggJTAq0Wk
Zpft7O16iOJE39QarpkvysDB5K0Le0rP8tbgzC9BtG/pUGFOBazvKn3kQ866tq/7
nlQi64FJdATG4AKj5StctrsZlmqL/+2oJafPUaUNfLSdeUnatuoEjjcAA+CJKH1H
Wr8eH7w8y4ogzIP4JqCo4szY3VjI6qnLJcOJbVm58rgfqDmD6nCHiFczcADCcYak
n93Rev8Ce8ZFr81uszvJlUdyyKbW10ucZko0LCxEzEixQQbuDtcPgfJIu/mGN0VX
KYiKMlA/Mq8N6q6KMLv3niMFbzQZSaZU01A8JTkvVSUc3qc+Da5Gru2jnBuqAOju
hdkktBF0rMyj8CR6LuZ6IaCmBiJdg20AgnDWLm9q4iYGXeN92YxrMxqzMBAetT05
L+mqC5vLAorNFbaIKIxfLx1gSN8lZLiQMu+g6Rxf/ZyfyeePhO8IYlFeCJWMKife
VuKVj5GwbxMQNgQofYJyGYXdjNOAtHt1kJxBmDKcst920pwwr1DHPctyEHgNbYzH
Qs8q8eaMVSq1hQeW3hrZ1bAqoiZswYKGtMUxDI0hFjeKn1laUXTzwzerrwBW7E1a
frhxGBfiPZvB98sPTeBYkLprIpGAryV6yvCryI/NwQPH1oGjHq7T7KK0ftsqek3a
Nsb/MeYtg64A+tE1mdxFLYHfKqXNQeLr3TlrGN2tRmzHfonIoIelv2H76uudW9iw
GcILKs715tvL2wUm3OAiK7y2tEx2Odo4CPXnMiXOVFJyOHFJoQ0uRjGlYmrjaN1C
czzaImdmkruO4ZENw7IKhHgtqgjwnYC8VbjtdZFDZUJOAi62XrEoel+pW3usx9YA
jtaUATpExkG9ioPPaPhEsvH23RlddSm/x1JGN3FoxZP0yI+zgk9byCaCeb01SXJO
TvOOz4V/sTqYNz1Gyzc35FIqFatLyGitqBjaANKWDPK3pRCetxY5weGJuAlA6zOq
5hmJOMm8d+Kn2XFYUJ+Z4nOjkI42tFgKjl1Olt5dWl6GKjD5xWFSW2V/Z1ScEzM3
OGlC0LnSGZScmQG9BZ77T4+V8xEJiP8ZOVOEt81DW0ycI3yGGlPSPvbwNTK02rDZ
frG5TZIyjyKkwnR38y4XdT7mO4icMptL5YRAmOATyw0T4rA4U+0Spxb3F5SXG+cM
RNiRJWvJ1AQ3egmwcGADkpxhZsxx+AnRGSFenwRLCN+nT2Cy0vdMuspPQ5bIKP8r
n+Oxmf+hsoVty9MCDxaCFKUkWjMaEcaHqlLPPPBK5y/dzna8XrZ4sOo3daCwBUR4
ExiHzTrPVaVINK0mOVpayippaSvQXneTz7TNTOSMgRTsPpyZXBbuRpRK+NstNfDS
ZcoKT//Z3knMqg5SEzGQMzlhXfmLnZE/HYQuo6H82M9HyspfNjaHaOeejaYybu83
3XzFjDr4jj/Aa2zs9YA1RgYHy37p1zeMVXZgT/+kTdR5onnvihqUHPayYDdqzpzg
VcdK7IydA1xe/rnNIOlpDbR8y7ia3zm4FoMC5o3Wbsi9PNfEUrBYb4A+nwA7GXts
dQAZ+WDmnUMoTsaCRLqk+OBsFBwa6JP9WHcL2KRFGq1ziZiIn7JuY7wVTh700XOu
iV5ov/wQ5Oio1Pl8HKe9uBNodXh3qBPPhdoQbfOl10zLf8gr6REVJD6MHgxVyvDX
FQChMOQJ8ipo8SM8xoFSx9yZNg+aDw1azd2dSZ4DbJfOuVK3XF+87Uih3e337Gsl
6h5uTk4xJBzHIJW51v6SgvDnPCwn3V1JDuouglha4gFQCQGA7t1fKLuCDb4Hx0DW
J/uoIMGZn6loJPNPreRz0AAPUJ7dm3ZqaA0J8eEeyU21zHDACb7HwAqIcHEavicC
QsawMDktzoQRxJp1b1cbSRN4GU4npii1SWmc2EwnjOLFmknAVhvoDS32vrhMErkJ
Bd/ZFK01br3ejakCODW43jPKnnERrTC2YrTRFS9lpCMK2+lrVKTRvb+l49yUVr5A
3P3d083Dm50iqWNBYmd87K2itS5M26yq6Bnk2F7O6Upw64n5VGB/bMJLDqwgUBNk
j+COugH1gQRMXgIHYQIJYsE0DxwLGpvJJBSxnHV8tGLknQNInGGik7Fc2ip0SpoK
4LCGffo2McRW1JaUCP0K8Ij11/UqkLBgC910XMGFCwHtcq2ri1w22Z5wqUbWflkN
g5HrS4U271HnQAYtysYTzpp6++xlSHWRAced6u7I+GymuSjdpLdSF26VLg+swM7C
11A/dNAdzs1uA1mp+eS6LrcsavyM6q5a0m0JXXeAbYPt5gzzjzsRaX1P4SOKJ/aQ
0qell2w6X+Ah93xVpTKvYAzc0vxrbrs4wmqqoMNSl7gNGRNPgFmBnx9b7gvZE7Iq
bNHs3peUXrKhUNyU3lxUrBQWuZZt5ixlDzCFAm35ZrKqvW+X8PqsTDK8AW3cXaD6
jFenRRjbVIr9aQWacqR7ciGgorLjqMzAmQG1oco3IlXmj/cvyeNH1wQx52RNYN+0
FiwYW3+Sa7zsZd6soOTvNT2y2M6MZAYuZFTJRCsk9LbuDqpgvBuO6vPeBduaq4SF
KlOaljyiww5nJeRs3G8I1TeGGUKLXk3rbJjROAA2kBzUIKZ8NLp04+oYIm6zliTw
vRVFvra1hyRD6Av2O9Zung/jRidEBgy/PVlXwR/0ZhCF3ThnhYYJSn7ia8gzsBfv
o18UtEMzsEf9TjgRQ9/K1PVY2MaftZhwAYemKuRhgLNlJ5jVHamNiYu5LUIzaAKt
fWtHC8nrbcL1nrwXy0RmLqn0p2zoTackijV0Y7kUB/fA+9krrwH3Z7BOg5ZVZ67m
zR2HTRXNmAL5LUW1NGSvIdmrUjiPnqSX7uFLHte8hSo0gNQQwuYxTa6qiDw/jWiu
rqCNJVZMvoBczZsE7ldTVoTlvVTvImpvm4GHMxqkWCviWECiwiMlWRgzbSGdIh5A
akJBVTvm0oncK+fN0AMh3vmVw2psa1gf7PIKS+FiT3lE/aZd66rsXO07kkNorFB5
CPB0Yc9/OBh5V3WCrw4BidamUw44qPqBEY1IiXgkpJliN9cHlCsCrNvo8s+0o/d2
myxPUd/hGRisgmDqBKtR6OsKU+NmLHJp2hRk71+xLENV/ysPH7AxHibMGrXYjeAY
sp1Nc/Vb0ooMRfjXU8/4sGd2pVB5CLk2DAPTdjQM0Vif1j1mGd2r4Q7yiSn38XkU
LEJOL5evxJyVx6lKVS2hMukbcIxt1z+kzf2ss73Ta3XkRDkDj/5SL8PG8ClFSsTb
38t9ThASgKrz0VSiJaRzaCAZ+VujqCDTh43gF54a/gTzR4YUgFgpxV3LP+6s1W6Z
EhhiUNlW0T+IDjqwe7/D01KVtlfxgcvQQhanjr/iE5zswv2X2NHWMMocwgzaAoWU
J7M9peJwSimV20EgoZU1EdcXAT0PuqYer37G7FnbltD6j1KpDoIZ9uIaZg4UJAAX
Esa9/2vG5pwmRRFngyC84Eq7tez52ztW7pfuIyK7Z79HI0ony7PoGRZwTNKOwZ4D
Ksi6l0SUqZ9a5W7t1BVNkQ7+mxn3VSVhDaF2ils5mLF7NcRBGQMsEiX893/S5hSz
K+uBGw6peY3dIDHE3zlDcLKYHhyZZZNewzcBOC+a1Ko2A1xvu/FJfBSBSWoEtDCd
kCb4Ecq3ofWiUNzQhWDT+/x8hXkv0/1I2p9eDx9+ZaL3OPfSpEoJHxmzm4VVJWWc
Pp0C4RdyNIR9ZatwnnPpGLbxideCp7WFnzRBr1SK6vxJN9IoqwQzZCbfqcoZUUHD
tsIn65volNPkT8wslxYU6jFTT3IL+kbFj5F9qP4ShOcF6nwgP6AFGNSA2zXwfgZo
Koc+NBbQb5/uRZCiWCTnKjlnoC3JWMS4hpRX3Pk0RAx5DJh9HlCDdtBfrsxXqOi4
KmOs7SDixVWego8Y00O2rGEMp19qyQZXnfm9+/HmyhKI1WzDws0bNvziMckXlVED
OdSgC3A3eySpA8lV6DJfzGvVyvyC7YWI6VYT0My3o7A8mfbR526SH2VhNpWHElQF
svxGTNmETa0/kQbHBaRq74cwtzcduYUR63OIKGFMiCghjlBA3+kad6aaEFuiCZV5
VD7T5aL0c8uw+Ck4gVWQtLEoZRG6vPhlOo9mj9kLnho3sRZEizz0fgbTdeZNk6mm
4cvFBy+nDkmM7nTNLJGWFdWmIxco9AThrXzQ0GtVCbYQ4KDQ7fs60gWGox5BIju+
vsgcrsyPCFv24xDTOZr0KVMFmd5ZB8ZDM3Qi80rny1dkRp48KbqqzRh+s4rbLLS0
xckEKVx9roAcJ6doowNv07wLfm8+K4f1gP01+0DSRxLColk4u99cJC9na9A884us
NNX7kF4z+60bg1uZa2zpboGm5GGxGxzVmfjiSRW8e4v6gr3Cm2/eYlxH5aF29tX+
c/r8DZ7/Kf/gjw1TcgegpKBtoOTlvfLr/oRoa0oiKzn7YebopXaZ0X6PtWRmFMMu
alj4fNn8CPcZcrI/JgtSlD2rLRuTr0fOc8jgofmXVPjDI3pfHIezwK5e1u5a+dtQ
3cgMoLPp70oPAXWsSkjeje7rR3GppQzacbu6ohwHNfSvpnNUma8Oo0SMmo1ZanOW
t/yHowaUsPMmcw/6voVPbAUTEGulOu3U4Ck0NFEZUuVZ7q7jeoyPnvVWeQnLUPj0
AoeqxZqkNLdtLq42oh8Cf9Gb6b/P8QBw77iQVg+KfWAHwMbrdYXYao1HFmEzXe0o
rXiHoVHD9s3ag6inU8970BHSp0y2l/yymIWzTEHBSnKh0G6avejGv7EsKxut7mRK
TLM1kPyyQD5KjaF04FPt0jFVWkRKWcQO1aYvfpqbRMwjXFty2kMi6vaKzD/Ragrs
WkQDQ93OxhndV1bhJwSBQ3PDJthasiPplvKGzYQMwXEMIkI2XD//59F5M4GhQAl5
jqvnR1OHnE18mhxbRJMB5RDIMneRuzJWveoWv5zhdDhAHFmf7EUdC6LAyrS1RJgb
skzJhLsxUCJawpSoR07fJ+3vtzH8jrmvrSNzMlmbgrpayrl+mp2qTRFJOZCIESw6
ZKs/UDq8knUs6P/D8YiSNFnWtM2sZgkvayaRMz4RdraL27hCYsYyK19E2myTJ97P
DlCirazuyGRW9D5sNhJlvCQ0cUXbbRlQFfS9hx7/bNc+fnflL119p04yUTK32YT+
5RkpCdmEQDzVCndueEwLGHraQms9kKrKvCEMNCSDyX7OFXTpnqQmLLrAvxPRr0u/
/ymSL7k7pX6DW3LdV7hYlUUAU3T1ESakPPOjiTGpxAPAD8pD0o5fLHzBth2QrAAo
uBy/a5VHjRWv6cGBtL/XTECvD1kdhBc5zMRL04rmuxlM9Lv8IxZK1wC0gw2LINht
dD8FrAoElbcQvSaN1l4Dqsbg60kExFaHzqsdo5KbCwAU5hKbkFd6aYHmliETiPvl
GLhIuJFShznuPyujqnxIY6gRq6aNcepoOpazJP2Gkd/pLgBEXY+cVtiQGaxRU10E
cZIDmPL9Ndd2mIMq2tWvA6+oevHKSnG+G8p93k/Xcq1SMbXKEJrkJ/hWnn3sQbpa
3TVXIR7XiO7YZO3utSG+ENDigAGS/73XUbrv5pQO2NNK3OKzpFXMJV7nLlAEgIMr
iPrY/7QwPOSWin/M5oj47jdv+F2VG99ipM7MlRLrSQrrPXiPsEjmh3Swy+CJUA/N
CuwqoH1drfkye6AkFJKNP+9BMnsD7tZEJUVeU6KJdbLR9X6dTchhBiVgkzohruq9
soPd15fixpfbJqzDwMGFXp5U7Sx1yVfpVu6aJ2YBhdqejQ5EUfMzjEWL98+RXY33
zbmaGwt9QtNlhZccNneSYKTnpjpfUVGIbpUuNb0jcWuYFiNP0be5UEThUowB+evl
ZDS0pqQbsqp1RgZSZYKgOk2aTTy+45JOJlkiqI2ETbusR4rlzyQH8AWzel8W7HcP
3RRqBpCc52gJRlYeI0s3ijqvlwf3fJ5DG3I73DD1t/2GOF0cT462xbr9EQfm/1oN
AJJojSMLwVubW1ypSkhtMHfMtVFu8zboI81AfItbQEYmIwh4d/cxMzVKV2FO8fxz
F3Q5qTT21Tcfgo7JtR+8e+FhG8KHVh++DTkKdI2FbIWqBNHZyAVlK0UBLLwivQuS
DMqsfTAQgi3uFBReaF9lWfS3Dt1IT4dFCspm5D7JcsAB6nol41SHW+5txkCJAmq3
5cOm9ZrvO3OpkEEZj8BlDFPMejFfdpQEZwm19twluPb28l6WO5hIwL065JtRZtR7
4UXiU8tisW9G7WmUI6VO4Dx6XaUNVVfwqWeZaMK2FIsKNqFtx5imrUhtdOQgXjSH
mg1fN/qJ5n0dpDu7OEBekJygqgvCme+p77hGKQxODu9OKV9nFxiW9w9efvbaeMxh
lmXaQfCXASIym6kBGKgpdATr9FIK7uJPzFUpA0vawHx82mgav5AZ1/rdE+eE+8A/
9JDQpacQ60gkgqWrQmQir2Bp+lPrr32XWvOCLtDiQnoZlhcYHhEIxPdUGJZimUa8
97oCdwu0vj8I4x+Qc0ikXfZo3k+8ANygP2JhQ+8pzRHx6HJSILyALLBb4hqMq8Ok
UktW5VbDLPknfBmpw0+Ld/LmfRfRatXIKgApWBavuDFs6Ui0mDVuaDO78JxUiLF3
/k8Q3DGBSwLfklkdIg5A8TzX0L3I+sogvxvOMQVGw72AVJvx241F/w18UhEhMlI+
lzgUHP3CxyaJDzTRdUGZJ1n89dMwOYL7/5HGRpPh/17uH22Xt1z9T5QTGGaJnq62
G+Zs9ni090lUr0mRnqCfj6/ETbitycdhD0ZoqW/Km7auujEdYElTVroHeCDMMhmn
uFNvbEx4T3bREsmjC4TKoXhEYsZUfhNKsbOhD6E8G9RUFPq7M8DA2qS5bOpIfWyk
WxkKqmpUSW1t1ri2aGbs++JmB6W/SgyuNuBbYU0ufj3YOosQQLAxyxUNUIfPR3Ks
YY6tmzGQIJr1t3eferyv2vbjxZ1YpEGs5c6TDji5cI5/MKHOxzmMUEQwkXDfHcZo
DUQXFMuoNwkDQwjA7qpD4/ULyXKXYkkj7LaHL62RGfkv2Xn8P6vkNPBlogqotK/P
TDBGKTeXgj6IXi+Vc+SOh0NKvN9sgtQPb6Ova7Y/mvwIR1+GZgwSG20QAHef8MJl
gMC2pTFyToKFJJyAmeW3FIujtxvNHfNXenRMd73zHBR3GaCkpLC4sFI5e8P6XrH3
QSA3+RLAlaEUtOosS+pXOD/35bbUA7nBZM+UQ7t9OCvC3dmWQpkhnAnkM/Gf98eb
bqG/XnFfqLx2pyktIyPLb+VZAiLTXvJhLdgEhQ/OtH40jmd1sMnc/bFojf3JHxLu
4FDNN04EpDCmavcoobt/GywT5ZnoXJ6dtNPZ8vVuvP/4/9G3YkiYtcoL+WFvhux1
ZLUxcCEUzAwe7GgO4yCxGzZBKWv79dqxk4yGFbHuRf7B0qvmEXMxAAOiqoJUyosi
P3FdHwxP8YKCRSCCswOlY/xoKQPUkP1sJS7BsZi/hXtwEArZgK7OMkWz6RGrYZux
LZOZgsXdnp6m7Dhe+diwVdRSVtVPQAV9aix8/FyxlLNu+AEFg4CoEQeil3MirnQ0
H32NRyXWRiFSlsNmLiKKLLPXqEtGXhph24wAYG1kVLnRzQVpD55EsObQmxAI3POz
Zaizm08OwxgwDCYNrMqFEszQOZpX3EFFwbJxe+Rnbo8NegQnIbsz8hgcDlhcJENg
Lvf/1LsJNf75mawGbVQKVVvTCZ5VyvtCE6Q8ABhJIHYJqMX9TpnyVkp7JKHg7MGk
DBsKxjDe0r6PrEBjwj2a+D8Ha6OgSWFQysIQ74JTXXxoQ/8Z4i4sE4bOxEINU2jX
bSTs2s9sY8Afcxa/oAwbcA4UQ5UQ4VI0phzpozqxe8CjRKZsOW/NM5iERHWRabNx
Ncl9l8zH2XxNW5cqSoQrrryDHJICtA4t/pNZ1MlQcPiKGChZ4hB93qnCKBXIUq44
/DzQb6NjJw3gdOkS2hWTnKD97pAgmIz8GANemwfzYTAyTK7c4nnYAp8+iVLjsxZq
J1Jj1+6xbodLG+OYj/z6xMeaYgrxdjJUw8IhtDMx+McS4+pXYB6B2hDHG4GE984a
zJU6QdW6cHH+6UqyabXYJXAeULYjiBXc/MnsEux30+VIUU8IU+vdKi2cT2LIuXKs
DoG/jJb9CLvhOPoL2VOr6pSosCbcVpNhOk+DnsOaP49dOtxZrnaCYJtIf1uWVMqv
b8je8dh4AOWJ6UK0BkTF9SE9uQ8rSZW8MLMPUvZaoBgWjeflv3WQAdwPxAZiyIAN
JjAWo7p5UvXwRE6cITHIkfeLb1ausv/bTsAmWtuAWjbwxiqiJsKX71dz7CyzyL8H
SvpdATW0MmenEZNGqkBJyAOFgjTUzvmaufA5b7PzuwlVjfEjSZ5HZW46+h1Z+CRi
lfG9Dc0oQ3NxQ3uJ4VNsrC3oo5OPq0+otrVR8RkcHowjRntrIDB1SBT57vQVo9wH
FRdLBB+93MMewYY42il7Sx3Vb/QLBLBeZp8AzKEGDTfzwrzEuw2wAvPZzzGFYIsv
gZta2hR8N1uKVMRjM9T+wgtfV1124Msy9KtFM21pdEHUGTL351W3KgvTZbY7C5cS
zjvRcwSKvFv/+3zENkF/buVSzUiahtxVgdruzpyP5OgBJOxJAz0DsYjvki7l3kRG
ENKvD4DVr49jPPcuQo+7Tb493Ues1GcgGsm1/qKbVCHgo/CU3r4wRVoEMB1d+sM7
c8c6Pe+SOTs8FBeE8UM+96L3m5fRJgjTsqbZfRz/RDHK1jX4igVfXQHwZQZE55Wi
MQ9msyaiPqVDeHiW4Do1Ih15wfaBnJe9+Eh24CN5XGhMXxk17F29k6SgE2Ghovo+
bOiwiD9sumrtQuDB+nzIlCvG1IDNYnoHGchOakG6tcu6QpXQOx6hWxqPBVxKyImD
Wq6wREDXNMf+z38prQgLCZH1SQCYasYlyby/msP0uRYEc0slyG6Pek4vRLQNdM6m
PAoO6DY114n4CBiJR+DAMThbYyiQfEi+SKh9ThH6HRxrQMqVM75DrEV0w78jIAgY
gxgDS7PPXUAy+UEK9lezWoBVjVbQ45i7jW3UTW/jIk2DiVd6DZC137h//wqc0hyi
W4z1+QyBfJ9sxuTC/05nq3EIdK+aRiWj9sSxVNr7ZTAvXlncg5IcLldeuWLmTfSm
JnVKpBkJEKAfkII6gBS7TkGhU3sIROTZ+nnsKoOFzoceciBZw0lWCubQNImcLHgg
Y1iviJxaaQdsHUiqOwBcFDGRnh2mZEWxQ4vrovcMYBhOlegKXCTa8Bl3jjmg/XI9
G0FpOtsJXfeFpJfogv0A7W5IkbJuvvXJ2RyPou9t5C2nEoLGxAUOPu+GvtnupicS
/pu0Dl/Mr9xIBW2hEL/02ea0rZ7iOyiP+GVRTuqmCuIRN4Jh9vKrR2HC64mBiYYo
elSFjkQekG8JUCU+gclQWdAi0Ya5HmHGpVCpf088sF8KDTHXBwZidyyOCf0sivga
c4CrddFC2VyY8CEUKgdMafGZoQE4LYcJneGuXrlg+v2xD/6cJxPsugICiBuE1Q1m
Xss9Z9og09+IwXQH5GlVtbzqdp9drlXNiImOYVJx9CYGCEnAii9HEux7mGWsvCIY
lv+rr5yi7n1wc/ivqU+3Gbqd1b7MrPrAsvE8AUjq0NV0hDz5oTlcmtFj5efKKO/Z
0n584LMEto+e28fQFDJdBfDyFRelQUGMjLOzODeqbQj6vZT9SU6oy3Ix38ed8Wya
WRE80tUf1g6FfEfy5B5uXxAzcGNTTtNX6fcr7hBR9ddaCPKiVkl+02Tcv/qQN3U2
CwTOJOXfRbSpMnRuFPtyRfi6JDVIGUY2rfA0pu0HHnXxGM205DD7WoPTSk4AJVmV
/FVmgFIRItBXROLApWQECB3LKmqoXWYILW45XNbxMj9NQPxWShhQr5mw8NCGd+77
ALyxhppyuNSajPjOibkNEUjqM7PcxbpbRMsWc2Stw6WQ7zZknSRZ7tTRVDuOqJbC
SPU4acvlxAZ/bhP7K+jCzrVdNtwJh8Vlaz0CQMG95lWHse2IuJLuA+rDjPJfF2l4
yfaBlTx0/1Qi/+1HqUDWWTWy7Epf+ohxxLMg96tDGOcUF03c+Estpq9Qd4KRlUio
DzSYpF+bf8yH9LYFqz+hR2/W4jrrObZqsS12joyL6vxJverK2ZMq3B3OdhpyJC1n
lUhME4dGCxT3WKv/YFMlYqADWXZKHSwLIpXsHFNxQ83jR8mOCcvBQHmt2NFCMJhZ
8lTxu3zHApDslipO618II5qm2OAgrZ55KFfFiM7VadQm0mJOwrynluRwWwmXPBFW
V/NsMhvN0jSI99GiLCWh8FpjCqPfXz927HS0+l2kMRJkm3UMDAxKdvKaIf2OU/Zz
e8F0V/FtaJKoWeeGxiw1xnKfUZENoVxw1LKkgupQhgczp8h9W+lghJtMhrhThMsr
ebkoommibnFndIa8p+3YVVD4fAi6uJA6MFXeHggyGNPgWe+eDG1ZbxNaf8t0fh6I
x3P1YkeY+U3niiCdSj8NNy+lNaEG3y2CWcIPALsBrzD8nWbIt9rM0qZoWavZ+Y+I
vLD8myAfNmp3AZs1yqSlskQNAVipv9iBgy8jLOs8gGxhaWrknwWLrc4S9ZT7v09k
1P7WBSePXXCxshJ0SYDZmPoTYhMKkJOw8VLuAa2fP4IINoDke/rABauJSKEg233A
v+f8XGHgSn1iH8BplXMedPldjT8xIqWgYGaAn5Z+rWcV32+zrMQ5ihCSWlpzOFrL
jbD2yNuTnlMA3f5GId6ZOPk9qmwjP5zj1mLci0AbNJlNkFCSd0Na4/sjUD4hrIuC
7WxY+7OxvAnHdyQvE2mBW82HqF8T5AqNz6RMCyUz7tVrZ+UPN0mCOqO6i2rhyPR0
k2NNnoW5tJTUdO55HLbpO6nsbsUhHeLyFRmXIZ3iRQOxsgAqXumTMM7I+gYXEgV2
MiGp5j2UUk+IsO5hyGGChyQ4BZUlWstrY4m6VVGQMVBGcjLQmZTeR3Ztd2HjVofA
aXmgn9JunCnVDhF1vLsWekcAw6cmxIEZ/180QNu9JLs2MNYdShiS9RiSMdw0xD84
hlDCxcKE/KOSnMbfvUWkQbfzsU10Q/hQuYKT8MIYKFE/MhiXiPxnKegZUmRV57l5
a9RWYP8AObDBstWRzL7/2e3/p6K014SfuLbmIIv5PemER7ghUeT4LlPBqBYHOJ2s
rzmskM1dqoSdqd1JXxZ58vzWwuxbCALbc5ktlgapJglu/OXiz2EvLFebZXbSpq8e
unh6yREJYop5MR4hVAzJiNuDSz1z6bdc7qoQlqZWnHKqdzeGRQ+LLO4wnqkNOofa
RDseAWogxyoSrScEIdI/TA6109VkBPtRhS0eA8As1UHIVEQC9/e+kpn5ibTuX6GS
5FJ6C44/RMN7sYg4mhiTW+aVgwrKAtVV7RAgHJ29Yo87tGd86ef2CmukE9lKlskB
MoKUSgkQk9u5gqxB7/htjc0DSPhA5zcjxaVjl0kRdCVUUz5GqtPmkJ0hX2Ikg36/
8V0Su2LeXec4kKOkR6f5Iv2TvSXtGBaUAAqr6nHsxG8EaFGqYVtB7Mt0/wteFbm9
brlIjLsYaaOQsBLRon5G6fhfo9f5AzumWzoWypoCpq8sHVF/4312hVVzh1R8mGwH
eQBaHh/D62J0y3atbk1FtcPogjhi3kmgXC1jwqQjfJyZ5BnX4jygqbKgE4/Ayean
VcRaAUiJrcQvwMEE2L9Y3JIaij0yCwedqivg0Iazi5tyhtCwPDXLnDh96FuWEbJE
3oCCZ05hsH1pz1Dlw7baA8uDq9BftxJQzIvkJxUZt87Cch7ww0SfScSfxfBzZSOP
OF7Gh9dBNPzvk6v7TVl1q/x63YGBtp7aRL9jWrGHbtXr0wVekKNG5IPvwQufcuF3
rbvb36Fk+hbzEpetyYBLMLnxWGOMCRA6GJzjdKmBzGDX/044+ng9F0J8XbN7+ewb
8gW6Td0j1rnb8SxlEbg22WgCeqLwFEprNMT8wStYLZx8+4svaMhl4Pat+jLYaJV3
ZVF5Na12ZT5SYzAIxIQ3kyDhaP26JlqHO2GH5GsiRBTeN93UYNFDkgoPTQ25+Nuv
UAfRAKsW2yO3bS11f+QZyN40tOTbXwPfoXhA3ViGLd57Cg9RYXlZ6JYKixLEG2qL
1pxg9AGi8YBbkvsUymKVwEN2olThYQp5TrxF1czHR0qMb0JFCvs0kLGlqU3jrNUR
6lioU+xihGbh7lRZXDmGkJFa3R11GqLtwmiTIRCazmgbZbhkdNis/1aMXuonRf4+
s8XgcKjtHXSf1n3kiie5p+nvSgpPC65vdygYUslXlfsC7SeKcjmGjXsgbbgnoLMS
cAVzH7P1r0lTMC7MvE/musjobORRh2dStlPpNcyjp/TUEIJz0jbvlXotq28AG2yn
FMsvmHmIECJqEszmdKf/mnqCCkFrLqCrAVfaWDr6UrKS+vx5yaa8imoFrfsxVB3B
JIbmzvB1DHoOj8xuX3YTS8VyKYUlozDwIraC3a8Qx/vVY2ZTz1rzOUPE6AseDd/M
mbD7g2jY06kjOuyML39r8LdKoshHNrlQvT6HBygWPoJEToiq/yZTISs/+OOqA2nW
ldGrLuHB/FpjidEUML5OvS+STk57GGPZ7vCQTz670g7jXqRrbBzxAfQhWMhVIiG3
r8Z7iMPJb2uudHltSGiWhhZtKq1bCx61eYNT8NtSmoBFget/HGAtgQWDUpf1f8+1
a2+DIqZh0bvX1y42qbCBdUAFysO7JJ81FceVOKJkViCp+Lw/5lPPRabhIRu5sh81
3ukFrsa00UmU0G7dHjBJQ4D+AFBL5OVMgt5iJ1H1PNZRX359FSPqXMWVMLIXlDAb
cfXmijayaMX4ssoZyxG/Lgl3+jrj7frSn93BUMH+Vt3Sog6D3xM/S5bncxTlcdxX
jJvBxu+ovGPsq0xMjLUGO5y9jrWZD5JnhuXPS/T8OPrY+INxYzJCwZuTMFduOyoR
pDoVzx+NermvXGIPSUQ7ZG431Lv52NNKUNBWGBP43YvzjR0jgPeR+dX+qFReCML4
6q4OXwBjuMHKZEJkMXmcviKzdi3FNT9DnpxnFAVLEExMqzg+BrrZuJotUaLEiVS6
hK0pc9Gl7W5dun64n9tuc1lLs9QUXjV1OFQ+4lCaHWqRbIrA2DgAVlXCZmwLOFxH
UraVuLKWZ7bW04ASyCNd6v5HqzFxrMRgqJbP+XxyPevOx9FKcMGvU9QaSlWDFewv
GU7ZeEmKdV/0dV2KhSsuaveUji7MjXWAS54AdM3ANTTrH23QhqXlMCriwDhIoYIZ
v4Ux6FiWVOXye6PolELtc74G/r0HBUGhgIxHyZaBiXa7PShSZUfbREQvQoEgwVeV
j7WPc5n3ZrJS7xqemo+4DqxJ9tRmKZBpl/BAPBKbl6r+t5d98u839edAoAQo2rO0
MBaqSRSXfxBxjQ7cCx8AuKtUipzgOqje5c4E2783HQ9rM14zV+QLgu8I2jox27JA
+K+WlOGAdlmumFOynm9LRxOeFeFsDA+/iZJLX7uCsTKpyafYrYr2QM2KJFkBgAGr
vXD/pP/z1hmxJbOJaMze6Vu8cMhyyc5/WysTGCufqOp/l80XAWS9VqaM7bLIPUev
WJ6gYeXBCx8h1x4cusmchEX/GR4TqAYz99KGmKuLKbt5ie1bzk3xgntWdtoD5t/1
mztTAutwO9o8p1yeOhqvjvLmhkAVu3LGFj6vbr3iDBw4eSyZYhUSH4VDilQGl/Yl
vZMQrRvwtHqyxt3iEfC+Eqz2OOYzjyFsWwuRi6Hvl1Eh86kNn471oiVysE3vGxJF
7skqOwC49qheDrfV6i2Byfjb+kxrMP3BELLGKi2F340zhjw8bymHxlCxIitLAUqe
Mhxy7s/em7HWS+Qdqs6HCpO6JLC7Fs8Nm/F0i4wfkO0TLFYxsEi6oIlREJxSwS4W
8wv2fWkQNAkVMkW7mhAvJ6olvxyfU/YWubbhyZnkREfikNxZSnF/VsDgMa1e3tyb
WuQFmFHhX8qAyL4Jj3HGQEAPcxmymWU8xDWP6irhs7QtiJ8h8tzPs7W20Llr91XN
WBYwK8jAvHQPmIVJ22dublbv5ZEARNnr1IsPGc5bwG/IqcRkyApeN8YyhLGW/1V2
rWn8FbWMbpMCYr35QNUKd4LOC4vyGxcBJFziCZeweI77IFAnk0D5Rr49fOi2KZ1Y
8BKYQBejrg5rIJ48R2GZuvuWVOatadySrBLOiOj8QHwbsurRkmqu+GqgVpJBakZK
Tn2HuOvIfAU8wYdJ6ZVUgR4ZNwMnLl67CBSc13/kPw65csR3//m7bCPGeqCFcKyK
x2GDSG0ilU81n5LPZU1PKxNaINyklLSoRevxa8Grse2ZRlQoS0wJuPwyXt/XjyBz
tLjzBIo1zHELVm1DJWx2IMvGasQVFdBVa0JdovIsmhswhrEzsS+pHsgPy1mTQ5Vf
D5otiEgjmuue9ENo7kMRq70crhQ1Fw1Z+KJoenjJOmxm1GhVcSOPHvbkwh83GiTP
6Er3QCXAQtApN3pvNT5oiKEaeMVn90wGDHnI1pBw3MoAzq7Xwv9SCpBC78cLhMm/
0AnWYRMO3D9C5/sgNIOiyiWaJkEUU2F/6wDXhmkJagyIxSDuT5pWyDQ1sinUUm6f
ApvqVHTYt6kaVZIuPDRDEKOFXRqTkVkrbc7ntduagTRlTOjavwGRXAoZsu6NZf+u
gDzDFL2SHei1VaBp7yxXS5ERsjCzL2KEjB+7TobP4gl52jPLUK7fYDpxxwYb513c
qZkMWbE5CwB1m2uFZrnSkU8TIr5NtqjJ9vcJHPZfpP83z4SwgA9TNglL9VW+mL6t
AobrPztK/38mouIDovawLcZyEcTUEwHpHFuNDWWp5c0LBCMndxxakFxq8pdE0iwk
2ogGkzd8xNbjanuKojYahz4U5HyoWNzkDVdSPtMzHY4szsfFQfB85bKJBQxcZalf
UxWH0SJ6skhO8PLc9c+cuj5SMW8M5rCBFyK0/wQ7qo2pep/zxnrdqXSSpee+uZmb
oXeB66mg3j2/mRP79UJK2D+Sorw2lIo4M6b2d7GEuyJEvXqmiA+OuB9XG83eQ+R6
Y4YTnx/KZHyneiXR1JNv8h7p258J5Z+x6g40GpaPs5lRmzN4w49H9PzqCUJ3Pqaj
zSEfS7uVul9d0KzKbQyANlbWFycGO2L/HfBsm5JVBrJpIanQGuZTDlVILciKnhQN
l2qIJZmDH1P441tlvJ0i4/V+ybgIPqBCNQYWnwiZfMGXb2akaU887y5qt7WH9pTG
UWRY/pXM2c8VFapPXC5mhvCtt1EsWlFzzpwc/EF56AZMrH/ESA2j4CBKdYqrreoz
Wgx4UduCF166rs5sZxVEv95BEqLaCPzQcWdhV/3yG0ixhYs8eVAuvthPEttKEX+4
zyq6I2fplDgWcioKqvekBNXjYRv6p6RWIxR/xnr51zerxjGsxdi2vfdbs4hEWU2C
PNl4C83Dan7eAe9wRKAhVCgWSxiPjJs8U0fvg+tR1TUQz71Jdw+GnOsXojPw7W+M
NTnRGbH5dw1BkqLytUnjh9H96bCHRroRNPM6zJV/BZbp+beu0O7E28CPOcpc3vA/
7g2l8dk23wGQ8l9UhKjGkviQcMFCLhEfC2oI0afVTxsFtZStDr6nIwASCqxQgV0z
kPeDWvyQqrfBDEnkurMFgOnaxpr5jluQXlBmMtzThSsEECujuNf3sZNhP0Qa+9nK
lBKuvLtxUUWVos1XFBTjmRWuAT0eOIOD40U5+K5CEUjNXpwLDv7hQEphwuQx3f5G
T+G145XsbwaDddi0jXEiBMvyh3ty9geg3yahP3nGZXirII2N1MHQsrSzRtICIaUK
g2qYBEd4utWxnApFyIJzoUd35yyUmIt9cCXDIGio91K3CsvbbpC0k5zw8mnmKLBj
rzdNr8PuewlCDYgEQmEK89Xj0u5SJdpc+V/IuTcSzJXusVY0CFyFdgUwmTd9wjOd
bMVpjV1GNQ6ClmRRPYM/MFx6mXo58+1ypO5jVP10GmzR2kVbNZY4kL0Ad1FYHu44
8leZrB/loVGpwLQgDwn67VzyOfv8l5FekoPLE2FV4MPsIbd37+kPeEYX62cWvlEP
d4RCvOfP7dK1Y9SP+ioxxRlAO7JIJblwIJjxfVeB42xz6EIhn5TTT7O/CT1qZAMM
IALiPRKE/OJOUWrksvhS/v5kZnj2mFeQluKrlXCoIGv3LQgzJHxJp4q98jD8pQFo
fou5fRPNjBjRBXthAQiPjEy3wbMdlG3SgDqhB1Hou4QxcCwWYvmvvz7+kw5CfbWH
I8+AuyuFB/p5aCVyOvprD8Z7e3rwbUJwWAykRPbxula5GmBgghxIkQjcioOIHuZd
jHwIOS8q0SApX3HRqxSKwWu9beUNMZmXh1nU+IRaZU5HOu/1VW9fmGZbRzx9efhp
Li35X6iwDcXa9yuHABJ0gUk6IxzdU77qFLI6AYfi0CRIp3lAfUqX53ffA6jZDaAl
Jw+mwxrfHaimzvZp1rkcm3n1Dz+oFvTvW17DWX/KhO/Shh3YVof3X8RJnmXjHIlW
nyCZWPmzILf1JGYFJVQNXR1S7jpaJ8170a2MH/7KUE9+rAcbuYuNewcwx0bhB9D9
ZVeRlatYegWvs1O1W6PndY1SBsaebnB54q/UVPo2EIyroxeFj7/5+61c/kXlW5hY
mKBFfEJiMTOVN3G2dKaCiLkbQQLH896fhiR7BaGkw4aRt+7dvS3fS9YQZIQ3TzBX
thyyT1bUPooMfYSvJIaxNrtqm6fHp41Pq/vAU3terWKRcPzioNnbv0B9HqtaEsfH
xBkEP3Abr3J+bzWaHrkBqio93gUiGGUFryR1cELq3XkG+ZBIMAJVcfQqhQYd25dg
+LG2YFF4BmvsnYK3wduIlOO90VRAyK3qqHSDJBkJg6FfgfD927k6yfiYZIUMym9w
c4pLSVYZSjH2oDEg9rRT3816FxdVQSqKJ1Z70IdoEAD/VywTVMKAeQ6+49bW5SOX
8v32KZfAXBXtJto9M02QFam4IafHoJ+2saPQp6o2DHkEaXT9QKpqyNBWy9Zej37s
oithJjMTNBevCjW7KRPJVcDAT3i0xqLHpqk1Uf0/n2jKx3RkNaN5XDp8z+OUNm+4
8rsAV2cIpZwxbGJec1FT0lkFvVYpl/xa8f0MN3QtQWswIP1V9P55OUXnxpIBTQAl
2gsHgdaTayMppZhNHh3EFJs9dk3icGgQnoe8vYevgvU9eiTB8buFjgEIUlOqRpmy
b5K2teazK49RVV1U1Xzph6IV7Rf7gSZfNfpVSn6KdKp0E842zgizoY8g8slCXP0Q
/LYvmHChYaBC9YvrgFY0B43atxPXPxfAALYr/w/b5AWrA9y8g0n2TnyczRse2cDq
DjgKco0Es2ecmIxUxQ3ccVWc/fpwPwp/a9EFjD+2qLKV5CdfyXNJMdRbF7vgFui3
uzQQJpznXCaTMdc0pwfCvpfciWpLV34w3JdpU64u/2OOS/ez+CH7Z03/BgEU7/Ig
SNGtqEIRpk7VSabSJ33OJ6v9Mv5IE6URkwcNuhZc0B4cRtfwBdi/OzgvKkkcZOnU
4RfyMbaufBJ//viKsgRnRyAeinU8nxvU3XHUaZu4jI2hnLJkpT42ZVbBlY3BPqzM
c5AIHMIPES3ubcMt6EBHOVlstHW0e93Z+ttOVeUWdQlRoHaFUqLwCWCg7gODmt2M
QQuaP328DRrlFtnGd6jqjM5V5KHKdRD1nTWftIgtSlkn8movTrjEWgYPnXcgG8Cx
Iyp3SdWSIclS/b9uIguxhZdsU/qmKu8jkaMtysLpeDO3ILW/FxFxAiGhgVQSNTGr
DRM6uE2tnH+gg50QDVm80+jlnPX2vvVDwSqzSKBw803mBG2unvwR8v0Nv+pHE3iW
D3h1USFLcpYbW12wf/xeRzu2XydHXxiMLP4qbp8Ax5cFo8gPPm6+ejYYxExIS2XA
SARn6CprY1tnp5u/zqYAptecyg9us9EtFoiCbhZG2NsNqpQ2VHeSfe6IKFRp4jTi
3vESE5/aso+nocrriLAULdvGWEpuw8dtUmv6X6RI3lDfPIYb3E7Wl5ZBLZPDkyxt
IZvQmNDaC3pmTlec/wHUc/7hBF9MDOWPyzDKakqdPfsPNMRRK0o6ITlo2LLVDto4
i4kwhXpvmagHYsbGz0m8rgKYd1Wu3Iri/Szg05cPePklcXZ9KfdIE1G1uSpyS7uu
Sj2ckbxaqwRJ7z9e/A9uxJ+ZcrPchaqc44BhobN4djew3D/1kLs8EsdRf0Y+5xYq
fXTcGx1w9RoefmkYH+lstbIRi163r7cTaI5sMrZSbUcvQNUo1MmQdskSXqGfFXpO
BH1RfZvgyRYKYQsDVVgxVDUqVSYSaQejpo9pHO0sKbm/RSNIn/u3mpy2CzrSpRet
R66WuSf0QO5aZUjnYnbpkzOq8oD9jPsgXfdvOMDTl4QM9T3MGI7s7+1TcQsXcVve
u8rxHiBTUUG2mDXxQJre6KbWamE2I8QUH4uTA1nvi4cOlwFIiS2VQpuqr39SBzrY
Tx4wiLwpevCDs/UpMcbtFhToiM9BeyavXAd97Gj7U7hbPOB+llLrD0xtLtxVXNSP
rnlzQLKy//Wls5ljcxl13UewQcpJfYXR8qTS2DM7Frv3aYJq61fD9xOkCGD26LNS
8GA/daKKU5/e1nFyc/Ssu+RDLAgzqwCquOo37EV9J5LHGiDOux2tnRNFDNTJugF8
igbn911XHo2HlyCNKyuC9Oqk37c7cBeyg0Kr4rWaIb2xFwBLxBwO/DU+WvhAb4o1
rAj6+XqZAckUePMb4Y0Ay3AFoqKHVp5dvrxQpBFHACSkPrwOttjeYmuki2cM6vkK
77bWJKzKDoqZ7Y9kpet1EPfjCjWS3KLbzhbKJnk1jvdlJAjTqWJnkT6kr39F781s
rRqgT1d2An8WRFtoF5/ofmKOyxRMhhcLIQ6Rtgk+HXK9stZaW0flvYPEHfP2CqE1
WhbNuAcxmCnrwAj6r9IybpjMMUSk2Kj1h9ktoW0+7mlZvYiDehkmtUK2FfdEN8Sz
CximF4WODtW/SviFnNgR6Q07BCYQM9HdwxjFWisyeF7iH3fb4LobcTl4aaPSZkpO
tDIypdL4HNe1f9YIt1FEEaOmgojUO/bbpK4a7w/8Eaq7MNAeik+Y/jzMm9v0A5O6
I6EMqUpC1qKYweh4m1TR9lGpx7rhQk5n0b+Tw4n/MRT5k/hZ+ig99BgFxd4JYKm+
QXio167RhaP249eGU3j5izgQ75FfBATonOtcCV35cqQa64nAgqx0lP8kB7V9ZR7P
lQXOybWqTsFQ48ibUVRot+6roNYqf+MNcdttTnhiZ75RCuoZ3UBq7F1hxNeBAdpY
FgcI/g/5Q8+2MsjwaRjaeBFw54m8qkW+lQ5WKxIwQXTvLzMEONPuvZGDQ+/Ubp9E
Sp5t4XBu8qY1Xq6XzDVkSk45R6B4CiJQMFDKsm2lJv2R5YLW+BdYzE4PKgP/Kt8w
QyJRJoOqaH/xZ+Rj1Z39cBHef4iG2qHng6Nk7mKtki4QIEP5zAUH2sVOR9FSS5ky
KQ4Pp0CG89+eQ2fWnGxe99LrfPc85RwG2PsLF2BqObOKzl9To06eqMNQPmoMi5OX
ece9Q2ouQZ72KcIB6ka3ZJylZHrasGlgexqNsGkdsVWUwc0DSfWrK9sZIcHu2SiO
uDTNRYSpo5GyLO7SLdcgM/i3s1dhoO7IzSRBhFtHLroROqBUiIaoWvdNufqcGNHt
U7TrQnYaqM0RV/7VQgGPrtZ+q5B+1O6PQuoTWv7jFylVu7RTapksbN2+QrYJA8jZ
55VAfWZVYwvhTlLdpdOEY4K4fI8QzI89KWy8jlm9EMbQ2IVx9NomphG6KEQ2muzN
EAJpXqWdRRPgOT4Wv73fM17aUBw+lIVU2GnSSF7atkKc3WW6aAB6yGP+M3nccMFo
PgTxlZSq1jWg6MohRcTQ9XKV3IGeloiwDFtMGRtYZ88WVEpy0Xepc8A5vCW2TPvn
4pQz1JZRi57D1E35/8RfOd/ygM3DCE53CX1SWKnY7hsbB28D9dlkox5OOE9IGGN2
L0oE3CND6X/3uDO/vSVr/3uOxQobu2laZWT39JVyFxFF9RvMtxu3SZvllMcc8LU8
+TjJmcJS3Qe7lmNXP4xzaEF8gWpRzwRgXrIEpETiiySmuKqvzCwB+PNqoYfXUc0F
lxUNeF/OYlXAu78R0yWd6Crsoqfscq5axbIshzyhXESG4DB3NDI2pc1SpS8AJrgh
u1XIU0cckKVVhXZd0ffEaOf201ZExjHuehjgZhBJCiilYpucEA/0FcE8UAaCm4Dk
MVfvaiaajahYhzyXZNXPjHimnnHSn9706g2Ely3vUTfYvuMgvYwboa/LsG73tiGm
lY1bYJ0giDH0OUEgJO5jWyNXftZsbvFWFJhY8RXswDqsGa4r8O8kHQh2AAdz19QS
S9Nr+T3QJJo1veNfXT05r4sQP+ZWDLd5x4wwRPi/BhMnk4c4vU0LUx1LzwLmMz0e
L978NaV25i8OV8MmvpBSZTiHDIOCfiB/AOZruGbYgWuNWd5TvNTFcM0Le6PMJcjW
MFHWdQ2Uupv6i/Ue9pcOcVEbQERSpbbKdLYcgHh8MeloebSr1xvhESN5tGEbZOtu
YqZm26Xwe0whvXb2vtT8pxZKb52ZeygKeUlK5kmpxteNpXrgVP4ZbyBIgydHeajd
pmHxcMUfOTDrp5vEQrwvLWDoBeXMz0k8lOWmls7ZCn8yd6gDnIJlhwDKz01z6LQN
kF/RGRGPHUNTiValkSi6OyVN4WGOvx7nWXiaubXeFwqPWp/3oAP3GTz74/+dQmrP
n0RoMaRSr75MaFtx+iYFPOT5ZCWoU0UKievjhJGEhncVIfv6faYtr93aneAZxkiO
1gdLnvyHCpl895iULntY1H3W/uandMZmbb92c4BeI8SChrQC01kwT3QZxoXPeAaX
lSpANKZVN1HULI7YoHQjZstej5IXJirAcgWByrTMlkg3bIi1KPynSXxF9rFTuYrp
ZwFyrnw5ZbA63ROfbCz2YWXGy3kWkY1LioEzzbxWjCk68ut5QQvtM03P7qHTx2zu
Y2e6xxeVw4UAdsdLODzF9rS/UhdRuujiq0jlZfujk774pAV6QOXJTj9iSNQ3ootJ
/6brOXcMOnPOQMUtWMbuT9D5fI91IOV/m+NP9Ikkk52nP3e9EvF3gvSMnLxqvHhJ
kxaXkkz1U87GOVlJy9vSsaTYK4H13hZtNtct/1yPbmvu4h/bA2CyR1BVxtA9BH2i
TMFY1HGXxS980ZzDq21l6iEEnxqxG11jImhh/haqOs5VWV03DNLWfGNl+QklFloI
5hPp6NM7z9CqIXL1QbigJdIXsJNJbu8e5411jf68d+Chk7lqMx4u3ZnDJQCpflPP
4Nhc1DsMikK4nc8a000ygN9v3ivEG/fP8uGU3tlWbctLhHDFCyZkag7RG8U/DUAi
rO1ue+w6SCMwR81Qp6WBo/4E0O3ZJZKedXVn+R2sbhjGychu90Mc+bkfaBV8uPF8
bSWurg4ILzYrq7nKaGegMTp+NGEYRzypqtpgsTunAVol2fA7WWXHTjQsNVs0y4vS
93Wj+Mj21nwAeqN+5rXkEZGrNkvf76a2CirkuMFmeqbKe4jCpl92A/7N1/GWwX4U
++RAlks9YQB2bbHXrvjrNhEuNT4FbvFUc1C+AvRWBgOtc1VTLTz44BsXVfSMUL+d
DJ8AMRHhoP0I+eUkuYABcts7NjoyYYaidIO79s4BcUV59JzDZZFrLJASGj/6VjbH
XFJ30SyIPz6Z1Dpnu4beM3zKayDS2r3jtbBjNmyTG/RDVcfQ6KWm0Jjy1bdfQR6l
0R6uJRQPSMTk5xDdusUEwNev7J8QUJoJMbRLepRqbSNxX7X8XUWuTqWjhzq3syGt
mgdBBOUIV3zFTz92D7LD3E6ulT2hWXcC37X7m3g8iHh319H2lRTYET/EsVpCKw6h
ylNjSTuE8tXoBotgL9dL6qSQuHrwbxfuAu35DJOGNgk8NGuJNwPDVqogCn1J78tC
atinw5BtzOT6MRdi3LAD2bjBl3GvNyMgXVm8QnPw6K1JurIlSEQoAAEtbmaYhw0h
bRN7u22fmTXaNIdKaIIGijHeJhaoofU+beC2OvoWhWFpbYIVIQjgNbagrk4kuHzY
J7uwN/0QdKrFomSQ4nqDCmDvh0gHlbvtwZ1zcKlNO8mTO5FMX5NrJcyYVExHygHd
PitIJynPR9x25tUgRBEisEU3hY1GZKesA4IkEiGkIt4mkkuRcwv6KvpopCX9kZWU
hN/oNJEfoYd1cqq1ooDRTbz+h6+XM0O9qgS2DpOuExaZEyms8q9Pktoy8r8EyDvx
kurPNl07ne7EzkcyJtwKpQ4X3v3o2E8i6nIijlcy/KDqZjc/kNQGBCA9qOCI3NLV
uBiAqVOvZwDmAHvlDJc/KF7Lq8M4wXtfARA+QgOwaj0wZcvqKvHjkdTZmP96sKrM
M80dvgk8/HqJ6yn0p9SX/arRvey4eHCxorZNcjdJ8NecYfZK+aymPrT/tQ/2xXga
OcvuBsEATu/FUvv8q4lqazANTWKPI+KPOJerqs++8ltIIlyL4LyMZTYgxkWdbkiM
bxX0ermKhtu7RsoyJJN+GyiGj00PaosBiOAeggOkgHfaEuvi9HFQEjhpwcxsfkAy
AxA3TE9OHRwfku6bETs8F9r0MitrhJ945v7v6gfKSVCFmc7i84vqe4rB8C8/evKb
wNWbJE0hRpfwZm2u1DVwD5kmm4LT5HTa5n5cbmFuk59oxWkk/UMwAZdvaD1r+0Fp
BUz6YzuWDiym16rxLEN1JJ8XioxRWKwaE0+FRFzStV9HSb2nh6nIbX2MhCdhwfa/
ihaeCl39FEfhvNKrUs8MhavEPLPdzQxnFOggcn44ghBbCNjZW0ue8/eL0H+9aegU
ovP+bp6FD0xEZDjE5ye7HNXZUircYOjbhsWM054oLW+M1ONu0tAGvLPHhafIYgd0
r74fblAaWXTFj6voYp1yUvo7UK8LsNsYfRBKg2JK5LNIKpOT3KNXWj2eos3nnyIv
KC7FaRPr7isy8Kw+/6plyRt30STaMLroUkg3f347aBA3GbkZlIH3TQAgVpFkAri5
Y8X70Tu4JHnjwofM2WPr2Wo27iS73TDPjoUXQ8HFs6qxVu+uJfK3i3eVlcEQqsqg
ur2iXA2117An/McwKYcJLMNbaHx2m9mkR/AwkZTZmbn13JkEjO45mGGKOXSE+Fyl
nLA2aePyDg2byxBsjlgi0q5/eDp95PCw/XdwqK9ZKQtnplLmpzQ+8WVApusisH5G
/H9ak17nThZSm3h5BvSG3+TTF59RMSxxWqeO8aDcLDhqyE/9euYYpyF1bkICDDiE
zWm0UByeBHo0L1xecnYIgCGefmJ0zDwP7oQ6CEZUjOSU3KsWnU5qfX4WAAUpbPrk
pG+4TMS0UnQk1ErGvyf+KfIhpCwoIquW6g7lEt3ljJFiZQr5MvyH8A66PxqahDhX
134pgn4vPXELWY891DyWGx5zU30qOl5ZfEgjo6fJEcsyCpax4bxkDuJoClJfSqS4
mnYesCZYmKO34w/0oeYZ4LrOb4+D42G4aS46kY5HlApZBj9SwCgyxCG9JNH/l2LX
ij66PLIR/4hTqHBihDFDQnYMPkA08D69BMNMpyEQlcepa4Ii4gdeoSZBQD15TB8u
/7/e457ZoamsjWeeKwfOxy9SgGYKkI9gTre4tnWZtD1VQRmx2ZvvC/7Wyk32OC2x
PUCA8x6JKFzcbtBS1thi1S0JdeNIUbgWfix0hexQOEw0+RYKsuhPTW7pBNqyqY8c
CPxgfBoxwKj6EjS/gGxeUy5nGIpEOWJBxPEc2G5oNFNY5GvnkG2lxpfrf3KMvqVa
IGDfqvuKcUY+VqGZIWNIFoSyZrC4LBobqq+iLXt4oNbNz//MMHugqwSVP4e4jPz1
6gSdMUn65uFtPfA/xh2rB/5uZGOn4NiPfoJulfXGrYqPLlcNYc79hf26vwgD0swl
BEE+l2+AB1spgENahjoPnGsnBUi3trnxRTofTBpAHiY5JLveFOKQs1Vc5m0vu7hI
gPl+9/58rvU9HAvXm8qJIH74D9Wmhk+8tbA8bPxOoobJljkDsSC3FKAV+INCNTuB
DM5MnDSrLYBxq4waKSvpeV5e91Bx15E/uNXfY+LcHgUD014JhLrlTs0kiMYzAmrn
fur3bI57lD2wSXsYNCNMrWrCgaytLPOIKcnNuX4ldW0EV1kBlYxLuGayB3dpjKuU
xGeIrefaZcXtz+gyB/q/Ei9zBgnZbPWNiEVFER7350Tkpp5klndqgzATL8qSZRD4
BOeX9zRYBYJOxpGaFiL/4wQDhW9cZnWZn/vNtRoSXF9sdRPtYjh8SEJj45WCo8a9
hAYZIp1HB4K+Teo48ZDF2HkGZJK+LKfFt2q60WS9gObAro9t7Wjl/3PuyHmOT8fe
Lx+QxmLJT2NCa80Ilih0z5hakADrLDSzjLPHbao+j9Avsw8+jyLb8tob8thkhvFY
qr0ttHsaSgQgbNsp0Os2Zvh2gsTXcOTMpqOQ134inhIXlMxx79/hwTDpSw+ppzTy
8oqbg3jgDyzOlSWD6tq+hBvZOiUidZByfzUd2WNUMuTiheJVBvkAKRQXwFNUhkmr
u8GjptS8tvkMREEMT+3DfBLC1ZbJCxFKWBz2pDThfVPKR6wiPPZHGLBI76a9beY+
s+mbg8Bti9SDJZChjuyh/2GZPIfsbuqwoVm0JqnG29jLfPyh7K/nBPaNWmhpCfRw
21TqIpG+4uAPZ6ey3G1d5VLW95xw0/abNXLbKW91AXFOemHlI6FRmZeLNmUTJ8Dx
1Dd7iKG1hr/ykBK9AaIYgkp0xdstQPFkNHxo+mTtYHunRHPDAY32Yr80EeHpKht+
cd8k6VYjXfYLCrP9aMHYgzSHPYIv1z+zURhOayEWidUM+QgXxeEW0UkzPk2M3wi5
+dbcSeJ1BD59vxyNrctlpUyLUlPDbFm/PuKN7jwTEuMTO8D5QHDn9qbtfFReRtRK
umXKt3cacgwpBQu7MyJbNDg76jwaCjzROp7+kDj0rF24F+07ZeR8BqsESgjyURIu
zlVczwi8aARxbDiWNuOEFtxJHjI3nsLcxaXaKg+p683DRd6pTJWlWiTESZdoVeMQ
+dmxZEO1hSf3hC6wRaMrgo0EcQx3uVqSe5eZNCKS2bczbRe7VLbuxiy+jtz84DoP
jcS692wTKr/Bpq5iJo8+47aQ/Lps2hU0VPdPH1nNtot21A6rnqtW/76Y3RTISdY4
xH+VI2IKtoNoEeBKvPc07KGBr22Q0CZFzywaiiPzQVdC+Ut+euTk69Vj8qJEYgHp
vD72cSGuDCYfC+e4aK+/h6NwjC1C7j1Ahuz3715kY+wVjNKOpehqQP/r9IYLhHgz
9cJ3aXj0bTzBvBcoPbKeQtSO/d2AJPEapz41KntCVc8rV30+x8aipe8sjTHRY30x
cei7CGd0liqpeAUhzIAgy6xeTDsfxYSvvYPSAuj3HDZIOufN4CB/a/b92MYV9QFA
xS1ZbnVbFA85yqX+WZ+TQY7NVSt1cWBKUl0ifjUJpd0H13GtX9rM/m6+ANzEklM4
HG7ScRxpl2dwFhXFZmWX1qHNjfop/Vfpe+QrEZAIxPjCbqMDC1HzOiCEzTJqcy5H
CEuhIsPaLwN8o3++EbYXlc9QWcn7oR/CedwgWNv7pqIPL3GMp4CpKPBL56+hH6XX
Fpd8CbXzBcY7Zw8TlT9i/pev1nOqBDZ9Bmc0HB3u+ALJgtmp6EZSgLIQ9Nrnjitf
d8VmSj0yUHmMGXqpBc3S+qdyiHjFYMvheoRrDJ31fdiQImkc8tEp96BGweYdzmPg
tMrodyVkcbpyBddYTqztBMJg55AyyB37uxMRCktcWeNNrqZyOS4q5MFmtNyHNlYA
i8u9attC8qIVRhnOavhsF6raqQvmGYdF7cMhx0MCPdDutnoSSiNkFFXLPBWrYOVi
ml/Uv6I6hLeQivROTs+2DUU32NEGujORoAp75qYoPeU4NBhuowI4pq929DMyIt2f
IH/eWTWvvgt4AbOETKcIMVpfiQNt9jxQ2nHr4AHV3JBBe8XabD/taVUJ0Q9Kh2E2
HorKlOr7bUHwbKZso1kBv6bp/Cb1WXp91N+app93KB4wNU6uzaWjXT3fr43yv7wV
1YDc/kxXOl/J4xkN5Kjxy1zu4J5+jnE3bIswqOc7cs2INWBAjGC4LNBZsiv4PZ9r
HkAM/U9x5UBcbPlwrnPtwuxpmXFmm1sUdsmExp4DL3EJszGnMiJ8v2OZjl8dM6VE
IF44CuocpjZCAA3rvMxojXDPS5tGg4kI5NyF1U3268Z6B9p4XyMPiR6Exx34t3Ln
B1rAjab9x62UJykKsS8nJYgFzP5xcfwryYADL9asn6bn3Y8hktoZ2Ya5foKwv34J
tBGDr17Sh7mB0zj4Vp3GZHPyD6fw62xyym8qSgLVJ8LnQCctgCbjhl8p4NFy1ii+
6/SNF/THVEuIDMxcPj4YP2EakZ1bQ5JZFQ8+zefJvgK2pXn78maO9mlZSEUDH8i5
d8XPGFM0ZIR9Vs4grwlz6TreXGso+qgAhprAVojlY0wLVYGxMLK/fHwlllGD7dho
i7XvJZko6B/7/X/coHE6EYD8EZ8wkpmBzScLBQXUFpg/mLiRQiI4/eyO4BMbbADe
2mhwwlvZnzNFtQSFQiuJp+OrG5jegGKtMKuYL1vb6Hb2/rAWFXQS8AG5lOr42mjy
pOdgZRMcvaNJAebgT/dv1IoDWNVRy1bv2H9bckRPUIbyw/A4bSYTNs/DAwu6bdFJ
8UuvKNImD9TVzJhlOSHTHd2WvkDUkPZgPrQ4S0J53iIDRFr1f66eNxRef3275eRo
t4K8X3GgofwGl3AFIo3vM/OBLl6A67vazZs7z7g0Pco5HyHTnEqF9SmNGAkpRjCJ
2ZEf6huhjPOwB0q0WMy8bX3gHCudqup7ZrnYP+QMXqqF5coR3RWS41FVNat3rdRM
jZ2astu02BSGeT4fhyNg5eFSpC6vPblCvHxxkqxWywBHyWrksSvlSPc5dTGUtheC
5nhjJJDhoFZWF5JvJslQ5LBqTapDQvzt1RMteZT1+70MzOWQLxa0BspQ7VThzR8v
jzSq70ZAdO7zTlIBvjSXA6XNRgSswnn1JkNxxFjTUZ4Wo6moJR/hw+ObQEgHpEAd
fmRJJRZvoXfCAYMMIUzebhaJIgFlb0ixkf/Pch0ayuJL7c8MXe0E8V1spg0H1TIr
vyEWD0lvIGjHTrR9cAzb1pHmMMeyUb2u/X9eLG/elp/uBu54B7q9mi3FnGNe0ypf
MTmJdkrNftiTGMC100CP0wIEIDt0mh4/1DQSNVIxdZMaMHmsITXvQv8rp1sj6tgi
DtL52vgrRwqqlvrQMzltwNnrpq3f6Us0/d0ojBFL7kBKgIFarFAlDKSkDAABiKno
9TfxybUNPUHDqcsyFpI+SjdCyNvgKqkw/UlWHyh3YduiN/Jr+BcpYjPaeXXwJfOl
FIOBl1s2ji+Mp3PVnxiUA+PEdJNb88cSIYR8pA7Pkb/AR+xsV7ieNhi7dxPeHYgz
l0xKoe9NBauc0pUIyOZHnFQZUxW/4387q6gbov5FJ3tNPewjXKgmaNOu33JNwceQ
Uy2GFmC81TO9TkYtAfzDyXs9RIP8ZnHRRo3uT01VtJv603G3MbF5owK0UDp4b6Cq
TRcl6Kj58pSm+d76eV2rRCp65egPDb93+zjSr9qqbynVG0MZRzCCdfpW3820JJLF
gkGXq/2QCAFt+alhEMFNppF60K0PVSD+ptw8QTdZ3C0VOcWm/J9stqvhOq/5cr6i
F7sh3hfi2JshIEQy3BCje6wvhA7FVr0HgyfHtOUYZlzUE/IdUoYNbjkfqarHQYB0
cSoDkWgJ7kod7Hq0LJgIk+fM45gttkc37n4R9d+jceSXFQKAOldk4YPrqL29P6+o
3i6OvZqta8lAksS8FttlfPWuhR45HtBsswlBd/AvHUCsV0Yq0Y7dS8+mnuCmiYAJ
SvZsRU0zkE5vqjUwEE5bph6zaB4GiYIohgIef+tsgvmfFk6mpBMpsN46z8bJt1+U
NVYpAHIjjMEFzu8L9LpeyVyOwzduxZhsEShnm8nWhrm8e4OmxecJBYQ4sSm82wQM
EGhGdrDTCrb4hALn1383MfebHNiDneBrDoRpaLl3L5pL1o1izEdj+igDUqcvv6Jf
ry7RkU2Itznq6KWtO6YpCScVr8ZUCTGdENaWKHJicn3o/38MZBdJ2ScR9RSjD1HP
w1ndW9/JUYDNWWsk4Bd1uVznze2Jz1Ukl7WXOhboMY5O76gl1duCMUFW5GGwYIum
GobNcZij14rHUVeOqz9RmmLrACKeFYHUm7AwECvG83nA+HrNEikDW0cg9AM5/HtH
bqZnqrk3Eja4WSq2WVxdhnzNQDoHOdvHHHA2nAN66xbAtqRBPJfKlH13eXUeM1KB
CK7m1L/d2pNQkMV6z27PpGcYiRTyBUEZtNQHjKnoyqpXr6dsDKUw8y/rzdJw01nT
SC0WkzFercEV3sLP31qVcvXd4YZ684rQ3bKsR5FTxspAK6hSJ23c4Hp9DBClOCte
8cOfooLw4Y3GcAjB49AA3wOoULiT/AL6G0eaC6nQ8uDj8JB1yeD1P0joY7D7kjRe
XyM+4JMRNlqnFYsBLMe/ThYFh6OfxB9XKMTrIezvtQT6aebebMvpryxvZjAYzxYV
k3Q61Pmv8KLGvyZqcbtGPLVOl87WAKVMt6AkQceE+NFEMOeqy1v4kp1s31D+318W
GkP0DeXAplrcG4yGjArjzLBLC44MUDzA3YplwJIVi1qNR0GxXQs03wOSJ1TN8GqT
HHQjW/tSb4ReV+66YEeiC9FI/GfEPAYd+vBkPWl/eDIUEKfXdOJwDtrLRrSlQHlm
NCi+7XvnBpXEzBLWo4TzPoKMSWt7HN+ufmMbVU2pDmvxDZegja+t3Zmcheu28hV0
bky6kcjLVP199oR+eoyLVP/boOupGHS852cAiBsf7M+9eMMMQivB94ZE/7S9c/ze
7O5jPIceQ7TsIkNWBOTA8xCMViwYV43vibf8aoXkaovY1j2fjlMljXLUwO6bk3gq
5xHoEOkudd/K0JZXRxWNsQDjnCaKeUB8R4/pBjT4IIG6pZTKsEKENZ4W/3p/i0W5
9dE//m5Ac+RQg5/L+FhBdu0QmFq9Rg6k+0N4o5iXrNhK0nPnc9PTOrVpCmGtiyGE
rrQMDYAciqqd4c5hPPDAxJGdU7aoWyY/Etc5oNtkZL7apqQU4N+xnONp/CCnY5BN
RQ/6ckCjRZisGw16t6DhrjdD6YPAv0CTlHJs149TSuWFAZK9cYH2GFJhI2szdxl/
sq1GCxO1eRgDFiHzb6xRzwLUmQRNw4DvxPPWBH9CByHVHCDVjgEJywG8kSydKJBp
Dq3I3Zw27fNeMG6y3fj6ngDdT69sE+QUS6dNkoEsOfqG7cDLpAaNlh7MSBQWbeIG
559JJUOnu2cMHzL1qrmX1GE+oyzFWlcFAmasgCx33FEDEITMgiESLWWd+amXZ3vD
ly2Fxne2PdyjGMj3QIKKxEbXnAGhRApZNNDZ+eYY00SdzUlPiozr7Ns0D+vwWejI
snwuzarjPcp1vooHeNOBqmwfxxMqfB9oOJxFz+FyPRnRxF4oszBhDgYoqzz3Jx0W
j7kajhwhZgyxB7RPku0gJDSdZy6MCCpt7TEzut3H31HePHVJwdOMMSlccTwczt+o
EpxTblDS7bGe39/UzOwFsY6NquNQB3qR4qjRNl7P/Pk5r+56I9+pSPQTLr3KCc9E
O5lBXJMn5MGaNjkbHNvQ4MCsDTim+XiBhoVPPXCsAgK6Pfp/0QAunMgj5LiCUl7f
yyYnzb2XdvozBmcJTfkvHc48ZhzD5RtDBfYsuwxMWSCZXk2oqdFgZwJqQCCP31EA
zOC0YRZ1HMQhPpd+XvJYURzt7Na8kIHPywZXFrrg/H9yUUMYREIy0H+MVSQ6dyd9
6XCdBXNSAadXBPNtduisI94hdSE3hEspNP28CeOAnegt3tmvHvLhfdHvakLfyGmr
Zm5zq81rO8otWa166F9Xc29AKkdp7EaKHTICTeSAjj3Dxt+N4yRm2Witv2LVWW0v
G5rMgbqXYcihsnfG0v8wRFS3zcJ1WAgL4Wn+t6/qTfo6HmxmNzT8+3gdEx+25GTL
Iy6V/vDKlNpqkP0/nAp9dQ6L4/2ZUWbhqpcQzjWI0yiOOqZz+tkkjeg7VOivgV2E
3oVCXk6RtclbXbvgKTWSoo1IAxHk/LjwJrdq32Tq7ucfyVg+pV9VG/PFbkCa859C
YL4TyCmEzsPBCs/uU+poVuAdzjXJVheLsTLNKHQjTOuAstOt19hCMtbbBMTZoow4
YsxecEvXch0fk8FOXwWqD/AMp05ivSP2rVM0F+r/VJf3bf/FwVmDZLb/RTUHOus4
4NHmHzN7vJKpEsDUaNMeG/I8PL+sDKcxMmNWTGrPhp/ZhxPJ8ndfAT/6MbkhxxbB
QC94DvB1fFZErCTeUFLI8kHNIfN2rYwko89sUNZO1rvQArX/G596pUlRQaVIzCeB
ddGUNOhC8hQaql4lB5aHoMRSlyZwXeqTnPwdMy5BupRPEXXLV1NXHRSFx1OdSabb
XBatuKD5fQOtRa6/0AdFL928nVCNbt0dqAFiQaKNPJmXtegeZ+HFoJJXp+en1rGC
e2fnkobYvcrTkpS3JAcx71cim4iNJVZAwSeRIhyiYdQBQmpiSQDkflQDSx82QS3z
yQurIy9+Ym7V6Ab71XGFuRMi/1q+Hvvyt0PBYtHX9Oa2qi9S3lOTmmq0AW0AdF+j
NfVjwSkq/rbGuDgmn/pYSM1C2K/IU1K9/GcV2rAL3XEa4HW/vDuUo5YS6tqrMusr
LabY3LnCULp2kRqMsSnxBdziIJ/cU6/Qrp2xs2psClTjvoglmfswiu78YoeHbXfR
CIsXFtkecCGLwjFWkmdMaffXKQTTiqLJO4v5fQUVXV3gFAZh36D+LiEi6rkxRpnt
/2z0mfSSDJ9Tu8s2jIhxJhx1pX08qUYtvEmCdsAquunDIHBmjw9KRYMIjTnuvPXw
bdExWGKUEUzMsHMCxXPpSejocMyYby8sO6K48c9fme4jgWC7kDIJJK31ydzMBjlA
8gmBu8IkMZLn1nHkwGzD9RZ+w8hpG7iXPG6RDS6xjxb9rgupPvHFoLVfd448wAx+
gYK9BV/+91R+ODYubrwnsap5y+coV1UDvkIUF9cskoFaYSno2DWiQ2gugKodJR3g
YMA5sK9+3kiPOHwDT7ElqzjFwxfdl6Vn8cy+UUeQbXpI1bIFp7nMT4wWJmIvZYwC
HeMZRWkSNKnpf+GT8wRNkPvWCCHC1JAlpzYtCmwhmRVYRgA9KFfhckfDXAVQm00e
/LtWSETIMo3Kke0fMDR4K/5NYmXPrNglIjgqhhXUoIsXb9yYdRjB+xBJHGZk9IO7
4lbLbI18THr5+8Ab1K/sc5vT3+4j3JrXiMY1xM/JjP4BRp0N2vkxv6o/unYpfPzw
+gZDdYGYMkxD9oTY3mpXgZ+Y2rJ9K1Ho+t8LCvlFFFpsHaKAKi8a0myzsp3zpM1W
2WWV2f1TQocoA1mJsftC3c5ICZdtq03UyBniDAa+csnEglemdTE67TX+E7nV5QeF
BbUzYffXkORpHyDQBQrbaXZmPERA+o+JIBGi6vMuF7SGNCb2eDn2nlRY4YBsXTbk
4khBlQjh0oMTXko9/SO0O9viuE0ZwcPCoc8zVYhnckylmRW7LgWTsN8w5VLtJrDO
buqnlwk9wWO1CP+2OuwKG+ydSnp04wXr/RRXBsmVzM4a5vr03nWCPkS/EZRXCJ+Q
YGN8DSaQUfMCvYDRKNpcbtctABDdlZxeQbDjmX0GfzTCt2vQUw1aHyQNK1cSIfxc
oygAbXZKjA/O0JXDdnxT9ej/QXMaqLg7etWDnsmuy/aT9U64Rm0RRo8lchCXd38s
IYgtzjLGZ4yed5aX8zTrl/kTa5ezloe0V7pNQqtm1dpqDRWQmez05KN+zWRWu2Ka
WXWQJgi3tjvb+3+yr53g5+ktUjfLbiCDG6hbrK2nAC0cdOyV8ZONbMUV5HqyCqpu
wm/NiTnOW7Qwu+7kQVxhjgDBkarWjoAsTjBdcg5CMTp65dskaY2E9FOoWscJ34cU
Zb9sN/mEwvmWSTHKw71t62TTkF+/cZGnsf15I3CRtqzX8g7hPdtK4vW/qmh6plv3
j0GvmN1HzuTglLvV9WXwOELSB7r8ScmDF5q6r2wYvgEBPLtdFjiN4QyV73ZsxCJR
SnoAeg/hi3eWlIvhvbCd7UJ1NMchVqpLkxqpg1AUE9FKFCmRKYdKoeNt2EOL3icX
Pc1HKTnTKQBYhOhfKcMsYywqSYZt1YA55ALbLDQT6BRd0DUW/atPXJSM+IxEr+2Z
1suwdTr/H0UUj6YUudidSVJmL1gdhwxgb906yiwZrC2lykQeEK89QEek26i5HYvN
nAgJNxFc9Xc3mw9K/Xcz6pyAHZ7rVZvqLxam02AdOmosdHatwV2m8B/BeFJs6b1L
nmis+FJQ63ZaEIC6R+RoTHIN5THXDSSH/sErPAWMlOwDYr9A2qXn+BEjm9kZ93Zd
+XlnCvNPfz7/TfF0rKYcXiE1t5aIdWvJ2Ir6E8j76kGkypo0rL8X0S31ZeHZmiNF
vLdoHBEWjXYY9nqQDKcAqkovQnT9JmgsEmKSh33f+QmBDv7LVvRVafXa9FQafgR2
+nnuqQGSysdCYPqNUAySC5/k0MOB8wAq4fY+hUBN4AvGXUqfvVfGHD55eReYqXzK
OvPYNi9DZEZkXl8dOQXBdUzQ/a8V4XIMRmOWD8N7QcN1mhEnVMaj5++GY0sMvv9u
763V7WCrW7Xeg7NCw0ZM/52zE/3/BnR6ZdCEMDsA6zk74FqbPOGd3pJIGeFn7TrA
O8Lex9Dto/agZwnc8r+zgEI0CeKpRu3jRr+cHSyIyZsplyn3sZAOCZNR8JcDD4bQ
EGvdrw8dKFVIXhWZ+IpBHJLO4T0lodc1hCpUisEzxrhDjsqUVfoRJNpbOUSgVOu5
Fbr92jEquHf3xN+CbbJiiFhtXxKntU7wYTqUnkJ7W/nswBjjTV0ROy7oH4rydqXW
+CzgZ4O+Rb33A+ur6uXrSqTaG1HQENLpDDgfvmB42Azf6y/IXFjB2gaviE9ytotx
qPKi9QHxYYT1ma/c2yP8trXhpdU+5bKKKCmC3ygpw1X3ajja1fnS5vwPR1kNOUVG
TlyggyAsrURxB8/3kGZ3oPC9+k4hThzYtwFieum19oFpRMW7MBMJXnQiBsDr38Zs
rdmpoorOURIvKvHuFffyiZlcOQojWWrV4bqulNiTGsPZ7/Cvs4q8ROTTp0Z+dMPk
2q6wR0ZCc8s7qThHNwFDZZLYOOdHh/5UgLtsAxtXXAAT3CN77Zk9QkLdeXTm5sJU
yh82jxjgTZ2bDu/pWRNxoi/HNRr4TBQzKlCkmPR3jtV85TOzDEWe26bs/0R47WiD
S1qns/A2xRqTTeKc4/yosdLwiovdADmneL6wIBA4OhwCGh0XDhBlqYYdaM83hyYZ
/y7dwy526hyBuqE5/wGEYwWkhk+390RqzYbvDkN80aLlUIITYcICpaPZ2rqfetT+
0gegYA47XTMlAznNm+p0uwb1IKrt2ic0oubph6pkPbU+9Xhxfb4h29XHAQocGnVh
nUv4tHSEOfmcGkY+Ns3oVbzh/FN+9HvxDFWph9E8Gu0abW7OGZaMKbSr7mKPHaCX
o9EIkJioy7J6PQNEzAm6uNaKJd9xQdcH+xabokDkKX+GVfPEyp0P0VdU3ycREF5q
tIg427Mogb4WXmgGJjWeOq+kuf4AAyz5it3DcjugtvsWrSOrBZgJRT5fuKgLWtTM
uCtfaYxvK+R0JIHRFvFAR4PVv/bsF1pd+K4JpwWu5WlKwPJIzzwqWVbGG/+dADMN
FTbtJEBCZhy+Zq4TxgUJcCzAFgo0QAVJw8ABLaj1LVYPvNqCkV6F5v3BeCEWHh7z
I8kcsh9z6W0CF3JZrFoFk+AaXEUX54n7l4UL3uJIg3PYOTztfqGZX/0czhJajFeu
n6Gm/JQwiF9sicrkqB7Thmp38+df0JUKkanECSl2xPrAFdqYMFiGfh4pkYK1RjUU
GfrCNHGWoqD+Vs7zzt3+LC+aWQ77CN1P3uz3C6htm6HyDiiZPZNc0T5RGtLrzOey
uJ0JLzeuohqTBBjF4dNlkajfRITtQyLoAQBAglubQYTGfcau5XAE/3x+vJjLGNDq
rwYWN1BFeKygN/n0XAygUma1aBZk+IlaT/DNSArXD5nMaCJ00R5EjeMFamzNRbhE
V/1ofnDI+t/hiXP+oCDDQT+pPoucT8ixqSmAI63s6YQcRpCpliqY/DnX0b992rIK
cAal1EZzPEVQfUkcvf4rim6yqSmio0U9bWEm1v3VESmRAfgNdBLo+FDrVepcqjhJ
1mgmFw2o8FzZftRYQjNsIaFpXpsaSiMviBHK39qGjpONFkGOp7ReqfySWvcA83yo
Hi9glO5TRfu5oLCymynT91m7b5MLwq/41foDe8wc22vsKpZ88NbtJ97lxBTtZzJv
rXQcQOrsv+EfuoNa4s6bajYm/iSmx5jqR/Hu+kK4NluTp75hjvFiHLTyikA2RyRv
8CAl49DFa8oitgzRkQLPCsndc4pYLgFeODsBWsaWjbw4xtRr+IiUwT/P/LqAmOci
IIESF4YiME5YQdzpAkHW6LV/SpzRe92jhZ+XIkT9+qFk/urMW+nOtlLJTprFAtTP
DFLYH8InEe8Gm1ngMH005/usxUDYONLl7mDlK6Y5C0kGqfuAbKnfej+7K94R/Xgs
sV+qezW4RAMYjziPQQV4QMQmFXh9tJ1aHGbXcHwMrwF4d9U0EvPtQ3G/0bK70loN
rgpsMiDOYbi3rRr65KMpcnCLYbnaqZDDFzZfT1zsPoAMmiUZUZmaY2mpJRQFOu/4
8abDln0tIrZQH8+wiFQSs7oG0wZ8dIXGv8JpB/Q/hzstzDZi2kRUiSrYMgbzYd9R
9yIOyD9iQ0+fndL95ytESabj9WeDBef+vTY1n4sH2keOIQjYN25lLBOfuzNMFQHx
3yUx/60/WAMvJVp5fbN36FNaRxNvAzs+zdmjkQipDOCYDdLyni84bwiqQEtP2LFy
5czSSTVwdMXTWzr/Jer8cm2gyHM52y9APzDChmIoAeg/C/w8qt93HfwDLdHAW4u/
uh4epSZ3eQMdJQ5wFGQ9ImMkadKSDtAB1UDNt/OkSBVklokHlWQiJX7Dxogj7Fwk
tMMwcQaziYkOOlFG9m/I5UVRHMIZe79dYQHzEDnOGElP8LtRcxRHtKvbsakrcYoP
BUlQeMmo/AJJm3OjdGhqFFgJfbRoAg0wOQN7A9W+EE4lbGSy9qaHw86KIbXHBN4Y
2G6dMVKk5QQd/djIU7gCI3+TGBtNIUp7i9SNqe2H6O0ZMvlKHluVEfnCNil0zKZ7
beDZs8I9KHKlCIx6G7quogfw+K906BgXAC3cJMQaNQrJZQ1Fh/WYSYkTsOgiOs6Z
V5q6X9NETHYA9OrrknomI/nB3gk1YEUzssQcKVPJqLHSHEDAaoWlmosReUUY1f3O
KNK6c6EEy/+hPmrCtki9Lm/VOkcUr3EvxNrtKHOjcjzSvsEB9Nr4yV24H21dYvAP
1gH0NCezfauSsqbH8EkeJ98/CNpcRXf8dpZb9WKzg7+vptTTECTnqnJzU5lidsTU
uFIQdH805b3Ztkz1qJK08NiLTT4GWFmjdLwhDDgN48i319PRSeqJt+lbPowrSAVM
BDUs+5B4Wr1ipomjCeBg9nGqs7lUKtqHDg1IME5SvZSwY/xYD7Om6bYeQQtNjde5
W4lobaHN8pxpnunwOCudg3mY01OUTCOP12C6QUMXiNt+84Y8zkhZWEs0tghr+zRA
Nq7QU5plzoS0hd49v8QEArEF45AcS1CW9kbtNlRvyRCyXgC/Z5ef0+rX+xwuhjpZ
p6r+0EJw0wWwd4sXQeFdYYJuhtilaamHmXeBvJEKyVwSNCWqbBIQgBuoHTuc4CuM
IJ5bwu+ojCzryCA9V7F4SKcBQAYb2dYhbIeBgJ+8OfUVYmSHj3sK4k+FujVG/rXi
4LpN32lJP2jlTUo9dsVVjj67GM9ZB3nQGfCkVCV2r7kGFm6WJdBYDUJqUMDwMxnm
gdMtSySGIg3DUfkOQuftRBDnR+ni+z6fXY6GH8HNCqNqgykE2HgOiHAdvHjZ1Ag1
0VmGpG5nCEso0vAcd/K5YAtVZjExfFaf+GMovj5g1e00GyYcEGyftmk7uzZbfrNB
m1FUN0fH3rAwkdpTzqSA3IJw1pltAToihjctrKpesWZTT9sMA0zXSdPDSVam3ZvF
fyZrnqVyLoL61KhS8ztcpyIAcNvaRIOtmhdhdyBPF8F3U6DcC6aJv3qgX09qb62w
IQAbHpHlWndcdOY8ZY/yjkPB3NpoMAFWaPNN0RGBUpaokZdJ70L8uWEh/4TNxZBS
C8VPX6Dymq0KvCMU8uL2qLjY2XDYKz6VJZKFelIH4nseHSh5BNB7CGFDSlxkKf2D
IUx1gVKxaUbYdKurggPeHVWgVSA/v4VsgVHD2Xr8eCmnKt+xcu+/gNRAKYLIiwIy
BMmI1BeGc5Sk6fBoMSqY5UyX3M1Ow8ObsZzC4HONM2uPe0dT3WtAF/EcGFQCD2+e
qKtmG54DvobOfEnpw86wyCKQpkM2p89PN9bEpJKT9loPCXYa3kLOphLF2eW+qh9B
GpEm9EnWPssuhiiwq+FcJh35ad0HUj2ueQ+/HDuZ0Z2UOXNEHRhscsawcsSC0See
9zcKrLdfvbWQaI9j1swVVG5F2ida5g4w2LyHRd+V7u3yXLCrk+1pknchOmb8woeF
XtOiuiV649oNAGeab2wZArkuwxTjYek445gRPCCkA1plyTlVf8zvEZrhpU3HFM3h
qAyG55sFrqoLmofxldxn4ASzKs+nCvJjHsQD2wqlumZJRxgntu1CnnSW1dtLFOPP
eUQ1DNB4ESVvpaag2xNi+eKA465a7By/tdF8kQBhOtcLuGsllK7NyIj/UFQEhLzk
JVSfnVYEgaSVEXt0yM/3OUL3TYegZhiHuJMxL0CH8axYamb6tMRGx5VQbR69sV1e
OfMuCAyNzIl/GpWNe2P4YvPNM33M7sbDZtj32e+PazOdJ6dx7dSkqtklcXuuLs7F
F2zSwHWaMv36VsfYnWeMcsqC7SaxXaad0ot5Kp/GxUFTui6H7ze+sAUHrcugcSaT
tPJEnBqIMShvHkaVxZ/NtK0OtzAj6qBqo4yoG0NI7N9q3uJeUCsj0BNm/JlY0Qmc
I4Neuf7Nfc5FvyNAZtOwl0+TH2E3A84wsx20AtkQIKWEQKrpcRB7GcfMj4G30FL+
PrHawFeZjad+PPOrJSzer2xJ36UHuZSo7aWl9pnVAZ5G66NzX7xNvTBNt2ux2ip9
DRLEPZCG2pp+29o6VYa5iwFoWogj1Z3mh8Qlc75VieXoNkjJS65+zoROf0u7G9Dc
yX9isz2geM/cTml6EVeq8RGB2CO9EmQjLsysmZY+KQ56svqBP8COItmRLXYKR9fM
e8K9Wu2y3ZWTaDiH0Tk1Po1Krz1YWHnA8gbkO46uTmBN+Le2Vw2fPDa+ABGk1yuB
h1fxv6+z+2Ur32/h59uZjnvjeWetLk5bux+g/nKyq7hFLxO3ppz/K2ai7HBVzRG0
FLbxrx3VOOEYQt1YeYMCmG/RE2QsGVQcQGKf1gJA7lozL4my4g4N0yypkO2bCirS
NStnN6HUE0sL2RaD+Df6851ugOMcodASSTPPFOqHjXhqDZ6voSvszTR3tRr8/DnA
EIkA2RCodS8ZVlxP2GrbwR2SjxWjKxYrngofLRPnRT2l7Mfsh/Q0ywBnmqR1moQq
AcbXGiSrqSZPgffIlxlga2k5VOHSXuM7QWb2xMMT2FHU91lwHB8MbKhu9IZ2pItX
HaBlmspyYPWew1qZu1thbr5fpUKXv82pFz5Pxhp8PBC/YLQR1zm8mVwOa1PCTe2G
7BBmPzTjjAIiRmxC9UCeGE4eSIxvRoZYjc0h66iAhfjlZVJ1GVm/UJ0eLPYagRk9
Pd99+ZNofsofquvzKBDq7uVCaesL3GqRuy/DXl3+0l8JmDfy7a/tS3OHgZYxYRMh
Bp8mG/fP+0CAbh3/n66FdsdOzXscbgBb3F8j6x1h26HLekFgJLD0ZcPldr5JloNg
//EwrJGN96bAT0OnOmTXFepBAb4qE3sUHzqMlBYpPNqurNUg4kqIzKhErWZwndPE
Hq+CsgBalr7yFf3XRgLAZfUXwMSqd6NpcgURzQMozjprC6AntvdUd8aXkSORzlPY
8p9MJMaIrpLXE+711RHnE8gMAnHdl1ywc2KwNjSx6dmlWtw57A9inE4cjhSED4yh
FPpwVXKj44LUYSNNYtscX1CxWZoH/M8OOa7Nai8p0TRoPYBoW6IWY4yv4H0HtHwE
00rwxgh0IWD2a3MR2yiLI494S+cidvZwORys9q3QBJFNdxlF4ZjCk5u+rHDbk8D/
kRk/mOTm48warX+msTblUW7I8Npd7pI8izDMepmzFk2YxMG6c5j31Ng7LyM86HSU
nYsyaeEPydGQUbXB0ljf/mBVpBrR5Fl/Nu/eAVihBjWuBwe9HPV9kfg50Jn0xfOx
nqZwhcTSCSw/SfX4VrK3dyZjRJQYbUJ2mWaWg5Y1e/8lSI/S+ER7CKu/avkIb5I+
S+cGpH6lb5PT++OsQ04KMPCH5Fgfno0zv7dinLG2b8hn4h9Dgo0O0VJ1hsQvSIjI
sTuaYNvbE1bZs2VkZuew+g9rcvoLGZb4FS8iBh5RVY9vncLS+M5/TkTR/4o6ePeo
LD4REaws5x+xu+jCnlnjlhEpvuNqpNfKBjXw2DTcO+9EabUBaa3mfltXLTBG0MAC
xfxqQKNzTLA0MQAq3AojWXWBFte1TWZGK1tBOdkRIi39oTafMUpSkKSXjhEYPu3d
o0jVtQUpzVwXnQukqrDys05vvpb10CUQptF282jwts1lPi7ZvygzwcZ5RfRwniFm
kV0WjdMOvyxb9Y8rva9kIXuuuZwvqtQhk4yTbUhx6je+XnBfSW4I8eD2mvzuEWhU
Eigj+CUdO34eostGxNXELkDEDCIKTPwwCHjZK9mJsuqXfA6UPi0CBfBlpqT+zsek
t6cb2Olnb0+qATawrmYi13I9VSl7wrmLUFv9XwVwh68XV+mp7eiIx7LhGfpk0GWw
R4hKA22EMuEI+MhJiuAOboTz+DfFOX4mWJuegrBDPv8NdY9pbtJm4gVGbvL5KZYb
XA7aqOiiOvCu5aHFFU+4Nkf0SyX0doIbqAY9HMT+w7Svzo3IvcZ84Mq4pOUFJcd/
qsVWi5Teh2OyTIiZa3YtPh4WSn2yREWfe7aw95CB8Oi0IALXlkcdssLbXs/bIyqz
uQWqJZKIhk3Ov+sikr7l7J0SI2p/KRXB6/YOsY+BxS/fUdIbY7xxEaDJ3mPICXci
vo+6VOUVeI7O6ER10vl+ObHQhPNEpD4ElerlmmBVigWtJBd6XL41vlUn/hh041zO
INUWD8kIdab1Eu6oqRbxL/zmzE7z15pNc5s8VyOoYQDI5xZKjeb4WGl3yItNKden
qHpzDdQDSYXyq6tNCeSSgU7rMQGFGt0WaU4twCAXBEQaC+fXb4gdH3e+sgvJ0PBa
NsKIMitWHzW0yZwWXvaXEpeaN03prbKqEpTW2oCb+/ZkHDplPfJdOep29/+teUNq
sXkxJ9c5CJV46XbQyK958rQFfqwFB9xvkDaM4yXMdHCHvliMOkg6q0UaqRjX11Ci
LoPozyx2I1haF73Yv0NbkgZBULdV3JgS/CHY/iwikL14f5s1tjzXZN471+w7G+3c
Cy0tVS+TOGmPJqSIDRV/1XQ+7cIsCB+L9sGv2OqudsS1+P2C7lhs09ezYGZoV/k9
4k35rxu5oTUqpDWBE9ggKT7gqryuUwvzzeLW0MFYHslIsSm8xyhispjoZaH+H9Vf
F8wmSwXL3VzVBHJ8vfybBFYIY8E1jixQFSD9YB/UxXy4n0beYOnQHVMxQzUolj1P
RshBfQuMJEWyuRnvi+83zR/WUgIkbmEUUhzFA7D1ZoFmOb6ZAbBI0z88t9uyzlVi
rDazb8HS2IuHQTYY8FtGXUjqIXPFK+OYTjLESp228v6SOlTWQaTp+m8haGhiLhDQ
YqPzKfjVigBJyxA0e2xozHdkCzsC5fcCFVCfxPRKWkcSUk7y08J3y+CuTx/ToDMe
uHmI/lA57siJ1Xp16DaZqHcpeJo81Plw5xnMu/IjTDgquA3AS17dquaGAWp6HZYZ
OqJp0RM5Si4XfEbRFpPn1f/ZyRbmpigqKJh6GzoGSzy3BxvDoh1oftVUiWZnFyz1
6W7hJuvyxLcwjDuyaHAbTPE2kmvWNq6egq5OeFNxMitM6aWd1Bkk8M+zsloJkekY
H/Fzz7LBUp/PWZ6dnHyH8itvwPXMuXxZ4mAV/jRl9Cepz4bv/Qs/7yk6x3hLhGss
1UnCJq/9IAdTdOEtkELPElfHrAhKyYOz41pAvwCQ5kR4+0vbsje9Fv2O6V8HVhyh
CF/axCfxYN6EY6Eh5FbXy4qVxiVt9le85wzG4oOCqkvI7Q1/369Da/syJH2mSijX
l0gJJI8/9wa2u4nG6BB4EmdYr/A8yhLbgLqzhUauLqA3s0Og7KIpe/uA4021rEW4
zqu5YFMLiZbWuVbmIhXXqMzsmFrqM4vfO/rPhZsEIhi2B4Ksw8lAqF0H+C1HSPKx
B/Xy13LprCiDHRaeFNbDm46diL31EWWhOVWvlM74aGGv43OKZQqz+gSBJ9o0yIK+
8WKN11a3vmsOPGYGQQT2rEEfW3kHftzXRd1wHx5QyWAyN4hRTUa07Pr+zXPCkFeH
zep1a3ZNIuT2RoD+rUfw/fYqdxGr0k3IW19oHOAcFvBR8kg0E2Vm+pW2tbuH1Cbk
4zdcYv98zueRT0/lS5hOm9k0dLkLbSsIqXMw0JKccpNX0wWPsGVyJdChMMjszOLG
KNAhGWq6/Aqw9XMK5+19gsB7x8k32Ca9o3Qh+BZr4BrVlXnujLmD8MdBEGjw40x7
pYGdXX9Jn5Us3EFq7wlAmpbYlAzReJqnAL1QhbAndiTJ7t9hKmqyAn1rLD+WUw0H
w+dnYw8+SMhOPDhqppfK3VK3Xk+Ihkzz3whWFKdTG5v/MPWugqEVfCAagram+mvd
NzA6VE2H5g0w0qX7askVae4DvX9nxV4NOHkpuekP+dce4nN3uavbkUsq/ZjMURDQ
e86Pr/LCPrN8bwtcZRD9ZB1WvSFDZ21BBALFsgrBl2OTk55tdGMbK+X313ukM5UJ
Lb7l2UhQwM97dxYiYZ7sPmqFZx95Iw59HPJieI1BJOOxcI9dkHLeePz0sygFOiw0
pd5/Z8jxUiZosZSmvxxOwxgfyGiJb0RQ3Ybjh019jxoxWVo4JnaHRmZcI019GvWO
K0tBe6zyBaeCCabKRE0c54zuygSB1nJQsMMTdSN98kF2nqDonwXcUBdfhu+8LlAw
NJMTGqFQb3tmuyrXDWZrRXECo8PuiB9E/6m6C6n3l/X3CdHFNZG4qwIcHaVZ/Ymw
MnIc4aELGMdW+TXP0ZY9ttx1CUzVfgYSX3FvnhyBDNerRMnl7xwXboVWL0uwx/Tm
rNa/JduYL5WZGmv92oM+Mv+zn62NQeMn+xYMYfStkea8VzpcbVJJ8EYYirUgVTF3
O2l8ekfrBsKKpARmuH2iZvNtUvaC88TwbXz90ein3MyFyNXGjJ5VMKnvqmoahk4H
bj8uvTl6I5N537NVf06WPEPVKXWjFdol8hCLG6LWgr661j0smvdkL0L+iEvqPORg
VYRsGR8ON9cDJmxjhwbR087aS6hQAV0akMsmL5UZtWtFspqqXTYv45mmvZUhR5xu
d2Fn3rU69O84GTWRG+ZMesn6ZqAAhj7u5Qwl4UlDMhUjSYnP297snirH3V4DTQXs
9bZCz1iRf4mdn7VZbHE2mV1yx8ebXJ3Kqqd3tw6dDrfsKcE2TqATHeQvukYvo6S3
AkGlVrZilI+nHDn5AlRXaUAhSVNRzLIAV8Eku1on1RKDzY0oO2w6YH07MK12l9Qk
VKp1SbZeZgn+s4vqfL+Uv5X23Hm2T5z4UEZcihte+pUGX2TIDFzyCiyVdPJNB4NV
d5L9I18HrRXyKBziaDnTqNapJPovDsG9aTt/oXO5nW6E57sZ9a5mukXVT6cVyzhh
MzZKD++QT9IktobmuVlWg+UNdiTC6EqwDibxWt4vl9+GKn1mHhNlzT4hx3IHwaP2
pzyYI6nW2FvdWaYKOHirNqohBlmbqvi1/E4q5yokX2UdfHnZmGk4jG4HEpqDDa2M
h51O/g5dqEcFfAn2br69FIgNiA8OKUTWRccUvvJvbcL1zSz5gs9R8gAV8T54Rstu
iAJAaOuDStFYkvIilu7LkYj6dRZPBntk9XAXsUS8tsSlWXieCUBDfMUe+90+WDKs
KZGtYN3/l12GKT/yLCP2ex5k9RMhFygY5gnSbEv7Tv6fkBJtkbHhHp0nXsj9/D8Y
R0F7UXOcBUMDNv/Ro6dXYK9a2WNSosGUK9E6b1Z5n4xWWZcbGZpNz7cJsnXWzVVt
oRyRhWZWp9aHocjGFA/lKIG1M9S04D2EVi2nkIrDqoD2zY1686AjqVjTZRCJ3LuK
iC9hGCu7e14fKq+8gOV7oH7N6WODLY4/ya05GuQp/OXbvO1bSBI/ZY0khsQMjg1m
LvUTBP/SX1eGHkzkIJDf1vlhDFMYgQRg0qL0Vwkf8qDunyx+mvAwKpZQorG4764F
10Oxa7eniISN3I0Swp62XxrU4uUvnD4uTmQULjnZoMaLYhIR8eUl/6oHQRKaJIUG
BLiT+FxkbiKJ87nAW98MzXDvlF4n4C40O/7XgMMsv2jP8F0FVrxb9y/m9q6ZEHOH
ZWRAWQkSQ4bB8VZ/r5RZQT0+0u1/i8tt7E8Xs6iECl3pBsNl/uRKfD/udRzSB8wb
N8wrzRs53ilckc/u2zUh6UIRn5/hfpKuilh+5CrcXJBe2c9wKoZU2ljpWVnAb5zI
9zN3UfXn4cBe1Babs6BOeQo/5AUVuwzC3wqh6VFfN26Ag3Vxdy63T6RN34Dx6K4X
8AJaufTNDm3bt9YZA5QzaaGklKqR1fyS1K4dUJpki7ERLq0KpE8vAtpuVaxb/Asi
gpDmcVrSdusdkKR5PIIC7cE5I1Fry2mP2UwpZtyIsQJx25WT86N0mUOsRrtGJ3ae
TjmcFMpSnBncxqwzJlDnUFN3iggBLgoJBdNFEc45+YfTqWvIOApKAFbD8yc+TVur
91D3Kazv90xY2G9y0wDBfWyKTK3ne9SO0mmmfWPooH7WmkAjvSzvUp1R+x0WDZ+n
JAKK0UDCpUHEYAuJifj9itD66SwVG9D2y2Eibp2UOzIOUx4W+8CLLoDA4q7X4R8z
CwwIw+kZTsE/7ctNx4b2N5tg+0Lkp1DBFcYW8N8tGEwyiwXAxTNqPZXBtP2kUHj+
qN4X5Yn8JPZ9LWQ/9yr9tkKTFdqiivGPPdQABpAifvW0C/1f3aUboulFu9JErv69
Gb47wmKMEw6tn4Bln+UFjH7itRyFoYMNKioAmDMFJDQnAYoNJulyggybC7TVR9V6
waFRL5dkZdCoPH3Z/gLSDIB9eVq2NU/gjbzTzv5c+cTIxhp8sl8BxgvMuojPtifk
7GJ3a+Z0OnAjzBIVD9IyH9npY/hvPqSUlKoHjMzl4CzguYOoKqfcSIsA+hTNEJJX
0aUgrgTKbWakIhv3T5LG1TVGNo9VlWQNOTOgEnBCG0wYvI0VqNiapZmeS8D4aiOx
OLRRXOYvWoVwFYBpYLK8eAkvPyF8t64Aj7Z3d8L2U3a32BJtorCrBUUHsjFCvKDk
a51dQQJ/0RlI49GawCA0ZWIyOyJYUx1Joj9kp3a3/wwItyC8gk9eB3p1oHBSsI2O
nsL+gBc5ymv6QctSd8hrLItR1KRmICyrIXHCatF9XmgxUZghJ98h8ppJG8AltJhR
ajUdEkp1H5AwdVfDuQ7weA6aJ3xruATQ6AOmhc+AVarItdjtDwO0fUYJjIHqBXgV
+pl6F3mFLztQbifKiSGnvhTcGZFaOMOBJ8YBVfm1j0aB9Ogp/MYMWl4L6ks+MNTF
qGzuRFeWnJTQAWZm9uc2ezd2Ijq3xsENJ8p4M0cZr8b+htTMmceiLM8RMrxVDUxP
O8shb5345Hc0e7fiYWzVFfE/rKIt3SWcdrJkKzSQTzDIdEyyDZ85ggvtYNQfns53
CamR5uUD0/IPwqVt+hyDlwIU1IbyB7byrHe8wLnxahdu5zgHWgQ0xO6ICUUsAyN7
0DBVyswAPIgCV4WqtBhQXKWC2T8mOddDJ0QPNxSu75Y/ILF1+HQElq2jw3/ThvTx
AoQSl7nDtSqC3bT9QttJHHhaPepBVUb7Vi2b6P+Qz8gPl+jyhWB2hwsMAcmjPK9e
VEWc/+vAJXTwmTgXx/qJG955gUcwpKagxsVZqSGkQA9jl7pgVDehtecmeBE8Ts2+
Oy1rlwmDLKfrSqQCQqmpKOqNpWLF3xQr2zfGNhCnfXaLjW6gAIneoZ+ecsYnXxsb
P8Rco1EuEbuRNWvITHTwG0aOqxPMATcRUYiBmuRYywZq8L60aSAGIKeG6MGX4d8w
QB8vpjl2urqKJHEkEPGm1VhZCwcjDQ4sE+bBMMgW/gvQmlnDLAkxmrSzfY7fsjEK
nZu9tjgjB8PgpuzD6W1fwButLkgYfZsIq1eDjC5onOvVhtiO0IZhnhBgfkjIDBt4
e862tQun72upVuZMsElxU5zdNEZvsj+/ceUWlfovmVbRG592mklheEubPqtDfcD9
K40DunueDfjQe5NJWW/iArFZYqYthKS8lQOtiqURUW0XPuVqWeD0jwZWZR5jcsqj
biQFu1ZM75mHkaqYWemfYsYqNMim/Imn7l62M5nyvlyqPC9O9HMtKLxBY+Ot/cl8
H5i/MPEWvTeahFTxSFYoEoDMOCQ8yobJr76i925pwsE2rn4i0E36szU9yX9CJeBC
nxUKT8HLyXmVlfQDVYlk9ltzrj5/lcmgIns5/VUL5YcgnZQX8EMS5wHK424rv/1N
YcNALzoP6N80JLXGKXzy6F0Sm1RNkVDtUkKUIRtCU/VXRI7XCXYNTcYQBM3Ir7CU
BQ7JBoTygjZUJbcUZUIn9KuitTKXZCrDsBZHlnzBOvhrdlu2mLkgrffxcbCiboYe
uGv9Q2Ral+lL74e3teWWCCf95IEnF/YjhPaZSQadWM3b5aLP+5NsWAeJQ93E5n+d
uIoX8W0TmijAabkmS7SHNIJC5VMucZcXhioWID1Ynp+gdBSjKfTYzo7TF9wEej2C
lICUanfBXdK1iJULu7nvqh217MUQCmDvsuGZ3Ylx16DAMTa1UEcJaYgbYhp5NmQg
l3QjorAupxKZhfapanBsSIfXbK80l5FL/Hr6sbQAi7H0lctHSLy10gVR0Ixir68b
gDUPEUDvL6SV8UAJT7jBIb2Y9qkCM9IZ53afu+hx3PtwpoehlahOOPyvPPlo3xHT
5DTcrRSboc8vIO0dW20Q8ASrsRQdZ/nP+y7qpo1Lrj6yZz5Z/I+vMXcqHNnSDyur
uZkqbaLyJpgd4UeZlo5Q5LaU/8dS7plBiGjcl0ME4K1yt+wsgX0FjOZXkab3PMg8
NuH02SkVABsT3Rh25SipjbpVISTzb9oK3ev4Im+QkFTDn/DTU903FaTY9nYuAxGi
XCeJewXMpW1W8JaRaePdViT1dDhWkNCvUxbHT3+NOdpLZo4fnr3JflMzgVlmg2/u
Lgy3lil/bnseVNc8MuopdXrWw33k2MOtRb0dYDNEDGeQBIxBqnznNMbtCSTuiyIa
LsrGr0M2Ypw+I8AWrmfmtyD2y/15qmvHoAcrqBBWpgWSkyI8ciNQnhuuD/PIfD7D
l6Y0qMxbrRDCFG2MGvQ7c9z5vUi4Wnc4Q2z8Cha/Zq/3HfoBtLEnfTwiY298Km+7
ZB/K6N0JTYG2z89f3ryKtTaszex8esr41ORu+ThZRCcGqpkUSZtlPEU0qsNH+95Z
o7Wnn4kQPtnI+pGE6Y/Nu9EfjsOXnCZ6b7794wa1KrjqZIe4ChdMz+HbX5XeGl9m
G7ua/juXva5ew66GmR+PzbeRraAZIE1JUK/CcLF2KGkb+BpDa+Z+5k/+oJmoyOU3
WeoiO5/EswiHNguBB9CuiR5Wfodtv9YICapjJ109dDO358ikUyMSW8mLmhA916hG
QCmDkOqlt8qFt96CkkqVHuYzFrOe95xnAyyRNOLdEuMhQqkW2emKFyeBW7KPKfGb
EdlPbRE8jORkeMxPx6IjTMGsEL3U/3BUdN4//Megd/B8aOCQRrb+c7WnAvXIoOcX
tzWUYNEiyvjaxomY4xBjuuIst3bHjlcbVcoNRQfpPSMR8gV5Na+UFmGl1nfs+0l9
xTM/CzmibYxSYd4E/RcT9zG3Xn73UZ10DVM/R9DOk2TiGV9oBsWxZ2inN2FKaMr2
UcO+Rh15M1oUa1i4hEbmHj+OBFBgX+2w9ix4NzKI1dJjYNk8RC3+jOSP8jqxonap
r2HB6XvADECjpxpTHL+4dG+FRcbAI8XACCkhgyg3D0BYQqDdjbMnYYbeOK39hkSi
Xh/y9KMZQecInLrfY82rSj9HxVmxTo5ead5A7rP9/8IOlCwsgqzrDEBOXzPai167
iB7POz+RoVxxYpTAGVlyFmt3S4xikM6/omk6GHpXcNIC9jytmU0ZgWlVPELGYXD2
n/lqBdxas09qg+mVbM7uE2NbL2GpL+NTPoyjveGoaCKvUJjFV7l8y7vQNy/c1+6s
vEl+H7mDefFFsmrU6AmyW6VAdPIhOpXHPomJIduJj2687K4uAeDmOJjBLhORxUbz
1MuJLKFszlPQ4DXUztIVKIan5dVups2kg8DNMhAYgiRWQJgG5+aSQjVwaE78uSVG
RpVTiJ8c+0+d3fcINvG7/Q/HS+O8R4q7x7sRU0zhsbImEKKecoR4a1riQ8fDh0fT
ogJQHBSQm7VOs9AVSJor1bv/seuozZBGl9xuNw7Vz5fRJqNJGCt/ciECkqRQP1ln
uywXl7Tm2xuDL/6HXyV/JW8klIoyocozTOuovawjgZgZX5d1LJ2C33cQA2o7N7KV
96lwomzR5E8kOEqt3BWfjYqw1dIpNVmD17z94Ft2AaoqjHHSuCyPJdeaTZs3OqNB
jTrki59bY7jSOsYuM4FosTL9w7pB9u0BpT76Q1sal42oHXLp4LGtQ79oYMDBHwBC
RrTJMe39Uuo/KjdchshqQuvah+fDJUvs3LoFgOwE8PISMc230rf6yDkRz69oV/Ng
PClMwzDT5mrc73ijsWDk7SNg5qVe/dYoVg4NKIIWN45GXBcpGIPK2aFc+nPaSvJO
v6eVcTZQw85qL+fRkG10TdMCfebkJzwO46nxZ7fZag2ero2Vgac2NxVHRRdjbD/o
QVsdB7FVaqb/Jx1y/yzkDCzqnjzO3gSoYqAYBXjmUp+6uftWW0z/zXiMHrOR03SD
KC7Ep+A5Y7/wEyHMKGHSLH6PAaiDHgN9qhBBzarUW6pKY0H76RGuhxY0A+satpdJ
jLiA8nEp618+/3PgGsFGvX1cbhofM5KlEUyZMFC2xPuqP5uzS1WtynmcLo/T6qDO
eKp/HBOZXVuh+1sfl8ksQiZKdbOP4M4YxCeiY+GL2jveU+5VkIKfjydEbc/6n9cd
OAHG9D4GTo4cnZucIKgUF4+0o19PQ25Dgn+ozTGVrtkwODeFdlQWFK5JpCSndcD2
ozMufAKyM1+gKWvEJ/7IonVD7Is+mJAx/d0KVXIOSo9I4+qISaYO7BVvutq/D7yL
hQK+OJrua5so4d+hhLSYYTwBXpxIuEJ2263UGYw+K8ezKe2tXMlbnd0htt2jmxZH
FL9/OgVrkwgUBtaXpLkk8honulord2yldONT1tCcZqgb43kba+JZHbapXLNPDV8w
T+QTTAkJUmwckmCAUEIv9G7ugBl63Nt4q+AwCeytJxKu7+HusxcD2RflgC4LtndM
36Hw6T5RFyxOpIGw4kn8Ge9XneEpLUw5mugzGrOPaWAv01DiPEhDJjPrkrly0Mrz
zEKPgca0jMBX763/BC3Ni6fysy9weTtfp0oVpjAvpknqlJtOMnRjGkK+1O2Gz9rn
LA/6/wcowbymLwNJ2ASZek6LbICBSnZ9b45ZZ1YCElNj4+xXDBDnzkIypqrt85/J
K2zP6cYKfasT17UOF3v3u4XbrW+arCreYgOZJE7GLTg2VLwU/Xm66Zfcxvp8CRov
HU3EjEJCfpvm25OkPE1+Q+QtXMgc7MfedJ/WYg15W8rsBo4y9bdmcc04FzJgFQnu
VKcOvs0DX7CojxOuUG5gIHKQfrCl24tDCwN4LlPbPtapeKJykgnhLwnSrtXYIr+z
JxX1hVUZpr3x9Awm49ez22pn3CXaC0iT4BqO3fGwEmxyo5lChwSb1XHZXwXGuNRD
UGZha/7g6NpHYw/kT1Gx933HFV2sOJyqHcgdD/NBtDC6j50FutjLHj+gjuTP4vPa
aoqD05FDxes/tk1sdRQ3Sv2PZ2mzdXf9EFtD5ggPAo+1UuG7bK1b30ZY2Z1mBpX2
Fseh3W57Gjpybiz5NwPw1pbnotQn9paUg2wrXFhn9r4UmBWIlMrT3jgnkalZwOGy
DdMWEY3KbrYtqq4/PWSs325htmxsloNmJR5IN5eTP3ldYTlLTmHG5eeBHotzXflz
2aYyupkzR3xNdnZdq2sOGGxjqWfjdeIKLU5IhX90irvqcRRfI/uxYlNDNlEhtoh5
5Qc5oJ04fX99TJJQXTuh+5Yr0iDUA8l6AabWAt4YaiV00/w/hEKPZbpWzYe8xusa
4mAJqMkCwmBCVpZM/731R7Bi+Ho5diTaCxe1iXhSRozZEO55umXoRu1pZDNxN3rG
8zkiALk9weGrpj0gV21dFDYFzUIk71bNkA7Kj7H0Tmj2o/YwQkrVZSYugVgowtrE
YMI2vMm6sK9pzkaERvYw2kSdrCF5NpXyWo8PTqorVYBvgjv0SKUXn+tJqyj3kqXt
6Kv8OyTfQc5WiXQZb97Wm6u2XbvM9yA0Pc3F/5CtmM7aYJVItXGcKLdIpEX2MFeX
bcqb1f+ERnrOuDGhxklXXrRlejXeYH1sbC9Nve9aKO1gxIXnbl6U9xvpiimtqaX9
U7HQ6bkblndfNr2CA5TaGIgC2hDVrsdvm/NSC5nOCwlNBpSxLfwYKKyFbUPKTPkv
pIgK5oR3Tv6fVx/sZmg9L7qsXZtGp6TxP6H60vm+kaOfsocEDEcyO4AB+KSb4UVQ
i/mNGrRr3S1V5npzi3WbArOFXsnVMu2GD2yzhwwN0L6lCPcUlnpt4kbkRF/CGs5g
qfmFOCuQodm7fsQ8h+izt0BvzrJYo9lN+jj6DJbxoVHJvPy8UVG7OhXpHKi70mxt
jLTVzUCHJZJ92OIWdZxph+4tbpKXor3YSwBzZGTPhOEsS6BxgiYxNemRxVYHsA+h
Ems9trkGvudqKwr97Mo/pM69/w5E1KKNEF3QmqRBRXLqQV00bTCKuw1a+GlXTlc6
B+oIJ8dc9rj9cZVDFNVCc3l1lTVbL5RwTNlwh4h+r9+JsqBMiQt3Fef76E83Ezmi
FMqBodzASnbnSfXuKNVwWz4RK9JnqeHxb/HrTtApnGmW5Au8/T0lReyzTJ4mKL9Z
tJL6JCU9rjSeGtWI7cHnNyZMKQ8qOHQtgCsM7x209jssLtBwlKjOU0kFojVNqmiB
vYrgRq0n8RLkWR7J0wZhlTzY8GObSpOOYaJ9fTssa3USlVXhrEmGUfXRd3fWqhGn
qK/OKu9WDLm92iXu4QhDW/HFTh6Xg0Uk3pmg9By/aQHudVjuXdagtI4NwUNyyu35
J/cr08SDWTYPe5bHUeozlBzUWNRYlCN3fyGRUXgoLf3Vm8+P96QjL7sAh0yPUxB4
6ahhjXX0ZuMDqJNPjBUZJFLSH2DM7e8ajg6B2ZVLmns146iyqvuhiqkm5S46HKWY
BnBCu5Ksfrdwkyztlbw/Wbo7CpO3tz/j0ChxcK8txSf8+sXHojMziEJaeRo3gUzN
sMK+8ebjLxzJLM+EG5UE4+NAR7MGhFAIIs3HMXEilhlP6R4AwmsUq5zk+7iVPocH
HirNYpYxFakkeW7eE00Y9gWXTfEaNrgbB4dOtG5QZ27N7jSSGOdMzQwSTe9YzF1v
/s7ahGelbkJFmiQSM9GjadhnY4D1+z6bxMa0SrRN86KIeY14+BfnZ/F8OOyIZMwx
qiFqxmoYkP0FtfshAK0IX1Eb1NcfUpDcahndFKwukY6eKTfzlpysiN3WtUH6pQKl
m0wcMnhfv/PjpbHMR8ny7t2goILvddDefSMdgQgUlFWsbtTRkDaazRHsR5ZBokp8
G0cRqFwtClpCak408PK4T4h5qWSiAPUMvwZSCRzN6jKrHnQz7LWQKxTqRjezutNX
O5r+8D88mNM+duEZYA3brjtmyt1GlFI5NXw30GYSvBsWg+l+KYMOBFLTIqf0a2kc
NZx1Ooe/H2ZXbccB54tf75d+acaWUp4XDcg2iwRY8m0uRLidbpIpWGX49vMzGVRe
3YULRNx8oHQLtG5Q7KgGyXgg6UFCnbwFaGbgtyHvZEimpp/0ljUFUjlZ/k1J1pno
gYNOehuo/g6nKeBBkZ3oj25naW2v2QP2J206Oa1hPHh8PYgFvkqwfVTDq3n4E6X0
oyq19NUwx5xT8VMHpOcAChpgWad7ChQM7pOeplIZ5YXHcPB2Td391WsJgHQsQ5Hv
gvkjul7bCtp/8CN9AX3ATtIamPbYS7Yf4R8wvncmEKZqsyLFde1IYKJn+KBolWlL
pHifRPiskk+TO0lg/rkYJW5OOUa8kaDWUlSV50flI1WRUeSleVhrq3M6U1nxcivP
E1sDiMIkNZgWhgy3HmvU34rB5xFyZRHEa0lKvnH94bneLSU7IYo7PESKWnkJHJLd
wWrEQzovSCuQq2oV4ebCkFxmwXjKNo4WR7lCJILghOfWUTeypIMJBsnv+j7OlXdH
gigKyTG1cAiMC/C1Vgny7/+nfScMDJpORTjCC4ClTIO16Se4PedLoF7Uv9Geelil
/2oHr2aEa5o1fSEA0ETDEwxuajyZqi9El9pQGYOZZ+8bR7XfpDN3PnijiCFDccLp
GIsTkaWTMcGUt99lwhfzPsK2R93cLgkbgIijXG1yicO7YkcWo0s+Ollsq2/uqSZl
XolOJERDVXZjv3bNw/J4RBAMBsFKNzw3OxieOTkp6JxrsE1tDxVTJI+MqWL+EJ1s
dGiD3julAndOfkGRN7Wo38BomaIMrNPPdTYhVW5EYZRr9gXWys2Gh1HGirX7CpV/
e0zD7eJlYpcR8t/cXJEbzWTUvLJ9IkIsnujcLrGihbxKqi32BnnNJCFpvdL2lC3Q
SfXI88rn+ywYy9Nn/gXcjlJ70lXkgsXi2Ydn5AcmDeyoO+JrDpxCHYmUQSVQyllf
4OQ1DRfghixkqTn7xPJL9F4OtF3axrtN4yj4ogpAkF/GW+id9vwuPGmK+eD7rqhq
Hhy/E6DAShVgwsOfBoOmgPA3G+MJzqygFZ1ivjCxJOgwAxUTxSzhfSbYUwkxsRky
A1UPt42dBF5vMa5j/gujRWTJsxAyOf5W3wLXXYUxGr/9VBctcssTIBCmTOLWytqG
bwzKLGu0NPV5idzmX9alxgotdXizDtIn4eZjacVlqVt3dCBhxy+zldMtZU9FHTzO
t0PMjhJb0HkZa2BoEf6lZ7UrMKNGed+Y+SQZz8V0ZInv4jz9SIcTbnFPPItd05sF
KMfyjrTbc9BIK9n2hne880RIdkThTRKpdoox161v2pZ3m2kmj1YHhrX/QUYZjmeb
T9DCyL/Vvt17yiNs+CQzHiwo3hVuQPwoEcdrF7cRovGKv1BINUBLKeOWdoa/UbB6
WKcxpmpOhJlHM2SIihxX5osgQOpn/GmDudS0s+vxfAoKUDhUgQYccgy0NoaFB0pj
nwh5rLWwrB44l8W/rEvq8++gP0rDIsC0DF32tjRFRlcjqYz6cGrbr85GkSRfjY6/
pMBczA4QU+xplVPaWCJeyPeBfqf3klhW5yZgHTZ67ZjwaR0g2oPJ3iY2rvAtsLR6
GYGEYhTOrWWj/EBt1Sm6xtlyyMp45cee1Zb/3eWrb2KGQLXXJgR/asSZMYMQl1db
2G0ZTfr701jUkjUHOJ3yKd5H/UMelyM7wTbOM/DSfCcFQVGDKIhyZJn0JKyhK7vd
XNNtds+INwnwQYgjh15zM4LOeSMUCYhHGxTFl2A55Oro9yNmEaJgZcwjuyvNJnb3
SjY9kwLOizD5uTwbKVqfN8Z0f/uWM5aQ7Wgtluc6/NxSpxPfffYZDPwZlK+xWrTo
8zGYJxUKVacl2C9W0O+vrssSHUvNqaKKCf9dpW6kpwsS/WrPXZ/DMoGMjxCF3Jjk
ZNGxwoCVr10XLmuXUzV1tWajRlGlpRgVYzvthchd5c1ANIaD/cKyfWRcYUYl7fmm
Rh0uJBCiv7FMbas8lzjwoPcJ3l1NyrIAovKC/dIKe+MtHhxBqrLsqRrWEAeGM0N1
t8r31WW7VXOSudlYnP9TayDIKwklmGeGAyDxR+KijnIOboOVfOA04DqgbyNOA1dJ
ZVxL1HImZiN3o9gCLxlUooKUZbVE/8Pv0GuVMk0+S8iVXDvOffcWKEWXNYwPdA61
ee3iTTpgjMp5A9SKR06t+ZMQmNBRqKmPWnHRMpi1vl4R2w48UCKlRQLEZWiUE4YS
L/iJMVVKYfDuEgkAvIh0EhMrzDCb/E3li69CjX6j98aopH5BdmkDt+52CPbENIyy
/qI7Zw4x2aq0KFrpTQq+R/Y0IG3WsDg9IFZegJayExRWNaND/gIEaOKdQ3jHXjom
m7ugiRcXRmMXCkEplpHowhAhRxQ8eCigvBXpiY1mksk5WNcMLSe32PwmrOPcvUtm
k22H78lhVUQ8N4xkSH9j04nygPEVBbIEvRaKs/WnhKU7K+FihU/Hvd6Tod55qC0Z
3EuvS/99Of4PkfSVzf0XMV8i1Qow8nxvidbKqLRw2VWNq5Pw3peCYP1/wAOfKo2Z
lUBHidLeIxPMJMisl2idDZwYb0hFhq848OO3Hj/W0R+MS3gCXJkmPKxDVOGIi2wb
Qoymduad/bFrE4WdStfapEszC0BWiUOPZjvtoeKx1VSe/E5D3d9JBtGF6zEFSWMk
Qsxi284fMJFNaOUdqP4RITi6VFpC5n6BddtGTduDuNzp6ZHhZSb4iu6g147UCnLu
UR34OU7fiaftV0RtKpK4zokIum6HlW85lP74IwUTlWOYlOJCdfymh0O8uDBt9DhR
5TGD2duk6VQjuNVS1ImtSjZ9yUu1CEa9p6ofNpEFaafxuLf00SRoj5hc/UrF2QyP
t7nhkMkE1/qXlVT8ZpnukH0wFRy/oSkKdw9gGN2U7eGBDCRu7Hwg+P6KbjZPN6bY
XrcH8ptJBGzMWHisxBvS99tGyJ9J7EaYhmTFz2LPxqgdXx07gir2A1SOt+f7vaUk
O+GdtiZM8MOo2+3O1mXtNq3Y5peB3weC1F0Bn99x8845cUVTV68TEZDR2M42Sbvg
n5qWWxhatffCRubSvvU/fqJjpXklIYmobwntr8DKGdCvP4vbOfblQf1bgZ4LaO5R
EjSRqX4XTBjHwHmPEQQSvec8Yi0usgqgxcojQad1xdR5Ora/5NP0bzby/TLuGZ9K
6ZB8DPaXXsRAY6elInu8QE58mc5snc/VDXfw/g0TuUZkDXw8Bk07xjoumjj9qumX
sAzYA4wE6L/VoGNBSbqHHovaepbonDEUu5n0TxDLoBcC5CVFxdKBw1DCgCJs2T01
4oYaLy3KtSYDVXNOtumtvo4/Gbk6U2sOg8RAyfBEMEodN+fHeVIfVQWdHmdqUD9K
ntkaObEqgKRiu0iDUtQBh1ZamozZQRUgbJrlW+uJ6+kraFm1r2eGiYzxxyBzF8Ye
CkNrLSaN1BJWrQUoyYIboEZb+Ff24rXzGDwdZZ0AEobu+c0UuXQSXTDHsIuTHbdW
vKH5niDhGiz8Goo3rrgjWYeOSaIJNmlCI8mneT2g5c1VF7/3YjeuRG0XFL0kd3js
5mPES7Oc1LXPXx7oVrLmDK8lKvWzF1gMVgpcD3fOhYdRo0o3ZrEustDyXhqvaNah
ngmfRQtof7J0/2rjWRLBztH44m7zhhKAHDC4jGMVodfkJA/8n+/Je3jprekhwVKw
YMmhuunZOPOm8OnzMSHHDrzyvha0qbZfFV5olUF9zrudarqBcTOxnF1Olbka5lG9
0DKc9EjsgqWObnWLCtx1a7zJLWfYGKdIe9MDlubkGxE/xv+O+fs0p3JB0gZGlg8u
/I9/t4SzCCZ44y4Qyfxge2XbKS1ELZaVOIfSzzY/mhBNOgt2bZz+hQrWqnpa2v+c
GamBM/zCBabBITWNf3WlPcb2f/ySrHxzYl5WRoTG88ZDKv1MprsasFXBF4JG7tA3
sDoS15Z+UwStDsEFuMzF+HNPjnQ6/FLEaQt5LqofQrGCB7eNLK/7NG8u1KKFlVR+
tP0H9os0KlYjNh3/DTxyIok+drBs9Tsl+iFuLuX6HDE9KAenDuDvBcOgLWe/aPsv
lnZBbUbnBUAqRwXkY9xAkkklU9M5+D711pTc/87SIZWvZGSYyWPWnz70bQszUi2U
M1n77QvvDU5Qw0rsaaMNkKaXhv7uicIQrtcGdFB3kq9bRkd5XZbYlcUjXa6RkpcI
e2FcMTpEn7oDDLHyP+6B/oPsEt0dKE1rZMA6JCwfYN6E/iQ10cC9frRuQLbLFJK6
6ahfIu41mb5Zx8lNkm+3VwKr/0m82ofRJpZ7oI9RirSAO5PTh0o8tGbs9ZZFvj5d
/0cPIF5WaPvpaOJPPSszLzyZz0pQY2McpC/p1xf8s3KiteZybTocvYiD1P7HJM6k
/mfZuoAltZthT9vm+P6i4izFV1rFerSCgvSHJwoAfyapPYzoWoRGI30Be1hD/Hcv
/YVvHN+ACezp3jfJ124DzEVcAiqvyhMaO/c+BiCmm5t9Ms0gqlTc2uJnLYBswE40
KJO7gzA0zv+dggbqLFsTu3pyVunKithwm8o4eadIRzNcuW2wp9BR6Dt5gp3efMb2
bzjmvqKMyymXWSzrYpvS/snaJBpXPAI6qQjISSewJIq0g4ys0I9k628Y9155d8FS
gs6sJt9zA9obq6kQBRUBy8yaMSN7YkUR3ylbRCmndMroH1J8V1l7NwuXYF9qkpA7
jt+Ho+yZwuInQwC2vyclSHkbEEKx8N+4fRSbc6HmlQrszi8AO2QhZM7mE9MsqZ/o
2QwrWKyLx7WCgposJc1gXHWg3QtB6V6UAnddXM50ALS1jdhLkcyMuDA42vvMVbcv
TmLS2w2u2nRKXF+pvBcQRtQ25Jy2f6ytjgEzRXm+hbOQP5b7gu9lOMEX6ZuHHiyi
js3XGBTuP06qZuXtmEywxldZLeU726vD/3pg9YdBeNc/FwIc74JpVZ9aECwC+37C
P3t5T8Pj2mJWwN558RWR8QNQaMeeVOtpbfFOJ08ta3cnKsmhC8yMt/83rP3vY1hd
yRbcNPtShL0IPuFEpRY+HX9PAVaRR3+7H4MfW6A8+NbZl03MK7n/ZgQ+N3uxcEY+
JvjEnxiehUabTBY2pAyrieABxB2WXLlSi3eMjOTtZBwgBC7oydwPzzwsCZhobik5
9Q63B4Z0UL2bWHlnORp5i0pSLtiDajeUxJtZjJE+RBySwbFJ9ZjwWJO9bNPOBK7J
k7KK9eOG95kc6RGBD3oBLcrb6zgV8c9Zxx375fJiF90A5boMpKitx9c1kB+gg1L3
Fw+H47jR3wcaj1NLaZu2uFDHQYTXJMZxzq0jpTdZlZfkF3jJMk20Pusk15vStc64
MMgiyljyEFJaEdrPntyufXkLXUGJlgobucHWyCclSw2XS3M7FjVktDl1zlcL2l6X
mG6NyaUM7zoCenocGn2Sa7Asg7Pb1z0Y7XgEblv2HBxrl8LChGok13bLC23VB31w
2EKYO7Cwsskqpnex2wmDb7kQROXEQ7feSwjkEgq0jcd+pC5lJluXvytM/qsuxl9A
CH8mphUwRTwH2a5NfwDVdvOhWX2ZQf36I/XKiqLzARzK/mW0bOA5yk7ST9+Pl6ol
ycpo7nRXw4EIYiG99VE0LBVBAO64OYriujzI2o9dPoqm3h0Uh/P7qNzp7yC3vo5J
IwZmdiEAWxXwnGvKtwS3wcb5djEUzJrBnsdFsrpMPz7p1N8qFmFyptYP2MBXp8nX
nA2NxjIEvJGsH1Yalr9YPdnBBATGNqC0h/XPUBNIVWOPS68b2kDaoVaqKi6MCYTd
4KlrProo0mBK1Cav3C+FD84gAxj8gvP3LxKgkLGr91qO3W/bAbFbK05KSPKs50LZ
1o1nzjXYmCfeXYpfrShJYxbF9YL3byw4LZKLGesH/loEkWL5dDp78U9Dod/+65dG
ekioBRgjE10vgXcgU1AowtjXosOFF7q+CkEyvLmc3ehV4oAjTTyDrBtKCnpkG3HR
QI8F4EzVIDlN//1kgZitXojJIAydv1biqjBIIuGbrTqMMCv7RYZaunDH4EfTe22A
IFoEz1beimGChEXD7zZl9tbyC3PGPeVPLJ4nfRWc4r440fL571H8qPimpimfxHWP
CD+hsYSYMc9bNLs8oG0M3DXxQf1DvJlKDi6mhBKMGdhatbgrCkWeEsRPoK9TEcvG
56EEGIA7QvC1zhMxYCnim/F6UTzFXWbuEF6REBvvMiBUwSgzUiZvPBxpP8r5K8Bx
MZ0Qmfi6emxXokPqqa53ZsysIEZ54TZ2Y3UqDbekGcINse+ZUDjHnCKDcQvbpk/w
mDtyRECXubbZ0DBFJ37gcvQ7OWf1s1GZvloXmOmdd1tJBZnM5jvHGlQcr4LWravr
mW97UKFaiTWrl1UrGXnHKDrO3oFVsNtj5FqJJTRwKrajhzHoo0YrVaFWh2SdPWHD
bwGSe/z9kHIw2osHKq7nGOQ+Ya+8E0rpJN04P5ZnVaZTlPs09iJrnzcjpwdPejVx
QbiuMQXdnSiteeWrYT/Dq6DWgoFaTf8f7Yyx2UVNDcczeRvMNI15advmYuY9EtWZ
UeXh0AOHD3M6J9/8PVSZlesZV9OPs4A7DuBsiSZ2o1gWMFiiI68p99ORyh0VE8Z2
hrZfQeTAFZY0bqpyiroWfRBwQ6zWXhhiCn69UKYvOZY98T8p1IR15Z8zX5vY+x87
1R3n9bEnNYRs+ZDd6bYA0f/+idXvDrVlQeIJGq2wC5eJM9yuB+LAtITBQQ5gU/yN
lSbZupLG6CH9FND6dRTStjOQFZKub8sllRChx6xGrGxRGqQnM1LWNoHS6X6yeq3i
dyLkMqcXgI0Uiq29L2UkUPH4JlomC10Ct6xzrmQRvqWQ+cKpB1JUAKa5bR+ATEzE
Pm0IvoUb/ifk0Em9/Jfdydvot+RiFEX2WYR2FECYvGx/qVmqbuit9ApCMF1LRaXn
G6UKuOMgl73L0iuxN+gAi6BP2VfKkq6ElCjCVuWmT0P+VrQuEoQtUOxvPnHCZ7/1
ZGd6aJl4wrpkPzC+GfJWg8dwaJBmutnhckxHpea+At4/qnHE2aGb07a3hXNLr6k5
ZHKhCL1eRNoYnbdGnbuoLsJ8oPGRWXn34UgELLMIUmLUs4oPWTIR6rXWtudRsOT1
r+0cKPz5VaaW/Nri3hJGcHKPEWcUyXOnAtxdjMK+L6pYmiLRTcYiA5d0Yv6O1F9l
EL63effm5kuXUt9Jm2pWmuoZoqHcAX6JOzPRm4S/+ZCSwa1Er+ruF3p5r6pbWSg3
hDMHXk8Uw0RFojJYgVGzdgydMjrOUStwBatzrFGH7K6RTS3/iWsGO9is2joANAXS
X2LM9WZnYc6hRJYOYSCoTip0lmHPPwYhTZTUBj4sJI5m/+X4aMWIZcNCdJhIqrLM
9rVaGj+853os3AuIhJW9a7kV2hNaSzk3m3bgfLO+3MenlsBvA1AAs/j6ATjTkJlP
oXUlRhvKdMbgHzLT+VLQ9StfUh19nnfvxu/tZ1fFWS0tFa5yVib3YEf8JLMNgx8M
JvL+Wfwkc6Qw+put5cve2v/Sv+Ex0q9QykV2pnecF0j8ocduy6xqu0qBhDG5WLcC
4gnFxNDljxdOVxReS5w6+jNsyLU9Wun5aoZst+vF4oeinb7H4V7jkKYn6egwBTYj
kJum6JMkp10fvE1CSDm2iyE0V76ZSdKHeL+XuzWvNIntIEzCFYsnV+01fBWZkPYV
SyMLGAklzp/IISBAnZI80a6gXqI4iFJnUDhZQJs4TtBZFxrmh1zsrYzv3YYwkZCA
EuL1wI/1UDWE0P843DlIjBi2iB8t5O36Np5SC0K4vwsKn0xOthbXMxPSHzxaMNFB
SswlmJHtOIe/yr2cxTypqD8NdcTZBa7ZYD2TSxds4GeW0LnzkDg5mp2KXTFkqEj0
/OhuiMzWWpFu9h/x7G6Aqqt+yw6fOIKqzyphhVkZYEPfQy39KFUk28j2FQZDi0v4
J+yGNIV2HODJAlAHgcyIpIw4V4zvMWc0/CJcMskN1GlOthTwS6StQskmavc7zA/D
YtXXD4eJZar4AgzOfFMbI4R+YGEWdOtyhkxIOdfmC8FdM2cjfe/YXp1hcQJVM2Nw
/J8b6pSw892ygX8W3gTHCkC0usqljYlHCZ2LdgMZYeP3jaZoevD2EwdR1Nx6k5C7
U2wDDZOA3C/VorDFdABz7KQgL3QBUbpBYlNDvL0Dih208Pi2jziufGTibYB9Y1XB
+CpXUA/CooRQP9VscsdkQ9tAY6q+YXY1lkCKG+ogfkHCXfJGHJG4w3kh76fmwAQJ
2KY6UEeQhruEVfjY0ag3hJKEI7OJRg3Lw/RdWwZGaag1nC1gOQQwDNmXOeYDS+j9
hM3Zs+cdTL/7V5UVOCG/Iay/5kHyYYG04t3Db+B/N1pEMA8SJ+CrkHeEEAMOeGwC
5R6cTeXI6PI8Or3CXksuW9a7ZCRNf/aOoQ0ZZx1Frkf8JI1Y4argx48YvV929yof
prohPkC8V3ze9AfSed9ekGgj4PfGFKMGwqPaW55ilVliJ42tNNCNP2+QHn3wgBGj
gdGgI0bAPnAK8XP9ZzUcOy5GWJHz+V3KxDg1RwBjRPpTygLQ3I9usVrUwTqQJjn3
+mp7SepotrGoXNd4zP2/5Y0zIwtNaY+YeZ2vdawITrrubB/ID3hSWwN5CTk0Yq0N
PZUla3DH2pEWNMWbbKQThQoB7re/MqnsUBl4SXOwVCfbw6rxv+9kqMxnqupBsjrE
94kuJVV59ljeYjhAkYmOTAAEbL7K771zOvvLgq3TkNbk4OLwFReMlbRXymrkMfPr
Yrg8sAM1vrqWjLyTjdsMrUb8rKm/IEVY7FKNgdhOUgohX0LmwM/YSanRnAwwLMDF
CdsJKuJ/UR8SUwdirtCy/EHAjigVTEymkyg5E1/Aojf0Lw8M/+p1i/8Tkzn7eJZa
v3Gm5rsp8zeUly9KHDPg7YNuxEyrruweun6mPoIcBEXdurfbVXBWctgnFCn+xj52
1iTu1p3xcCTzsY2a3qSu2p726NP/h4hpngdjeOFymoyX/nyaSDzNTSH5upb42I6D
7trVB/KBY8nmdT80c5L6FXSOVttsr5qpph+qo8Z/TQ7h2OnGCjAuoaU3WQMkCWXN
t6myQO5pVz3s1KTS36OdVlXCNOE9YI8/WkbSjTKiNhAa4khiMU6h9/B9og+s2Cfr
wE09Jxa8jV/t05VxuCMPCpxY2ryKbbZ3DW2QuN+WpxJVTFQbusjIHLeOlP2RzpBm
TyRraDSBZw0NMysayanMaXFwGSTP+zQfO1I7G5mweboJexbSa/8tamdz+MzFwBVt
j0UN9619niH/ym1t2uAmd1kpvPSEdm6ckHQ31Qa6IWMibMGQeBPnX7dMSWZu6R+s
l+CnwmYJWMSciW9kI9DOwzkTdvd/d8dqB3DCR/otMrFNLlIuueCvI5vTN283w+rk
+GdBUBovd61btI7o2PIrug6mIp8M8ynwFEgQLd0e+VePUmNcNq3QKxIw3TF/tTh1
PcEflsrM10lcNWNjpe4bHoAANBFlS9MDYMvC9zwnYDqne/b6IDtzeCMfZBI9OMAH
PmVQPcijbaPnjYMnqKyP2hutfI6bL0SgWwcvOIHgqHgmaAoybxFJbNts4Y7lWkxg
NpLlmbl98ieZiC+PFOholu9+5PFj27V0poi6DQ16ZM8ehG5lBnCo1Fu6wDg+zJkf
Lt6N7ncVPFoHO/k3Ln/GWgA+5RYYKKiMOz5ZjzTxz1k//L/R7geXLxUHxlMOLWlS
lgn6oR+eSKxV03B/hGu27OXq6LlSQ744WrCicQPTphjxnu0/vjkYNB8+3HdIKt7m
l1OuSvd+2zk/sf44kBItMSsornhQjJflPLunSOqn5DDJuz2Ot7csLC90e2l6Zqbb
JKfXdjxPDqPTWActU/T9tc0bGGms+ACBzujQooA8UaSUQ/2ZZtCdQtCyhMsWULs8
mEEbTogZeA258q4LfdSu82NmOhzI3Z5+Se3sKxEgXeWZ2lM/rfrv3vzNjiUuImtG
cZjuSmSe10ZhRS/0ubYSdZA0SDKuyKw324aTmyzBU5FLSVLtnSEDv6TUHa/UNcaJ
nEEvuvD7xg6kI8Dg1/H2kJXwe5A6zu8Msp39diAxwdKC7nPowsMpG8/FqhMqOiTy
y2YcP6rof14tklszQr0iNkcgdsO4kGYkafWLXD6p7ZhaA2so9VvU3hmVjsT+4X8V
7xLiRc0Mci/GSbfVy30Nl4s/meaFE4a/jzlDCx/6GHigyb9bL504mHZqj7BMFVh3
pKwtRkVHDO+kMCTSajDdzDXqgGJT7ygPqq95aVoq4CgTQPkjtQT2fLogBb+KXG5i
DMw5KmmfT/mgoXN0OCRPYctqmbwCgNh/arrlXgSO6DZAexa+OfPtgRYu3fVUYQog
TBYLabeQ2wTL6lhQN8ElZiSifa0ldbSw6Hatmfe1k0dfu1UvTBTSuPfJRNpVmRr0
ZCJYBt6MFHlcmZipSqb8cBYFS0EKN0z/1UXkiP651VrtjHTtCCRoDcDeFconOccd
uix0WK7rr3qRMzeLTMwOej5zt0zpEPTYKq8d3Fqsol92hRqXV7qVQt87Ynbpg3bT
GSebUhdI52S0Oimqj3egR8Cs5CMNOIcprfO78wTSvHCuXQci3eVpPaRK65jg+du2
L7HgM6zLYlKGdpr5gLcCOmkvrQrSgyUBvkBT5LcGTvfVI3sn2xTkRqdSCvtMCszj
sD5/Dm6AVLQfdhq5sYwIQJ0VG0Q2249tA2pCM+k2ebr9buM3Tp3w6wHWaHN0bgcP
GyQ5VdnyWCdoUY/KxLlUYTsvewEZFHN7SxbAOvvCKfquLKQwniFuj0yqPu0PwyaK
pDofftzAAG9y9IDYo4x2Sx0cnK5yf09O30pgPywbzb3TWSOuQqUaN+zyJd6daP1v
o9VsMiwdTSgX9H9DNAIwCijG6JJUmsczxEoo/ok2Q5fvevrSpBWIjw+WywK0esM6
39N8JP3VEJvGULxWqYSBshhujHKAM6G162NzcG86mVbuLfySEl2vgqZneoxc0VCG
LBzkLq5CL9lCPqAwpaoe7rfyo+0loIxjQfLOQDi2NnEMU7fC2p8wRRLadVG9fQyb
PhbeQiTrWZiE7iTWmtu+4wlgLCmSuQL/cTTjtt1XCuv5+A+H2Z3pyRT+AeZV5iJw
yz5sZ/LkzJCbVI7OlzutrVBUa6GoD9eSRYV4H0lRtdwAoVj3ZC+h/ig5hmpHW/5o
Y2lZpYMsVQfThDJoS5gMesA/UfXXJQ0yLJelYgRLdhWprb/ypnbtxG1GAcYjt1iC
XWDV+4w/+566kKz8JUKWwLdZqanhZumKWdrw6rH/LwIprhtCG8gscaOO1ehuxmMK
W3wknF2WozNIfrAw1+2GFhVQNYvYGd+vi9FO5v+u7bhujmYzUgvySNM4bZ+hkkIL
6jBrhpO9Nphv8soOzXkRxCPerSgKBwFflxnm76J885T8ZbmsVaF3G0qOEx+zjB/3
KqseN70zPOVFzUtUSxTB2O/MLCEWxEn3RqRAJCgHV1LBnHY0cgDnAWzNdwFF7HR0
4ztQjgfJWesEUMQLf3DhIjtSZOW99fTygDQhMXpG8sEX3pmxCeyYNWQoflimMEGO
KtjGJazEt9oH5h9Hn4iJa9YczfsmibwdDJExL5oXLZ2/MgbMMv0JUJG4E+VxFzWT
BH6bRkT822uCrJP6iBwLlJeV+WLz5qnFs6G7X+sefJ7tQhbzOezCcyuFgDv26uvg
dU1RjsZ0mBT/BL2/LSorjMhFlcmDF6l1msm9tyJEq+EcejpUFE9EXbenduBgmznj
/6AhTvxZXi2yVkGln4359EHCLQ3WhctyUF3GVs9XdPMPHppO0bnXC9HUQCnoB6kN
fZUNrVvkISp6ISYCdlwP5BDi6jgc84x0BVVYwSezF9Vd7INSkk/IyUH8yTXqH0fp
W2SpaoykyOH3zdSwajEsGMrPAxZK13XNzEx2baPCIgk1iCv2JpqSxkEbGWVXNp1b
zIwP6UwK1RN7QZWzPH+cSH+PWOc3/OTqiWE4LW0psVjVuwF5PmY73RB8t32mqtBh
JZ3Myl/N6S7gVKAV87o0LJpMUYSowLDOg4HysyGVeg+ZoSE9vPjy/y26qx3iBjiq
Vwk2oy8J/uvnoYpO0KZdIpLYSrWHZ9nJD3SPqCM+ju4/55pCw7wjdK1qGZFtvk09
pXhIgOGZI+fzMhrLtnSukKNQWwBG7I8LFD+eggFMGKhIBV8WRNKA+C5e5ogWRGex
viE4axR8BTLAUlJhRA28HAIihgEW6wbhVckkwwbej7WJk8Yd1e0nEsvsttW8CHNN
ONQk4neILWpH84YMI/c5123NT74qnKfbyoSt8GDHEWYzqT74lVYUwv4y5mYL+xr2
7pWw3NYdRtZIyT7FYySlLg/Nb7QVeZzMEUzxHoL8DBNi3ArruVk/w+oh1sKOwoW9
LovtTKg4FklkIR6nQUpWs4w2seRbsz/Hwg5x3XLPjl4YEaAGzUGCCflusU4/on25
WHY8DARpm6fILinesNzlxBcu+Aqr0rRqXyDZj7WFP+0hv2sau3Jre5HXtc+f3rbL
R8cSjmuNVMAsug9VAdoj1kaW3Pb4HvjNimF7P5gENOYycYd/2EL69ln7USsnsY1x
uHdhhwdMtHauY4OXl2xFHFb20DQsN9XTUckc2JYpi9htm2BMm6/GtA4YlS6k5sf0
tU4LZZWM/NE4f6aq178VolFTUNUNEgTmXvyrKiIo3LAIGlK3C5enx9Ij8U4tNE+r
JVNWU2rS0BVUEuwCyEthAGGrTo3F9LhCevVRj8QjQjG4HD1YKRBlQOpSkKIOrtcM
L/UNS8pOM86f3cOGgPYV+cDAfm2qiVZar3wFhEl5y5Qe971uOYG0RRwhllA8ux8Q
qIifJk5v7AwBCux6k5G89VMiOG7At/TyTohWt2ZbA6EQZuKrxecVjL4Wlt/JaNlb
pAk9Ka6b6VFvfC4AaumgPK5O47ovvibYXmfXaDeWoQwQgKMdGuABA3U4AATDLUxP
MVsOI0KEr3fbjx/Zru6CQBiuY0R1VleHH2uFke9ut9clecfXTEBohZGM2zMIMBWC
dym0zxj8PhJxX90/hg5dg9+Go3moPKRR5Twmb9F7qPvcu/9fR6SE8DEYK6aToJ65
PDzXx2kRn6NkhxzlKaDRgJgxfgYwvtMNZeoJjncqX6AYxIpaeBwt2DtUxIWKHyiq
kWfudPpIAcOK0RSs5PNGTXTFVM+7HVusuJ591gLl/Ac0UL4m7CKaoRbAkdVKpRis
81DuVH16TtXiu7G8FmhA0fQyDA4ZymMZ/9PdNMUtRN5Pw4mgZJM0+qkn2wcnQANw
BqUtw4BO5vllgBshu0sX2NpAwY/5mPqBJxIK2eyyUAcYT+YKXk21qbHajbV3xpOS
c4Mq8zzV+UjQ8Hn5B3bngyM/ec+fIuc+dwBWfBiDasu47YC/TlYqw13/XgQ/0n5i
HqVAFxZ3Sv9ELmWy0i6oIdZfMyKaMfTUpe9vU+7Y/mCV3tZD+bRiYpk20+kBTv6h
elbOWKw5UPCTdpO4d0pBhv2gYk98S1GYnSHBarb5yMXoJdWjLssd9AQnXZvP0EJr
vqvjJpjP8Vtm1bJopGVXkT7+gH31TIy8nTZVGpOrQSMqLwy8fg9pdddfZ7NKvYfH
PoHtaf70Zj69HcC0UD0ZK7wQ73fbrPbCi24Q5DxJXsvEyKaTu2x1rTrSPZel82Rd
g1cheEKLO0Vhi0V+jsVj+37VFpRkT6gvEcN0ssoKK4V5t9qpSQQAAigimMewPo6s
VXEkFXz+nQt2LSXQTwCA19+cziin/kmcR3iHQmIP2QgLKQAOaUBMazq6ihBI3LZ8
zeMWxex89KrkiRxUZLOo5SVeifiWjnM9+LLw5DffZLvYckxmo0c3mMz8ZWP4Q7Ls
1to1fu71p8+OpQlp2XQRNqs8PYGEx1+uV6zU6NpwS94u+6qw94xBYRbrJm3r5y69
Bu40n9JfTPqck2VJ36TVYA/MFfcOLOy/60CXFDuQnGy/iHgMjYSZ6jUE8fxZ8czN
hhrHWeuiQdBhnihWUU5XVnh9adJLWma/PdGTvqWj7dQkTIxsAFa8F/HbIw1gwx94
/Y9zbi780+0ysCwnnMfdOczi4IJopK+n+nW6OvidA5oj0GamfQABLKKHOLcjRBQ3
Vtk2S1uCCYx89n9W57JwDzEv/V0VeYTpTVD7raRuTV08qoTw3yslas+8B/cTkg+K
oiRqInS+GDaXFuVjHnuyIxlF6ttrPyr50fy4IixKASWHslNWNbwBIfAKxlBK8eGo
eDBDqDOUQz4y3zkplb+3zuC1WeJpaXgxVVHfUKPPvVQX5UL7X3SY+KDQdaaY18yh
gNqa9LKt1D+RTDrdxvyvgSKUQvMo6sx2/ZttZvq8arUstcZ7WwgQZ8U4VNU8qjr/
vStv9Tsx+Z37+p3tLl6v9I6Z5/BLQFMMkAaHModMIKhyBRiXKcP7yJd3ts5bsbsL
HKMiO+IN342WnOLeF+LzTZpYRGh3o0grlOYaKegJK9qwUZxu9D6lNGw0lR8aBgPm
BU/h9BAjVmDGre7BcMYjZt2z4OCJto+6gr8teMsj1GUWZwnIHq5psNBDzIXdU4Gk
Bs4U+rsesy/+h4XeMiKzQU49efCWMI53nRgfRrkGIyleHjAdyWVxomtpXU2zY3UX
LM/h5pBUlSjB8Dsg8cbRthuQFz5C141wTRIhu6L6j9r1Eo+I5jfEMzRzPfqKZN26
YhmhKgeMD88EBlqvU+FC96ByCUXo7GxB/r6plheLe5YGHLQKLl8eR8l3ZrPtygkL
FYS+MIkd/SB0rPeTJjGDCGzHh78+699FAPy7IidBBq8lyyc7NlVdMRcLYRi+14Bc
zeRezKL0QoZQzD6cIKUu+y2z9zJDYCuZIZok/1FWO1feNMOhBqY8zPJ+ItA5OaNJ
gdjTvaLmOm8lbti6TW5x8vSwt4ipxwU3jyHUehEZUfXBVvFRNOglKGqPAZLj6gzh
82zvOhT5xAlwE1K6th/tvOcddbtOftBJn3FAqBcjsT8hzKr77/fiYWWLvsPbHVUd
n6i5TMngYcBZ8WgeCBw3y0O3dDamAf+6KuOsN0i2zwEhVpp8iclp/UZgmMmoyLih
8jN0lZrsNBbHGpZR07YQZKIk9iWgoUc7wDP0z3nf/ZLGOsWj0nvf94ZUUQC6B15X
igz9MephkU/XwXAQYxkk7hdhzv84xoWkN+3HlffmwuyqT5b+C3dH2DfPX+R9cmFK
QeVFdqKRGfYwPqfPEfotrFKX0xNVfiuUHgThUSLxtzcfYMryu3gFvwbzRNAzKFOX
CgCmIPY2+xotSkXo8Iq4JCGNNJlH2tRi3S1ZLZbcgsl1VEGcSoKU6q5Wegp+zMS8
kqhE1czfIMPc1Mh1yWDX4Ob0EDkY0wfJrW9UoEYIh6BlBWdkjiJY7LfTQE3X1Ghg
F5JJOrlMlkmnj0SCa4IuSQ3wuGSRKwwNDCCfI81Z3U6q7FBzR1yjjl/vmocV5gBs
T4LxqSpcGplJ2cnzgWbSsbf3UZfScUGPG9DmJkoglvv0NHuMp8k8WWXIknuCT+hq
K2/hGCTTUB3CwCFqRQh0AkNXz+n6TxT3dN9WMOYWsAiy8TuWLz46h9mPK+wkSMSj
57sk75F4sCdXaB/QtneqJ5VOT/KU4UPi/Hl8glQZO52Knh55VanzEr2uebJ6tOiN
z09gifkcvo0yZBUCeaV7CbFxPoI3n3dhdpeqdvXMxOUTfv4klYlFP/YxqtA682QY
V/nwNQpTakB6Hk9i3czZ7GPBY30EA8ungywlTfqINu6CfbMXMfnj/UFow8BLPLp9
viJMsiEXSdM3rusYKjrsLVTg0Oj8sLGc/E7G5WliVG5g+TrCr4+KbcxRt/K8j8rP
QUQm+JJWZcBq8MAbq+27U1728iIbPS3Vs/0JEPtD7cygsfmPRU2ObFmqlTeje3XJ
O3nkKXAn78NJiiXi8caEeZj60w8+DNkEDCvcmklp116v3b5qPMHPfC9F8VTm9Zbv
cCN44yDhtvaBQfQ5coohuVLactzATCovJKXYxuj9+bC3uUpOQOB31kSkjXjoBU47
SqsjdyUNmYgJB8KMq119kvtt2EWP9+Ah36NCskMT6LkWq/GNo+v3wJsF34Ti36DT
2lLPRkpOu7QpmXXKWJf0Gmf8DW0N8/xJEXMe+cCiJe1i5o6TEVKSG7rOsR2w4zxI
tyXh2M3B0HJ8TGPTCkLua7bqwHIFR6I25JdO781bNRz/+jbzL4pA4Jh1vzRDXI97
nvtE0WSHOQ0FUL5zQbYMNJDjT0srkTpaywGB8FkzZAZf1xVq++1/OnX+8xCDH93s
KIQArbuC+QoHfrqn6+91eT+h1xozXNfZ+LhSKXf9USB2rPImePQ7xMDiRwVT2/r/
IBcFqqpoQOX8tpIWH7qQfU/IoH87Q19QeW0Vl/5qi9gStfnkhYVeojMnGEKS9Dl2
1wrDOfF2qOiDoPlWfLfRkixQCeGchhg6bxdzoGZwSKHLvuhFZ8C2o9Krth+3YZdw
m18Acv9q3mTCDI3+3nkCbgXmi3OJdkoWBeMcJXepsAkj7b2kziSMNXD10h1N6HjH
HfX41Q1gIOrwAUkY3k6mcaH/UMTWIo58GbBFkpIEorc9v2J8YSaOq2rtN4KRL15I
yepB+k5ksH5C9vBxDfDziqf1cdyT7ioQJ4VIsMWUlMsf+MXn9i5hs+phlkVCbGto
LHYFiWrTdJtcws+kQiix+J+9i1z/JSzzI4x2/2iQaKZLon2DTgtEMBPjgCive57V
TAtwWzHx76C1ml1SkoJ3xfcaiOJV7VVfZ8Hd6oy537V2vso+/QHdxXXe8T8aBbh5
uGmgILOaTd53Z6ghANj+vq+rD8awGL9UY3wQPH0bZAs6KMXHtcEzXrqesBivQw5G
T0HPyBZV/mBNpEULqCB8XG9weemB6Xz01UXudBYWmhwicxUWk3wadHk/QM+99aV9
S/5UmMZbtj7ygoyj+FzTUTxnwY+UCBD1In4YXFbya4TO8mpnvIUw9egOmBdindfM
5BIzD7oMp84Y5fpyGtwGlb7ei9sEhRCJWE9Gg9YobfhVI7QlXiFecNcWqTzHEiQ3
F3n2rD3fTAkLvWmKb51CUbaQcRIigxvN9NAkVykTuua18oFxmWwjTOlcuaJZlXuL
YC++BoU6XvLQqMKxIKOYe8HD1yML07goYFkrClKXT2b7WAXCiwqjxOCbgAtQyho6
2VlTlLI3tYNL672fuOCiOfdggKFqFZ/DTWDjjCEfuZ8zzeGaJbqhT/UbrWtx7aBW
5pSZbJqUSCVVXdxA/+/yVZAHFOup/PhU62nv0nuHkmwkPk2S8FVnRb+X3xjg3T66
BGJsGXjHjG7otKeKlrXtHqH9XbWAWN3OQxeWplzrKIe/Rl4sKucvqe1z6E4FEOML
v3RJWTcNNjiwt9tQTyvcC0BCMu5QxyOx4now0BmoWS3RgY5ZNsrfCWVyi4PptEjM
h3/1i9PpdaPjg/y1xcgsA7onOKCLwX9+3EVtCqI/TGeov+nvdKk4glFUxD0OTORh
OLEUgWLFUVXEiAYgMYagJJXcy7qB4RTwHDBP5VUMFj3W/uBdVE5T11a+NifnyrFQ
vfiSK0GAqevj+RvxzGg4/2tk3ijxSaEo7QdKA659tqCVaOSVKyeasKm43pCLkjlI
aGSGv1UfUC+oZcwSebA55XijRusBaKrmsy5OH10Uo011VZ2YcReLi+Lpw06ypxTW
arobAHTROHn2WqS+ypk7GIHHrOjpN6HSaXOon+EztOMGiPSj27A9rwOj2uAtg3Kr
GAt9vf3Ikzxrnmwet9oCxvzH4OahhB8wqYXEUuQQ2bO5xBV4bh9Jg5ygAr/5xYjX
nz6g1ukosZ0pZL2vUasBmfe51hL5W/qORBYtJwuxf/g6IBn4Frz33ftmqh1hUcCi
oL1Ko8wjYTf+MPv7Ejr4YhvCnNsoC94wx1IUwhKZ79lEZMtif0iP+4JpQxYxbKba
5SSqh4pkz0lhULIP+Cg+PxhQm/9+an42iOKuwXI5wc9vwIZlQf9ROUV82RLrU6Xh
jvArL5NLE4vsJ2/vo9VZNV9ITis97+JUY6WsbqwmYp4ATwFE8ZlkOix9HnPyhP/K
tbFJM6aM9bVC+RmGElkOqUQiFVNRZSxeEXK0+uFjCcrIphbxzwb0F0eBHbQjrtZV
eA/mDKYX/Zw9wkYwi0Ol9TFx9Hbp5rSqob6mp0wjj5DWGa4fp7cmuJkzsUonGlde
EK8zdwkIes9hW0kevEVPLKUKcvbeS820f8+33KvG4AcS8lR2kQ2IBj02gAY6BybJ
HOwlIYx3NkcHc3rIcJbtBHh0QOaOcg5lhGLjr9f43y2IV6Yh+d7KzTQcLTeeQPnl
iOCIjZpdIObHZcGJODvgyrk2jfOxesxG5N5O3egCZFR/hRl4jEIMCWtACnhiKX5G
TSZKwIZoTqbsf9YxpCBmhyEKXr708ceS4FjiFXww3RpUJ7M4RDVczUWl1QhjcJ21
zw9dLwDFkaAhc8RhBF3pJeYE6/1I7V58ZMF+q2BCre455s103wv0m3YPJDvWeBvc
R3V1TzGnuasrjv4ApicAPQ1CVl+H5gLo5UqWYStGAlRgBeTfSBpdG1GW64C0KI7i
kI9/y5mPA5FhFGFWLqAph9wSLymX/KTKiAVxAVl9w1WIfbk26gg0vv1neKtD62m+
Gqp3kSE7zhRNnYqmlDvQSQdEXxnB0dyOj6ckfgY3TKfPA326EkfnNnkotHInNqXr
irmoyQFkVXqlLEtX9n+9+xdbb57Rpxx+21vHROzZfICocLheUZCd2OKTQBiSO9eR
rdUz0JjKYhYs5bDl326ZhWkkP+DrJbTblziKr2o9i4LiWRjT87Foz/6AyQvdDwyC
P+tzm7KJBTDkhMrkVEX3x4PW3yVxYi82jv3XHBHtYhAaNNR+v1oEH/ec9Fxit4eE
feXqakOoSC6Veaydu1RkZHYozheEPWOndsma/BJmPFPY1j+gLbXMSw6gZom8rljF
1S+XndG1Vve0T/PI64sUscmB1YUNANFXLqupMqpEKJNldVGORqCZnL7328JGHb/p
uPSDfnYzwDoVIih0+MEE89uedFMYFX0qOGk0rLzzJKJsQ1MYcQrqLi7ueAPOeHtQ
9dYDGdKhwAV99wp9sqMi9sBI/I6iKkA5DYG2BdpetzDFhsdfsdXGjhbjCeLkSQa0
PNrm7ok2AUxrwp64i6ePlGEuT3NhRaMidPVZBY7J87eEZnXB3DcAxLQRHoK8RR9p
7hJlYKMFq59vPpHCMTr2XyZrZCj9XyDkNzzRSNslcYCrkt6CrDPbeirMiJvjlIYY
I8K0VBoW/YJhhnxDzJ8cOR5rVBoiu/HIWY/hU3vQBWX6Ypeh5vAMxIFUst1wqNud
6SmFNpaTlpLCuEBqvkZC8Um9AELju2kkxJS4HjF4LXRbKFEMf/1zpjCe/P4jO2oB
UNLmAidYMF0iyIw7d/vA9hZRmRo3OVt12R5UaGeaw9ZMridpzwwDkfhuo10o6M/p
U/fsPXcweFYk0nFBjPQN+sKnCDfZBWCL4ag7K07RHz6UG0o9jThzUJxFASVbZ0eF
5izpJS9uVUfr593sLNfkgPIzVs/W/kQCRcBbbMNCd/yzzSdqeIZ+HluliS7vjxz+
ug57qBOHqt4Sxr6F8kUm3A3wPdYQbdMClcndO5yR2gVTTaMEou2l0w9QjuqPEsAZ
cQN83RcBHFL9wFDrAQWLCt+CaLY1nln1JFfuavlUiuNo6Dq8lf4FWWNJ09oalaFk
J3UGiQ6vpSXfKX6/z1yXvrB01cdRD2QLlYSGPU9hxfQ/zjgjniABytB0XCpQdiA6
JSkcTRSbhEL/IMuGxxDktV1yIquFtLuleSnN2tcbJcCq6uVw019If3o5zPL3KDfl
MBdaLZrr0caywW2Ld9QN82NC37XUogBQpAhMH0qUETETMuere2mf05PlxPYbHILK
G1gb1rwb41MiY1mpkTgf7BLW7ZcONx1Zrz7Lh6FeL3VKCwewe4NDSeop4J7KbwR4
O7FkS0OL6gGn9AWa06AWt39iHIOh83Cej1dfG2yQDxlA4V/atCrVzh/m9RytmC0l
6qaTthn5pHHwgIScgLXtK6sT5uhXp7w32Id2Hkvkm9vZuJQWvGKzA3ltXyfhVdAN
vJf28v5JjOek/0+aV6OhT/vFQ0s+xFi50PdGZk8CEQdQOMnoCPIDctozu4XyDWtE
Q1+F+FgIf1bBe307dIIkDAj2xpL8UG4/DkILR2DrLOtxNs3wVAR+i/c4eBkq2VAb
jZlvkeo308eNPguVEN7yAMor1TcgaS19uxFdfVrRs1PqSTim+pS/XdrikA4tqLDh
eenQqNva/AwPshUJJTQxtPzFgEY0xMlvgVjDGwHV1shVazgwL+qqkkueGxmH5zlZ
uXGEGjFviEObwiBVGIBpYlJFslUraSSZoMA9PY4gn/eq5tqP9T9Lfd1EQh6kEcp7
Ek8qdW7w84uE0NZVazJGA5RuDG9KmLE/4Z1x3KExqhQRGjTMSZEqaS1rpfAjFj/A
+qmeYSp7l6TGXA171Hv/1laOLIwLDn5IPWMLLX3dwNzOVly2SpkVq8OHOhFidP54
dvRP4J5zxPpmVh4XQdD6Cy0KrSqqAFmgaJOnVF/ul0HZDNa3omIjMFzobawMnIci
AmT3LEEgdWj9lKZGnLTJVxTrO0JIBJQs0EgEHcYDlqBsvyraY2/lKP83zaTEXHiY
ApZbxhNPWIPZCV5LqWY57N4GoAhEp1+/DJ9irYoveUlcD6/wbYcWQQkUe8Uf5NCO
L0jTkxNToP5rR9n7VxHYz/A5dspxyuTgvlATGXQ1E5nA+a4uvITGhR+Wvy7101+l
EtbTSgea1ZTjXzMTCvHQzFF2CFTSqfZhf8jMK0M/wgHMwwoqsIV0R+v+4LrnCn7I
hkuyjcX4QUfEH9Tm+W8BTNjNDFK8rUduB8imYrnEH8bGddR6XZ1nN5vI4bcjQad9
ObzqGmPXxqeonxzzUQEe4873ethwdCrZU8qyJozTQ41jsNwPu6oHn18doGub4yiy
82EoLMiS67vv6Y+zfgJZa3dDMva760OElebAaHi8i/FbKrFOEp/89Jz/sJg/kN4i
aTneSDBi5g3U0fYfnMcOjDNuy/Lnvc4q0ixc3u8joOjRqcqRlI6OV7br1KCTSC1e
47KbSRqh90Fn4XFL5mre5uYLsRWyaLH1PZFE/2+lkhhYNdR9t3aX9XTyjYA3nNeg
L9NPVBTt5v8OCwmTyHQkqAyIgy5hzi4s/CWa0AWApmkYbH3dsm4Rb9Y5Ga1uJNc2
x8Sf/c/Ye6zTZohwqMVTllH+YanlCwQTfcMEWU1NWPVefAq0+vIyFLbVPfx8gS62
/qFk4+1R3mSgcsG3BGftrwwJ7J55fm+d1sYkVyK5L1XvU4/L3esaypjIPnjMTw7h
GAdGKLmRxHLWB/JDgczPf6fgxXLkUOMrz8wdu2N3NrJoxn1ZrSQroE+bhdVrlxGw
6AQ/ZepTjlU9gRf/5v8i5mHOMiUrZBgpmtm3y/NXNvLDCFZqO/ngXD+yVwdk10t9
nsgbMy20yNU+NqKoZoIIKTNbHIdS1nCTXx6IjsHfb6tpZLonjquz56LSkA3OTD0e
8z79NodS0N4exE5Yh4S0NGPAPnD9WaIOaR1yX3I1NXIhDqTJKJYBu7hGgV8SkSSk
zvCCTUJMX7Ph7Qw/Kml1bML9XErgDfHgwWhUe0w2XgiWOCjrGMvsp1w1XlwX4IM1
9qK6sBH2a6YWNyEtuP7rirqsyFIniSEhE2BMDfGTxBFwGFVwoiFBQYqCgOp4meb8
a2uHpCxTyYel75YCu6rZDUbXVTg6QGJ75F55xUsTmfeKQXsj5jjOX+Q0a84E611k
ZOM+WtEoYdWKt4wHb4sb0FtGbpWQYdftr7JYpgZe530ao7G9aNY0uEP0UUGapzby
5zh2Sh94n4HmUMQNmmOjezy05H4F37P5nkwlZSzrPJWkItfJseqXeFAQ68KHovAe
JbYaFxWwxxDh/paCzhlm/CNd9kzW8DOFyzRMOGnAAQJfFLLDB9MGVFwugHxjPlX7
QR+h2QG4RkwPI+7nrghbxgGYzn8TF3fODRWnJS2q+g0wzbUEW2iCeEbM7Vvi03GS
WryxcZ2Dxohy5aorObQYIyV6dbm0GdB37XCPiEH/82xYM1Auofoa8J7NSTJkjaXE
jycNGT77vuHDogllR6TM9mWSD2WbdUVhnlnNy3TYUF7LfOoeNwNO7cKqW3PDBAIC
W5eVIyFQVQX/qCsRUrrVYP3MCIOyayMp1GwlhSMf6ShV95QcSXErsNIYzBgfCIDt
/BbUYGlQa0U1R0dqiU+TrACUkhuvpH0WVQjYN3WeTgf9v3O2pBRnPZRP/NCqmjcX
yO9kRO465HggaYNiYg6KfJxoPF2hFFA8EHqH2+SGlIbCVyszgWi0i+xMqA4iKxJG
8Cxp0uLcJMzhVXaXI6HvFIJgLpvgR0Cjqr9o3J0nbavYO3Q0M8rKsL94Hkc/p91Y
okADAui5WOzaTuR57uGfvHt2h+wELiog8WB5EmFWxpL1q3Kx0sSpc/y8zOWgIFrp
71Ak0AScyWyZclqGdSetRcYpxtog2M8vokqsBHGTS+YYXQFlmihTyQ+/itKCStMu
wlrgOmVNab7MhAwxZMwvZmunLEMv7zeTSExDmQJIs7UzInm8K9J6FHZuFhBuJRHZ
izOn9jCcsRY/a2qfD3teRaGtR8ua+pD1RB/bkxu9TPaSBYcsj1WTEGKcefFzERaC
izXF1hdSP8Y6yzNCxanmCo5XU1RWeJS7Qg6oatH+4nqDnlUE+Ba/cIYfGU/5csDV
FvQVI9745kyf28ZSG7iVMaFN818dBBLkNe+sxOzD+PjVWcD47vR2/FxDNkLHfqJQ
+J3cENc4wdCzJpvl0Kf+FnF39TK/f8RdLk0P389rjlF7ZITTgdp0Yhio91iXDldZ
uVkFz4+e0No3Iv/FmHzZ3ls8NdZ1H7S0WzhxDPyS1SJj9JiU0XyThU2D6PExBhI8
EcBR6f9q2QFzWDd/SrmQhGWHjihU5fF6bNxYOKDUmWJncMLwiaWayuxai3IULUR5
+Q1k4fcvuJCQ0HdgWmJkQKK5ZvxdcH5nByGhWpddYjw9322/THiIMRdy74F++J07
t2wR3nRWe0xOG1am/K7wjZW92ko44rUw/CgRqRhwcjH20qWSaiD6kIZuQM8dU+yK
SBvkQGWJaDOYavpja5aQiOd8Y4BbLfpvDlvBXw0WTWGd4ieo/8Goc/29SxFeejb8
kLkTdAG/8PrPXeUXWhhTFF3RieUnGj7PZSgQeCXHfd8B1B/Ac7IdISYqiTaoZB3i
VzI61rH8aVMCHNIJtdmfJ9FYhuzaGrt/ZzSHOUp/gxamOLwgwLwd9Xd2PjOSxdwE
t7wR8yz6LwAkxpQ6bDDj5C6EIBmOyS3Lj5RjZSToyYt9o28m0qxIAigO0xaH5LjT
zNabO7Wg81tXUMm3dJqnBI/6XOhQUzDVsqL0xlg/EMZmi9FP+52rmtRuUV3uBnT2
PuqXDG/5XJJgKbkh2qWulxtEnImlKpkwb4dv0Ia/Nwb37/7udLhRfi4Qsmq+aWcI
NAV2p3SsDp4hORaLcRD7Hx1EzWjNDCG0gbtFCDdNeTTTnCsEDGQzPQiC/GuUmm4U
iSvC3T7eA/59pORzp2X1BQVTiM8GbHBOvKhc6SVYTho9gNhUgZETD2EbOPTBdAch
rzU+5L+RwbEu/L+fEOQkZRUFM2JsjOnfJpBjtZauXOw7iwfHP9MI4D1MKfiQjjcP
9SLtSWpRQtM0SB6/fSHLOfBJAOb1r/5okJRlM29hmKWa7cfK1vyseMvnO/IzuMub
8CiV9dtanubtcAMt75n9UTdW93n8wsNcsiMFWPAD7hj0xrX+mXO+e1JEsysZMLRt
RMbd0JWsePjkLBpF/m1pLP6bx4++TIxI8124Eh99S2tNUsaPkGXLzW9ZkR7QDKDb
KuP8eKNpWEz2NyxIuq60xeJCAYeVkXy7fTZ1Ty75oDnxuD9LfPMO05Lmjf0PQ/k4
JzXeGRyBY1KgbCOBL5pByTgpio9E52lLS8mcSmySwDoQGMSnkJ3SxybZvCbCuqOg
N7Fnmqy4BPdmMxeyKJo05VVkmLtONZeBj+jvtxlCBsik+cHwt5eY6B2L4xBwWMk7
qFjJfywTkAa5rUT4TtXn2tiPB3KOiHIayR08EBrtAJ1CzcA37H5fgxekbf/HX3Ba
qq+32GxiX8goM0Lbr3QtYuwFS6Ny+ZhPz5w0mkFC6OupwpfKc3QsylpwNhT8ddts
0KRmk2BeBhrP6JZdaiWcTt0D5H+7bdjtg5c4ZAcmzuer4kcMnofLkK8PToHL9hse
/zKpnCBo28iGygUzsvyFbiR+y3qoJoeCbkeA+rTldaPnElWUenX4ASLki+qXCU3Z
d4oD0eHJlbzGN5UGi+slNH4qc1vu+n18T2JCAiLjG6siCj61GOSbzFvuKSimhBim
w+jd/exTCMOB4+0sqWh1axi9BTNgCo9WFJDiR+jvRtvZLcw6Ymg/mhZqQdD2qsus
U9KmCGj2KxMLjwNNBTcJZ+kn8R8iBHnymJIEdKdkgVvEAyjwufhVqDYfJ/ErnYfu
FbRwNpWqcejHAwP6axjP0+fEQYC/J7hZ2Rs6APpY16ZoYesBz/L509GA//QmmV0a
MWpmyySowCTcM4u4iJdu2ZWldZSN4yB5leEMrirA1aKW8kGv/uh4uB3CSFUk4JYp
/oQ1XpuxfmuwRTvYCxeZh2wIQo2lNT2/u82SYWmDBlkpzdKf4tknGL040zhMvvGr
yykLrUZyXVMJTBfgpdjkpA3YG83ycY9LFGclAsvz5Jzip6J5qHMYNlEmWd12aJoG
0/FZB+C2shIJZDscOGorXGkmC0ZlaeNUyk2QguUrqmdz2iTGixN2wfuA22B/jWsY
OpaV0jo/I3lls/9gB0fmJXcumGxbdAHeBO65Sd1wSD7k1i0rpg1inGxIOKaIGxaq
UjVcTOZqneBhOyLD/TMborlUwWhUNCKzkgvbcuDsFz7tpWJH5D5ZvWoXw0zvH3Jg
Ynpy1jYtSubwrm+QD1GtH1lb1MUUMYQ8ivN7g7BjvXwb5dt43g+PuDNSD9tkwLs0
4raXwhGZvc76nRzFcaqt+Fg7qf5fyEHXCjeGXr0TgQqWVUWyDzaKDf+HpXX4lgze
4cOZvqnmx58B9FXnT/O9YbW+Fb93gSs1SzYlEe7z4FcvS8JMQjByJJ4fbzLPbv14
XGuJvAGnmIM/kXaugvy+l0lPFJcLzkChiX5UWMmHuFmyrqjTEl7hfWX0MH0Vsib/
bumpTBWCisjZFkMoDwb/zPYD7s2pIEVAFS70HvqM2Pzarkfqxl9vSk5sd5hhHnRi
UaZIguTGMgUGw5KOFZBGl9ZWEUiWXXQanLT+aSnalxJS++oT+kE5AFFIZ6f6UP2D
MgHUPOiIs4dtNNdT1R0olDcBCi6l+BEFCiPgQWxVM8z4AwV9urqy80vRmPuxo95r
jamM9A6YGgZIzDSj6KZhWR8SXB78xtyVv3Wr9iTI8NgFHdjeaYUzeSl9vd9e9yDR
hR01ukIlAVrcZJMERgcByoACRYrimn4O8ARo39fePN1mSyGHij73pvBlXOZh7k5A
jyjvY1t86fYmHHDlrWyHUQpam4bvjhQr3hH/hCl9gat5LJCblu75g0AEZta7+wZi
oZc+t6aY4kfKKIWkz6PcwPhQbLirlkXPQpLEvvU+d0PpW/j/TF7CB430mGxsTI3d
nxlrjxz+l6fz/0GpbM+4IAMhX4tfS53BcyKKPaeqQmONS9N11QloJZL/YF5d80W6
R+jJURcQ5xv2GyCDONQ8H4viS4K6woV5zwqTwqp1P1SEo2HOTueql8BMSUXdrw8n
yPa4ytuLzfZ6FI/zgDdIrNuXlHiQC/0K8m4gNZQWWh6OMhfvRhm+QgJ/ncCCZfrE
UjSBcd0G/bacRZkOWRvU2hghfE7YURtFPNs4xzBLMqRl5c0p+9W8SohXbLNe1u+M
9TKefPhpekNe5IdUBiO9Hr45FkN6i3WiaQTE9ekiy1WwMJFrq2QxfuCE60VVG7EU
3x1PUTz28jLVUz4tdfTfP8WBpa+gBQ2oQoIALnteFVsGmzm1ZWz1hd23/vOD0xlp
wuDwAlWWBX25+ELQfaoVoIoO6EbziFTL6UjxYjTbF+zf+fFYLLlxUlWR3h3jLVWg
6Mvcc/CSHgOcP7yxu2P19UDErjAZW+hSMLeES8q43roEnx4la06C0rbbRK8lKCRR
qlixVoLkgUSZ5RNBvm1oWTqZAyhcwNS7eLymTRZTs9peq/gf5akxbpp0qFWLzefp
5YG3p90G9xB3qINlA9RJK3tBo2SNtNW7l0DlFfEU/VlTlVMM2VXPhsIHM4s5OLfm
85uaTD1IrYJERHUJa7W9vT7FbR/6wMn6FOerslkrUuEobHzJ0/8IZI0MapTInjHQ
f1DBYgLQXsdLPQml/mfWNUaUy7ldliCAUrZbhe2BFXx81HSGjEyfZPvtlgvLsM+E
PSE6iof6cKkWKo6VDp7hV8tYJdu4Po5AAwEUqMGiY14WJRlaIwtU20C7SakjKFb6
HkxQgvJEG5Y5wuQcu5FVRXxAtAobZuzqZNdmhl5XadTDGHDHptn2Ehry+TLqmL2O
LXdNdG+PLsGzzcOIWqGNCA2jdItyNiJIkTmuPqUzmbhsWU4uGjVdMaGIQdVDQ/92
MM1dBo/LevkdpIxYNTimEokSJvgt1gTf7eM7lr5Nxyzm7gOATyMoWJDLX/VYHzZr
ZocdgqLWFR1MIvke8T7I+55WHEhmVt0+6f7FfcdrQtvJk4KbNiHv39psZY138Rdr
PlXmwAxEqlTiYaKK/Pr5dyPdx0qzWv30CEBcSvJlEaxGatfnzuz4dqPf7qDipzPf
24LoYPk6aBruzLokZPqTNquK3ReL4l1RI/KWywhj60wYFPScEpreQBoiOAHba5Cl
nFsrYbRFvApqf9eGQqxaGQTnil5MnZECFRgJWaOM2EC0kj+mZNgTGh4zVRoxt5VR
UT+CbJZp/t/x4wF/GXnrPeq044PDsnxV1MMDdRE966/jI9D1HsBSJil72HFjfFal
m8jLlVbCvfBofc4O/Scym3WCcJiXjTV3DOhQcBkA5MYLo2TqteonsgDJ+NE5Bebd
JszGjQj9AP8PfnmaKLY60wQhxv7JSi3/2Qq73v/UoAiujLCmlB0Y/n+O0Bmt3f7v
g58pzPlmpUkOvT1SJqvsSt4kBSeNsa2knyXnEfN1nP6B/i5PsG9ErupWfhBm3eYY
5OFA6Zh5Q0ruabMU4zOwzi1OnwaqzSIIe0Ucl2oVwyA9Oyc4VrrggE3uwv8/ab5V
fTkmZpZtEpjLVThmUdWzpdf4dTTcovFcpbcBPUj+FAaIrNwK/l4mAMO8sW7jCXp2
K7+XFMY5nnQe5GASin7/1kmciyotyJjqU8z9OnBHlHWec8yXbpG/9ycQNJQrGoWp
iH7jjRIaRMC5bxixutTCMp1XujBmjwmO5viIthCyfxp6X+dw3epsEOL8OBRjs/dt
P3BnkSJO/g7OqlEx/r0740ATObRIE1eSgLBnpCr7BXT0a+VbCAo/yMNRXo5XZu+Z
CK1bDVYz3f6C7QN0yqQ26podGdPF/usvWSwcmh7ycrrjeUp2XoiJAYmsT6zcgg5k
CWtYE4di+qGsSKqmNytqiAPylQHDZyxOJ7yMIcuzjvFQwMLjHDkl/FQFmjZwdSTs
9PdgoD7l8MTCuZXVkt8A5v9S7+pqNIbBJWSYTN7j4VkH30Poa0cqbY0QrZKwdwB3
W1CnzfhcKkXGBQEFkAkS6fNPNPw9dbaIkvB9U0lrYt1b6BNZQuy8AeftwyhcGnLQ
OEPuFCAzcf1o25GZPEA98MTN//WzemThed9v9zXrGzG9sy78ZX5b53uxfKWr62Kz
56GIr4Kf+7vQNKrNbXPZbS8L59xnL3uHRIR24yxa8BmsJjZTyQHY6/IM1KyNLP7j
lKr4RpXCWWmsfZKEtLxnVkOwNYX0NLEDPj6LEw5WZTvVDwXbuMqvK61MBkY0NCoA
U53QFB+hJ20iIgyQI+1bRbZ0MnvKBq4ybuEKpWioDEAbPhx4tiuJk6gvDYcy9JsY
NipQ39/lgeSPVNzsjAFQ3fT+4q9kXkzi1GY3eHTMc+L6TVIFS2S9T89be8osPK47
XHHEheJU4N/AcXorHC2tiE13D0pGDSODdcJeVKNg0qb+4ykjAZVTPpqfstY+Ngja
r8AJxDmoEgKoai2E3y8zQ63vC24v9qEVm7tV0xn11KnawJ88ieKwdgDOI+rblLYR
/MsDXAc2reoEX0RaukpN36gzz3QGerrq0jP7UMrs3N4nrIMTfSwqDibWrh4FpraV
YPF05vX27ZXLYDUB/3Tql70EA4KCoNUvxjg30o5QSZX4NyQrIOwWSzwCfAI/aCfe
JdN7phGQfKaW8JvOD19IrEzHFTB2Aj0C2cr9MDN4hRiPzYhczyQCcf3JdKwUTxu3
H7GWgcYsdvWh38czbd3/diFPtH9Qmlh6O/Jf5KLHZ2uU6GrpAqRZbRBjGLRwE+u9
CrNrzeIbgcfkEcUciuHrQ9U212JdB0D9MrgHi0jRRf2Q24azRIteF0QsWcWfrRbs
NRBw2BqdALZgSBMfg30mXt2Zij0NIfTTMQikysRGtBXjZZBtCJ0l1t9PYZyFw4fb
jUiijkqPexqcdu7idcJVLg112VA7MYTUm2spKUSZU1FGrch9YH2JEFthB1xTjovH
G2gLL9yYYCBl/uhL0l2bwzdqx/R5xCN/8G9X4RLwoP/NJ24LguEyd8XqwE3C52wv
q5q5Xr8zCeYz3pn+RqMRlhIg39TpTWgyTmOaDfSJ7R06i2RWReZfSSNg/imxAa4G
m3M/t2EDOOr3iZOnSKXD9eG2R6FVBYLBrCT77+b1AMx/bqwd2PXaPPCFipoMJVie
U7dCl1kkT66lvcOkiAgzFpmeOQFas7/KKd1XMJcPKC8qTYlr9c8+4rREC1SjIboK
ik/MFX2SzEWWvdYp1oE924WmXCu5yDXy5F421vNgQzTTBj4WfR7dwWLhsscvxQ6S
ILbahtEXpznddmvC6Q8AaUcln2fjm5UEMZOea7rr+5yClrX0B9PKetKApeaDdDJ9
GsgGo/XbL7rS6g9+ZIN349wdrsE044noaNZtkIr8Gje1OMWnPYpuTbOMSSV45yM7
ewoCXlwSK+9FsoHUzlQM2EsAshNBEw2Q8lo1wYE/kkym1RCEodC8rnPpRSU3fdBf
O2sfZYt6rHUTxjiw/YfAFsaSSnu3e+kYJvtlKQzbHrSbOoK2SxGyLTGevTTKyudH
6XlAkc4hKiYBc/gCRxhE3ZMLqyJV4DQVv9cPe+jBX/FWm/5RItp8xfU41Sif9apj
j/HuhcAcgz8NFaZNJW6mFyauAWiqi0GfkIxBjC8V4saFaiRfatEaFgCfD1BrE75E
JshjiHxhXJz3Y3NvJAVND0rC3GGQYzm4ZDBcNuEOF6L9XI9/txfYz+yHe7CIPw9H
NvdO1/GbvcUwWXxJiKs3NiBDIgDCtUUymPP9VP7q7b2IY5fkBmMRPkbbI8n2oRRI
hjMTvHAGMtHeOdQzUsWDw/JxHMBCw6c7RtEZaYF5teMPkXpUCVhA6WoWWBHseNtv
ztqZdyGNeAJF229bDyu8pQRDFMURTrtYeA6JjoZvxId2EnWCD50M4/yWtbFlZfRi
nEmnLOayzMe7qHKlLdP9F/HDOfAODUtz+ZvftwUTQPy2Jlc/mEfrhwdoeucEocFC
lDMtK1YxsGF5DeWT9Bgi73du+pASZODkRw/r0brh+gdQMrb9i/+O1ZHDf78pHP++
0oYYktevOj+x7Y3yFXsIagy3sEO9IY6Kc6cD2l/A7i2yFE7PEiHMIiywohZTC7tD
9iHKxvw8/Wg2hF6EixdeoHUJNqhqkY98xTJaM1vVDcH3YeSgJNlnPqoqsbdHEaaK
3HpDv0lNrgqFIt/jBhECYpmJbpPwqOmOEtzU/d+68EzofliaOL1BOXrozIjFfMvk
pD4Iqdrs1Nq9z+7xOHOb44NxLC3OdNv4p8a0H5jx2NWqW3vz2pO+BhS3hXjj3kjr
nJscWjcFQPx3OxY6OQXvUy02VMM/2sSar6iHQ5/72ULFUqfIZ27jnuPTY235YRxy
Rha/WjjlUOVZUEZjXnuzNaexqak0k/Rk/wQcj8FIqnky3ynRUS8uRbHjaBi48Isw
SbtUURszIsu8S8NxK/7HN6fE8Hjg+cWu/lFEwXjrPBcXhBPs8lP6YyFSKwDkwTfx
J4I1B/NZiXglqaCv/UH1iBIZ2vYjNwREhkhe9T9G5FvdGPFLEheBU392bZLvX004
HDBSnMGMfYE1X/lzWIwGkkJKfPj4eQEWq64fSn0fhSLkIW8Xj/F3QtD76kvuhbka
qm1XOFtVfGLsJRAa1YJ0e/8sB++sAQSKyHII3ZVjDB+ePxPziljnb7m+RFka+OZO
tAQujSug1FPzQACx+Oi1RdyHYBo+/Z1bc0L0Rgji+5Kb9G0vIyTWBnOQaMDsg5m3
kUYzDnwZFn3rdRoRfb2/QTx+80YoMj/3UFInD6SYNftJpq4ecv4a4UqThvp/e/Zk
fn6qj1XVQQbq5GEio5U5dBUdUcI1j3tT4t/qlKLuv5LO7+i19L1atOAdg216U63b
9kOHEaNQy9Svs+EqCB6i7CYABoYv5SZYfoDkiLrUNkGKQOWm6/j2MM36qK774xol
Z/vPPutgT7glNk7dhT8AV2SxycE3Ds3F1SD5Wnvus7tjEmOOUvsJOVOJ+UWm6AYh
NvSJZjYpdzoruHtirr2MISUxOJxepOP0nwdb75vKcUDXJt0efNdS3c2OWPkuYu3y
m2LrzrgYVkQg0RQ3KtyXn50b1P7llDJN+m6g37qXJtyq+qa9DLA+xEc4giFyhZCB
qI+LExT7tn4V5JqVGYqsIfhRyJCJjJPh/bnpiPpLBLkTcP/K1nn1yhVpD+Jij8YX
9U4FP3uwGS9MH+bkHnUfTER98d4NZgGWSlsCxh617uVNkQhenJBZwIVwDsrhpqCK
iGfHatLMmmqcCLkaOq9B4AHAgpZZv8qbDAd6rBVWpv/VgR1sSEm++XChrRkj5dok
YiAvFLkFBvBR/h1Dg6WFmRPsafos/nM48QTsMjPs/gKiAC0gADZ5CYhWNdfHpYJ2
OkVqrI+Or66pQSlZ9K6mE0EsbDqxTO01mpRjuHeIqSQJBbq/kG+kSKJ7MC/nDwxK
gxbECjZ7E4bRnfdr3rpNIRREPhi8YJq6nwI9byNYfHIv2dbqF8RoCQoN7+rXZbFv
KXTEW2VScoe6h0QzxXUmhFjenXPvmeWFmKVFXLAWjtErCrC6GS5zmzTtbEK0yI/6
749wn7EXW1pcThchePciqHWjNRsdjhR2b30BS46DobFo5O11HP5gsXvWrgpYaFP9
POb/gEtJhSGOP1AEACYJEmZ3e4aBWv4ZJSY69URghdM1tVtvaVU3Ta8OIv4qNn9J
xHgloPKkhga/m4HoGIngJk/NzBk72/2mdG9qhCgSFCPy7Edz8bQOYCXivmMU7nAB
czem53ze0jm6vqLcLhLJkiFbA4bPtGTDatOtcL93qn46H47Ro/P+Rx6V/lNQ7POi
MF4dPBwFKLOCXRDpDDxN/rH+PgZ+iPd6FOjw6tYELV8i2lkcXjSGPvbl4HmVNOxP
LLHWAgnfdqTeyoFuBETeOGY76ejdsdyIMtsGWIR2o//lZLVC050PVtDWTvP2RUQf
WtAUk0loYJ2Shsghi1gorlzPjjUDphHZx2L5tcA4RF3wcQB769pufzSfW+vTiUu4
D+R4/Gj3QwOKGuLefFfQjupcFUDkiCetLRaEy58nPYR7ab446B8iNLh+CRMUiOuP
pDUp1jEAPuBLidxBSJXbNFqrgcEPJCyqF1eO2qkQaVGr4F+hsn0v62sXcV9SWCYA
2j4wVzhnLTEp5mKtZi3tmAlGVzEtSVZQP/b+6aIuS+a7gDuxyNXL+1UFnafa4TOD
njZtFODD2rIh3mz3tpdINGRT67ONtQCuHZBHRFUlEOTbcz99S58n0QUeyvmcXj7Z
l24St05ojH2cBnhWH6Wqv7QhYqUtvCAtZBdzsgiHo+5JpuPp9XGFjmxo2G249q7y
5S0PQCDYZ/1Djfwu+/H0bCbvXF3xp8+OqDeh/nVdAFOm1MjjPy6JAGkqGy6IRiBc
fmcDzu3+rvkDnXIGlzHgZA63j15E3BAMEIQ0ZcIFO2Kydsc50fEru3dZceO0W31R
nT5ueJGJcpN8U0BNsKQU+jqQNj/89vagewmuxi2tp9JW1z6xw69cfB+QzFofpiDi
6SWq89RSh3gd+zUfluh9bYLvxLNjmOIxmjuJxYEX2n8QWhaC5LnTI2ZEyhx2PUp/
VFrli6c9olKL00+UZtkftHcTQaiXGTHdnQQ+ibRtgcYWfnpVMPKWTQQJAO+9fnEb
xWI8gqzDJ+MlSjA1CkbstzyCEPhpmkZZCXqqYLicz3BC4qyEvA0dLcSHCEzIQYoj
b2SH6MBvpMmrR8VLfeH/Z0Qpu8dXFj7WSspawT842pDap9GFAINBNCAXXeB0AiKJ
ofLd4lh3dP0+0axh/sM7T0gpOkhEfbe03wFs60oObH0xGqXdsci8CdyRQ7rRadjA
j7tTznAAP4ol4QhvCfeakXwlXi9o3DSKDDGWjGrKdHIxGrsjW+OqG4KgIgL14NM9
D3zQDa6zLUL21xhVgnI4Bmy7t5vhn7DFbwU8dk0vXKOGMTTXCV3o38/TCBfhoMZV
LSx3wtMUGs9UcqiB8lPkgQOrbpmn/VQX5E4wkFthV39wUB2WBO0SjF/OmC6TWu7e
xKZl3D7JfmLgsd7DxcISQMcO6MutbEJxWWLWlinz1KjuOIvy8uwmGcnQOQIub+mg
s34jGFXVAzRfBMsyF5Uj+nIDd4jKvBFRI4pX726nt+bQUUDOVYdPBS+g0YRnlbqz
dwsduwafJ++6NXCttRQz6CY3lRgvLhKwsgLNe3tw0ZZ8LuraZ13Prz9S2bzKE2Ei
dy2wZNcevYwXKehPPJAqAZpEeRnwLWFUWSKUYATKh6sObGTPCtTAMxl9G8gAhshF
NN551GGPdw7GptLtOhbmbn99HulY3qkSptIQ9KefoB5xYdW888xkpHQt1fREGCvA
jkFiWscRiUG6xQtTxYK42S4sixr3jbKdlY5LRvlBs3ZA74Sq5mMyBgO3glVEiET8
DCCUWdA5CE5zUlGVyWTsjOzGOKLIpQptvNzsYf7VKxou3rWUwXDuFuCB98z7Plcn
3kbAvKWzzMIFqrX3pqfeEQseliwnMy8oK3si+08v/EBeH7wCSYYiMJFxeFk3ktGM
2R0uA7sCa3gJK9TBUsNorYictjEUnIF/1K2apsIuAHGFMh+wuPmVapGIckfDYTMR
16OkeNei/uYyt052AG65awQtIOKUhzkTBRT2pynGckmEhNtb3V2459WelPMV3VaL
CzGwMJCrGJBrkOq7lS1mryOgb62WRD03ShwWLH9vz1R75DFvWOkKgB5twgMS2Cjf
CbsIhEqVows4yKuuGG2pMpLachvEufamqUyJ/IRWFkVsPpVkRcOXK7jS0iuOac/S
dRGuzBL4gv7Nbj3ug8PcsREuvNZuVx7TdPAsrkkUdtRBf/ZiHxAtsvGJxqREPcfE
fjDxRU1FI3mPowUeNLLk0aGwEfzpzzCQt3W8MHMmxh8OEpCE91uTIr45TeZM7v2e
Jfl19Pdk9hmT+k6g7ZtJPA56oER1JDleoeZbIdC4vsYgIVXamlfRar6zWuo5pqqZ
JM0AZIvUgibRpTGpMXxa263BkgmwaGmxpIx3X9Zv8FcbWu0Ft0SURfySQm1mLIB4
tzlkP4bmB7FfWChZK1asqlN9POHUcWj8SW6KJDP4EdpwpMSsx+9XwpsT1BojBRLJ
/GG9mwIY3pgzvN3FAIct6HSobt0IRRGvUmqSeq179iUSkb+QiRqwbLbJ9szpxgs8
YX7dUBvwxz7Act+UVZ/Vo0IB5zIC9xsPDzabImbrf6xej7HLT2frBIMhHUqR1tq1
3TRA1RMt4az2QV9YizVco8SpJCgWVdIO9bUJ4FD5j5WMubcPzQDnMgWb9CtV4eoZ
E3f0s0jzTz1/Q1O/mVo5/J2y+9ESBfI6Bb/nFsrl8ybyrHhweSQEn9WAELsj9lGR
YU3t0UA2cppoPIm9QKMLXusr/4GDWGegUd7p80EHmk4/ltZcRxnSKvwmRfQOZfmU
WR5CBEIoSjfKGOroGiSSnVTaDXys/Fh1+BM3tK11yNY703L2/Z9+GJBgdd1+es8g
lidRxsXSqgpCwDxJM6ldcaGz6KG0yD4ykgzR/20V7f8PBeMWw7kz26huOStFjZQR
ktxEqQIPlQ+CNxjr+LANyjgVaVDMEm0x/0nqbm9WpLMfwSoR9MblQOblNEgtTZ2v
uqjTqXpemSKzz8ZIojohf+tWMNi6hpq8Q0fEhlSAdqHEqIsGDmUzY32qLF485Y9S
AumBgeLztj/0oxx85oqUh2nzndzjTpMUBsuKWctoT8geXxA2N1tZVaAgHTUMex/8
S4Pkr+Xh64Ledm2kf+AeeSxL00999ab10NyOY7EsGlYv6jMsxtrEjZsyuoBZucJW
KDZMtBaeyqJChN4T9x3ajV2qibehtnpje50XyKBSH3DxtNLIwK2NSUheZPkb4e5l
rayQ9kJK5rvK3LgdFK6LdHBPOD2dvdlXl2fm+zeWSTcCv3rkUD24e9V88rljT+0K
WWF3jZAXbBqe1mn2atHdYqR0pYrW+yqVdSgob7IpD+n3Pf0k0wUQcP1Vx19qsVc+
QYRg3k/I8dMNIzNIpV7Un3xYiRIyde5DBF8txcOW1qeLGLYVInyimBgFq8we2QH/
BN8NENvgTvynOFuM/FD5/7XTtPgiJy6Upz2scmcPBZtjLqPLKuc08iC9US80kwq+
ZBfIfQRL1wNN6adeOibhe7IeUGiYrXKyOfP/QNiedh9+/rfawwhSmCYusXv2nwZ6
lR31uM4fIJHIu6dgyBJ6WZRVF0w+vrfi68nxaeX2W4qDClUzjprNgFvCfwruA0tc
vO7W8QQQ7BilMliQ7uhH6pIQfU7qaJeSDO36Po5sR5dRq/WoqnRtHqUdOXtD05ni
IyHWYpV0jw8pOOqHUiRDlzzgNgVjdHi+mRAI9+EVxjAp0ZnDbz/r0mWRCzNa8ifs
8hmNH4uTobr1KrhxNyUCjc8BFNGOTGZF2Q7Bk+LvE1dWykyL2ABO6L1iKDWa5Tc4
AG+bus9MamB+f9ilzwFho78KB4v6BxN1LBBTgBsz9vlOC4t8zhy15ayayTbvwCGG
DZvpnXaLZ7IiaQGezbtp8v/lEDR6z5dm+XhXZG/L1DxH8gySca59CpZqlZzBctxK
dIArERDPMTrzcL6lBvVqrE6uKmYtUTNNaIP4G28J4sabNn2hpW+3RhtAblJwAOEd
65t8kjyfRHAFxXUfDWd9zqXtPIa3nV63NWSjuBzYp/M2VNBRMgu/a/hHhx3qQYj0
o/zulbQdM2BkCi+25M/+Q7mae6N/c16yVrm0r946aT37MXOXvynE/dXhC2NP0EMq
DfF3UWUUYMw8jKpx3dNt1+Cq86h+Yn3/5nM2aPx+McinEBKOEAkIc0qiVhekiZ4W
iYhPIwnKPPjYwTf4T1Na9JtRivZxLRoTOUnhqemh3kSfnK6/MVVpoDJGZ4KlTZex
8oqSJ5SAgbScm4Ajr0ZInpytIs+7Wd7UNHQ/kKDnMHmmzrpWfn4wR5+qAlXR+SaI
65KAhaTz9bkpQkP5xvbte2EpPoxF2+ei9jheIuUPlrmzlCZEWMZomFRNuFgg3zJB
+9TVSR6oFGcoohL9IUyJyMeoybKVdtZ5IxSXQbB8RYACGY7lbP/zJaurNaCWhLm+
8sUCDhC/mVDYDwaGgDUBgClMCEjDCxRKQJvduuStHdbD/hu21iTLqCPr+OSE+qk/
fjTOorARN0n9xf/xUYHyxaKoYGVQ2tTU6HyN0V7lTAb3wuPgdkx3cQbxAK2n8oi6
K+3iDQHxLOAT2Xo+9hqJJIM1cWqHTK6WmAEtX7GJvzZoVAEo1eRcoqEub0+cnCRz
4ye/Hx5FNjgxUS4jakB7c4TWCnGx+lV6EOrr76tCJXOieOI0RIOq1tpjPJKBR3If
XuGowDyvfv2u7cXPu/pu0YuXEs9WZpEzwX0TN8szr6N0OfT6yyTkdh6c76x036Z2
4j01cPhjIOBbaCJQTEq8wH/VqMPMj0iUE0qDV1gcU1FwnOSaD4NJRSdeJ3bXpkss
ppXENdEF1XiC0590EyN74jc6xZXQPbl3LvCzQ+HMAIDm96eI9lLrlfJccwGgZC+5
xZVfHQ20tD+adWF0aggkE53aUhtqMaxE3hmtf4j1Kd9jMOvgaHaE4qo16PTgAlCV
J9ilOVqKTFNFK1RjrcvHUgFoMPaq1O3xRSMxTUX96DYOClWh9PjSWTONO6qvrXy3
T+Wmkq4Xnm3gsvJgl+gl98WgGSgsjGoIS/M18cDyilNGwFUz55V6ZhplRnlE5hhV
7c+9J3UOBZluI7GWgoY+5i1S6BdOSbfuHfSP4JjXwM83aa/VaQLkfMGBMFcZvBB4
p44ys7eooQ9QWtIUmxDrxrJJGSRzRgLUwApxTFGTFo7dSp+jb8CQsvRQD/TnBeTQ
YLOgC+sRktic4uGHMfooTniyg43qXb28VvFG8b2uwkgSpkXWaSFHyJPtuT64vbgo
70MEL9+mcsnUtPIHYJ7g/uLmxLvW7IwtYT46zGt1JawZeIIA1V4UuzUpapagnkch
3MTrAwE/tgJ2xD2g0HCfpLDtYeF7HVq7J8bzqzUtc5cRglytBjCQKVjospOsbll2
dsw//vey7ZL8MI9MsAGuYgTpI36mZKf4UhemvKry510AIrtryhpWy8HCrRaSFzWk
Qqp4BqUxUpBOFcKDyeT4PGGyogwm1DPuYBsZxChuas/sTYRfJdUrpivYPszZ8Yy4
ttrYBXAdk+z8uov0v0QLCuIByYpoF/KuSV+dEkFEklLF8zvgnEHW/GmqRnexF2r7
v+Rl4WsheA8PuePDLZJUTayvF8wACdNKfFKn8NMI9zm5VP6RKZ03BYr/eaU19eQ6
y8XHZ4T33rYhXlj4WNO0y2HzTq9JgMkJhOLc0j/mdj7YKmn5RIG4dmdfbB+ciu58
p2vl9nxfaLatBkGQwolxVBTqT0/zU/ikbwbAsAjZ/FJu4plk0CPdEMC1ba4W09Qc
m+IpdZ7gRdvXAN5Ll/+hEEPwvAcjZ8G7vA544t7NY0lwUMOIbG2qGpJaA+Lw2nIR
nVzI9iWInVA2MxdHSRjR2JveGx8DU5SmofkGcNkZUJVnGuej7G+svmP4xnMqRYOJ
9q4ZQc8IeALAPFkQj1ZdOV0wBe3lGWpMtX2J0Z2GmNWRTirii/6ERYTwUlfXr483
bsegtzR+Fay/ocGyQvFFIZXuzqpVAfn7nfQe1/K7ZD5SsW1OXpY3GFTGoRDDgawD
95RXijES1Bqk1VgQBp9aDf9Nx1xuaKkUBOUH/q6zrQ+QzJqDhPTjn42jmFYkMk9G
lqiR2fIq36pmXvzRk53gY/qikU3EUsV8QsmBqrQXq7vmkNygUFAsv+2ZVThSkyM5
Kqf0jFLnJgkmOVoblZu+nXl7ZnRgdAL62EPNxcWztm/CZw/yZN7gverLbtC9Lylr
l47X7amQtSBkxhrvw8DWj8ghn2g9AV3YRQe7w7nxDgB4c82ageGVTOZ1JCy8NyZx
rP8vIe6rr/tYKzCFEAVc/6xFN8r9nom9dYWEJMVqngrJ9qM0AgRCQ3qSdxPWSTUf
tjmjWqSnN+awslc1apVaNbb+4S3opykw/gCRAQmRwz8YR9107zrMl2f9MFKkkcuC
KgPzFJmYSN4U6n0PDY6sBdPE9VwRw1ApT2mBayXxKIgfn56tai5M49ha4B72UE/N
1mBKlnppe28osS4szFAdaoka9SDNv11g4igGPKU1nDHbUNmiHX7wkKMiGqFJoKXN
3TeTWAVjJI5551ehwU++a7/eLq0O5FXo0r6pZdqxEmGQCUgSKd9+9/cgUK3WKl/i
z7kpKvK1DhTnIWuWOx2hdVq1k0ZU9sxPCHfbU8n+dNiGf/GFyDh+hM8i1+SrCDER
+c0RTQ+HnKS+750EEaVflaHBlc4LuN3n3IO9pwIQDFJiW0+PraL4Sz2BgWL2qVme
5vdmDWP2LW0TztOjwAHvWWKg8wmQgrS0B3CdxmSfXZbuj3qi6vDW8zGltxzs0S+Y
mUAjb2det1OOsZKNvgUXVS5EScNeTVHxCOy+S6PQXZ6u8g0ImtwHo0RM6lbhuWeV
xt3LF3UNXjhtP75CkZFnL8dj08ukyp1jUFHOCqLWGc32bNsGLi0sbohoIO/ZQn09
pBwhiuaVlU1ypdXnNlrIBd4tepjFgp0lij2Oy60hVA3mPMLgHqtEu4MCwSe9Einx
sr7sR3BwWT3SAQheR57eQjd/UNDbgeSq72TJ0wWAo4lbxAnUCOEOxU35/LVJyo3f
DxWRxVmTbYcMYXx0uNx9f9xxrLArjC1ST/Nk7pZ66WIQMMt760UDf+TUH69vPCZH
QFLk+SyCZHpwXWyqmBJbfGoMFHLstp4lWpTnClhh4KIsrcYhTDJovBvT1fjcHQxt
1hkyanj8kIEHfGY7BPAX92OunDWM+A5UwouusenIg8oo/8scJ1mQp2P/zz6y40nq
MQ/xidXfopBnoeS9oAZfw2uGRWG0JvxCe6e0UD1uTGgwLS5JTfEFV/wSSsvMMCkq
3zfgL7SRtZrgvIP+du+sdP6mfUthqI9R3kXQIR8umPOLoyHiIqNXUTbmut7RlP5i
FC3bMlquBjLmp/o4rnPcpty+4qyhzoOZMYF375NtRhNM8sDajMhCRN3cRgZYYxQc
h+kY7CYz3gTgYZWi8adwPaU9oFFR/deAVF0wy4lsT9PRudwv978i3qeVd/IwYSEh
PAdwGFBA8iVb52wgihIl4XKRN/wFyoZ1BxyLk5Z2inQsnAcLtDPXw+Kb2bGm/mhO
h2FWbAUCalZ/KhAK3ditOxfx89rBrqdXnWQkxPx6RdKo1TS3pxIFXoR/wursI5wz
E4Z/c+pM4VJKWDNuEBaoJXx3KOSP4+6G27B4I/elpfDWpUBGi3q8pW2IHzUYTA22
nt57McC+Ue3u9EIZElxOWYmZUj73HbavAVJSkE+7HNC35TPHuS9JJ2kyRmA51Kr9
dKow7UfqGOfJLRLL932dGj1hWpmMUPdLET2LoF58xD7bvfoSKPZWDaeL2pyvfRk1
or+bLcrCiqXcK7kZOMlD/mIInZpZjhOu+P1kZGIp6/M99UeGan2IIJWTlXXqMyRp
Rzzs9oQb0OjDESP6B7zv0xMS2JN+jD2n4XCNUMZ59UPm0DOwnTnHLwX6f3yN1jpX
UmDv6z7yFHCN1W7bR6u/MNDrAvfy3T3HbhIUgJZNbayvyIaC5okqERoFZaX/0cnu
rp1VxYEYB51rQ++1KJfaDfW0b1X0U7OhUfmMeznCL9tOS3wAGWDL8ffBjEhw8J6p
2YjKkfViVslI5p7EPaKm2c885mA3fIc0vgzjbB23XQg3w8AfoFtiRo7ltRtleKy1
fRMm5idtHsmlXwKVGUT13YHV8h6AN6R4VXoN3q7FGJhz0RAePfAhfRMiJK3IPrDn
lkF971SDJaCQWU4V1EsssXxXmH7+nScsZWH6Cb16lJSax7h7TNPAhujAeC+cdq2d
3qA4pLxqropiFeLvaJLFtcONOMPd4vHPjY6c3XnTjcQmTkMox373Clyup9t7kqPh
ceTAMI0zMxkH6a1zDO/DpLlrmzsSOqzfoe893MWCva8PCciU/2WnyyMXsMj78MJN
5YcG11U22nITMaqF6ID0uO4LabDGRkxIvV3ZxyBBG5dS4Jd/mEDBuD/jYh84cgNg
3Bs6R9/e6QxJptrSA6MeS6cKPrjhtzAuWunnzZvDH/wVgmpFngmBhaUW1ILoMmRO
eBe+rkaxRuHfOAYAnnwnmDo/+Yir4G6SqJydneDWqcZD7APAdqgpJ3b1DHU8DQxZ
+B0Ks22dARTrE5XX+E8wHoukvDJu7yDUaKg/YUcsDJUEpgfb+fAw1kKA3zYCf7rG
0ZegbBzU+2KIm0mOT57rcsP1pwzP5Ue6dQehRL1P99a3wENhzYIjmmXkdyDLSCF8
IQtanBQ8oZx3YRA2hPGiAZuQ3C67oLVNcIsNJPHoljK23mwvc6cZNLwWli4vmUcZ
GtBL62BeAhQEwSPFXvu+PAT7bVz5W0yTm2bMp+CNSVonyel1Kvumecu1DkLVCh+d
2XdTyZRJt3Kd/wFyc1o6UCOk4vLfvp9VkUpPxPGVMDI49AYVY5oSMNWgaY/KV+Vu
6/xhbs+ye4jK6rMoKCFwWHmIlR0GK5V4MHGkDxEj28GAcwTUSrFVPA9odpv5D3Ra
Wi/wE8o5jCoHiRMtf3jKDSMql2XsplmWU46jWvmSIqgXiwS46k9xnjLQE9KWeZvw
KpoFIi67vqtZ7azXAAegFRwP61mTIpKYM3Fl+u215nR/FOwLjxbowPLZA57W2q2s
9Vv3OfUpD3Q2Ht7p9uk0tLRfVWkSWbq9EiknEf4BEevIklNhysJ2p93/WPQmSdrL
fAvy4b2md2AE8ncQxnViL/VcrTWjoAB3UP3CUS78J2QYrWYYp4qLWZ5ftiWnD/ZN
cEmfidqBIuxJuXB/7IrhVxVxWhJjdDelIRkQXVDMqwDkxlMy9gJc8MrhM96l96K9
xgxPDopLC/KHniSzGlf7K+Vg8YZZT2hYecQAaxjeI+HtlaVlFEz7DWeIIx4JCLrJ
XGlezLYISU2j3FfXBKU9FgifVaE6s1Y1SExwFIs2pwvdcIfdSprphfbFIsBRo3QK
Ltl1K+xkIWzFRV7Sfo+D+lny7MAUCuAw3MSlHDCUOKZ0qYjFtffAlihrxUXWuVqI
XAcWX2MQSBiksFz+He8W/ae4ljjPlFNJVcbn8q3sdXMiYqUHvPIZf+76ut3KLdMP
h/KV1n/qQtMY5euufJzEmIGWM2LuCm2yrviN/sopUaORIhEf7lK0qufJ59W6aJKK
Kl5kJv5JN6CjIxfMlGPeiubdjdlGwEbPNvVK5K/3lvve1QqqcJba5PVRXdo79srA
2PsvGcDsxpDAFHgUBfxS5dDZ46AukoENBBSaTy/ScNgmMtoJlBbzCgnV2ztTpoqn
1VkVADusNPKFXJ0s/DfYmxbsL83meQXNJX/rXShucl3EqXN4jWpJw6dBUFYLwdyg
eOs3Alz+KOWSg7z+6QIU261EHwTG2J4pBiw9PzxivI7zcEcQuZo5nr/dxn0PcHLc
/Zv88z0CgVKWXcdShTXd3gqbRU8QGUJHgj2qRtUgtnE8fhIgGimRRm9tmN5m6jM7
6w5EwDKWO/8/C+Gh4wdJ+G8oLCT9Sf69mp2ppQ2Z26lPGcSuNcoFs1AqVBlXsulL
ZxnPlOb/M/hsmB32lJR+okYWYFQnyTDTUTcevXiOgIWJLqwDU/CX67qv8Cnf/GM7
BzJjK1wOtVFHxjwmL2+3IjNnj6tojJ6Z/CNRCtKOi/BSy/VaKCkw4cH9dCJHRnYj
yTRMORGRy2HwQHuFWinVTwXLa6fUJdnIO6jwVoPBeIav9l8ZVaE62v9wiOJQBf8m
xsWW/kirJ9pTFpt65XQ/TyznsFXiPdCiYNcVJIglG7pJogK1yIx2T3QpsmG264ux
YsPA3bz3lzTKy4d3XCKgqTTpzdbbKkYcYLZsJd9QYRklFvMmi6imkK4d1txL/ynp
xyxBTxPp4QQpAf/bPLivxk9oTBkvK6EvmTPmtkk7HxcwzGBvA+HWaLNPBx2vNWZ/
KxygDm/6Kj9/NRUcUWK1xE5Fh4M+txtUPItqAD3FgsrjSBamFnJfo70yat5ufZ8z
IsZMLIQjzFsP9P2+FFxwa8JfBWJmM2juFhyV3cYGSAfOUsDLZ5em+O/kR+5u2K+A
bftfCf9wsheuCer+TajtHhnQ5k9AJ6uualmTRXFb8LhO7i8/RRMdZ8QG1r5Y7bju
coOop1uLAbmC5LBYI45mJGbRUagY332A0Zn+Hame4HdMoxcXpkiWDAeEpo4aiUhr
TH2CjS0h5QoQ9AO0KymUm+DOq5CRmUAp+VAwAYTSixZygU8K+nyyTE8Mxpfs/JIM
8NetC4ZCpy8eJb0mxwVEc/0vt0bQHUHd6jxXKsfXHb69rQCI/t77jQXWTO+QnAgL
pkwtvIma5To1uo3sZ7OVbnZZnTgQ7qZpmqfQ/PoFUAATHBUq86jsXPAEjqktg8wp
5dBZ/CxhshLy25nr9T7UrqggyGDjC289UrMK6Z9CYlKGBXBvY054GR/nuJ4F/Mas
w9h0dlWhfgNggW76zwz6BnqZvRBpnaRwqR0YXZhjMP9TrOCPknxQkPYXWb3p4K0y
PWd4sixyQKCuyeRyiZqcCcinLQkbEkq5bENsUPWXoimBOI7bz66KAx0o97QP7n1m
WD7ZEBngwX4kl3xttirBJ3d42pNlmX+AfrtN7iXwnaCiQhwLcbVe69ptab430ico
Mv2nVS87YxyNNu8qfIPKJnj7vDFWSvwtvRSFguaXewvCMz8rPPM1Ep3iAfjbZkVC
uOQ0oYz+a/e/KpLExMA/MuaiA/0VK0ylkniB2sCYQtH72OaCC1RbgXoNx1TXCD0N
7QaGiY4S6XSNSqIC2wipmaAQzKsZX6cnIm50SyywAhkM8c0by/zvuZPW/paG9tur
n4WtCJ/VcIFDVc0IdRE8AxsHSKPPFL5xcl820l6oNti0/kJo6Mr8nzt3EApO4whD
Yv3zQZSt6PoXK8lJMfbxmC1dxkebEJZ4XQyELDXOOAyaqsR8ors+OCcDxyiQY5Ia
RGFD9QHW8QgZCvYfU+A6Nwl+FeRH3pIFcIA4rGdwLLQ6OibfsuuhksVjTY5mQ65e
QHOlTbf8adV3gfnSRv4QBem60Ff4gbS7mLElpafqN6k8Wr00ku7T062HbaberRoI
ieCQV+RZ6zc80kkgbQeBkycZDpdqZbPd1PA/4HL2Uu7rckFGLY+aZZxMA8gOZ6r0
hS/Zl+Fgo0jiDZWE4DpiX+5JA041++a4iGrQJrVuIND2ZlSLS+kL8kUPXk5MAxhF
UCbjhSCv8IYnm0mflTpeA309YRaZRgqNvQ0FsoZ9Au/0zeDywuyDHnAVwxBYeyWH
nVVgt45YNofQKLo8qc7lpX+HeGnZsmpyREv5DZa9TnmWkc2djkS2crXvPKNUds6x
7CgnGtJsmw5uXbxspqf/uD6UWTVkRAyCPcgIDXHIM6VS6e0ss83qA+trrmgMgl2Y
iwbodN/WWVC8uBRQ1cQHOXnMiMHDtjLYXZOdy+t5r75IB1Fj0uFh0OsZJpDtjYtN
UxA0tbWqZ6tZ9i2Ta1VicQ+ZZW4zrdNnkAQVouspwtZGdpXk68m6XQ0zekJwPJhS
jtUKEnKLhluJImzKhttLPFPICuH0jy+9mahErd2JSOFKTdlYxWnNA5ThUy02595c
QBQyiM3IYPPW69jx43KtUN29AtfWBfFEkbY5SFSPuRHeaT5xXmukvr6ZryG0OB3T
ee7Rhp0sMTUZQyLAPiWzZ+Lh3ep2xfIf2qDYfcpmF2/JgtoMKBKL807TpQWWrY03
PyNacw3iCXnfGapWzpGteAoDA3X8qou8nEF9McavLVhWoSgQwH3fRekl8wDMzcFg
JK9vyFpRB/5yDvMcpgHQoTqK2YUVt2jH5CrcryM156CeOA7YFFlYqp+V/Tb/oBGD
I64xGITCcMYFGE+4t+QMHl82dywude3VmdEMJmkoIzLX2yhDM7d2AGqdafcA209i
p0+UaCN+PFt4fBOtZBR+ZFTCkmbVJNzTAlZY7KL3tbdqrTCBlRQxIyN4v6Fk7snP
+mUqca9OVwKc5/vceFJsODBGnIKh3xlQllWv4CM7tWEs7sRAVoN9eDsVKphtk5nn
dsg7vgAPvv+x99cFNl4/G5JhPtmhp8XfHcuUIXhgdRkwI1+u6zKQy/ABFcM9QtbB
9iYmVxJcQufA9FEuiZyKsmtz8v9sdqZKq2I0R2G4xeyQgVgKkzKWAOI0Lm91TARy
5Hair4FxCJyOo5y2q5tx/r4p8vc4UgBpBky9PgFbBA5mch+Fjs2SVsm4M4hQnFhS
dj8NhgQBmPkT9sHOvKau1hZGZxVWMxiZiDeKiyoLyQWreBjGbTl6Xcz4YEl2dp2Y
QMxCLMG2dibAoedpJEBXoysFWMN4vyvPeRND+aGPtDG/sUIT2JNRKWkeh4GWAoGb
gIbhJcQpx2OCtQwcq5LZdcvJ71nc3KPlODHWrrktJd0xSREJUwGMABeQrcjxfPXv
pbe4MwsLgikCns3o1ixfZq18ZR7yPbtxGrgGvY8IIwegQ6VQZ/a52hHOm9RfWlAr
L8R8a7uK4H0O9qy02hs2kd5jW/OjK8TPbD+RoKMfqRNMAf2K1Uyo0zevRn75Af78
ihTaEwfeTiQUk/mZQoqHkAMrj6n9BVoSj024o0SYx1NE5QNpNoVvanBMRWAP3gDI
qkeYykalb1beKhfqPRqVwFkZYdmq4e7kpWhQzFsfGWpOPQYdxiR2q+D55RMmaVP7
Tt+PgenQUbxu00UOjGAV8gduWijzr9ZkfTagd4rCXcMlxs/dLHS2TyagdVJQ4THu
g5U2XpypoeScpPaVCbIbkuQp192HO/ajbit70LaNoAJJsF55qEbbyEFsrnBHmDa8
aDY4yVc+qJfVlErRbIiyalJGVOeXl86xh0vn9VCmOlMGaB/mmLcLnmu9U2pEIXH3
2oNZobaYyC5gzKPzIvwY+xp/47fWRGze6kvbBc+iy/Q5uqqcfxDNWjVuWtEPC4Dm
qEx5IrJpF3LR9Fcr0qs70UcdvHEZ3HZL9ZUDlfGUjvgr4JJ/FwQw/C8sri0L/wpy
djLjQ/KN/9yykCbjhtvFlngDNvsXDUqBmuk+mpXhOc651xO1lIrnEwA+Ql7B+QDY
Jh5MqJQD0580jivCM7OHlQwvm6QIm3Qw/7Giq8KLgCWVoMluMP3cyLWyqx1vVej5
DphD9DZgFz9nHTnsn0g1Cd3Fi6myzTPsMqVyqUtCbyOWC8B6FEm/HY+jMUGqnIhI
IGmE6RGyV83XhRAI/39a92IMNQznbuxhz8iZvHh8g0qpBgHdICwnDlnPM18C4wkW
287E3bbhJO2y9qMs6WHAbYGI5mqMZgMKsss23dd1ajJFrVSx+N8LatdJp+p8HiTl
dxgRg/zY8nIe0ADLQM4fFt8qqV/jq15hMVDGIyUEmFKcpLXnKgQnT+cTYVI5oEgB
m9brvUQukcEx4/55G95u2TSr5gQcVcBhQ4znl6QBNoXmFwrJI+8NIWzO3Qdf9zMK
9j3pfJeGOuzxQzftO5NY4PtCZLv4RAoh9+q03ggMako0lRqnzeD/8T3Vc4dZeB6r
oMF1pDEvX1lF7Q8oVDDgiUM6QsVEmiJ3T9rgaLmSml9KPV4vLsgLxHPoXlNi3p59
nSQq7oHfIIlxXlj9uPJYN1AuC4jhNB7yntMz5oQRa2y6piwEaDbGxlCp9f8bxzjF
mwueyAIcGpzWBet6Cssadq67ja81rzkRVAIO5hof6V2vZhg+wZ3smOKVEP0dbLk3
sfpytjFFtRD/W7LWpCJNagF8HNnwrfzL0xww7qls7H5EEnsTkeWPN25u/I7EcdOv
3OHK7as2utKALl91apsG+0zjxRcgNW+pIId4GE2FgRqzQ0YXQXiVpbMwdNbroPYs
WUdiYwvRs1jXPiNgM2sOOWwq0n1Df59O/OJ33mBexaaF+t+QHhQ9amRiw2uFdhVT
Yx7pcb3vCS1oSBvDkIxG8hvV3Fd7mibMW08vZptqrUVd0T5r3TQ49ePONEvF+Ghy
nCoPtYRqO4/DemiGY/BuJcX62KFdHX8SGFvEEo59mXG+J0RUwlCahsGABDeVozLI
wzNNQGZy0lB0DWo2Ub/NttCiovVy94oiSbFAcUar9HeP0nkvn55Msx3+9IWzf5ju
tvLNPnflhkfFzm8eG8+1p3XF5TyZ94Qphj3OHsSd6KoMXXPnMNGNxunFcGYGhoIF
D02ZLJSSKpTgOPBWAI9ZTGE/K/TwX/Kwqod5pORtweVDyj8ST7mqa66qjgN4OM9r
Aa0RhWfLvA0+C++OaYT6RRrR736xvOz2VDUavIBoV/5hcrLw/2Zp1gzUsPPQchGw
/zYOXv21mQbyUOuF1QBzqDZufUitc9R6wiGzH0pRuXIEC4HML8+VclyQjufA9l7Q
YK1p+ovng4CTHLbnSXSY2oTM6Ypy5RMgIIfXS5fHZsM3gEueva6tN2OL+vPkWI0H
BW9P5nllC8lKagKF4Ia7Q/6rwSKYUMGWzl0awkJZa9LS/9TPKQYrEPKotciDNCLI
YjOeAIzdGo7l8r7iHPB+YpbvrVYeXuAj1nuTK6hGjJrKQuMZqAELPgSHvLQC9q2b
gQ/j4/D+dTHRPxDaomcLTPNq48hZti2MQllc39NuuUSL1kele/KmINxFQZJDGcRm
zLnq0AsriuoBuIl3RJ+TQeR5RYGp3zsliZ82tBJfn+Sx65HiuFHzAz+gb6nakHkS
eRYp/zOZkOveFvoMSE9oRB7R9iA3Jzp1f+PI3oFOpsSDtihMqqVbToWurGVgZmx+
qUG/rxyKlLIlGpq2wsPiM5r+oqjq5cq8eGkX0HarTsgrAbc61I61ajWSHCxPose7
4zpGK4D1H6MLdsBJF7kzchufxNePddC4Kg+TbSIk1CCD70wuaB1ZdfFggE4D+MHo
8hSvQ3kemQHmN3jpzB4H54VTjtW7HlOyedu/00SboFOwv600LcLR7X/vLbWvVyTN
6ECC8M2lq3ryOSZFQuuSZCA8PKDKJnqiXcZ9BeG9F9NfpXqvoyRCbXqStnsrRnz/
zS7bapS3h0BOVSwWilPw3KWHfLpRySbXV/vDM3wahRs2ZwRXr7thhgHDVGa+Ak4x
QCdRb8fybo/TB2RiklZZPxW5sCZTA5rFAB+HljWTeYvwmBpi6UaqIN9DwoKdJ9rp
37wEhuyWhhp3jIPGyPqUyLH4JThqYIkYO8238jP3qVdQFi4dSQqdbkw2PtuXvsgt
FD/GrGu6Ak3EPJCHJ5qYFMabttaOBOCIn++0eH9hY+MRksHI2tT6rCtzEwdFSGQt
U7meEhWd5+5440jWHhO66VV4zzxVQedJSF0/CVeHHiRPKQn/rQr20c40tungcHhZ
3YJzur3ZmYhiVUFEp/1K+tkXUcLrtSarYJJWwn5PeqvuBlWp492Evq6ky+78epN4
5oWi1C1ZbI1uuB+f8PglOm5YWFQdCXttQ3X9DAvLcK+G6p8i2uhEjL62Ds+fZCAU
6fImj9HN7Ncse2ChdXdfjlWULDk0PQHk6wwUY1w8fq9T4L46wB/B00wZRVqjk3JB
4QUMat0pLWDj/FRF95iMDMYPQ9bMnE30SDQmApu5qB8wB6NTiMDLGGW0Uka+dgmX
PAOyONdqONJa/xa1eXQ27GhdWMLq0ozpzpZ+T69jAMlEfStYNMb4mURn4sN/Ag+t
yGjj769w/axGLm+UJOj0cTUCR7oMks2Mrd6eW5iSJkkkRkjzxKlhRj4EAP17dJTg
ijLGWLVuo1KOdl4qzb8pbgcnzI7ho412rBc3w21BXiBnXAzFDl7DVPuqpZRfBTME
3Kbgfya+11/Uan1jpyD00K40ubtOVD4/vLqFq0EPvAp81fo9P4KJdQ4F0Nac993T
40CMY+l9QRjcJ+CWZNkf3iW5X79yDHEIhrcaaAMQ4O0CGQJBywSXjXa/PnyhTnTL
jBKjF7o0ci5F/bVEOMTH1qq4lOlNMjb6o8wNTH/kw6WrXYLmILzvFjrD7c8+eD+T
ohZf6uGaC1L6guqmgAA6WrKzX6IwaB0XGUNudCmvlOqr4F/DfTZFOlVeoum8wIKh
ra0x6lMFpd7d+mJ/YBmZ/NLRCrITncEGwZ/Sgv/o1JtDJetedQPMvnpjG0weH4co
hBP9nsJABfVlCsLA0AWRqZ93yLTwsTPZ6ZtjkwcBPL/U6ArOe1lieNFGJDe/3q5I
ZwdWu5Y7DNtwiUzhBtpDDLfTrR8T5MCW5SRZt2y00znQwbLRQqzivNswoqAYWN+L
/dUpTHHjocFt8u33DvwK88UNzHo73JCYSl6ZeXGe3nJU0SaWVJoCb/CdWQrwrrvu
6attnhMVtH9XpNt2HhwqQ/Ndb/LhjKcP3TXZjLZiF0fECcgCs1GU7V/94oQ8IrLK
iu2SCoE/Kl1kH+iCHGc88r6h6bJrN8L1k2gJ0XBQ3KBVENcC6K7NEvmLTIgqV1aV
GDlODbuCBG+pYHxuP98PMSabrz0nEjhoscy9DVSXw2M7mjLEtpRkKZz8ascx0cLd
Jun/MpNtYYdp2fmoLFsXZAvsX+gKjfNJyIBi9cPJBX5kVh3hNi85K13ac3RrK6YF
cPbIfDTs36y7UWfN6lIg3BtA/jBIqofohGHY/vF1DStzpvd6Flie9kJCtAosKEOj
JQ9oUzMR4GPoiEev6AgKXgoLTasexrMxChnVZhYwk4gvuJIsYWLtQafkNJ9znMaD
YOi6yMcKOtH+sNR200Gr2I5oNRaYNHWQnG/MD4Ux3wHbNvk66iJ+vaE/wuRL7TCc
Uqj7zAm6H1wUHnEH4Af6vttPf4zKQCE04lb1XJz5kXrIcE2PLndHmQg+VUXjaSsE
Txx+8KE6kv+rVmdTUDCudXOtfmqZnNpM5OYnkgCXk+marzVIBWoGC9nrD9IFSG85
p1AQxd7fFfDJGQlQhhKyHjSKXox+qOAWKZmun3KGEEQZsoK8rGWFVgHu3jVxOpw5
tPKWMMEuSHU85bxFjHX5xm0T4YWeuGZYzk/sIgN6M0uHmQNHZZnEtkFbhXFXBU7I
YL3mpTxFZzs1g/C2LMH0gKTKFw4mb68Tn8ij1phcLzB6hVuWj82EsyoGO1xEyva3
74vAhDDGByYMT5VVsOIj5CO4PXdMgn4LB0n8NR5Ke9+o5fyKLSqpFdL3X7/225Lh
eRH5Pq5x3sdNlOfLPDGi+Reg4aOaZTbsp3CCrIy2rz4DPT33QKzErGihm5D4Ffs5
VfFuolMoNn+2iES51un0AjJQvA41+RfhL9SGkMbdGMRzvNbvRUgV8a6277ffhrt4
I7JWzl/4n0vEBVHqTDLOtO71T08IQz4g+VrxnRDQUA4oEVZ2kuxuWVTZ6OZcRH77
iozoDcFpcM+OX3tqjvzAplJJF3vnwxZCPnljhS6oqwo3SpZ8v11pnpaN8sBFOHir
LMNvRmyCD1BrQYNGd1E19Y8RtwntXYvidldcKRNLPKL64p6GoQZe116N7zfboFqT
HKqNyY9Q++Oxc7MI3AbYnsT61O1oMfLB0b+Zbia4JMp7+1cfNdOFA4F8ADVr82HB
/yWUyi6nBUtzhP2thhh9JUGyCAtcbhdMu8q4tU+evK+6l4nc7GOXv25tv9nJ14SD
QgzsLzjEzcGxRW9LmOixdSSCpnA1VHTNuqNaIQXOM/HXDkHw4EmKZHKwUx29B1sk
f8sxsg42hhZat8FiYfXpn7u7+a2yfC1hudpA5U4JKzdHVzNRW3BgYQA4yjBZqGap
ejtOLre5YkdZO84DiWrbYNX5jRrtdT4P2nJIYtb1IFmFie/YEvG4PgCemlUxL1ru
zLO6HC3/kmmAwa9PX/SXwVa0E6Q3kyxijIhJqd6RlH1LDm7ZU3REMZg4u/cO+Bi+
cNs3yIADEOq8AHHF1Myml+dCJ5pXN6wTAo0vd0ZdyT3gVpKu/5MoRPsF0Ahl8geB
EstCgnmgKfUPpTD6YW/uv3/5Q2NFzlcITkcpdG3F9RcqIM7pwQLur+wyjUg7iyZX
ccdnBojYJGahA4eBOmWBfelc8g+KnZxHU+VgAXtjZkua5v02PCkbL71JmEEy9F36
KmHRVTkHS5Qoj5IW1xPn378HJ6ywAV1lWoNn2F6TEZ2+l2lwdTBo5KNqpM6Gro2U
O/oMbtzrPRVg8NyB9zwjCGY8DsSWzg6Uow/AXsQLpTC2sUewPb5pbWpOIFYnLain
SvhFysuNjpszwAfmaw2r18RkEjnwJDlVDIGZsqIwprZWTozM+5qwwwo2nrQ+apIc
78va275MJG38zuBX3a/q2B+CihejMlJ7hG0fw6f6igpztob0RIvHcbV3sccfIua0
383Uab67VAloQdQ99pNUXYK6+29+qrZSalzUEYyhAKC3sIuVSxSwiHH6yXYOhEDW
J/2Z5QZvs6fp284CnIqXQKmhZNZrJHR+/iI9wofGjoKh6fIbpbthKqTzg+dl1z4R
YfrGNWh0+ozba/84t5pTqYbsJx3VhkjU7CgElc5/kTpu7QN+CdRcN+yneauGNWQS
iCoUWLOwLOap5+il+D6hkWRlssTXBstlYrsVMBODMTvCZ7g66u/h3xPfMceLu0m2
5w3L7uzE+756lE7Ynoz+oIovgcEaUhUhWNd/h3C6GLr8eX/dYfUXkHj1CQs+IDMj
AF6zFfsQazIOuqda1pWzBZgB60JzLEvMy1/gU5roc/pve3nTbW9HKQcX8z8UASWT
fj/UuVj0x1LrslfOvT/4y7S7tgFwDVOJ/Ep1YFXf8p1Kdj7UDH/mugjFrCyIAs2Q
HyHpSEL3Kyb5gRGM+2kE1w1plyY7ETpae+WrdiQC+M+pqavwk7oUceY4qz8XYKoB
3FMIv2wdz9Y4rBzEt1U2gjSIQsCuN2KpjkeEW9ejGZIFxQIiXPhB5tcNGFeSEdpR
iHYrADRgmLhlCRUW0qGUxrNVlPNpqk1ae6XyPZnwMySf/fFuotxOzG7W/1NQIok8
Un9EU6WbNc+zOHB1Ru32iyEk5txl625+v+HDe/CGnfIdSwi7iZECOn0OkH319Aim
Q38J8ELyhc2o7VEXP0XurXVJFbZAjH3prKztkvOyda8NSY61qwk/MX7j1slWIDil
Du+qD1bT+2qJNRXb2jxhx7Hhd+R/uYOu2KtNOdHS06FhMJ920u+gZ6Kj8/7pI2lt
K5nLWxAXUuY25ibTTeyW972WsKWL2y0vz60gaXdIiAUtpNx2K9MuRnd/fS7jqj9p
WzIY/Ca+hxOovu90QkaDChJCYTDmXtS38T0yzgBFlX0GJqJlwELWpnKT2tAjXfC+
e9SXra5/9HtVn4+5T8xOEkxWMhfo6aTT5K/DGWxYGXl6NgqIHs5WXSgJEaqUsSWS
viHwJfX7zoXGMvGxdG7A2EQEDdOlCYu1dsHBrXbjWnU5Bbirs5MGTCwRIEqNBxSC
rBo+MX6QNE40VJSDXv9JrSQzYf5VtMhuS60mvTu7IjgA/S9WOkpDiJLgzzHBDHyx
/Kr6orLRHhn7UxwFqyGzvvOT1GFYdBCfOXXWi0impmXctGRcIafRhT/DGydbS6U4
CUHTkmVLoRhiP4VzMh3asjFgYvClP3OkyVEcYcv/RwHjuhZ2joRH33XcyJMsjb1L
ieTY3oFKnwR3pcUKXgOsFCKh6k/XiLZUd01EXw1LJ9Q4cUX+vAaB2yGa+XQWWS4R
sqzMiAYpT3NnEco0b7h26KuVaDzGJf+pqW79iignEGb3YmRNczSksnGuPFfepeLK
CIbljDtfiZI4YdF49MrhG5CYP4CcsZDZJrnKjKO6pCsVYFW1QKRSjlZ9XjekfhPs
VuXlMpakBfYIzr2Nyf4hmlTP5QbZwZwL4Tovbu34f2R7S1fkKznZHIlnMQk7svyY
6uJ7/7Jh5gFH5jZ6FZhcjQTbg/RVgcJLtohhDJgHSZuAxYYsUz3Yjn6FmppVaNpJ
iiAszNLH2bm0ISLmEAdJ6f/OHVSNi8xtoTefgagQ9n3Yr9iG1ortoWwQWgZBXEx3
EsSTB0i12c9+OIMVrLhETwJZ2kb8y+azkOQJxUmej0E3rcI6h9aBlhMHbZXkKbow
NHLYdFJUmm3UIbOaJT+K3SAqsW44cBdkcj8TsLByPZyrJfDrE8ZjIrFcKD9XOSgm
nPGpPzZhFII4z5lJvyO5FxbwCLNmJlbbi+r/aKttwnzpgjlIFMsz9ZQUB7y0TA65
PIjwscQhRSnPnr/eVlThjge+XQVCMnHGI6wGXv/26K4CVVg8Ums9nen5WMCd6Cnx
ixy7vg9aeT0WXEP7kb+UEL+j9wP3E39Xb6Fo+eoTub211aijgFs+Pw6DPdYuZ+dv
lE5uE6NFxo5wRaYmXef181bwdk9VxxnOiUNnIbeQuU3nleSCkB3EW21vNGVkCQBu
d7seUGppzilSRoxh7jrhJbSaQxM+hKbX7YT+54K1ezz+efb3TIP1niPMN2dOUqyh
7KyVZzcWok3T2abNHuscqCDGFHNMSid1sMxeZP8HylSZc5WG7by72tUjmbtaiJF5
wDN7ZZJIyYY7AeaAFCd0M4O/WX/4NCBsph+WrtLCGK3BM2AkoXGQy0qMe4Zx9cWm
OleEHSwBqPsQYnbdDhQ8e5pMgzI5+t3Bl/2V5RmsGAkSCQnAtl5ZYPJsmlYprsfh
VkrUTMWlD6w8eM0IEAuqF8o3NiEJoq9JVp6BZSlhrJoaswIkLK3pToaFsfdE3Fry
vs2kqTqaZhSkjm26eNCHRxIzr3LbEx6TdCvjYNU6oDtb4piaNkJQLIscLfr5y+hc
xPNt3Q/oHdSlSBB52FUVGeCOwsdCFhnRFD9tbMpqQPuxSD8kzluXahqp/oqW5gRz
zPNIhUhCVqmJQ6RGCJI0Qk8PmwCOEtOLgwvPq0vOp/gPcPe80WRiYZF2rN2vaxdH
sCB9DH1l8dWwJaZHgyQBUVQH3fgZFbkZIeAlb0wwUvo21OozFJHeN12xSKlTrO6H
16aqvd2EJvlOQbgwQ4KV9OwMP+Bf58KJzHrT6SO5QPtn+RDjDYvIFrkLDseXNrLw
H5iOVEHy4z5UI6S4809hyUs1nsIZ0v31I/V+kr30IZFgmE0RXgnBjUAHG8PRcPks
gaIV665Dvb0zShWhRsfswOFzhd9NRyaQzyBsuKrBF1hi8/aCxKXiQVUCZKS8lIrf
+dRtBMrnw2wkta49ZnNqVrKX9dNhcxEoX86qb2cncY3PGBce/mFvjdlxRr4wj0XV
hGer22Xc73Umcnx8aSO3k7INj+GnUSLCp74zbZeGsfTILkmvGVKi1FWX40++gtZF
6nl1mXpGIe0NtUSATXFgE9dnebFcl5CwHeybMLmLmqAl5QnUk+WKEpbXOfAJVh9P
8Eb0oavSxNrHk7W8+xTLUlCBx4vmxAltK9HU8BYYRuKTd3nPWKzIFb9ZVUVNs8iG
T6UgZFLWNJFyHC7kalU5WfeyX7J43x/qVZgYhPaar8q2AUScnBLkSkhNUcRbSZUF
+tBr7oRFpWIigyGAmheWngjyBkrQHEbzPFewy+AijvOi2cDZWA6sGnsUenjx+5+x
ZU6yCtRbjMjKatVI1bAzitO8IxVS8ZAFcX7C980NArOStmrDeTDJ09ozkNtU6HvT
KINJmG9PbmTXjIXv9DYkyVhjecSqhoK29iBgV3EmZvA1l7Zky62w/vXgdKIknRXZ
dTFTTfhFOlrHxcpcTXqyVP3jPMHIbhiWyMJuccgIxz4rOXP6N6VSs1tJHBZlrt2m
JYG5I6MRn6Dr6ntoKsNX74vMu+jqHqmOubDu/xa+JomuU+K0xPLFC3cQybsabV9n
AKU48VUzh+RcC2ctVfbGRbEaJmjlmHCsiusTcB6ABU+sad0T/v+qMDOd7lemFFUZ
x6sJetiCe08fdG9Cxxnp2czNDEBLvsY5MoC+Exok/XkQUaL1c7uwvZiqoSxF4Z6W
9Rcicd7s1dHFlRU2zVmUqcK40UJzjGZvceEdFG2zOICb5WsY8wiD5lsIC6OyeXl+
Fe3lITzqHNayFWg0b6LlhJ91n+ehkIi138YViINemJ3/SY74ZDD8sMt9mMn/9Dey
XewHsPKSC6kHsTo24mWVRQyiXxMvtRr2PqIK8JTgHfO96mXkoKhmDBfL5qO/jzLB
izyy48j3GK8QimDZ9fAnbFkphm2at1pS/JxiFmynlraNliOYqODU/I//qj228J79
GGTz5TnPiBAP7ZTNUkgYF64yMfyCvhu7ZCsLWFzYknQPE4r/xYedlw/So19em+jH
MP7SBZAi+ZD5qWk6LhEB0WRo5wMBqtvDYi+1B5eEMo9QdxG+QB6LnjaCvx6Wk+L8
BRkZ5gawoe9HCRZyEhq7elbPEWaHu7dAa/8uhAegRgV5ktnwcGtHjfZQodI6XPJA
PihKafJORcOywsaAetNYL+EguRBwLkwJwhzFvcT2mlZ7LoWfBajs2XviyKoSwpWX
Uf5mQWKLgxj0CVevH13a0phlkCKqtApkm8QNJVhY4d2gpPkfFbShRwZUI7pcoLz5
vx+r3gPEuz+zYA8zgqR97Kf/tIpWFOdcFiKV1ReFtmi0wPnb5yg7n+lrTVOtdDnE
S+OB0iHQSJG9/9Wm0ZLrRWvi6PpUZ+pLtZLj1SR95UIH0FdaXHsU0tcTBkeoKFwN
YEM8Y3dTLGHQHPoDjzvUBKO1y2iR+x83dDTbX+W0LuwIfD67CbB+QqwYYIT+LbSf
YAEE+Wl3FLdOJjUChvkO4UCxB7o82/0/XcuhBgSXB+aOzduqEAeLZjk75bE2Ft6w
N6rYXYt5MqnqjQsiRDRXmLysfqKr/oFGzBIlE0XeMWQKKYrRS3Fh95iXHGYc/m/4
IvmmKTK6D5Jjiq+i7akNr+pDgXVi2Mej9rn9jJhlr9swCWcVIMSKLCnLSoDal0zg
JqSbsdpL67qLsaTZN3Of7mBuR4QXPDmBPfbzEFoyMeqaaKQ7em9172+T1jNQHqDq
k7NlO6o8m5U3gwrkcDQW5QCsSSRWYrcPv6/ncrANvfmmJF7R2nLfnWa6xGf2ej9X
mjsKhc2XEMZBUTThs8ea4xqISC+/HebHFhzDagVFtC13BUP3bZBwe0qKEsjaS11A
UMn4qSjvP6MgSynvqvOrR+SpTRcZ/mZJGQIzQuymfnrTny1ZR61d3WH2P2O0fhu5
oayQU+i8TDd/eDjTFfuoBUdKhrv57xfA7pd+FjSh8H68aAbHt7MRBVDogk7yZrQX
2oyyCsF50BafZdZMvAyaWeplT6ckYN93wSWTwNgjs2/yxKX64gXMuYgUw5y3S4AK
C98fEAQ/v+m458qG/pr5aK6bhdhP+o2WKa64CcFC/cnnhUiQ72vQMj4uKGurd01O
tfbosDLDo2T1oldi9jvWHySVt4vb8qzztrEHYaVHcuntwDtUi1S9BdBiXRm0R38c
4m5mlk5BkbhlN6NLTLoG83CME/xGRYyKSY4bn/imdLDygkhkKKQcmvsW33vmaxHD
YMDwyb/M1uQieL4aS7lNx6LoL3jT/oP4e40FFxcrkQeb3dqpC8MuapFj7raH6qpX
QXr4OnKo2MFgbSUUAHsSf8pPiamXnsoGecR2MO+VbLikTvKMVYJSxoK6jpx2uIcJ
HR8j1cc/HarxTTLE8Z82Z9CpCY9Q3mj4Ubes5LLoeUygZwQ9I4k91PkwXZejaQT/
IOVVMskTRjmi/xXlExQwhMWlaKvN6t9sft1hJdyL3VspsfnMMSMkS1ltwL1jWf3l
NRQ2vIzezIa8I9XHWQD9apYZLZGW9ymjVddrBc6A9Tp33h36KKTRrjrRq4+da0F3
83ilXmuZtqmxIk4MwseXRMP+BEb/C32v0JzwsA+BvMct0Qq4co2d/BDtGkZ5z9Yb
07syAjmUDWhhkPDPn6FRJBpRI9FZJ3BhXMC/SXpdtQ/0GFX0GqDp74MPyolUqkvD
JaLs/+pAp9X+wR5MMcDlj8lg5MADQZUuZIAcFvY/J4jtDVWdUbiWfBBC9nl2c+x4
5uZy7sI1f8nmx/Dd0HoKLmyShaG4+5OHr8yU0nHQX6EGLHUrgKwRhe/nQrrrjQFv
zSmeBIr9zHOpR7bs2JVxOAOAAYIH+GYXeg14SekI/4RIm1dqzHog6OusVdDBmq9X
AzvvsR+QSKAV3z7TpHDEUzq+aeNsAsJw1EUhDBc4wZH/j5/JFYaQ9X3bhyBqU0mo
0mImuudY6siv1ImpnnZg6eubAsGyEa1yNy13ODdhLB9HBHH5WwB+KjekLlEkxW2c
o3DlO6GUkIbMMR0TXNsGF2Kmt3ViyY6Q5o4gS3x3jByJUBJRUrdYbeo/L0KyH6Mc
nIOZ1NQ8FccSI/OsG/LCgK/S++e8KbXbPyuiCuZkSTW9fOJKlGCPusU8vfTAJrqg
7IzsVabFIhgslG00+e3TGD8Kr+hWOTcLMB5cuf1GnUGH2NVe+gVYgAtPhHrPwBnj
t2O56kUdnz0iFw9nvcbnrA0DtmWV2S25gzI0dtyNwXm85c8LaWd+Xlm497VhJ6nZ
hy464QGJF5Zt93aPx5/D/XWruhViJ8vbwuBfnC13YyvtmF1dUCUzwDJdqLl/JNHr
SqcflpTeCRidwWqzt/As/ZwFycHyFxLCx8YWOBjocmW+jwqY3fJpShlqygzc221+
OAxyYSeJE920zRhz63VgKKJ8e8E9bgWUSnwJTYKjdZshoAKAS+RZh+BJs4wLLlpd
pugdskoCur0h9c5uZqfjqnuOq9ueKr1psLr3EZqTCQlKcxlWihNxntYpA04EFMW3
by5wLcxeql6f9CS8rA8CmtC3cYGdbQi3p4lXtP0WaTwG2oA93E5wlEEP8l/3T+Dr
q1CeMuuLE9JFyUONNbCfpNEOmPL6kS3rZz055RuZB/U508deVoJYJHlzkd7EQKGm
dlhKxUV9b2be2zKawC7GFqfWHKtGrKWWir6uEvqdmMG5RvmClZOpyoJnj2aPrP31
O2HW/SlI2MKdMbJGOrT0/r5lCka0CgOTVjaDzrUqOZfvTcClMejoQchHafZTmwue
1IFeV5grCWBhTnJfMDkHZ927RGqctHFs3blD3HuMr702rnFNras1dSC59aMMjW4P
ub+MJZgKgI+TKhWQd8MVjAaS3P1Dl5EkpEPzz1klHOl5VzJSNktwz1rNqKGnulcV
557Vy7czLsDZg/Jm7DGbpAx6hNMwTVnFPeJYj1HKMl8kN+IbTVUYmaSVpkZ1LJY1
ka4eC4l/IEZCUZPi9W8wt2n9GfbKAvmBmLu3xz9TPJB7QYVAJI6b63jFE5aWnTKx
LaJ3/DjHF5ZXdD8Bj8rg01gSnSgCZqTBVnKDV8Dd7Zo+U5M1T49H6hRr+fmAmF9C
qUxRRvsqM+jnwJUc+30dpHqUJ0kktGHQlc1fT5CKjghSFaOqEn4OSv85NQz89ZeD
iQv4ntRVFcR7uoiWROE9Z+EEeLVtq5fQgo58INsEkcgXmAtNpSIfon0HPHIPhRUF
ufkeAj1+vtDaxCU59Y1GEdoB8SwZHTyLHqERRQhUev0vXnNxQ0yQbCTNJ8Ga9quD
g+zZKigkUc8dIYUQ61ypLRdowvrV88a3IIu7OBY29nLMvMw1tnUwO9kLt4hAyivi
ge07HMqV+2E2Vljh/zswuerOg/aZ3JU3hBq0WQ7PyHfSVjAHQ5ZJnM/PLe4llame
tCsz3oH+I3zdmQPOFKB0dHGZlgPw+7iDR/+bKqVk25+UqMJtYGbGypcmkPk0Gs5J
BZGa+AEmj+PHg9Ja9Hv/xjPkOtAAR1LEz4a8HAfWJHJZTmQXGPR/XvTo04UMjsjJ
IPHlbqJEAK9gTI6w7w33awCXOSKN18uqf1JDZxiHrJsIMCxKaPzkcw3gMptZ85F8
PZVIIsAmsvx9DaUwD//phzo5J6kuwdWXvBg3zU6UOdyZPMLY8zJbgNIL0oQrwnxl
/yDj3D8QnQGoHesDmvL0NtZdKYnJUXbqG8BV30GEEjt0NTCPtiafkGM7YbXdArR1
SrmyGmC0HCc1WQoHuFzYiyfTjnh4e1ytkNnH6F5EY5TEUaSVTfzi+BdK/Xu+lBbv
M7g/Xm04YEbfbuTBEK0OD+R6o/4XrcynE2AYAgRH4+ZP6HuOplSQ61LKWp5R0s45
GFhDs7tr6EONWA4rRItv84k0q1fNnNeyggBp9v3UOKcrHcyR6/Y93k4C7GCScN7G
WB3J/DfPGm0z5aj2j/3zA4Op+NjjMCukYpHjkYhXCLD8pISNCA3KrzhrCLsQCDsx
05zl/nmPnC2m1Nk8CrZT6A7JBFZhLeAG7wZlsFQhBK70Al2vxi6zVgyWIuh2dtcx
+s3f8B6K6xg1xfpn4tkfLHoRQKF36YxOhP4TE1dmOCnJkMrImb9pMLQQCIN9ZJf3
+faYVeaM3U2eFA4wEFddX/t/HorEgpklCysWSg/GCN4RAtI7dO8Hd5X5RzKmV4XF
wWHSyWB6pYHTUBopATtkBEmla4ZUQiKkF3i6+zScgd8eqRS/BF4sWLFrqeHTBnvN
9bJcxnlfJP/7IJ54JKnttuynRQByfTQDLAHjd4RBajZYuEOlj+1UYgxXh4XRb5es
mulpi6XebsXtXzfDomJf/F+Fqly4JT90NjayCjV1ZeX4NwlJqUpL5HqTKXkN/vAC
XJlsWlv138GIRO45p4Kg6d0181KXYYZ38hhtuCzz7/kocHC8bFJ8lTD2eYW8vPl1
Bech7qq4KZZv9YlaYgbFhT559BBERx6kgYuEJaTCUlpHvN7Z/hLOalGqps88GVC8
2ahAIX0/nmwWw3/fNJZ5nPiov0+NL8t8rq1SC9FGriGPQB9L3Fp5UuRM7zsYD+i2
DdUeiyjTW/IAq/7LlPTlwwNWEWqCaga+/A5aFDyIK2JJ3/oW22qYjGJNY6oOYEee
mjlTME/22xh7aFHQ8hubrR95OVrY+ZStRFWDZ9jkwMloptABO4wBA39b48BmNrfQ
2YZ8jEGLtSvQT7nloOum2mj5O0bgjsiQyxTcopy6UjEIbUG2EOYyOYH9slSX/FrS
DRZn4heraow3L9wB1A/JT6xf/hh/lCuyTuWe71VTV7Za0uff/GoslinAqV8vxIEg
lIYNgwxTwAFJUXJVknq4pdy4xLZOA8Grj+wxSw3mjgtKe77QakDHfYT3iTKKC5Z9
wYgouLWFCxMhDtyuxu14XQiffC3XeBiDpAXMcyUNdQ7py5FlDaO9hjr9kspzKt93
r/g/KNbRykHOXGYwDPU62InPb5BA86qgTjbesvgno+IfYCdLhPZROEuiXNB61sgj
BicFrlWiG00imK/HUocRo/H9FyO59WayKP7FF8eWkHJQuP4pbhFLUcid8vrNoCUc
CtEtCLUBQwgg0LbIstfPxF4pKoibSigN5YJ/6+az/hmiAFLSDiQO00lJivANUZhN
GOEwRwlMzihAvAlLdtm7bn+tTfiXfkynV/TuTHO9kWhn8mI/fs6tzaTG7vvUQ++8
i0ZLzLX9xGszwf2MpNEaXM+4pBDz3FOWacP4ki3JrCg8Ff8cnYdcCYVms6jIMRHU
2o9r9rx1gMt+nuzB6wNUf+tSD25yugA4XBT6KPrBNzWhqXXOoosUWjeI1YiZ8p/E
y1M0r+aJQ2XCba2fE/Lbj1tyzKjU8PudVYYBK+bkK3LRGnFN0vAYAA/165ms3wE4
595On1IgNX6arQp5SLtup0oJT5yTWKweccyZB+cEIE4+wtIxA3xSb/5LUpLCDV/n
CUsmfdh4TNwOsH5lkoa+YO4Eyd+b0deOqLI7yOtc9go6r5ymk9Pb0dnGjGhRIzsm
SYUa/6weSN9cILz5HVIyh8goGoirzECY1Ok+ZvsuhmYeRTBbDVb0+7UD83RbnRi3
iKSR8VGgtbOqBD6o5+wNCDjk9/D76J/3D6u9iKJcjXUm874JssQ7mcStlXT7Y3ce
JNbCQj29Kcg9MvZDuTU80h+i9E9r9dmKAASJWa38dCMiWKdkzc2dQ8XP0+X/Ympz
zMglZODs61UNhOll83AOPretOteUvzEoWKhUydSjt7wQ/v1KU6BGMV+QmQSsif0k
GycGQ3ku6tP+wS0btM49l9weO8JYASIMlH2dzvBRNTSh5aEZPzfO8L4+EFF9H6jG
8f/KQ3IeJxizdHVPBOwsKiOaVodgiHh2Bv0TwSvaN3H1X8z+aUahEW/uCYJ7ea5G
2WZa+l57GdU+lKlTxbr41G7nqNkQaWNELrrX5zXLmEZSyZ6mHBkabgyM/8Oiyx13
BhRy5MojsnQYSskETTTwHGz9sI4NndNQSqoxjTla6VYuaBiXTNDeV7sG5taUGSPN
Y0pWsyhU37kq92p816oSEuNUV8JkkhhGCojtAxKxgQAomBgfL7IRkoE4IGuUnl91
0wiiPFHBEGnaw1sju+2Zk3iC583vRmIZXGqk8Sqous+i6VFG3rGcpb1+kfjsWbyY
8BY+0e0lRXQB44O8ReELq/M6dBYIO7FjwUc2iAIrdMTqWfq4Tm0vb/hjTCCiJMAw
yuvCyh27zVpasfB2Le690BIA26RKLheqV+k2qH4l/P87I13nmtO0hyWgcpRULGA4
YYHaOZ+m1h4CzJx3B4gpDTmHomieSwfrxZXFHej27x7AYm4sNd8uCLK1gD9rrg/s
ddGSQ3FUH2pnNwBJll8wPs8NV+F+sM3kEzW+BCaVEU+f1o35E3EBc/CD9qk9An3v
gX04FSR/Y+LeVv7TiFteAdlj9GmBoaUh03oagBG31UGi0vehESZA7GyvGLAxRJJr
gA35TWzcD9Y0clNvZVB9NuIVbOEQcZB7PyCiH8GD+Gp3skHhfA7mKFe7QEEejM+F
Lixjek7V3+kmSzCcP4aywV7DiF6Jhx1U+/6UQIKL6F0IevKPWbV1lWVOz4NRwkMq
bzbEbT2BSgICJEc2VcqFta1eXs5DI1fCgbzXgP+PkI00V/Q2AmPvR28norgmBePO
BLximWgmuevoqEGIrX2xPHKxDe2gkGLFcEKXc5RENKEggPpH/odrFeG5GV1fzLEb
gYFeqC8hS597nqMqTSszRhwwTlQ+FrboUFcuxyIQ1LHVZou68W+XWV6cpA8i3HTX
FOJBvY0wXNEBqQSvGDXzz6dbhRXsehMGwp6wEaZDkZ9t5QF4H867rO+CS+DpUAYx
76hpZJiGdHI3KmfKfHKz8M2BSZucglbTnaeug/k4DlnL/s5C3LXcuwsD5K5pwomh
bnR8a7pMxSvC7rB+Xn4U9pwq1v9nHy1hR3G1+MG5jKmFo57io9osMxk8g6vOBLnv
jjf0WlAAdqcZzhDE7yhbkWo8YuRtVMh90BpIjPUNKgR9bHRPxFUuQl1dkiOpUuqn
fEaE0bznEIPOcgDkk+wqLfxk3zjbjK3kgOcf7inoOqLFNIKChiRPq91IxURvi3XG
TiH8MxLdtS48U+ZByG9nMFXmHukeWDvRQatrOm6x5mrZwxQYUw0BlHRg4YR2UYa8
gEfKQt6JRXndO9V7jRCk0z5ke1WVWmWOMq5TsXvGQOUQtUD8zRWUsW4RCuiolKN4
T2g8yhCnUtXhFDTllKFUuyaSRt6r37YzBw4+vNfnlgbe0t00FAlqNGj+cs6XzTnt
rnQyt3xbnEAzRhXeMoJ6OyBrBfqlTtL7PG5nCWy+l93fVBy4hnrWCYaKYGgn1xFr
0epjugRzf3vRryHifU31LrpUd6e32oIVBVyHjXFFY0ezpFxa++BGZK/CaPkJkALK
kXrvx4OFqDLQ10aQSW7Am+Gnq74JTcWIbXydpQgx5CDb/jQZMFcahilYGhieEnfg
e0Vj4Bwsnhyo0hP5N5YuEp4Is92RBaBsE3TsW7kAQa43N0jZcRMMLmcCQx8Ci6SF
ClA1zBf4bZZHHZX7wRB7fHRmu1HBypEouBPjfNmwE2pA4Ife8eV3aq0L2gh7lQ7A
TI6A5hlygJNnuYFfBWFaQ1/FZz04R8bVULDQhQ+vTdVCAbpg8AZiNHe71SgWfqsZ
WJm4rQevaZZhVRlkL6vjICMzvD6E45wv9/MIE519F88ZMgwLrK50VYlvmF8GY0Vh
C/cZfleRk7FMyQ8OhNWPkqU5XNSJzcAZ3gCu02RC3aq+FunG1j4jVm80djZkDCZB
8iVBn9FUy6ooljeFBV2kpcuD8eNjmE6/oEObkESLVnUNgKGQp9RSNRGxjOWlvPib
KV1tzLHbxnLA28/Z5EXy32Hw8zIn7arE2ymzsHCSjSfsdQ4W8nM48cfFORtTEASq
aVe6baOVHOer5AlIHK2ZegkgzD7rFTFC4/0zb2MB99AcxU2fcuSGHpjYYyxTTdQa
PkDvHOU16rjmVWHXgFOhBgP3Ity/jdt2NtGQa1Vifv/WYy//e6eHw79wwOEvIs/Y
Lqm0NTRh/5mXd87NEeMfnt6z+381Th8ATCDtOuDKgrnTyeDEggR/bfCy94M9QUW8
zJe9Nbp7SU1tNCPZNh/N0hCDMWa7Dzn/KIc3aJUv9lCt81ncAfO/4Og1WakJ8Xuc
8KS1CH6sisCss4tHsYBRZcDIpjeI8juUGB4fs2ISLnWqNnOHcs4O8KaYZjyQp4iL
i4VdJkyCppF+wYd2bKqDz2RZLhwHPUf3PMOG7wjnNN1+I6vnwdvFoWlgY+5LZUV2
WC+Sdze6UPr9nAfu44axjRm+qyQjdApz2r18vwmDOiVHZMeveuMbrp+Io6OTxMs9
mI6i6uWnMRhhY1l5a/lIQFW1xnybILccxBA/Ny4ifLcpKIdE9CdsPtqjjrz9Ovcf
VTwZ88ntnSW/kdQ7I9OUYchGjCrMlEfw331kY/CElDUtQRDDbSwDB1WPzBKFE/cO
gfDvvxVMQ0gE2WXpQmjN+z1NrUsxEpaKVwbK7x/QNuvp+g0ChE57akydoKFU65Vw
OqZtMFDRuRcidvBwa+rb17rF/aD/ASu7QQRlNFchXmVQ7GO+tQCg34Oag+24X9mR
VQdK7m0t5EJVTnJSMJF5GaJx+rkRn5IOnnauTB9Ou3Nn2l5p8r4YZzCVjprfa3/2
5ms92B9Kcj6n9EkYQoq+3Vyq18Xm/ed1Kv6OnTCtgAjLGremRbzQmfV3m8KYYIPt
TCwwc+WpfIr6A1HQzo7CeCt2mizRseDUN9bBQrKKJ2H7ovumXjk30HK78coPNg/D
IvbY5+W7C1WSFKItqkjht1mLkp3u4gXL/W4WkI9tLMl8C2vf653q8fd6K5nb0EEm
JjLtb1+vZtQmtc47RrfXz22qXCkxAJoWw/wUIjlHsrENONltUjyzWcoot6lk8CVy
LeCdTBAfJ8tG69R2aIykHqMQKMf0rd4rGafPVxuRiUSXK1Mfhun4S91hlgaGaBRq
B7SXsbsST/0S9bBJEJGStrKhaW8nMjZrgv8de8h8oMqLLOjUD8phHLiPhJ/RJKbW
frXwx2wzJQjN4zxvyF7xpWRRZXAz5/PHat6xKORw8zZbMcWiIQ8pF29oTgfclNqk
Y8YTu4/+Ewk6MClcuMuHaByxEYX0QOilMfkxUluAvYQD4I57rQXntnx3Ut+FN3k1
MarDIH5KN6kEZ04fs9+DQ9RzhakovYI/VuQaKSlsFD8d/QZaUrhhCNeAwbJ20KYg
KEIYw9XUVnId73fo+rotReJU9W0WQSKBe9IF66GZBoponlYt/h98LEHPrAGrNsVe
IVmN/yp99y/NuiVM9fRftqHeYNcOrmeLSapbSr/6Zv4MzvAG+yWJSNcDU/adOXQ2
t1i2CfY3WWueSTxREE/OPdXjL6NVP8jhu0oOpql6+vb7L78VqgXslY6T57whFQHq
qah9wk1oFsiAH6qWIbczcf+HzncUgrUOumNG/FeSNSxdKzLHD5H9SfsG31P1bF+C
pXMCFKOZGZtnAZPaUiG5gJZ1xryFuzhysXsU3JF6RPqjPY23r9VO6ZZ6aGUBjmDM
M5SWRXwu/9tC+k0/qSSEI+CkCkHqG0QRppocDmoKFWBUh726urjdEtnaLiFpSr+6
guPV8on4c8/3CFLerm9dNJO5h74whPaxrRqWKnFMQEt+x7X5kKRMOzN4VXoSLpQS
5FZa2KMd23IzWE4mAJ1QxwxSjadETfUwzE1Gyas+/HF7rJj7t0Z1VhqBj2ES8ubD
sjz1ZH07zVgmLT3sQK4ce2/4e80TSsmV91uWoTan6fdEha0pr3pwTf7zdvKaIfsJ
4D/ZkYZ9QDLR+t/Wu7nKzBM1TEdkJk8rFoKLSK1v+2ogJIvdmbytB9silAxBJ46K
uSJ2yn3lsB7t/oHyVn7D/npkvdiUpIkJn9kIiUtKNG01U1uxt5cI1GiWk8KYV3pP
QMRbxnkc6yIsd5bkCgvXZ/3GNBnOtw6HAhr0ebCf5q6v/7bAgHY2rUV29BDsM4DL
BKs2KyNHXjb+ZMwswpecRv6rOuskqzSLDRt2OEeAtw/DM8lHA19TZ0N5VEML/Jy3
6hW0rLid6IiVa8UimdftX4Ku/NYF4AQ61XzUQ1+/bs0KW4GKx0OQvbarhB9uy1T9
wRHtwOsMJHWqyKG6nlnzSFAz13IkdRRCGccV68qxXR30+gepuQicjyvLCREHUioJ
1OAlzSuGvQuqqRiJKf4m5TePVlCowb9d+UwuWmX7Xio7caaBMcXXfAPNRLZFhi/m
x/KznmpV5janVOHYZf/uZj/OU1V6d3mo6086i02t8QfLw5vn/Pc3LMGx6tjBWO33
nrrczKk4pYMd2TdWW8hsPTjdbQl1qvAStQf2vNtBC7y1cThS+Rwg5jmwcAuAWOKJ
mE+/UdJFOISyh4wBaFsZFlDiUazEeJywUH31QshvGONCjt0wGQCwDHgMV3OqjxK6
bv/zOht2+8wVGR2H+b8dzjhTpuECpE2RE0MKqBO2trh29HfcIjqsjnba/VUMq4VG
nP2EUffyEO0PUQ+we/TDFS3FEK4lmLXSLbGFZMkQqwYM8c6k8AUJ3Ka4pxXWWzvq
jtqelpKKzQPpqOCKDbzLnFr2Hs2LCaKwXbd9L8fXMT67Vm3Dtv0ZCikyRIT1XjOx
dIvwrQgSLmLLGk++6RTVojsLtgegdxnTJAahcSxshiLV9FAZOIvac7orTMMFx5m+
vKW7V2k67B9yMrhh9VAzxziN/u6e3ihPb8cuGz+2JaHAxMFMnvbHr7dJeo0IsntA
lAiTZVy2EweRHJfysbh2Hr4gcn7iDyYvp3xGNbRGbGX0DlieYJ+AMpQs/YWMxa9G
9phA5FI45uP0Lr6gaJKBhqEbD3Gd5nPIUqDIJTj2hF9p3vhm8tIgFOCygTUcTLd3
f9l0Vu/9oka5CWbHQW7/47Fon6UvnjvjTcQTY5rLuhI5dYKk5+aZIGhhgBVqosuf
cke/lbu5t/q9p19ws1F6tWwqFO/pvMpXtBH1LQO9xHgkIqFIoJuKawwqFuRgMYIz
BCgxTa8Ur/QKCCwbs7KoXOZ9tmNsRJRMB1TLnY7yIFeqgsXwg0r8uRPiHH/F+ZaV
iGtbyNsl8QbcFY6zLzzhdTwjxQItVxz/q9hdMOCewH4nBvFhuMJ6n+cCpFH8ro2D
lR4/PsNU+fvkHQcmCrOGl5IfCOQu+KAx0tw/pC8bQCpqHpxLYBsrgd8k26UV9Rys
L1mGs37T27OGeYIu9IsFvdN3M9AuC5pTYu0+1fMZpZO7S5N2mfSYmw+d6NzsG0MP
9h+uRE2LbRghwus/bd7NbTKXqWxaDSsRDE41aq55uK7idmABh50RWDmC/ndE9Kck
8YwcX/lozEKZbMlevogHGqh+OVrGH8IooOAw0bDm25X1xVR2e5/lMNHGbIkPMtfm
whpvMPYk4XtfQ3xTVnmFhhCKmZRG0RgpmQwp4RbM77PrWRW9mSjpJGuBCsSA6+WD
VLXxA1ebR5ecIX5FiIEXa6neXJxUqPKXZZiSOitvgafe843HERaD9rvspb+ftFi9
3y+FRK6bKu349d5usw5Xm1pQU0CCe2cov0v9Tvv7WJCI41NQOn5RskHzvmbK+qJ8
MsNk6YCPlj1FWcX4DmRdw/4ubMV04hMVPP7RX45Z9Lua/52KjxVcDsoOAJ2nmjQR
FGVKt/n6Ch7aUtLhM9ud13SBE25kybAlQo+jqqUnjBWLBWgmGoPPbD4ugoVEkOmh
KLfMxW644FkH687cvBw5BFuTjx39I1W2tib24OoGuxxPhVqoelq4QhWKuzBajQWz
5urQCcCTfBZKq+HvroF7ICDXFbLBv3NQsfGoNNEBFt02zAUxX79CMZpvehFUj/k3
QHv3cLpj9bNGRSTyc0rQJ6Qykja2Wvj2pTrJUQGa+KhjioHPGl4gwXlduqQ+Xf0b
PSe9VnhFuLZjLoVclvXZ7G1VtaeHnvV3oR022/TkEuZz1jQQbuLMH5Qo2i34g1KY
NhRvBClLY8H97oPCJDgedNSouPmVFTVL061/QAOvPKRrvEeO4y+B06H0/1atRcZO
sPz6mQrBfoRvKPXh9QQ6UGKZOMlG0+Mu2Wu2CCLSiAKMHIfqBafmruUHZ2aat+sD
w09pI0zMtERVpQQ8Rnvkb7mDOJMGsJCnns51jmkTSWxwRiowBeEUEuimI11VpAGE
vXwdRF9q3IUi/tMOslwuv6W63x9D5CRbkMwfBSWJKQ32RSU3SgOcbBxfRso7W5nY
B/znNmRfBWbWBFPPl3zsn1EFr2rFZjUPOaZ1ZpKaxSdrxCUv6LwnZN9VXKdZRIik
hUK58exTq33HItxqxgPI/MAhW7eRBoZQjrKYPJIPE/+a6tbafgf1A44i1bgoR9xL
r8DCvuGFDcZHAVW0LqfczMyh6Li2d7p3psQC9r/lRSuH5Cogp1LO0JcLKbp7ARJ4
NTjcEVdCKRomQXoa0Iq9VxG/l2eiQIXWtYK8umtRTV5rVOKyQZ+txSHC+8ibZxGj
63xb40jwNRRVxhemNQT5FsNMqCdUtWbEQ6bArFPdGc/C8SGiJpl8y2nwdE6lQpfP
rJcPXo2WZkksYZvB3QvAYWVu9IfzFbjjC3puOp4JI8LP5QFsAHh+Fw+A6039Gl0x
Hzts4DhyGlW8Gd30rPPGXxGx7Dg8473F0eZmtEQnl1in93Rv0NgsXKmmHp1PVEz/
Ks48oV7/TZVSCr6jSJeDsiX17C6ohalVb5g/aUQzBVLX8A66qS90VL2/YZ/Vgr1Z
CR+Nb0+0mlB+b8ILJrIXj4xv9NiSfiyYl3y+1MBv8Ur8NPoG3a8jZ8200VeUxwUY
j7C5/cJG4dBgfCAHlpPdToG8vfjY/+W3baGKJK3Hcqj17CUNiVQN6NjmR5ku3Puw
ja85h5mzfMxDHOSMXWokwV8Bv7gg+2s1yiHCnrgMDEor0Zk6L17oNN/UsgF/NEwJ
OtYl05cDMyKUiyMpd7BbP9jv2rDxFmAyipzB964E89nOI3AcsE1SVhIVMQWWutg4
N8l/BtPnBPR0ygnqlK4NcoPMKXQy1lHtMcOW8UWGxyXh5uNl57knQurkgIHLxxSk
Klhk64LbFg9K2a4NraCYODjZWSevbIdnLVJjD2EWhYr+jDugc3pSmseyU/EF0zYV
6GbS0hyiMzXnX9KBWSXdLXCxvLwF62gRYJg3+3mtY9fw31Tdieb1r3J53yM2aysK
5urKd5jwy2jxRY7P7qTdVrZGtWIkeiuZ0q+doEZ8+OkkLgmKt+wNogEn7mu2ME+c
4hX19Bd/C6+7Nm5MQCtJ4zOXXdLQhrHRIlRVgVbRst6QvVmbwIzTztvEIQ0lBvH3
9ry66eF9+nS3a0vyZAOLJUwhmojl3hVLuWqGzIs3U3hCRVgaHTZ6TwO/VHGN9eT+
CGaUaNab+WncFSgZQ9F3g+vXim8/FrRSA+8cbSOq+hYkEy+wg78xanISmuQUlOh4
4ttoSP8NoqANZjM4mRaSl8rRYuxiy+c4m2RpR9WheFonudwhlLjtXbhgPtXAeGnW
0DAwV8RoLptpX+ViotPZNC22ZIq08vnsVxEAEm+Wz/PI6yPlLP2FDLWiErePXDY1
JWLV70HAX0S8RTj4FhuqaMYyBo8lhyZsQJZiG5uR6Bs+HscQPB3npujVUwZbuHe1
/Y26AM7r7rkfJ/AwrByLEftJMetmRP+c5cGq+XNAF1RBpAUCaXbPAhEr5UeIC6qU
Msq714MuNKflAaDSokbD2iwyFNGxhDWbWtI3E83qWmoQWNvOBTyKNT701M/1LeC7
lx6kr0oGV5zjZy4SLAfmUF/tfw68jKpvuy52XsAtcqgYgpAi0OJhWqB20Va1cTG3
Zg44luxylDiIJchcfWR+aGNkR/1E+a9aj5BZ2FK81uEeTP03LMZdmk9APk9s0vhQ
DyiyPw95JjI2ggw3qmBMPwVI134yxAp5JpoBislhzGltEnNcLmDpymBjGedZmlDQ
CdTYlD36BXZi0P9M4NZtNO9XoVVR5TRUq7/NQvTVAJMgvXH+8voUYeZq3j0Bo01P
J6DmW6FiTAUNFQvFdSxYT6wjTSWqdEGFcx1oPTTknxzpdpBwRnmB44RJD3Z4tVHs
FXbcqFYOmNeoE46ZDmbsXao4Bj4fmrVLsugcO+DhhPXYnMvDaRPlCqqBSYKspDKT
AChyxU9i8fOJ9wlGvvyB05uZAmg80kgR+SSyxjjOOojdigDnkQlEDlVh5Mdhb6MT
Yo2/HDwgzyyVx9jU+nc2Ui4axso3NiEDsjc3mIIDfR1oeGaPaHZ3RLTK1LAuiUej
eIZRl5xXKKmqvAlsaVNuqJ9BjWjZcd9lZPz8tS4q6mBW2fAN/p5jc4i297eElwTd
2YypBTSRoAq/Cpkqui93DCOH6G7K4I5TmvpQT6S7Njs1tRt9nDC2juODjp1eX+zD
pGtNAg/Fi1jt/6b7UInDho7S7H55ISV1etuFyHuvGiMbj/2IDybYgII3j8WJaT/Z
aBgzGu1kuRgNWAI/UCFgW5aZLqo+T6DsKt+ymQYaO9onn2dDV63exRQmoj3LNO2e
x+YMgwPcexNkk6CwT3E4tmg90HMunUTiaqekHAwwMFsQ2+M2OS1XGFu1+dSl6YR6
evDvZGmcoPA0T/xxrnsBqP2ILoyhlZhfhEAVpHMU14wcMDAYWdXedps3wB2Tz/du
vZEwgzsc8Ekvo5nuvUq0naKrTdq7SwwSABRX9AfIrCRWgYx09JEZtjJFkpx8Su9q
kVe920BAc4GPMgT/vjwl4M1OAcidVX18iI0Q5+r/MBmpCagGZtdpHGnOo5aYyh8X
2ENvRfDB5OaoW2utZhF2YqNWL22lU2MobufXDjUhD47T+bczTuaNlG8qkrkQILfX
rKwwgPTmWxUdZaN67QkrClMLqmxOm4sdqdWhDgriO9ZXiQ/ks2uSTaqwZFQ3WLIf
g9s77YXZ11N8fmQBFSQ2Gz6vFoQSAzC17jzr/vSP/AFLwJxz+rAw2JCDwCsVT3tN
vQ8B86b4qmtpDk1cj78+wW+bBSDL6b7qxq4EGl0D/5fxrP18/3kvCU0GQvZ7P+sM
OH1TgYWPbo2AzYzShXoppYBYBv+VcRP6sWRSdq1mrA/5pupdty1pC0EjeYo6x9Zq
Ob+R2QTJGL0+K04+EzRVAJ1O7WjIN9wxwuA029stnxmVN8uTckdIdT01KtqjTfus
J9h+/BDzTWwituut1y5cIO4f1J5Ryd8ZD9C7E9dh+UbDQ0KR105ckcEwV8ceUejo
RkJql6Cwna+HFH53DRaCo3BQiJJEhr4z1kAV8U9nXM4sKhyMhf7/X/rThaXRaM7v
3rkwhQJ46eRfP4GsV1MXzivzSuMwZuonBCjEYQS27PWORro8L19Kb763PtTzSKYn
xvx6ZouwOBMgqGRDKaTlz+TLmrcP3fytvGLhrjXT3lqvUV/mpsjaUvQ3oJHSG1hP
dXlcWPpmMmnPz7mZJ1Hrn8Eu+O9UywPRpOVCXbVHc2yv2VLWI0fc4bgqGfLXpP3E
kVs2pM//1ieEwJFRfmu7KkA+W20Sr/4k1b8M+Ey0ulhJsLLqsc6o4ukGIiB3dxz0
1GnnliR35kvuhQj3moaiaKsr4vfB32P+/jcUPZ75amjoEUqmOmxrZGHfQJCGMP/W
h2zOVPxfpMzFyCJRw3DxdZD87osrnxTGniXSnSf2XRwQ8CFcKVNqIwVhNai/DUOJ
VY+ImWMVtDXVDpuIp9mFW1xBmVl1idcAn9t2htM9LTrciYJPBJbekQhJVGDTTlGb
urZekz73AorEr20JaMaHaNG9+nkY7WfJe12tOVDdrWOLXuLDz12BT8X9TxhZAX4/
HhtQ4dmsc92DqDBZ+J2NNU9+SL3VGd5uQ3ZqRyBJiOmz1fYrip+RndpQaqSRXZiO
kecsqxZbiDmr+SGRTc4GePIkobwPRProPK6koGVhgZRXHKk4smM2pk9tegZrLG+L
e5bmYmv3w4GcOwqx4cv4Izl+smL+8yvWXY4rDzMLvmJts6V5czfAhqwRI2Qav8N0
3ct3CxRDazrCB0m/EKe2uBVj951jxDNc33ZRF2CEHPUCJUx1mNaSXPCpSaOzbjjS
9j0mxxsVbTfLBqb495IBXGHhdmDB2rg6fFmmvgwziE8PpIz15eCinRk9nnwo/N4n
xOutRg+hiTujVFhG+xvI877kFtmarw6C9SbErQGQKKt6/amFpo4Z39NatPHP+92u
gNHE1jWTX7twAnIHDhuXCYg0t26PQCUyZF+bM1aFnWvuQSWIDn5d7YOEjoMRqGLA
BzFVk2TTXTFynMZ8LyLDW3yHDiEnRT8xvXSOV1pHGsCzlAo9sFX3FPP7B/xWVl98
MRiI8nQd53/yA5RB9IjdSuIRxHPvxz9nG6XiqWc4f4fGYj+fCFbZ9MKT7AQAE4GG
iHP7sgloLMcINwYIsO5Mlv1X6vCK8I9AXQaJnwroNXVI27+J7Os/DNCm334FcBQ/
hkaykFPNfWUOTLE8YazjfBmiy/4+uRabrenKt9oBjdMuWkiHQl2BbOcCA7xyzVTq
JPTr1V/Jy25nHFFmPfy559vIcIn2cfAl6e0Oqk86gfSkE1TJIRyQrM7Ux2+4sScz
Wxjf8MG3QU7VLAcLRAx0XuNpTriyUrkZ7iHcr48FMV1qth6k8339JFAYxaqU7dy6
2UrH9g8XN9ixpbz6cld8Ksv+OSVrkO2ioTKRVCV8ggp8jkZCTeRsjXIUNVCH1P6v
qK8oXf6mkvaQrtWSRzkySdAJu8N+RUN/ZQQGL8ynjM/DepIkgrBYygDdtcQI2lLg
WyQtV6B1f5yABggryGBWH5nueqHPZ6WAG83lfiC034sb1tTxGoJd7hTykcWvWlb7
JnsYF/IdiKU2cc3KLhZ6+bA3OeR3QfAzMYrsmM7Na1D46vZeMzil/oMaUmGGdtiQ
dqSQsXKtjAzx6sCvBJ86nNgBGE16r8UFNBD/KHxkqL2qbk2mi9SNLh3rFWE7avpz
TaOhgkbfemV3H0HY9pEIK2G2ykf6HYqaPYtb+Ndwt4WWjvQQ5/U/x9oICe2RQgBA
0d3I4V3ilMpTou4BRxN1Uyqb4AbDr3BMfUgEVlQ3Wnd4uSNd/5I2ZwW5rBNUhAIw
5cbMnAR8RcjsIu6KzFetq3gYjZDEfRdU8fqcSgzawFfH+R/xcIDKB4/3qi6sUaOT
edQHnB7U6+e9wxHMF6rVjI1F8m8n9+pjIs2q9gGrSK9VKscfW4UmhpDtbCGSmIpX
qtKlFvX95U30E91JMgJM8lMuYC1ffyBjHUQ66OXLK3qBkebVMtMebBrKRA2mnX1/
QyF5Z2gbXih416p2DXf+TAiq9xrUgxMT0ZGhKrlZWgiRYZjyhhATjRNJYJZ096oH
y4I50MykPf0ywEEEyKQGxsXhpWy4cS9Pj/HVhFmq2fFghQfizOB15t19OJwflWE5
786DIdrJyFR4C/z+7QShuVwI3apvyvtH7/BI7n4GTZ7nWzJUA0MkBINNaDoiQBMV
iujVC3KBDqubcJUBurv7fT9zNQ+Fgtjti/lPih8Zskvl7aHIbKEM3wLWmXKyC59+
mRRigBCrZ0unkqq9HIjid9pw8xmSzD29apMk8EsYi5Jn7cv1CqN5LBkQwejq95Vj
H9+ZubPjr+OmOjtwN/a45A7A6jrCvKX0TAfMb8XuVls4UntGknjBr5XvCN7qdr2T
QBEi5wd6fh8AvrOU8si/LoFDjN714t4391x8aPNXd1f70YvL2gTSy4AJs8Umqa0E
8aG/Yq98eNvAhkNfMgJDgGddosFeSRo0f4wVl16YgEJ/wbc/wCgnmKVwtARZCeDS
KieegA/48ssrhxN1n1nafxnUK2lK5hJNK7fvtrvDV138zbhxrpzmAJLLmmPImYcW
kvEQc2VqyvprSYGz3yIrwJPat1oj0HL3OibW+bF/46D/uoR5MR2TO6RqynN5iADK
0lh0Dw8R4T/C3o7AI4qqo7Fr6+LSlbJk5vNM4aXZpbA+Ae8SDKFelnJVtN/If39l
e+TjwjyhKTbFTd5T8e1PvqsIFF2YtR38YtD7KAMIr6vLsZlrQwNztC/cuYVlwMH/
pMqfTmFCUGwVJsh3pVdJmie7tVx4yfAfkTtZuXWNdlYJgxbyXLeU6JH8gXSzBLKs
/iCiaz+K6SHmu5fACteeetCIDFCdOvZDRHUIY+SdTSJAn4MNWE8enpoym3bAEZlS
/GyqAgsnKY1WXuk/c5SPNewTCCVKi2N4bXetdR4aL2mbWRQZTX/X8dJDp+Q38PWP
KMZDTLGolVn/d/Mmqc3Iv6o8zFvCJeLUewUxJfjd25O0CacrXJN4r7HhPDPQZSmH
cq3x4ZN9yzTcIuZ1ti/3v0YAklhTvYJ+rsxRs0dGQkB4bgytPyX9qHdG4CVousby
EhqRJTKvZ4NdcTHv1E/U4yXaBgP2Abb7SPx67d4SyNtgs6U0fwv/d7fslse+E0g4
KoQ4suP4Nr58XzrcIp1xxrpaTR1k1vBa6vLih1CdH/F/ldzoTGBS+p0JpwxGmvnZ
DLZKas0lA8Ic7QM6rfInaaAy2gFJaTPrNKQRYiedJlpRW+XpEWgCW/IU3qTP5y9m
3imkCFPHdoSuWH0wUKXprXOCIjbZ4Ld6O1cU/tAs1vh3J9S8Y2AI/+1eu58DrmPE
uEv5VkNLTKR4z3YpKCd6IDpB+KFLawzsisitaUO5Oc5tNufZaKZnI0dh0K8zMsu/
3Z39YUWIDY1FtNnTyEtCU4PvQi58Nck/RA81c7N08p2G2Zea80ZW/kK5qYYd+4Yv
/2NzMu4HmRg9NOgxuRe9gayl95LP2s9S4ZN2qYxK9p+RyRJvY1ggDKyihXaqFxcU
b/RHs3j1bRgA2+jcBZS9qlHJGDEOwdL7NGK+yX0C7b8patSE9vD/MNOxVyMccdU/
8DsUgNp8cIOAM73dVlkJMdACcFv7Dl5Fsh/kclmrCym/N3NP8jK9IFjQ70JwT49w
N1tMtM3TV987VaoZ7/ZzwNdPPNEb3h+chR8tCdOkFhwJjh1Qk+Zwy5r29VJmIOv6
WK9URuu6O/8+AXmJNr98GFdJbfCTcaa2k+xGQ6REpVelkNcGLfMVk8KFgZOHl0YS
MAKlMMAvnw/zS8gWmgJxDPvrNtgc4no7/tbtxNID5PLMTVEpjMNQqBbpd+7maUTP
p8mEZZj5+o6mMssnYZE9bHxa77tr5ha3Tzlz8cKk8HS7TQBTkC/+/wmOWgAGRL6U
jWm0xdZ8aofaKGMFOPUKDucH3oXpmVEje7mZqGuPLOA0mxtgW6cL986sjPuninTK
vrm8Vy4f/XrDDT0o9SXvRQDfQ5OBVblBhgKfONXaTk63w9EJ25uKXstTcW1dBmUB
+AfeSpauaIW5ApqGZiIKU2979u6sjpmpfNh/F2JDpnp85lVcRsNpAUBqENsFI6/Y
jD4bJaoabMfGaWcqCYLbHCH+vhF4HaurszOJt1gM4RGAFT4GenfPvMpRIwMhSnCo
hHuiEmK412t6KymEmfouKi+bJGeWx8ZLOKCjHL/RfuyBJv8zDRqbGISK9PlB/s0k
ICfXHqHRB7lb22Qg04Y9hRjSip++w2p7rl9VONI34kr7X4eL0XGodaeG4YT+In09
HJATtybAB6VtWRZdrpNYsgKIv1IR4YkK1jY0IRJ98MY2/QSVnsvl8ekZiJOuSGAn
1RZtgJ1wienmTCR+/6rctJZQX0LTQTplgqs0AtYJIPtP0Hbishir4T+C8qRAqpGU
B586RnCLWu4bC6Z1W/RsBP35kycTxJHGshsUKR/UHiM3C5AaAxvyrZJn8B+UJXiw
3Fy74wIfYXZIR5jhMVJpwOtUE1LHsxO7UQv+DiM1TZ9Zf41Ip+/ChehGI+Tf4M3e
oPMEvJs30n7kNYwmlW+wM1WvK3UZd33nJgXc0ypRTeo4U0OVlXBNzAVBRIUXk+yb
PV1m9onbRFO/2HhVd1fjhPyWs/fGxlUQBQYmbdNmYN81HDv2g42SXf/GZGYKiyv6
9iXystrL2vLdkjhwdjWav1RGNI1+HpbDB/4TPpHExepojVLsKBYuKSReapAWufO0
O58iT+EtuUV+wOg1KGEV0pzrzbev6NV2dAJWBvfU7T99fpipfTk4JwjHdMi3ypSz
DlNB3vh3alVBX7Ohaqe0xff22+0SgCJTtkxXRp1w0lzezpfCUukmE3WiVgNTOaVW
f1lDZaoodTEnMuRc7elNQhl85nrO+X+VMv4mKpQ/+gQ71KdefwLlZWvOvHoEJXK/
fcrwDicZu4pP0MnBW3IzVb63ia5pqF/0rCG2p6gcDeiEqcdXXKGp7XbYBP/RtNet
MFMhPOvP3gLuENw96DU61GKUHKm9Urx9bx/jtuaTzWw7WztsfMg1A27rpCxZeUaT
K9smScfmygW3FnsoPcP5u0FULLnzBrKQd+/jENcUzStAKq/BaUDILuZv5ktjf3++
9OOoHWnnJG77KHUMHpH9ur0+Y1vpkFM8WpKoV0lApZCc5tIlfp49QHzZXywweRLD
G2t5LONQL0HUsuGfphC0SfNAcYDmnblzR398912KuKRZ5IpLfEyI0En9LLAfuCLC
rJD5HUw2p2b/oJt5ILHYwHjSc3qucQ1iGRnbX4RNr5eEvNVSXf1uPHqBMsccLTGH
9a4JRtBSHjI3iPbv+RkaIAZSF/muGmG/OGKlN4IPLhY/6mCeH8YDGhBE66ECsUtq
q5CzFbZhrLXCNbgDqP6zTkiA2+csA7xsLk+XvNe6y3dZncLyy9ITupyEQiORsYkE
wwSW+0v6l3lopqx1PGOAjrZemwuZyTQH/bsVarnvEj+4RKDMIiF7SSucxXDWRnnd
npW9Q8QayzohfyBJPYqSLDAJRUZVvj5R7iDN0Qy/tHzPxms85PNbELnzsYh/Bbzw
MXzZVSUr7Hl0t/8qSVyz0MTh/eS9eKqYpvZxLYh7j8JntEG6lRKWm8NeTvmpYtkl
3BfaZIGCDieoy/iRE11LDK78ECO3HNyywy2o1nOUwIo6F47tluTdjzrRYbOPtFkZ
0hjh9FDydAiA1r4+g70kheh0bh4+WH206aXf0tjq1rttbOeqd/kwzVPRq6XpSV6X
tL1HHAM/UKAn/sdFWMaHQtnsfiyv1GIZsbeIUYDr0O96mWbbI8OqJ/Mvhsll4E7G
25fLU/O+XsdAvhpv7X4gQqpDVmEcmhAEIWs3nwkXdsYUHqXwzzgsQjwzpXyPsc/7
NsKcX08qtGDBrCLd+uCQuKkZ1mxtoMlwSX5CJ2WopfKppwjqmuJqPTiBXQI+t9m3
aHXHUbuWmM+Kyo2CyTVQl2QpEqlYZ4378m7CPmTwfyzmf8z5yjKGcS4CoBQXrpHv
GYgBnL1gAKFYd7gEgPfreaSeagSb6Era2S/FXvP3iR3WbLLeUBnzKWIviz9F0sLI
UHKe5ZFzStJ+y3R7MaE1GYxbZEaz0sDLEhfvcQnPeD+nBaCaJyvZNhHk3h6w8MQn
c3ZMjA2x5EljFgg1x7dmZ7ay1Jyhr/QGax2r6TvrjLHvEALTfbGIxA6DcnicEUWv
dCxHiwcfLSr10W7RoZDvgHqB/DvwPu6j7XjQIEnAFKvWPozZyg9NWXeF6x6P7zIl
/mrc0ZO5vIsAyX+zyL3TreyEIp5cnVAZFRvgj6J9iAliGz3Lxqv0tz64noso8xyF
Nka7ZWBf72IOWFrmPQf0RO9qYtQR/d6a9cKbDG8o6DY0E7AhX/JHdUhsKo+aMdMf
KvcrmHeOgI2GsJQq3q6nvwTXebGduaHkbMNMtDTky8pmxbzeFgXTM55gsw4GqkJF
GrvJA57oK+joi7SIa8pV0ojet6/VzpiHrmatCtDZ+/2LNgxptdHDZgh7n5YA9sg9
a39s359q+kQ7sQtjijS3b1AA9tEnzBvUojWqGW5TQM6bjZUe2qoSR2ULZ5ikC3Qb
vnAegJMYR061Y8u7jvEgGpZEc329CltPpXWmbDA0Nc5lPzLiQlX/TGJOL/LtzXSy
fhk/akmnePxbELruB2ZMPdjO8KDTqmfA5n/ZLcrdUtArpiVMrGy16YyIGYro+6WO
9KHOFWHdN5pCgptpenNR8JZSy452j7S4AQT8PzVnCc6SjcXXyGDoNlu3PDf1SSZy
sLZod7z+u+9E9JSwRJHV4Ps5vNJltEFVhHrXS9/LwhIAm8G1IpPh/y+YIwBCNUv3
c2hNEJc2RTCs3wLKdJHoDOl14TJvsVvDtw1Aib7nS/5KimHH4hAE8Mox63zt+Qgk
AWRMychluyg6owN+1d0+TCHF6qUQldz163mEvDfmv3IuIm+EjAPf39N45J5VtNAW
UgynFvREUaR+F7wES+N5sUPFfoGZHdmKk91ah8jFvpPkXtZHovt+/Ajfa4ZfD2sw
S0t06op7PbYs73+CIAB1/IODo98H9LKziKO1DoI+94QT1CE7qe5XCvmIYAE6efSc
go2ikE+d12elplR+5V1ale1GW/VhFR9XIlhtj2VmyeNRhys4yRT3gCcLJD90SAPX
M0mrn4ti3luDHwt/ug0hBEHchaYWfI1qBf8xARYCTUVFBaw+h/JtugDczfL/o7nG
SChFX6W1EED2opem+1Wy2Gm8IHJJ8hoEul/9LJUKCoQJAm9Fecwl+AFstaYUwVDq
Fmin+6jGQqUhj2ySCwtpXBln1vVmkqqMko2xejTdAwFgv1h+5zIXH1BvEjWv7hvV
Awp3RCb4T4tPbz82IY8SgOaVQNV8+8Pj96PE06loYJQVvZgtzKGp+zN1hvC3mM3z
2EJ15apYctrt+4GUWBVE+eyf2egqQ7HkoV+SVxqQKr+58BAeH7r8mtivMZl31vD5
kkyIkx83g8g6fjOAjeUEnjEQ/PGwNWbylbkxUWGuS31cw/1ULa9j+mRynQrBP7Pf
YKIaF7zjeamTSIpQAR8GM36/R9GArE0K+dxKHr0b0FnFWCtey8Es4jizjwjJjfNe
PS+F+vd/dkTXJ7a5O7aINoMDh/X27L8B44hNFiHzTCzq/EeCnuVBMBUwiY8i7X7J
vZZC85rTLRl6Wifyskt/u0XkbJvP9oKuiNEnb0FeCmq0ygPBvLWTUt042VotzUdR
wgn2zN/FmGUlT4w5wHsGWQKmUvIt0o8nPocXnklTcesljJcD/4++ur1rMSS6Wtd+
PUOKf5JfRPrpohoTS7abN/yGIpsw08Duj9TWd2Z7rJx69yW6W0FS8qJOd15Gbl7x
t5u6zZXZfW8h53tQkKUjcr/pc4KRjoUBR6lnRN45731l8QV/uCHdVAlcDWOv0x96
1tpPv3BPVJQI7nq2pxE//4tKQZCN/jeDt97zmi3UYYt8MjyF9BCaAC1FYbE5U7a8
RzWaAIVZcwnQmZNyPY1CkEGr7saJf1ySU6OfbyEfAyFSpJT/8ydVOY21ECYhs0Qh
gdiY8W3a2Mnn/noDR13qBFjFv56axEaep3ZX5s+NLDmrVH6ZVe2wfHuPpMGXPYHQ
vmRLIk7wwPVE6VgwpzblybLxVDRfiiQn43mBJB9YNhrb4ZALIP4RFaztw0X2fC8i
vj/sBFYjBVazrkKlvOIrDXKCf1y0mDHJEnzpUA9NRNuJ3dv47rFZP/K9LZy5RR8B
9DEr4LqUKO/5r9lWo66X5D1AYl9+/QKuSSLUPK9kLlN0Jc2bZSVLS6NeqSOoP+1B
4KIu2HW0NDROoF/+5guVc8hRV6P5pq4tCEhJCCtG+sD5KUeS0QEIzA5zfy4/BWP7
/0Jfr25MzAbjqBb9yFXhY6t887OumABs6Ijz2WVv55zteARTtcgYRNsUckMhC+B6
eC8WfBL9l9YlNP1I9RZtpWFsl3j11zrIPGFOm1xC1MKG7o2Sh0WIzy5CPNoOQtZV
kBsDZSzkF2FgNNENnIFOh42eecLFkVd6RBfYg+Qqbx+Rv1w+fsd4Z2DYEyXErEeW
Fc13W4bnxD+K3C/OTEvJ25Gxu8WKqaTffCLS0jXmKtTD8nCoBgk3NwRXw0k8r+sG
8Bh9dOssJ8LWt1xJCmgFrJ3AzUgzAz53XJilD4HxA/ddXHuNaMLI62J6XMa9df7v
9IltsIosggjZnLPAEFDKhMy2EjpFK/5JRuMJ51tjdXAoO11enpUZYoeeJz0zimfR
tw3DKo0la/ECZUHEfBtlC8VTb9QtuaIUT9pVwaleIwUD/xeF9Fe/65oVRB2IABAO
fUhAlXOoLGRk88aNuEHbxCVtsbOkJTqfcV3zS4tZ+eoDyjn+W928p283o8vH010K
eZCC0AUHjNk27cjIRKB+t0oatUZGs+vQobE85gwc5GYA/zFkIt6A3YMalWwO8AtO
zeqXT9Z6zLsWAvRxmQaHW0o1yI+J9qrdYTGGdFv2eRXTrnWXO55YcaTUIkbWzSyG
i2qn9+vXe8evJzEY4iVMCg4Uq4kSjrO+xqbwW0vT6r7bl+RbqmCfD91G+kTvAgjF
4rt1EmTSkgL2BJ+1rjQGjlXoc2jBosrPeFRu18SuH3bi8gD0EHd1RF/mgnyvh5OM
neZ5CbR24dQxZb/f/BdePMvyuKlaHeqbbJDsJBXn707vpX2xjViyH06bLztCTf6H
1YPnCkcm1N+VtgaelAjIpu65Iwyud06L4Vht65oULezxBCcKKSvjdc+WqrTt4RuB
veSyhvYtvdsWcMIF7tdUbvojuRpAD45AWM4H8o7OSCd1jXRDzJDIdwPUsTibGCMC
3Ft9yWFDzHqYJKeCNH9+8wNZWgcBwmY1/49psfdgEMcx/bzVB6bo3Ho7QlUASuTj
6xZsrr8QxanmP4EjbRaLBS4u+4jmrBKItMvFWLgDc2WYykHGvMv0+2YfHxoO37re
mNJotURV+XfQ5gc50aBLpNsQZa6QklZ+Tf+fEjLAptqxTuU0CTNykrGq9LhYFYOS
oH+sk8B+C5PjLIbcwpHHAa1H4gRysWga7b7fEMcUJu/1tXU6xUYdUaER6S1JPDwb
+NSLryYOWZbBg4ngevHICCWRjBlNhPJ/7OLEbjEftmXDn1/a56LbKaw+m6s5li+O
g6FjCo+9crxtet1+OU4m2urxxeKBr7DPkivqk1NNxijCNONVAlWKp/uiDt4BZWCu
GFYfcRUsiE+tUmxJRc4wI28Irq4Zj1odKdU+HcTc8AUWQxuvS5BERPDGUjJQbSsQ
tPW2pTGHyFHVnqw4yB+4hOx2s3Rpi9tmV2+aIPlxtR/QtRDI/A9ORNITXct6uwsX
qLtfMKQtc+jR7JBrPRSQnvM2qb0WqzP+yU/zEIlAy0d9u9MuyF9QadoEvE5J70bn
pEtsRBwAcVO9JhQB6ZzLPKa3/qfe6kfVWy5it3oqCUMXeJ2bE2jEUmVvZfhn2Ptr
Iqf0ULQagCwawrVnbdaVSTCpNocBhaZ5+NeL1CFBtq9HWlVmwBnXV7eenZXx+U5u
VNEpYuFYZix9BOSuKpdGByWm3x+ahN+xVW3GC8oKgbhrzXpJHs3x+znvOHTQkUhP
Ndc6AUz8h+CiyvFR+HTP+y9yi1TAarWGddAWRnOQcctEKhN0I0jwvCo3Dgf9+uqN
7Fy6jRXh9CXxkLBasmLwx7tFgszNVs+z69DKBkZOkuuxErfJIJWFeppI9/JnBGPq
ubTMbRJhmNvVfV/CGgzgX7Yw7pcslndyAqQaol/mRLdVBNBu7GjaOVQTJ0Sss0qS
Vz/mxAZBf+gJ8JJ2bQ/9GTbBHUa4Fl9kHJTI9XMZxvD1W84xGL9A0kusz8cPzYiz
/NsLEMpvahzgg/aV7aw4uJYEDlxLoZ2NBsCPw2LEHirkyk2+p8f/DHIpbT88TFys
zmY6ncdqxoSU/vVJho+pz7wXbi6Su/fSfpHqYgkuupMSN3AvUv5f3Gx6XL3BFGQY
D3RIUnnTcRWK+h49GLc1hjbUWPog9+F2TF9xMqSxb3OyVCHn92/UscO62+ukNHSZ
VwCGGXLCpJ9UhkHY4nJFxkHkQRvyc0SkzH761IcnsPDMQm4Kbif05+j3scSvSjOr
CnzGfxUYw6PYbJIRzQFB7N8zXaie1heGs4wvgQicBGNoCI09YSfT4XrniH35l07f
H7QXGFwF0XC3kHoubGN4/h8UmLMYxjMI3ylFtAt2b0aCggpPMHl/KkdlBiT4bM4f
i4Uh0BqMhwP51e2SHTMluvjnY9U6OxZvovvMs1AnMtObl+hOEuyUlqtxJS+u8/GK
cdS6KsIZcVjn0FbknlEjn07LE+P4fa+A8hJ2Gf72OY5PwGTK0TynDDtVFnA4izqL
lrcwPhvMNyJo6/a9mB4dcP3tQWb2EWUnZLHwU/8b2nqN2haX102mJWo+L3ZR9V32
+duYfbUBLzbMTkXRWZyNm0z8WfVlyS/xctfW3ykYwfzf8nlPR29Bi0Iyof4Zay8P
EZkcYEmB6l7MmuvEPlLviqlmFl6nW9MslmXQD39ssMGOdK4YRHiOTjyu+2g+oFTB
aR8w6CBqQiicwnhijjUjdluCTph63aht1uLpu6cTTtdmiKtI8zzamBaItGZ3jy6i
xzlsIMgirTzH3nZ3jrH4afURuB15KO+M++44od35OAD/aja18Rg1hPeH46vbLH8d
Me2lgddwa7UrCt3m+LcAVBfJKL/N/jxz1CbwMSXN4zZDBFTnu2jooQFIN6cXYfxi
GvbaBxy5FuFv2X7B1Uo8mfTtojlXUafh/thfMkFl+oIUqzKwEZUJVoSvd1tkkrFA
uNVliiNSXFDug2tFlSuI7yuFIlHECAgBOmliwAJM2WAK5gPyZio3ljGPZVK2uCDt
mgFAu3cHKhC/p7WqRNUJMiiRLR4zOVch7JY8edSlvLFwIftD8grxPEpwEgvbQMcN
80+0+ccAdppIxvpDGjl/x/e6iNA0RCIlRPGCdhuNm14FjhDLtNMZBZE9ncHgjuwP
HNHGwgyCLF2s1FR89d7vYReLYkEPp/cdxesV0k66uewxlUXAWi/1eK9i7kFq0p/Z
4cnwXM/TpB6McM+l6gQJ4Ek+a9cGbYLS2qkVBCb1DJ0VfMysYSvBqm8X0yGVPn69
KQIwnM/ZJfeprnwsvRj4sbDgW4OimMql4rFZVVuUBu/9SsCXppmQhfGoLy54utzs
V9e7GfL1ur1UoiLrQWhT/50h23qz0lcK0g1dOUQF+cx6PwgVA60d18YR4273MzWt
O1mywWXF5xTNmbma40tYOIDximQ0BFvflDRFK6tTraFiOi34CLwoqNTN7HUT5CwL
vqitooFg6SfvmlH5cY32BBsqqQPgeLva5Pfwy5E2Ml7hBFjsyghNULX+u55GwIS6
slGX8YzEM8KoJ9mXsS8bJv1sQLh9mbU9QH8AoYhYLk/cQV3tllh/k3v2ME6Gyk2s
c4NOtVcxOQWJx1+mT+YEkekGLitjpbMczjvKuSBGkIXR61YsluI8HwxbDoxIXfM/
yiqSUqlCZ4Ii7J2YOLHQ+1gcjMVUfYZeyo2nlKZlburDjfb/8aseZhfVjJgNlIbA
2Z3T3gR7nacAEyv4CJMzRhguOBqDESzuZLN9qRowtFw6LwuCd0e7/ehrKd/Sehfd
1zQWfBlCs6T1z42QLB0KREHf2bTwFH/jFiZFOZV5nkRP8WTB1lVcZMW4xdVAvWIl
o7YzzGQOHkJkS0bO1NpYrFZfmdEUQltwbP4evHSljybf+taXIetL8Kh2/B6IA1ly
eCTfuKfVvGZ/ryXaAC94Rynx0DrNpt/Sbw8NxrCV2D46HKI8G3f79EVbtIyZxV8K
JWBwCAM0S+kf3kJEqdrPpF5au4ZJNiAE5AffqNHv5DfPuAGf4xU+XvMrggLud+Q9
wbTW7r0I2mwBp+CFF2iMub4yXSff6KnibZvZC0Xm1LbTVGgzsr8VqzBkNkk05xgv
NeZrmJ1kMlrfK+zc4S4gRc0gRcWp44UzFY9P9n7r4P9f/fixL4hYjuHMzo3PJ0+v
hN1QSPyGdGTBEAY9UEHnqvQytSoWQxKFlIzGh/sWL7mCm8mUEPW+Ltx5JtOvWJ9z
HGfFACDAJ079mkJjODe3S62dBu6jY82T11cfegQw51du6HX8K12htlvkk344F0Ct
UeLN4BrQB2ueFgpN3D5/g3xC4iC2C7vi2AzuU8ED/r6gIBTe3PJdfg5CdNnuKtzr
0dQwfk0yEiT3urgiV5B/9CDZIplKa040UU1SBcceL4KqoYuf78h5M9YhVGfR1+36
U82JzOqFhagn3BAX+wOLb7zINgSgWtKL3pYDYIaVdQdUI+fyEtsocjbPONpGGxbx
WoB1+nPolk6rDz3C5U8Dm7MM1OJ3NyII0//mKR8CAHnxKBHTZyjIWvRQD3wHD7v3
BNElB9G02lF5qR+yZj5cEW/Rdsalchl7UYZ/vCRKWHzXa4+XWnlCpk7QNhdUanUV
smjt29AxAQXPClG9TOFaMe/z+tsI4y6/K8PVSYjLRIHu/tHaHxJSGKA8g8KeHN0T
co+uriK8Xg8tkajwZYwf4AQgIhIBNgmOIPyFFxxLBFRogsAr7/dYZ3S4+Q+pHk5q
T1yMqgNww2tbQ7jECm+4oL9cfkV6TKchKWJhaiIVY6+wja2i/Tdw+vvdz6lw0ijt
YBZDXcGK7zg7JOWw+9BIBVwKHDwGfLiQba+CGgtZiGjfdGn+IPcT2HP/YSZ18JHm
Y+aRIwmzsiw9cEwASDK6asQNoIvbkebPudkFv7Z2MAFpFDJtZ38e1gDaavHLl9ro
zJg6PPRjNbnHof/PyPNnbYWNrxtMhLF76YY02HbIpbhEqyZ4FvXJrFDSU5omexqQ
baKcy3tjeoInrOPRQCcvBWIrsjbrAR8C1Dyz4YuI1VqSdBlSGmWXVJJ1qwSCgjvk
dQ0IJ8Bm/kDwDUWp3yRnHXnimbUdst3/yIwIpL0koWFQmHeSH93sphZ9ftkHh7xq
eTPjTZxNH3jwlhJDC04NvSS2ml7xZ8kYx8zGZAQg3oVhHhDa78zY6hoOfu1p5y0t
jAt92p3dJq6hOWQdhXdvXopakXJaPeP7dB4N51s7nPsStPVXxV/aj0jdrldNMmdw
bsEbPY8A4UPS4ZEptqrrOC64fWpD0CMoMcpRfYuVOb482DJ1Y4qf46ErxTMVDW/M
BUgZ1Y4kfp6nTCS8h6JTYQ4m9Nu6RQsYmmoiBrdSKcCG7PrZBq01DSzdJ5HdAcbX
O7P6g2eYfJ76Wv8yBqToZVkrCFfHHtrk2U2A1zlDfPozoAmqZTKR4zSjnDipUKE+
l57r1UsD/qyr+DAV3ERPXqkiwuDGQLNE/HB9tt7trseWaVCNsoxl1cR2gY6QIGpB
nYP6aWv7kySEiHJFKIczuxWRFUAHaDPKj02FiD0cKHtZYBV9r2Cl598uejdA+wep
liz+APcEni0bxNdnr/gAgD0AdUhiNKfjzU8hkE0c3NxDCzVEXajvpj86IazpT9Hb
Ye2dM7N3GIOGgXKu7SUeAJtys6gBshwJw3uIP58yzuzk002HQ5TR1Ijr2UL3Xcpa
4gP9jdMbxJLVRF9gVGk/em+JGatLMP7qQQ15AAHEMoeknbdGwNOAEdLiFZgMiH2E
bNIF8u1qXtCoq+wpbIxXVLCZ0jqHewqMWtIWdLsAT5PvdBnrrdvtf0zHjI1J7Ik3
boy7mgRD5eaRMSROqpARHo26GnAwnOXrShH3vHKrQBSVGinDptu4F2SAQHZfMl2J
acQyuv304nZ4M1ajCCEq6z8fjIAIkCj5jZzzXB9ZRNYrJDy7nLdNaSVWpXlEgIqQ
mIlweH3+2+8KtxlrRg/uFitadBsIHNfm8PAWr7v96iOep/SzWSaA+9VRhbyPBQ8L
Fe2U8CKfMJJuUZdgxZTA1eSqBMZK2XV0woiGOu1tGmf5vCbMQt1OB3yqpiYU8r2p
mxs9CnKdgprzqh7iy35sgM9vAEPEOeiNwEu+wZvwq0Jlu7IpM9iBgInmCO7D4DWf
RLPfCkAdiH7R8WxMjBEVOgo0g3ABWPFnuweY2wCv9hdcYeVpUOn/H4vIxdeH8iGG
CVTFv2V8KT32Gao3+Ei2PSKZLPcgMcizinvfvLqyl7qndxBb9o3rqpG2oEG1ywx2
cC4Uo9e2jwGO/OBy/bJg9/cAGJ2SVo0kZVlG4DHhlmFNFeVyDkQfMU1NTJvXZiAb
PhEo4vU7+NAy9GyWBGb2eXIK6g/C6IuyKA+rlX/JTzqecdtWQ0KDrdOFcdCsP8OP
fBV5EeOd/uG0ktFHAawVEYZy3/NaQBRJDbsufw0Tp7goQ4XVK63Svpmb0W+tVwkk
LLOLkUT4UVlINxIPqw5whiY9CxE0CwGCamXAnRGrDzJHf8MOWNHn0dOvUOpqCqEe
CxdxIOQvfZFuJykUfdPCtQNSMDdIpXWhdGnG3l1CvZQGg9su+PdEqJI2QNfS9kqd
Q8dCJmJ2IL5j+GJf9O6NDL8pEA7WF1PBOBgn0NvlBah1yoTspV+/EyyfJup1vZup
mMR6UumGELNhJUnUJDPOY/2bewywVsLF1atYUTstVWhzgm33rDKZr9UpeJZu+rFL
N7D4m5ND8Thxixii8iMvky4Tp+fYXhnlG7ycepRPFs3qWOo24meAZ7XBBUAABWCW
2Gb8JTP7uXMNA510I4LnBv/IkNCwgPKhhi7qEBR4AlamhqF8QXcApHo60Zsi5C+i
xwRx6FpCGlP/e8PN7rRhTLQNFQPTqjalzXAl7RYvGvF+kndt+LJwdQfYJSrfT8DE
270iSFiVS7RAQSmCwZGE1nfePc0liYcO0wVAMpTOaAFvVTW0nsmzDuhvRQUXib2x
0Gnzw+f/RtKzhScIDFigYsLdyE5yuQc/wNIZFaP08AmvTDq55+dLLFfJjS1DMiOE
s+zgU6n9RYKBpZEcwRLfK5RUj1uTnqEZlINMMdLlfPptP9zSuydyJt4qX3lMLgBZ
H02nrxeKFa+nXTpUFk5ysv8ZnIAzh2XwQkSclch/xO1Xj6766H58FlwaBzezzTSo
FE+dV8SdRIZwt55dgNN6Zp3HCCSQMibZQXNsYm9hDa28AKRlmx82GcyQ2TmDh1rL
suZSrcBs4rqy9hlfg+Mr7ldKTWgbbwcsFWBdF8WJAuqiAIeqK0esJ0HjNo5rTxFM
o6R4shTg9GBJlrA4aNAvYBNmT+ddZEaubvh8aT6eh9u1wz40yl6VXCJVO6547hOk
UaVZq3DeQXWq5v56tea8uKQuVEDfZMOIv0jDIdGM4WLPiMGEKTNf1CkJyj7/alu8
T5y3OpgsGO/prxPtAYf6/nRIFW3wLCMtQQpjk4XmpPPPTJrH7RJDheWW68WY+5hW
aaK4URCiBIXv7oUWtJMj21y8RNYmRDaJQI8VSP1oVI7jPb+hgeKBi2Gkl2ZZIUK8
IIxig8k/KwNY11PKi5wA3ul0UAXZSB0PF6pPzfTEbyqRlVpEzjzZtUkrBtnVfwJN
gly4AitqpejQbna2QYjbQR08Rl+BIFYtzTwwda/KVuvuEKEtLlMUtolErR4zfRFe
oKiO1l9Bjc/au3qSMiq2byCSYTJjK1hAmIxej/UQ7X0bDDVgY13iEe97Ph2MJK9/
Uiu/gHCRlx3bHpfA6T918A4PZKURPopXVCEkAxtHRyEXwn2nM2zVnXfbAcv2kkGe
EbLURIDzrFv87ojgd1CcLCPLmvXBFlThcIErAmDveCoh4EySvJWrz+Aa6E7APb6N
0iX6RiCtURpNzU7VyTXtARai6HYhhv6zsv+V3aK2mNJ+LGH4Q7szb5TjUcqm15/N
0AuWBEgxJr/k4OYNO8lJ8oTvrF0D9hjEghTVgpzJolIMnZdYrETTUgKBuPo8+ESy
bSOoubNPDw3froGFHCE6nyfXhjJEjKGvRm6A0TjdFEZ4Ru9E7nYpIQ8/U4Kps6WR
9dEaiqMmNG44DHtarfgUx8OJBrgOmB9R+M4jQFcinHYsSS13NvT0ZtoslCKt8mSd
PR2F/MdvWdjt1BTqTbEgtDma0DW9erOVfHjhOFJweX4Gpj0CsFK2v8XPvrdpGKBY
zAkPbb43uZEc+cVc0UxznYmaXz4vOeFNbHfvFFIhiPgujVvU5fiS0dS2+eJWqamc
04cYawsuSpSM7bxRsRXZ3EMVonqpAReWRNwI2UX8z2Jr3CLE0zTudIXgouMWjtA9
9sqMTrv2+0QJErDEzkbV9zc4YEF5QTM+qE2N7FK3SbaCdkUNMRulesDmf11Y3kC9
PEDMFFsW24DjG0Zv7tLly0gEIX5tSGLUmSSYjwmP+O8eHwIBybYjRLiF9AcZBrgZ
sCeVywP9vfR8hqzb62YcNQ5SA9jPbP0ynoXAXTLV6ENh+dZpq+p6B5rAEk8Y9tjd
hModfueWlhJI5R4t+wp3JaDdVIW+XVbr4aR6g5owdiM7B1y8b2BnucELayot7gc9
Xbq4YqrqxL4fucZiW8UibkOaUu1sUvTv1OHWlcOdYtltBVKQcTp+O84fY7X/4KLJ
J8Z5p/6Xq28ybtLMqqT5jxqKCtQv9buW2OHncSugjyKJhA1o0S/3nJ5ItC2FKdax
jVcXy/LuZA98ne2fUY0P21jU+a6R/7XxLEOL4nCH3w+B3Vsy3trV5l+YLaIkMS7W
pA5+xP5KbDcuOYqzPYwEI4e4fqyX4fhkoEbXmOxfkNXGirdlCCwTGpAza29QjnTx
8As+i4+AAxOjZm82dqVb3VX0Qek05chOwb4FD/yzY26C7uNzSojnA2rzpcqj73tp
+R5ckDMoAlYJlZCSdUAv7bjuCtCQbapGYSL5+00JMUNPK0IKg68z4Er+Xr/uYduG
2rG+2TNaRUFdvg78iO5RmSnyT/ppqgN88YHtRGj17oem4cmgxsonkvrAIhoBqyiq
15WPl7Tx/HDNduATcMgYXiSqQlme9mzp2u0yyEIffb4JydFQj4NONo7usnz1fVKn
1O/S9FFXJHeVi3lLqGZfxMD5lZLcOVWr9mxX0v3bq9Jd/m3kBXeTOdj369I78ikT
PDOn1nVs9JllUNP113neZPFjYxc+tnO9k5HOhLzU+0SDKoccFPej3fNdbOxkVAqU
VW7JzCKBQie6UZ1JXaaI4LG7qohOQ+IZB45NRVmcqrnNbnaKlfOHrQVSvVTbLCVy
CEyJRyVEwms+fbhemawWHgGG5tqdq2G0yFrfLLeUGtnPr3iBNvwIq/x7QuTfxVWG
dFQ24YJgPUeMaSHdnNe8/AWLvi3GM2JAsPKHTVsB/1TF+6GtGrDkb9cAVjeoWI2e
07e/tKYNPn4YIXj8xoe30GnL9AcPdcAXhN4PpWf2qGJ9EU0QONnWdueg8dS+JIZJ
rKKG6ybQlqsAevEKyVMQTHDIDCn8A+R70a6hhQtDuz81csswdZ05M+9qL9ClC/dt
ox+FCnbIYcxfSoAbRzSzu2Yv1dcnsg0JT2qGbIWdYJMWfxJKvgwuOHJ/VGV1ZYhP
bFeImI4qW+4ICUj6E8wbyqr9HivNGoDBc/8W3Ft7n/6wnM4eBvfZLW6X8UIJghfQ
sHL21hPwElbzNwC4lOgzhPWHzOJnF6bwNogGqO0ZvW4KAlOgUF6pYXoziKUvSlKa
DfZZ/350Z6IjB7fOW3EQjkSA7bt/4wvXGb7wVsDGrwuE4GvqdYI4yBb1AsDsHkXH
ebzL2EokH3rnM57HtdumlOJgWM/cPw1pZrp00vToRagVSoqr3/TJ8P5Pmdsg8f/L
T+6TXrM+cDo0I/ygMbeiMqFO8F5kLBU9li/vF/rt7vLXlrBapgE5Qliv2rUqPwab
sBx+AbwP+YIfok0guClltVAimzHLcZp0miEm/A4thvqOYz6u5fcki+2nUI0W7zoI
Y8LBQnTRxcwHNFhWH6cuX4O703mMg91RGYnJGmIDM2jxGGPFH4Xmhir2Nd0FlzLY
wofz3WbeE2xq0UmLusFBIFQlzGwZPzIXBGff9drqYNLCTzKRv9aa1/0Zx8X2YwyE
jjkkNL15lQW/ciQFlGnvNQU+RIsxmtyMRoSXkRYLaJh2qBCq4SAbHqJ5b0SoBhUg
LDCKBwomIUypIRppYbhCd9HCtAOSLs1yerx99t3s99wIUj8l15D6gZ62VXkSLcXJ
nWe0RyruE+YqDD0+1f/cYPJiE+ZJ0fFe57vA2+gBMQwZJz2v2x4c2JCIaJnn0IS2
LLuPaoibAZQC/aT8TgFkirn3BsDDnEg89Klxy3yQv8z+HAwJGaCa19u0PMMku2E1
GVJ0bkeE1qGl2o0VPbpwxDJVrT+sY9OPO2i0RMmtD8ZQDE+PuRRU5nJVwWI0njw/
ZUtA4gpP/Guwt2gsFI+/aJb3Dr40vbyk/KG+ZBvuICsWUAro8C3uh0rDUzJZvE5+
ulvrRkocEo2K4QiL+6n5JOYzI6Ab6kByeyOxRHlATHr8rr+m3/BdakuQBmGph/O1
jn+iZ+vNunT7pRRe1jxoUjIaPt8LXrz2N9xRS1EuPiTC3AUT0/1yc0YPHwFluUW5
DSGZdoq4qeHiq0ZLLZFaAfpFov3a8l2JhMMq07nbbSyN0IQK2oC7LbbNZfBGt5CA
kb7qG3bjxtAwMSlfRiTmgCLIM2NuQcydGJNTRzyJtgB7950mXNXggIpexbn8UcLy
g2LTI/ViIFL8RJcdb7QXPSwwRV6h8SGD2Egwp61ONRodVJ6bj6MtjuWJi5oWFXdd
n1TnImTLwNmezRI/ksMasIhbP1akc9e5how2RPc0TTdgnm1eYvPT8i4G5ELDM6Fj
5owOQXMn6aDtM0bB0xPoIJD5yXd1Vc3CMVyV8KXt9Knc6vY1NI2SvM2/sTLhIA+8
cOHSH/VZvx/GyalAr3jZPjsYnoFWHmRV3I8hpYywX7kbCy5IQKEEieAaLyPyjDuP
o5Ubm2IBWHXaiXxZWRIa39r0Om7oJ3zWKhgDIWYpkCvjzqG2LWGzExYRQnZWJZka
pIXM4Gscs0NV4HZxAvU6y/T4LZMWWxc9X4zOnRE/jtxxIwtABII2zfVrVMcgTrOz
/jKQNYLq3sR8BVvf2z6WOAeOSKwEsrnQD58qMiiUSZ/y/sUv2oAgcQ8DN6HX/DnY
yGdi4r3NFqkd5Wj68/P72IsccobZaL0kBE9dU0jKOnI+aC6T9numUs5W+IZ32m7M
CyoGLu2wejH3AAOA6VBjRsA4VUTu6IllEJsXnls8lzEDskuK4A8+Yk3tNge4F4zm
jwzivKKe79rdmT0JIByO/Qk1EkuyxdTOZ5vACJeY+jBnSw1W2/XPbY3tSi7D9N6j
1WGlp4oLsU2vv85JnQUfgXy9NHjQeSzStAs1752v7ZjbOW8iLbbaV1Q1Z1R2B7g4
X8JNBZEIiD9Zlh32UW7s5IUOrKCDxV8A7VrsFlsfuBCK2AQhLctAvOL+r6NPVFrP
Ki5oUuSCVZlBU/fHL7lv5C0s6KYeVYw4Zn58yRa+HOLIWDzchqg4q+TGYAvrk6WM
BvQ531H2gfrLC9pDSjFEn+8PTMEcTCXw2OhkpXDVAS7aUNCuZUZBhLGwOnsOvbB3
q/5iNYtTYygzOo2RK7XGgWRApLK++bWNPWq5UMxWwDmY6OfBm965VGbCvX0lKpU1
LiPHTQKpiVeGEzJ0xidREJWjXNOjff0bxwIzF9agxG2ksl2YjI9TNLvrSuNkuo8+
2XCPuWzsYIu5sMTEpNKFTLQBogzeYAY6BS3JqPi3d1PLh5naduHwwtoOiY98gQRS
89h1RDHzn39+PeGjRTLlfXXpJY8sXPVCDp49Ru+ct72oH/AA+R3I1m6vZq/Y8Qmn
o/hlN4ixy8wzdBcRUIfwL85aYqM+EPZXjFIJYvOugpFG1abddKJemp7Z/xp3gPKO
cjpGPlvE7XEiSvG8T+9vvIpBG1wvkUSjnX08lBEkTSSizncrUcDoUUBhXziqC90i
CuaRInMBJHt4WarH8qKE3u/gvW1pilz7yyAEK4B/TJpEE7kg4fa+FOsbg2wX7aps
H69jqgp+9Nb54M2speTJG6uBWcfPf7rBcTD3nxA8FYOqtt57XWnAWtarRAykk8z2
zVyA1fC8Hk018aCCZpthjzi/yn5WOX0pClMWdU+Q2K9DPHIj2fUZZmRkdaiDUviN
4rRvWAYNKLE/6YOiDciMPorZhKi/mEQeUGQWJ23RM0xkQvNN6MPzl/DEJBeTUAXb
2zM+/yuaHgdvVw+ym0OQQyq31PRO14oMyrBLLl9FXz54/wbHgPu5rVozreEJNzH8
T5bHGnOaPYs9BxvD4GgzFdXntJiIcl2ecMgStmM/f1910jKKV8JukSqE86P/5aoX
Y26Sbn6ZWY5W5VkVWwMTHI1wUXTTPqK6wb65r7wlNnS995ELkqlW5RPoBPwomkOE
0RDJmpHox/Klhc67aXs6+Ug0Wj5cT5m6MxOt+hjMR8Rx5tdGWOTwixoTop1cNlUR
C4AmI8miE0VUP6KWcr5P/Fpflbhj7I7aAvLRBiYP23lCh5145IpPb+GXM9JLvR2m
dP/b17WxJwXG+XeLCbRmXDROSJMjeSUnAr9jPCUISI/H2zYx66eWJ1sufLHTfp1a
XgVGnAvRYYqlCtUy6WMnpTz8GjrvviY87D7CcIB9+wbGrG/P9LtekOHp6K1u51hu
j22QKQGDWVQDDwhPD5Hc3A7soH8izC3jOL6bX+Na9CDCNffvIsrXywj7EkxL5Nov
yMoSb8ZJNnoz+b4o+YoqwDA7VqcCf8S4dr67ojZ1rHhEcWTNMGnSXaiABCIspkqo
NUZInbJbZUrcy2vFxINsXoRHO0LV2PdALAp862dESGIrcVRdZsiGA0CU9WEg22fg
Y9w1KvySq4ZRA33o3VySsVywfK6ffRArwDt1KSoIzhJ0cfPbbtt7TOIg4Yr0QA50
ExC6h8ifTp6OU7tJlCGGzzLk9G951mXlQQEG4UNx5rAqljMIRYTL58zWx2GXUbdb
YdMawFb2fHB3dXjh7aiGpNCFlXKc/GVRVed66vgOQ/mVw0lkjbCsiUqTkrg9M4J7
MaxQf7PBU5IrZuLVFo/n05v+hvF3F2CYZj3uG4RuMwhBjP7foA/HaRPgMbWmTIsy
235YPgYn2HY73pVT019AURae42KFJDEI92M3kgdRwDibu34qeQFxNrDYVNogOKF2
+TbBnoQ05Q4TarUTRXiHIUnai62v3np41hlwdHMP243Syoq5w/RGK1DoWGiionBI
5OVSlgP3eJCnGr4qtAm12A33PNJ0NTXKMy0MJa3kJJRQOtT5Cw8ERJZCAU9YFwI+
3bKMYjxvN8o1ZP18k5HxU2LhpK4jPp2qP2GYqz0ho+iY4+KvOVP8pApZO5twd3K+
3tTI2PBYZCHg3oIAVFrHVhDP308Ba+qsQxONUWICsA1S3kSVDsUYvN1XT1jV7Byj
fv7MMntbB/3awOb2TWdoH98yqeV/4woYvbdzQ8giN3HAmmPyIjUCwKkgjQe7yH04
lJE0I1XSlvsmQIr7mmbiVll8CWTl0lTl2vaxbgWFbRRBLasCxVV/AFmQMohE5h/9
3SEEsPew6vnZlBaXNfzSziq1ENsqblyCai6p1/3S5iNdqJLVHpcIs8dMjf+u5OtE
QcFVGe9uf/2wMrgkhOrQjmZ6+N3Rt7i8Fjw1FMgo6EgrlN/9IJxTYjNiGtLppNsk
2iqTLBBn1Jvjq7rS/0hGCG+c4V6NZMYuc3Ylk/P9TwbYMZelarpKzTyaFBae5vEf
QFjeQl3/TnEJMkgKGcdCWXp8tjFqHYbE5oz3gVR/T6AljiReqlB8mrKZUXzMjUzE
N7ENbdyakj8NStbmNLm0j0j58taW/Pu/5YGab5FYpPmpm/vKnF9Jld6edQtPYJTl
PdAI/OiVxNwm8pcvBDhwagm2EbHQo6ldN/uCiCoDQVDiYFYh5F4jRi8Tr7TEhTrR
GPWoAVdUGpeNQ+rda8c0g7HFMbAXzXbXv6BSJ+my7A90bKlWlF7du83Rqt7N6/bL
Vg3Fn0I5MSoEqgk4CdPX0m2lvtTzRvJY9NppYLvJDLPsBBV8fFx0vrdR5JVoOzVY
rGM3l0uTgG6sXq/FE/xIGutqGBhWVfjqzFCY7cknqxuSTU7vp2ZroNrJtppnb7sl
wG/hBJXbgZs0cIPvePPE7+lWC8DFB8BpFtNRLLjUAzCulbNsxba8wLmE372rFjYe
jMtv7yfpTNZ5cJV/p/Ole4jL0jMjapKh9neTWe/TPR/BnVJ8M4338iNjvJy9oqmc
0/JWQl9pqF06iQfLUvK6C5/6omc5dhLHt42euzbLGukkyjzNPwL98+jdD/IoJJml
I8N1Hu8XPMAJZ/4fsIoYqejRQfxV1oEQBCKQ5MOVbSCvphFSzfaeFmUs2rVxwAm9
yOky99hft7vjXtHbRPknXFXnODzcTKTEKqGIO4f+IoNV22myRtXygW+LUYC/2bgD
Sz6QOtIpekQvPej2m8DWsK6ljhded5DAv/BDGkaP/71owKNC3SjZedZ6Liui0f/J
kaFp9lyqQI1F9eB8zfQebXPqYF8HKOMZ6WTXiTfJ1vGrG3ck2iRj0OomHEsPxiZ3
/wSVW3o2nqJa/8exHRAO6f/r1VQ/Eg519+RDQdqYHLeUGSQ1ruv69WmqhDETpf3+
myRhm7m50JFN8+TUmEUkecHn2kzh1UWCHK5LOPH8RT4b3rt+Nvvg7LN5FaBlekzf
aG2T6nHglH32puGfiKqumoRycNGRhxI2BfcHDep0XvD7NWQxEkm/L5A90C3aIJs5
+jFBO5FtOf/A64HEi0btVpKa9QQE0sfqOSSEl+lSFFjndnWQUR98+iniu77pe2xc
v4Aoccwa4Usf8ku0UUF1DyEN98cIzErlRmYewUp+4B315ALdlhRpiPMfmQRMPv6D
2N1XYQrRjHlwYTanoikmrQCBkcfrfIB1OjlVqLOnL/fxqJyj6qHZSAy/gPECRSYx
+EJhnrufMDIEipfGd55pMnkO4cjHp9g4sMRlosDD4h8tU6eMEJrg85+5DtuDQQRb
jAk1z/lVcp2VIhkI8eJisKq/JbNC++tnOqb7o80yPArZAd5mMDTexSlO57dnBre/
TieOPLKlf+uP0um7/SIGFbTDm4FH6jvEx1y/me7IHxOIP80v7tVNr5iCDAzeWvVQ
IKwDDaElGUSBZKXnV4XlLY15Afy++CsLpV3BoHJU4Y75vvSwR2IQG9csR6bXjjWC
Y5DQHv9pyfNOozyGlKmEtBWUQ5QMlNGethXj8wo5tCWmCGIf6iFbHbgEf8u6KFZ5
ih//+EqC7puytiooz4r1S2QqNZNGnf1d/Vn/UEDOoOiXSGKLbJobH1nhG6WCBVHU
epTjkpq+a1BXS6LND4VaPWoy+oERAWrbM+OI59FMv3nSyH+anEJ54SBjM2mHVe7h
e57/qaTl5jIzAV5bBT3NJZKQCrF8k0v84mv1+7h2nF+efpFeuu4QW1EH3aqhu5Pt
2hMPgRtvyiRUE2MvAI7KwOsbQwZozSDbSPaTHuEWzVgE/hTu7onwceAb+n+7IdZ2
2fZf7FGtGvpZo7hU0Nl5xxBamWvRtATTQCbdNFcL7FLUdwcJZvqJHVKbq06UDDm4
j33o0XN/17qbAnBTOHTUy/ZBsbQlH9hi6IYnCnFKydb8IlDwlgkvsvI2+6TaXfvy
djm4mxf0nQ5BVwEVhHaH2q5MDJznenoFoLw99xa00WyxVEa5j2u7ZpzhNwKV0aa5
mU0FnE1ePaFW6UIk7ux6JO9ptNhnoDoDXbvTdu/pPA2QGKn536ubHYaXVHKvUyG5
gGmWCA8fbwX1DlLOiCP7SqN1ZZNIXeKtIK/sk3EprMZVlJa94mSaMFDGHSg7OboV
ewS2ToqUzm5T2mBdsv4WC0pENBm+56ox7AMkPB/q5FfDFJw+ROfK2Uwa4ZO8uvK4
yXtk6/sNpBVwmWGvFTAPOSfAcf+V/Wzm6HegaLbbjTbaBlpowyVdJuZhhAthMNr/
LHeBA/nFSfCRB50xnd6nGJOgEdKjUqa9yZKbh7wQGy61lwqQusTznl5k3RdieeuK
CBk5lCslzvF6fpnDvpIU//2ur4SXm6Wwc4RR+vmOUnU2+jFtmHjpcg3hZhq6OGQ5
Zd2zi/oyxmmhaa81N8XMhlA3cWsWlYyTiiU2QvQkWKUrs6FDD1ALJF3DXEE3rJ1X
gnqrV85fqwWJuwoPqwhApqMHp52y2uNUQp4i8yZnak6KnXSEJLxVte6B2Xde2go4
DXEDSN1rJWi8W4wOm5Lwk5lmE+kX+p8GqrNzR9aF71wecDv1jz0n//56FoRm7aZR
FcKCujTA8jEX/AOFyBzas0ROELmsFUQkhyEWHXQcNzIKppyQEZUsyImd8/CUvlqv
7wHDno/A7HGLtpn5wstXKGDB73Mikla5++uGlJ00jEzhplrQS7rsJWOcsMaakL5k
dxvFnG8wUQPTcj4CKPtHl0jRvhIgadRS6ZzCgZAGP9Ndx/8k6R5eN+2SMteUiwFU
B4wl3y/XLguvj8SAhS4Th1pqthTYOkdbKR8UAW0TH3eMAvC+fAV1cTSg5F3qoznh
qe2Nv0dXqkME6Uke41Xf7I+P1oU5/vuoVodmOqqey//Gs5vlVqj0Z/HwPOO/s8e5
sbWdlXjC4ItN8cCNa3Y8QYIEdHwgU6OLFP0fxar69KpiJqffskjp1GwhMvi2UL5q
Puy35oZIijExu6KoczpyrnUJK6C62NpIJwL7y4RPIrq1Xqw6VhTBoVgbMfGyQyaK
8u9MfhpDGuxKPpiyO+lIRDKaFcWmCZzSu07aq90c4FeC+LSPkU6oLHrf4Bpfm0D4
mLB2/59sJlSBKkpKH3xZDB16atY3CGIADOUyrj1WK49otLYG/nyNDlCXkdUecONc
p9RBnCup6wRrG0EIB1R29tdD1Vzhr/wH79CQcWb3rk3+AGcC6yDLdqNUeEA9cFT2
NMn0YLLAmaw03SrZbRPHuaygPyN14dkJL6TxRk7d/MuUj6IINjbKvc8+N56XmbcH
GHdjbseNElt+eNkA6/m7vOT64f1CI1ZCR5wqazo04wyKZlkk4lKqd9EDonwgbK8h
KP5Ldtl2fbDizRTgZ/nZ5q+iLGghfxQCmfPCcXN/V/I5eTHrCVJYhSVHUCOBDgLv
BT3UU7oaw+GrL+z7qD4bzIhVh4p0YI6BGdAhAUcTMFi3daTLhnAKBngMypof1x4I
kuhLaoa2GwCBfElr2/lZPjKrgGHflqBXeSCBF0cJLa4YAileZ5Fodwj7GiUbocPL
XYJnZbR7WiDp1lnFrFWOHcfMXMo6TvEYvwyqrNuw4QWde1AdMbs2FKgDJ//5XIeG
QDvDAjziN6+dZXQOXh6NJ87BJF6hL1bY2Lg4wXsWkzgJIj+TnIatm2B5V4B37F64
iL3RIeaqT9FMI9SNe+OSnvt8ztwEkpNS0UhZE/3u76sLs1+QqgFfela0LDwUrznF
lnzF+NILH5EBoJQgz2EM5Gh8O13YqsKhfyw5aGJLG17VcBKAiC1ox4kQ8SdO42iG
bdkifl/WwpUc5IjjCyV0jq1yKHitIgvnINF/w6IcMCBThVB5/WhpRrPHwsl37TgK
oOCWEqoGWbJmRQcFWnr2OAIzChaUebIEFAKxjes5/zwa/fBiG1d1GkqlEfxEaRCN
mZ78hL4Sm8eYDSt8JuNtF1Oi1dKsOkdwh5z/MEmrfTK7SPXuQ5dhSQ0CPb1X5QRD
bs4XD1PKV+SFxghnaxNx9CopR4tAYX/w7JziR/Klqi5WbEtacuXcjfAWGgM5+9OU
HRFMLDWQgWjoxdFeL90xrHl6PyzW0vhPukrZG4YO+CwLSOLy4EuI92TL4vdsBFWW
/d/JSjVw2G8i0ONrLW7cmlHREywcf4OH9PYYP5126WUEwogl3d/Ei9vRkJQzhaqB
PJMDh7D1syHlcKg4tOjriweOArBLfCd7rds+tX9RFRQrVpbOt6bTJ+uCACHJ3FeE
2DB5SUvJL8hG2NPvAl6MADaGrNsKY4Sz4b+14C5vMpZnKdbhuNEtYivzw9xgK4lw
ZciN6K9f1peqHUEfBlsvMDEe3I0VQnaCha9+/V4+L1mIAD1lTlK9pTJjBtcCtPHc
ELDd1W1lDQg0i8rqVR7VpF6CB5chGt8DSLjwKup77zcE8lbSAUG7vSI+0PL9pp3d
dAzlzBsbkWADWiPQrQxQOuvfgLu0COX3YoSVG6rzSGH9meQPwGrfjrtwBrshORJd
CEKZ1jjwaboAVwRUqDxIOPAlzQmKHTcK2L6ZPqv2zKDq7IcxuxX0gltRlt9HW/iH
aY7VVw3m7eXAoVkHULMstWijDrHxZJmGlGtd5nBtNGZqhTVc4kP9Zve+23PzdNzm
avjF+6KalnWB17p31aVi1tEFzHhGUsdXLcxye4pX3OtSKTI5J5tAacZwySafwlZz
VFgEJHSJYlnlydNDxB2pl2bgB/TEbEnuBryAVhgCvXb6aDMITj9WxDEu9FCPIdW1
VI1wBbK+IUuCHvkSIjqo25hW1/5010t/zr36XTHw4CAKCUEQhbfG45xbQLuPyghb
/rCM0BBUrsgGvMEDbY5AO9cfAhGyfxM88OYUzLnxu98mTEYjuHr7omXYWxiiGQuZ
Q7fhGkNaGoAfvYbcBIP5Lh3A6d5cqmQizg84u+e9k+aVAt9ODzEo88t3QUmZcFBq
+6FLXrG97QjQ5rdHdcqGIpO0ay6/qFp/6s2OQ5L2dKlmX+ihFRAtN7aP7ZFNsoxq
fsd9v1XCSDOTUs5pLw7wmfh3KdltNZNUyUBW7PGLYJJj/OwQlB55r6UX37EULtAS
96zp80XEKXq9S+wvmrEuB8wvsIyaC4Ney2kkGU5YhrNxHlmKPlmrNiZgFX0AavAn
Q1noTDUuEvhqvKBMXlMAg5BoN3myXLU3wtIFjedxCyodwhfkw/poQEjJvWrmFb9Y
ZsLfNfm8spQ4aGkiAU6ETpKFYa+iesGq3RDpCGWU2sk70s9CLWC8qctzkiryJhiy
kgQhSqK5JWc37Osbg6Q/K6Oy/6FbVLGGcNrsILaViYNS4Q+uDePJDMiOv9dQ5U7v
4F38OC+8s35qWu0O3VVEoiu3TONcry8BHc6GrqQJ3PvrNbeydU5x8nagdwd9UQBt
E8dCN/shgNfkcsC40aR9Q8efnniro+pEePV2yKA0Mhzd9HAzK8D0ZSrq+TjUrjXG
57+5TC6fh3knDBfBWycW+yZ5NbqGOS1XjvEpo7u0xNJQAZkgsS/fZknDQ/RXuZnT
mX6s8vzKsKw1G/8p+C01c8S6pALDM6uJzTzznl/Yi6WwLEpczBBPN7jU5eOMqA0H
mDsaI0vnCZVfZ9GS0KUAGgxhy50q/yFf0uiPW6Jc4t/wODUyWFVPpmYmPjHSKtlk
/0EQmJMoP4RUxVH58m9V/uOWEnsojhFl7bUAvWI0c8/9JpWtg7Dz6R2rzvLHrHGe
t+twfH4GErWk+Ck7zzIheWpQbSpyMdZtuKur7Pktmk4ohTF8G7PPMNgTwngy3h9W
m1Z1vyD17SSmjdX+l5ZHRXcRj8h7mRxLZ9YdxHYZgyYP+2cNrSQwz64z2AuXvtZy
Nb+I3UfKSTUM6CJT2PIv60l1W3ag5bEpI9b4q863FV97N03XHlVZJKui15Yl2uVY
laPMFtfzH6f7kDNbHK+GxT4XK1hlIV0+ARvcZY6eB9AMEgmXqLl2jWrX6mCCes+U
UV+KULIHiY6QXMlpQx7R7DQyt/wrJQ9fK7r5ZpvK4mRtD8O8TkCyA/Jlz576Kdve
4I0U98G+CtUkdqj2+foWStEyuAi2w0/Z8s3C54nX8ygGOiIJLjMvGgnzeY5cKMhk
SWrDAZShq1AYtvPpUfpktevgZRO/yVJ7Qci+8p5GF7HWt7ulAlgxA6E6a0PfpFMG
75zTUTNJlDF2UJx4ksgPvjVqtppYgWqG2EI1Wf8tS3s5u+rh0Wm9E3alQIrty+yc
6sZIjV690mEAgOYsCHI/IAc1SRgu41MYCyaQ3rpktxH8Ag81PHPhu2nHSpWrZ2eR
3S95Ig6TPDpb7jPw83gzGPpi0kzFx1arVMh37vvQK40MG6QWx3OjhOi2j/777jYi
nhS2qZzA4nd3upTEVqJMX9oj9l1dX552qBYC4Agmg+mXXyNdTEZQiee9RxM31Jdi
IbH5t47z2050LxEFrkO+3dsTBP2dbCdRnRG4T8NcRpOY0aRLWOsGKY07+UDUMZuU
bPQIe0hKOf9DG2sagKwCqFPOJrCXBJnAHE7/+1eYsncBOG26S5qcUzLkEClkP/vR
qiiA86gvtvcpI5JOCO9m6dhH13wSTMkB8QsItdWIappI9Gj7RJRDHQwjl17nfyPB
EALdoGvpgZsDWKcJ8toWYKa+jn0rKXV6eUJxnW7Sk46DsS7YliFoE543zsdH5BIA
gq8q2O70/3arQHSzgGLSCZuEpsgt1yJPUC/+vxp8cK8jKWLJVIB4QEQJQZ5sbvYQ
S65drIB9EzqIr4Ti5OjuIj9ylMJtofFQyd+CBTWWOS5RbtXoa2ZZXBNHYiOm4za1
OWVkF3VNBGvfjc2walkJN1huKhCrLzxs3G49LW4+6SSxZxE8gNRNNs51LoiqZNFj
06aMtLNjZz5+8TiKHBEQP1eE8hZIRVkLQbFDT+ebubS17oaXZbS79TB/iubPC4DV
ryrK9tTVPw5pNSeU2RoKsBTOuqSxdqam9pPTPqopzjgKb2IhKsYLSnWFJLKv9Axc
ncSPCMZUiImw9JSpFei7nI1zaqetzCKo5Gv8m8MnI13/exvPJoU2P0SFgMpxTye/
xAxbrRQLCCRSDpWyF3O/c98f+Nv0FzJK0EGRV89Ce6lUNaE2b90NgeAOdi8uFtH0
+wjbKkvam56tThp0zvrOu32k6lZTfpfEgynYS6gItNsI/JGsrY+2blzG5J6weoCY
4Fv+S5CGN5AkwUo9l4ZpS0ZixIEJF1ulgS7y+pNGdXX6G5sge0GToBBw7dWRe3q1
Vpr6Mh/ayGv45BInmD+d777ju8GuHiKRb+uHVRIPhx+bGBzch1RZIzoVCoOjzfi2
NyVYFsCAjwW/MTmhI5N6i9BsdEF4HCmdrDW35KEYAsUGpr7MZecL6H0jE2I7kaMV
BoYT3elIL9HjysJKEia4gFfD76aZzFnsOS5poaWgmzznUqH8++FlvvW5W6+uqRyI
SccdoOIriFYH4uVa0bTmCqCk9ncrfVfGePWqxtxA3qyUp3Vbkt99kxYbNzUsfRQq
GtBXrUpfq0+V9W0reNbIbauLVgxKJVZrHUgeKPTaeVOfo/msO497GERtPnybP2g6
KbxesrvIomRmKWCV7KJ4k0d50rNS2gooOsQgY7/2sPiwaL1/ee5FyG+Row/q0ame
YC4c1M5JVlnfRg3NVEYyFSES/qwOgOzvDsQwVXJjcQvgLFqJxEMd0xCfdvNb/gJ0
jzS39njHqU/bXZGSk4HOCmYLEp/kSuzyHgNJb4DBqHwmOv+UvHwiga/dGG7bO9hU
FJss2XuK6meOTcgqgvdL3EXZ0KkQScmhL6ArGKSaIcoB58M/NCErTQWeIbcyxlnw
DOFfrYEjMsenAU7xYOkInN2L9QW6Dcjn3SJHPBM7S/fe3VCdYhtgIaK9JupyIFkR
RY5jl6O4AQWUufrF1ShYJhqPjoj9Nx1ZLhLSAOlf/boxxlAmPrI9Osz7Ln9N8ISu
KDsPWb+lx1NC4JrIJqwBY3b/R61hGjoq2R8NUI6Rme4sZRH1VUmjd9y0Pq5gzquH
ZUSvxIAhLvPESTXhU4acUKGzF3ekXisx1YKpF36yzJUmt73kb9XVgAAn99tMCjSv
4cKyM0HRrpafk66t8YbKv1Xu+PXs/UQfXINcHocvb7CWgWrE0jz8gRRmAnmd0PSA
zOh/snMDrJ+VeIfK1cup/ONmr7TXI2cJM2NkUmyAXLIwaris4Nk+u6+YMB4k8XX3
870noEg1RPVTyWOLn2V7Wm+GlluazF0xPTZ3fKfQT3BxFKEAi435wL16FR169O24
QzeFoThZZANdINMbltN8oXB0ujQqpzQSCZwE2YTPGq9+SNCK2D1symq1BlIqeIrh
7hEAVkCpkcvBld97xe3Jf5z25bDwSyZYVfNTIEGDYbYeBScJZCGMRxYoqvg9SCLY
RAmmRCm82ymvnle7DVdpW2Q1eXqgPkBEkTLIwzBn1iXtiVXc0OFqEmQmpsePSPpv
3jAmkGHfJ49eKZPUCzs4EdWLqusoKjY5zXM4LarF0qrtPOOixynTFh0RGEs3MXsh
OKRlcIiGDSzTllW2nO5dc63P/axpUauTaGg1rKpYb3NO2w/CBi9x7QC22pHI2FuP
YiqsZEAl6W8JLs4fak7h/z/kiIOL+MLgmHqQsrALChbAOiYn0iRYqsQJaG7YKBDX
oawZVAV+Hx7SWN8i3totSMgYRmYOPdg7q/Nurw8Rj5PaKNFmy+KGBQzjJiqAzFVn
E0zdn56w34sw+/NHBDdiuCSibRgLmFqzSKdUTkVoXp1LIsV9P+CF1kd4xH0dwrGP
cmCNczMa2QP6+PXPO5SXNDMNfZxuiWYHgBuVpZ0g5VeB0zElQfmhxa6E76WFd1XZ
RNVz91LK4vOBt9xDh2qTKDtPJdAPJ8GGpx02DAWZh8fbxXQ3LDEH/sPhqkntlmGe
UsdnH8QV3A6wqQO7Evir0FjlqP2mXjqufFFsmhZwvhD3nUJAtuiWOTEBpv4kr8q5
smhPSf/nEe0L2+ZUxJjI3RZO2KNo27eJHARbweAVf0JQj53MpidPS+y9QCwSVv2Z
Zw0shwTXUihCcJR8F8TF1fCE7tDEJ1ofc9hrrvdBHDOKE5Pl7knBmW7FRDlJk6FH
Okq1ztT9pFg6AbEG8cuszYA3un6YUbaYWl5o60p6pU933hziRZke8l5ToqITAguv
nIWy+FSa5YzOtgzmlvdiyCMk4pXxIbsHgLESSbKswUmLr1EfaBmhd4TqfRlVjo38
KqE9gNG277QB+xcgpfl7nTTDKmB1BXFRbzgvLg261N8DBDizIYZofnRFHrDSSHvc
6F0snTJsT4cw9NPsaz7xaA6z8JzGzvApQ3W0L4kuHDQVEkjIIYIFw7gjN9VqCcqX
XfGPvDZ3tD2eg+s9y4q+/c94imt66cdDTXFUUwR9DdaykFEgrFOa1UhSBWs7htxN
eBaGRBEyt1Lvxcxeoc39nGpstESB/19mMZFuLbLqEEH0EMHmZXJcqXm2wtLtUgi5
kX//vPzOZVq/9vPf8VfaIRr4f3AmychCDxZgNys0VFp7PyNV7VhD5qcQbsI9c701
6+lVUlyJ7DFNtjuC1+vy7yvIFbxL9k0a8hplGMwdc6xdreUq2m2kcfn4ZJZoLjN1
5SHG/tpO/4aHsBXWC0cnx9ea/lhBCNXzJa+6BPj1g7U7ioh7ywDiOUVn4WfTHMaQ
sWev4yVlTEBha8cHSaKZvuDbv8ThmqMUSja5Zvb7BdlwfoHuYnFvUz5Iu+Td1fwy
JYjk2Rd5M90dQLKJXW+4cAU7aIVkfI4Z60BeiaNTmPTkTGRkpcQWqDFJe8JpkRM6
Dn55rm/cXJzNLrsIY3IV6YHz2skEs6JnuaGXM9dPKi3QHlCsw7k6JXzSTO4fYNxp
ruYQvFLNtyVwc3iy7WmcVgEoO82gxGLmpUrcuAn8rDI5fLHkj0hRcOfW8fBYXZI0
Mf7tMzyTWEUv0w5rJ4/EzsIP84Wr+sRzRJUcI/NJkXnBe7awQTtvA3J++nvftPWC
lleuKrHWvxqlX1sAZKQdWA2THDphg46A3kQWMIU75DZPKjfz9PPttNJOIMcaZW3/
wdMbn2x5j6DRYQJMhordNrlch3vVNZ+eKjbX8+kjwy1ptlUhtG1jpAo0M4W9bw4j
TT5DD/rISo7Wr3f5DBNRtq5SqdESdOIqdmqkozz4skSUIXWOkv9+36uzauAXZWj0
rULI1AE1kuUe2q5sU/6SWaobH1LDnaZqCv4tWlSWx/9xh2aSkEnGRiV84zHNY9R2
tefibw1FTedu10VaHzam8x2nH41z4vVg5UiUee6WPBiEE5yvw//iWtshLJUoeoBO
JCZ9KmaF7BW8ZiV5ch3sDsKm7DydVWMwB0SWhnZnwi9a/N9B1Kibd/F5p0vu2OfX
VZbipGzKuW6qvcCjzVOGGM8qA0u9LBSZPevQRqGy15m8SmsPEq04y+1CqiCoL4VR
lboJ3UWiHdF6b/7A2E7HdBXNmxR3s16rbJgTjyla/gDplEs8drbQZfs5Z3tw/z7S
r09n5pX50CHrvo2lbB4/OZhg7+0UcUWRYrVxwJoylWezxDSak+YSqFGNVX8yqVgr
QQwkXbB6EUMnbMG4w16opSuIMKAPBJ/rtXhC4F8XdhdqC3A1fvJpb3294RYWFiA4
6brBdmJjAlKvsMeYm+ueYDHp86fTd+47QJ/vNKnBAY3tAX5rJ+QzNGRU4oO99eTM
aR0EkniOiQ+tm8UxqJ1eQX17xeElKbT9ujx362XPAVzpQZsEvvDOKJpvl2g4Q7w3
X88vjJhVoY6MVGW6J6uH3iYHLS/mkmcPAbDolcvQkNCPNkSChGpgCL0jcAKyd6Qd
yNa1X5lAU3vxZFvK1ArFz3vmFPRh7g5hYOSeoiKMEt0oCdrEKocMLkbIqI6bXUm8
R1t9jovSJc48Jg9k1Hk8C9WMmu1ct2ywNQdY/lzvnqzjbabceajj5PdlVwVhh6Qn
BjrXyoQpD8EQCZeJJmkg8z3ewtFOAQjp6wVBcO2WGd0MXwqHSs3y4Pr6OFqtJMDU
8q9hOrRCbsyXZJTOejW8xw9AMwIoQtnmrUFYWCg4C5wC4c6HmLPsR+NutIAVZyKX
MLTj1Xw/03zYIpOeL8I6W1qVeqddK04DSvNt5UCk/td6XFhbRJlI3ShXDSwf4FbF
bgI7jqbkZrk5bVXKgjD9C/50EMEs78gD7o4UuB7S34Cc6/xnxldG6NAA5TxwlO0a
VHBaWnISAjAN0vpWl4kzH5G3chG4m8dQ5w9AzM0Z/3F9puSNTjIjST7inRAs4/wO
vaCdrRsgC+sNpzRxK+LBwRGHFXEhf6p7SsVX/sywLe6e4NES9LZeh8sa1MnnWwbJ
AvYdo7tEFrUFP8YDHbbSWxvrwyFrQ5VLZ0uK70rLSSb8zTPjaOEyy/CUorPB2N4X
eiUHKrvYD7Xom2y24Nm2puC2cG2CbpiqHxpHqNs/+5U7VJmeGezfp1amH5LgncA0
8nypEgWKEaisyinOo0PznEXxEwcDeStKOvftx3RMbVusidgIsTyLl/UxDXe5s3HV
Ch7PqtbEsUf1OwFYarwwCBo5zZtqbu+LbTVtQEGi0BgZW+Ky8UGavQ24W15R8v9a
kFfkFf2ldDm0TmXEXi67G5jMnHlXvjVxYGuYYJacPcczQLnFqzidRubQjf1x8QtR
IrGNG3F2lT0aIpfzAuoMhoUVfRY3Ni4+rRSIVlcvloyKaTi5QWRLQ9LlGYXKD7cL
SKcSnLcj9zLmYOkgfVMOcsvFrlEhrH3a9bEp2M8f5ld5IfTkpGgQMoMDBoLDAMjT
3v7MiZBAv45n3S/WzUQSUeKOSxXof7rUBKgyS/FzQDn/CigYywALhYO/eApP+xks
/d8FZ8ZZJE3QguNBKlcf3XXVJxBStlwffNRHqVxTYVOnGUPqEiayeR0ZNAKpz8df
6t+0kkTzcZC09vTdDRxA9y0ymbEcnhK6erj3hdq2RUqxYdm338rtAH3+5HRsXLIZ
7iDvI/xqRMS66UtOpC1Cb3px2ne0jibyN4X/NlmTN/Tu0dN/Qy2UWzfNbBJGW8sd
aIIx7YY5K5w0oqCD5O2li8n6q3HUhlRAE0QjHZoCGHN+2nJoKMKIzfQYq5VXhcU8
Z/5WJhxJg5OyrMSZ0PXgPKo7cmXBY1dinAspF4m6m+bs+n6QuYxScItrJrHHij0P
dfhazJnc52z6m4tv7DuOqmBgI/yP71sbhMzel8X3Emo9LdrdFsgVPXMq162AQP8Y
OO5aVSdMjo7obI4RjU9ONGKu2JVxu9lp+H2Dwc9TAMHdkyZlp5LFlEIddRRukPc8
iuJ+AiYUc5KoCWSYzCDBwOEjmh757ZKkIly4Kd0H1rUUNylUdvhBKXXkh6JEHOSJ
kDjKFVfmM0NDIF27RGorPQC/W+2RsfSr07Y0tSB9KMv9zOSHIW4jD+bSSzWJvhBb
2dQ4cPQWqZ7Imq6V4JJiWqbzk5GOJ1CFp5Ov0QCwp69ck4B71dVHaDRfqVg3WalZ
HEWrXcN7p4GamlLCDleTydkbciKvnegamvoclrRU1YydeNrCWZN7+LJS2J4icQQ/
hJ66jigVc5H64w3HkWmefGcCbyO41DYo9IjW7yBt+T101hmMS7Cg88tejAomH7fA
lxL3hfVIhA8q9NJeZMXJUgvNh4Aaq1w9tPxSHDbPJmkn2cEgCAtQbbQqBszMY7MN
hME9qpWfm5yqaehxMHPo2MMupdqXjCC2Z7XE+z2cDR2RnIBD8uojum4kCxZipErD
ZpzMGp/m9JsFPwoKvjH61WpR9X/GF0CUG+eAsa84hRkjlW7WzSVRnWk5DlabKMW5
YDN4zRqNiGlYWpGe/kDiauYMKVnGTs1Ue4SH7UImI82FFNY1JK0N6r+GS7J6SkY0
Qo/pSPY6vyG0c+VuS/Qx69J5BDUfmePT7rtvCoEa59651djXgPPQp6+OpppX6pSx
OpAFHiu81bzUI7m83q2fY3J3q+Bs1o1GFghCaNMJaXoKOvaf41GauJ/hoiCVxk2Y
Tap43EPp/M5I9xlV6Q7Mq2MH32fM4IdX4m67Us76rsZ07iAq8M6klQCjJxO5wQiJ
j+fW9C+BHBLlE8ZbU0zzMcm5NBsS/6Dsd39UduzfHdW3iOxC32Oq+wEPsPjgnXSf
PCEptkBhWEwiKuqoLAi0n36qToWnucE4vk6uGITEI5GUrbtcpLj/fZoB52wT7lvO
ktoZvyPdjPJe0B//eo5CJ+WajwlbOW94mCteZVYd34QVfFn6DcwEgigaTxR+CDHT
BZVzFC4o6IAp60wRsUiU/USUHKPs3tHEl9MAh3rHm0Scw0GA2tuiW+74D6FTqtQ5
h0F+wgmLKZogDcU5ja7qRLdZgioneOfMD7pm98qt3/wffwILHZm0s78PUVh+fqFM
njFCq0Lm5M2EtXL46vYxfhcIj5vqFrEcY2CInaXMHnMRd9FBusBgcjbk+5ldfXkj
7vz7itrPFLkmy0tsTZUIqGqP0kmHMD8tSbZLp7jBgpx0ZV9KjOVawlFqg4nCKsWx
VOfuCy8GcF9IMxxlpRgHH9M3ydOVZOJ+SHJaSZkbIzz8Ncj2g6Z2BykL93DaIrC4
rb8ykk5DrtpTSyt7Ol50DMAIaEW7jdX7VBjaP+Ya8yfugq2JujQNPQSDKAMsJ94r
Yv7Rz75K/EHYMeyT1ZIYkRTkUvSYnZDIO/rNs8+PYr+T9wcXAAQoAZzQo/ipTdyR
hULR7gvymJy58IjIAcPXzP2pPZgPqA2wQ0jriiUylWDgzvK6oIWHHUjYp9BHmSev
Bjo9/nWEgVNpdq5B7Y/0PbipzmdkEJFIU6bNn6M9uGEGM30fa+e4IFK0JY3GhJlc
tdLxvMlwuONUIxY9jst5jffYP1wgXt94Nd5qvF9R+ewMea2fo5/NXNC9NLz1WvLf
n/6XpRD/IYi4ijI1/d0mdm9EOyfw7eOSVn2DS2na+hMCIU5g2BqU2lDKYUgXVYAz
crbs99EwhBJpLow2nzL/pPZCD32/DOKo77jDYLCCyRZt36sOxZKiQ90vAiPj4+X9
EZoz51AyqVtrCZ0h2JbyRPVC/UspseDc+yq4rLm9JSsdlZ+51cF4xKkNUXdzTkuH
OJ9cbQ95/9mVH8rR41vBV0Ep1mQX2lY7LCs5HUz1uUzUeDWWrXnVWCsfkzEg3DHs
uG/hSfbgfZjitm5shVlKI0KTeBFx2GByjLVdRtvWcViCOyQNOct/RZvMZky35AiV
Vj500C5NU3ivJqLeij5DGTCnEreVeatD1nyQwaxMKeRKtH+Ue79d0i3r9uHGSOam
HrlvvMfDNiHPdX/4ZhN7qOi8tmKaK/vxRPrg5fdiLkMMYsq9Qmr6lpcjqKINUYvZ
9Sb59kA4NxNvbGtMgaxJqO4/Ww81eLO12WKUKB809xYqFh9MYu3EXMQxGNIdBFJs
ypJWeXYvHvWP4oExFKLBazLcZ/ux4psdxTA0OG4JAYlcvV28J+lJotrqXpL7545e
ULNJNT8CDJi2u0H4QCwvEJ2t4kcVPjDCpZwbMRu/LrfB9HqT0v6RmkccIrFdaOmL
gqBJYha3s3DKXZzkbtDl53qmcPo+bGQJuy7f2g9FQZpV4HjJYOOKpVkH/EGY8lNl
gYA4At/Eg6TOLheOHkTYJ9ylS4HpgtbsA3xRGbI9xZIXdMquBe5PctfYI2rMZSqe
9AeHE2dGjY4W+pBF/KP3PFCVMX/cQJc0NCpRqnz73lE1+G+r6AbgY+md9qENa0CQ
o+bbrGuGA1vF60u4/KbvxDctEIwnsp88uKy8YBfem5Wu1VvodZUT9Ikj/hgF/lfm
Q6xXAmZ01Htyi8Kl6GQmM4eUsHMe+Sb/upAkO1X6Rlhq1EOdWCom9lvuE+HH7E+C
D14IlOXXBBnuAREJ4dBO2D8WRgaSL/1sF4j+AZWHhorOz5+dthaY1/gVRjXxTDOp
p0u3R+2hx5sYxRS2/L3M0JKqocH25vHHp6F1/49URr+mnaBpqe5Rp1YjLEmMMkEa
A7rD6uXPh+GjFDnes54AaavAW4DncXczsUwEutwU+OrsDdSgoInWnYte+CRp2MvI
oNGUjAvQTbF1QJscP3olIbopNf7fyIIVs5uuil/ABXrCcoyVB46VRU9at/pvL7zM
IBurH0fn22i7EQaELkxnHHLoOnOuJbXKDDokXm5W2pfGwERePz3jnW12ggU+4fUL
MuDNpFDkNaAakNOiXIf2I1yrXGXWjCROAoSAHlgsYgru4wtaImsLa0h6DObTzrSi
zy+LrvfzOet+rVEI8iIhgnGmGPe7wbLGi7DsU+6TJVc5zuFvqG8kp3QI3eK9s9j/
c8114tRbkxAOqV3xp4Aso9qYBGrVT0WVW03+iL5VBQqwnuGfuomnaqQ9MA5WhSlQ
eDHajQitWHaImLiqRYGOGlkADLwkxUSfvjcvnOKhYGS1QZC5jcDeaIuW6xSZBZ05
hqyublRhGGbdG5fTK1cAsKGFirIJGwhVTLNrh9boD8Vz6s1jn9CwoKu87ERCKb+x
vLe7GL9npC6KLfZ1B0hJvpp9yMOWU0MOpRgM2/HL3LmusA90IA5HB8svmdApTBNp
PIwR1P5vQ93lrBvxWqLaf3kUH7utA6WY5dwuAm/ox26aHWLXnkGQgTWVEXmaOACQ
qNo8bjnn6u4pb5dshCGiOMhEDvqJiyGfa/G8Ry189LclzIyVJyxzDSyg5UR798ph
98zbwbxtH92GDMwh1ibmtY5jq7pwVWL9XX0PQLp+MRQEkb6eFCkcZ7+zpgGemTXJ
0qZzyNzP1+uLar3toVBxDPcIBgut0eORkXrTIuemDvVGgxfKWnHV/x7mGa2jkfdz
YMxweKZPgPHu3rOLWzfYqiPlhRbKLdNITA/bez40oORqqttsuPoURObQiNg/gO89
hRHY/1dK4QCMNhcI1QkYcSGo0XwgAuKOcCljpHj3ilLdYyAENQ9aio3mN6wYBrjB
HDZQhJqUbJe+cU8vORx1ANOh5mEbTMoSi1UVB7vMHqr/ua92Dh4YScfdC9VSwtDz
zjvV28kkF3EJfDQ/5X3d6qCeY1g4u7hpCaZeEDXe8Y2AekAL+MvSgrpZF5tGHi/z
25mVL30jIuRLB7ASlvUfOG3MCoqMEzSu70VdVPLAXQUKFoJgKb4h9wdTL/E9Llqk
f3v01zI+FjX3yOrryjRh83Ej/At/jG7GJc7LTvO6D0fxUnkal7Kg2FHt0FdhrA+9
HIqKkDmqFLhDMkDNQqCpcA6ZmaJJeS6QSmYZCkEovd6y77/jcMaKXDdMYbpEDeYt
Fe4oM0c6h5DXW7Bm8LQ5yPGMv90oMyX0PUNIsODElflbw7kSHmSGSbXNQd824kDA
35XB1uQXk8kdTZY+rPmiK+bkVHEq7BvbB07DTKd3IrijArWUgVVOdTH0iRLiZGlQ
1SzOMbuBohCc50/HONAh/vZFlKj0doV3xZ9HGl2/WWRc/C5WtinxjYjV0MBne93y
wM3J9ymyCV/ar2h9CQiwuMLGkgh/bwmdT4G9ZkEIk02hThUWb0QHV4075e3cION0
bA6CjWEOVyAMqlx/y9ncf5rKZaUcECk6BM05ZoVqg/UFnnFTVrFVvO6VhGdli2TL
A6fP0qFNrmcSb7Gw326m/PBfq2BVRYibF5RwoJehkg7Dj4T+wQX6hxsuDQcz1ox/
8oXcfSmUlq+doXlOQLDBIozOvwGvOr/eLnFTLIT307PwedHQcu/YfSBILfg+HWZ5
IzJ5DIAUxwiYoJ/4ZeyFIG7S8dCosiY+yP/nfy/So4Benc5IjuqepBmQBJybVevm
ZBf05sMfOCP61sLT5PGgKBhLlOIQRgdyLm7kt+0yvTUaJyCq2ZxpoY7LAB2NHmXR
17vp49rCbo3vAN6CSMEPsfFHiIUJyJOLpLNERDM7Kzk/q/CCwh0eRKVt7OFwOn81
WtMgOdHr0JDJPzGsSgBep5Hrn/iAkiwTI2sM0Jr2zrU6cToWBik8xot5z5J7PChh
6RfA4kFzJzSYLl1uNrIOh7lOMt6fSafl960dEJBY+xWzwxdrzrNtYOhKHihbjYa/
eX6vfqWe4kJOdFV6iJOmPOG1B5xK8Jpb8+Fe7YAAbSgMDMIb8CNWhmi6IWlFX5f9
Ha4Duo5ofHq1hRW/iznRcmnXK5NOA22IdknSVmYbeTLcgGP0635Qe63i0s6Nt/vK
0ZUvJwfsH2evDSw1Y0T5vTrgkzZ1CWBPovkMSJnEwtt7rk6yZ0Xfn3Gtu6aaY3rF
mfoAe8znkNQmlaCNYFw1r8TcDMyjpJKQarkYvKV3XxbYV7W7sBvlOV0UUP1Vn1zZ
Udk3ljX/QBDNWRsqSzW+zdGyYWruVqvvUHqtn9QAZMPw1I/RwCc2VIcg4bXGGaqK
W1HhBQhKQT6LAreDi4BR4deXwGWFDpC2NPhZb+syRQsXhet8W8w18yxLOHmNuDRY
Ch1pHgxtEkvUOdAfUybbN6ApY1Dmf45zmWTZVhm4Fs1BvrsDh88JrgfqU03HzyBb
CGAnmO4SC8TnVMsSQ6nOsvnYH7k1MsZPTJUQ9fVwDAnEq9OFbM0HpIGVf/72cwP1
2Ogw+Pu1DM+/UjQlF7QnGvgLPk7syPL0Xms4PjaACR0jAwEBwGO4tWT88bP4XL8F
CcCzXMdaChT7xQFC40m8fXqIttQpLfVQBqNhyD3wRXeI6yt0BlCyhNGQhU8K/qoT
/tBBrspYxSosTWhqmaCWjixM1jqsoLUeE6O+lbBA01HRTTT7YBf+6KbHwlP58CD1
FPN3y1G451M+l9uhBX+JQKXfRAxA/z3/3JvhSRunSkIjWzsL1BsH+1yMZoMUImkb
+TkjgxSDrz7A6JQ5/T+yjG5a02ZXbMUxGyGrG7DJknIH3BJrMWydv5V5Zytcximi
7Cc43FehQIGz+49vaa30mYbyO4VpjiG1GOKjUJ4ZwQ5eKmQw2BxJ24sE3m2HFqcW
mjdfmURKC3HYQUy9AOIq3We7Y8T0tMvMI7/H8GCt0cnir1AhX81Ytnck2Z/8B7KP
OSZDv6En1xPKbwacFu61jWCrVzAtW8Zv5FV69qqC9ENiP9CP2wz9Evpn4k1KXxLm
nCwuKzebj34dgA3D28KlnlXbaUFg48zEQbUCJJO39Kb6qPIue0nN9Jd7XnzerWRj
dBnjzBF0RHH7UtKynd63qVfWEnu7MdHJDKvO00utiWnyrxg/rwXjfAS9bJOkhsAm
4v0Z+XixKe68V9O/0OmIbmF3qIUNwnoR3V/ieG1gpbRzJNHXIz6wjCplUPf24vSQ
5PxqNs1rKOumROcvWDi0HWIKhdm6CtQoc7hYTC4m+wZAcUBSPwsV769rUytqkqYf
rlOaKYCW97PUljCrGPDw6cXNRExgwaqUr8yG/cRqE5zWJYzHrRGtMZxYqBuRdM0O
SXFWaFtjFM6fPORluqkv5SVueE4X7zRziff3romOS1ZMuSGWuBligHHy/oFN0xzq
t/zit9YsGTxA+B4wHnE2Xhyxc4JBCFjoaFCKvZmvKkC+glE+G+eZGxohe1bfW5F1
HOoPKuxDl/6hizm6nAOhMzoUJwvSO5oLb1gO6SMSi1A28StG0B98TK6pM+v3aCtI
T+E87uKb2HvDPJBUTwanQVuk8u2wj8VHd7tFKIEorDtr/hgWN9yIHmZAgcRj1/N0
OtXUdgsjte/54Zv4AvbTF0n4NBuCKiNpTpgUBuCzFwL4w+tS7ZL1cd1XPNtWAS2S
754B2wCtM1lVhEpwkRX7wFdyYcwONlSGg3KwXqyFcBgXr76n2bBeUHKi9Uv3oc7/
rEXjTGCeXyKrpu3B+qvrkEMEqzf5aW7ddeMdVdR3dKYVEpBG/uY9GVN7/1Jq751s
Q4uDkG4OsDRr3KBT8YiZbpCKgPjbJccZa9ED1pDjQ4GqrhuNvSqKMJSfjhRoStXW
2jBNXIIoC98oKGahi1N3jfk1oJ6OK8DHKUN0nCJK9DrlTkDmFsnld6Iu3YPDRAGZ
PIlR6XcSdNQRgMNUeSXN5MQejfEf73KFPH9Isk6ifduevFNa2ivT3OSmR2VEWhMA
wHagTPbHVxAffaXE9rvxCd5KL/U5mYUYOckfUXLRTuFtMwxM6LouWS5dOzooDZYB
HmcRg1Elf+rNma0RDOQaGVYO2h29Ks0V/AUyRgycGxNv4ke14heYQtKMJevvF7cq
cZiP+Eh+M6hDQNJuYrEu1Zrkd3SxAAsMjAf+OMs5XGREzJJ8H50xua7Ntdv2uYmS
fr5cIJHOPVrKQLMyDtHA7mGFurVwQ7STO837h2DNPS6fzwROTQSHpPNNg7/XNxF+
viv8IkoLgAWS/O1xplJmgE8bmur+LJt37PWWmGR/anMy8ZcJ9ZxdDQ+NKdKS5gHr
OfUDLMPS7kJDWINJlcvNZ3jPVTqm96RtYhAhHdrwsbdmThH1TnDyq1nUT6xuVJqS
rGbtIVY30OLVrtRQ68he01N8qRceyS/AwE/IWHDsE+L795RxaGBeRzkMsKk07qx9
YRf1R0KZRhYXYRN/7Gw+BS/jTfukHAnlIEmvLWv/xXQVVtaTlzeX8zpFRWoBV3RS
gd1hRCMW3fFe/+FUMiY75r5Wc0z8VzeTqkR4Jb3J+hHtqMwF/7mN1PoyB9C34hvH
zU+rLWTW//rOmya2Qn83GEzexKGzA9qA1tbusX9MFgsTQrA55eWTsRo0dQWP729f
SYIUMTDIs/5R0NVi1GWEA3PLtRFQDLeUl6vqaBbpAiVLGFqN5RI/UEQ3gsNfrihK
cncLIJaPkoR3inWphMlq1yX7sLnsAz8kLE4F0bo3DJiFyW5f2Sk1IWHsk3vrdPXy
Zp8ArL1qTQaBq5Jyc6DL0eYijgF4tofcV/HYNhknixqgDhwwKiIhOLpFepGeX0Ak
uKu3dFCg4PeVA8NmpZeP6/6SkGzQlPuYcb4z9iqAEFYazbvgYNKQP8YKXNX3jXln
m3T0/7HXQZ5yODJRUEIlClyJPAT99vFUtAF6RL/gV5RGfh4R+TahOJm5+zb5UnkQ
W0UIoW+b8yWn0A4PzoTxsz77wMDIPft4fxOuOaIShMoNOP9KzTXkbnq0HhbPhYOh
jozqiTbeeGNobV9GdJOwI5bcPondETWlArX9lvNDMToNtLixaxe4LJM4LDzeOi6P
angxtjcHdSzN2gu+gUqNwA8Kr8n/bpuJxIiFuJb9oUiT4wCaztP7BBHwcFPjkHRC
cxkb23/fHDdA4FzF/SxcRZePcKnGSMwRan57CAXzU/YJDdRUBckyB4pDW/ylF2IP
ik49/rpKoT7bKZGpk9wpflbo/+kHHc7Y5k8kmklh5OakOx6w6nTa95hBldfsvH7y
6oiLP3a+8hvSDEcpYIZ/9g8eiqkNh49cmg6ZLxM5WIDFdLBLA8fMvm+NluxrmC60
JswxzPbneqIu/Nr+lQeKM6mIzmILecXCeAKOm3SF7M4G4DzbTnV758Qg7LXrWV22
HH7jOoNdEHB/Ext1kdXa+6Ern3ubOtbVIeBuPeZWLmkLG4S9uJYwFHdyEYcbwJ4m
DImWP1dajKlDPZ2LQCnAsLdeT2DevX+y2lwaXcAhzniMigToBGW6ECN5hAD1gAtl
Ti9WUjht9x+jH0WIl27xyW8uXQog4CzUkJ55UFjyBUyJLXH9BYN2bfzuxPASMDVf
L14GB8Qj7kbJ6aXfQmO3+mKXJ1PGl2C+qr1c5OkN0l/PHJXSlktI/8FisBcxuKFd
21udYxoZgZuZbxK/X0BbnUYVIRGk7BEmHATMYtLRPYbcd0H8WX5HZfSBh1MrOO2u
s8Xnr40K8h4TsWWyqB4IZ2dcxDG3bGPgBR5owzdafH3t/ERTAO/EsSVOF5PwSerY
6JF/KsfQC/QU107sN7oDbzzWQwiaq7ZDLc+MAFsRPFnExij9ANK1PgaifIlocbfR
Vuw6RRo7Y5iYo8xgsLd4r6WJe/s7JQSpzZCy55uIOEi7xHpx/3Kjm8ez0G4l/z15
qs7yNiX+eyAGyKHmxc0ZlUePz6uSCEv8WaHSq8o8ieA+e8wFIoK7jmYfYoHbOSNL
TWZCwGXNXUMqVMDX3Y0/I5WEYJ26OArDS1fpdLIs/2WH20FRsnd+eFSphwlw8jup
e+E88WmQUTmXegKWwAuPTzwkQ7qTn2zbqXvHlBeNPCcVPusWAjRMRT4BJ+P4nKjs
DN/4K0XRosHXmCrDANxvdDeJJkj2bJ+xpFYkilCzCK2DON2ljtty+oQ1jcFmwmz6
+Td9F52NH34nXRrUZDS/QLcFiNL8/rOHZ3Hz3MlXqa0it7ZX/ijDiOC8C0us0Exl
7r5kT5e7QoF/+Ul4MQEvTjllf3GEE+rIGwYrBNECWCG/Z1slt7XKlHvaYkQQ9NRm
DNSHN3zhkK74we5yCOfN8dF0gBB3LTAy19IAk0WphCMVykSVYp8OtCkMjHREKhHu
jmQAyv7XgEhtHJs4vOEOb25jgcFUh2lyKzzVFQoWjOJSd5EDB5VTyJ/DCzVRX+7z
MZPh3ittUH0aLAnWwQFJttAe6Vamus/OYChDVf8wV1W1KbtS2OjnpTQ8s21qHW2V
nRTu8gi9/nvgD7igL27gXI2oSvVkDWGMLASG/rVqEh6m3GE19poBqSxvZK4Egnr7
tjYMRVjDnHxlhM7dVQ2Gda40CIv8doe4TuN8lxpoTj949UjIo5jJuS4yDkZfMBcR
ttZU/ewxS9zow6gAcCJls3O8UMxgUtvrmvJcPN9VM+ACrXaptwRTLcQPq7pooM9Q
0DmC8id8DKdbU9LUjv8W32+dcQ3J+0jUQypznN2O/gyT7Kqj5OM4J8p5CatazRuj
QItrP30YoyaDFGHwLJXoi8Hyb2+6knptqthe/5HKwJuRUELEIGGp6fWne0f8FCt4
5QMtrrpulDbEPgQHssUMoapQQxTtxdDZl5Nyj9mhrD8M+AKQPWypoTiVFLa4FVO7
/ylVozfyijiz6Wq0F8sdsr+lgcEp9SfydTPOrTEacQXwdwSRRulSQRuuNb33o6OB
H5X5Iz0h+KBU3wHVgafSbNFVkIZ9ccTRgtHHU2HaoixzYgARVuia2F+v8XRKdqxv
qlVLDfVXH/nlmPyQuUj9NyYFfT/iDbBmlmrJuJskGXgcTfSLYd16OdBT7WbcSj60
myK0Z4ASpIc31k/u4Zbft0qtK84a3IZ2cWiBE0shIfbYeYhi1IRRdgcivnfs3IiY
ssM5U9j8MpX/bTBiLiTnYQ4v8aqQf3AoDfLfJgCIaCvNjfpohrCbiOqidL/i9/sg
+d0dzCzFn+Ba+c3vqXz/luK8weMKJdlbwH3fTWkJuC3sWvaRaZVpwwCaA/+aKh6B
S9mN9PjNMrKPXTcIrciQlvXgfTvo4EB1itpCzkn1fB1bp9uP8H1PoYXqdjvlGhoe
8imkLiGaCjajpyrnwAf8GlRoXVPZ1SDLrgpyqhXlgVUB0FsqsOVm7SyOsLHrQ56O
89V6yZr9XTOG4hKxz2w1SLc5VpqcOdKxxlv5A8V3vkE53GxVuu6vnlArB09RWIRm
Ec4zsqY8LbMAXQN3PF3Aa8R0GJS0TBQEkE5njXJ4IiT0eg2T69CFFnet2fB449fj
b/AAWXL8lZcgipEouZ3dQeH148tJS+hmxeysFeykcnNJ9+vxC54mtMqjTi7dMIKA
2HSxgX69xj5rSy4MVlZ2lBUkhW2ZeiK1J2tZ/ep82aUcA9tK4Xcv+EG3Y/CccHgW
B6MOamnFoWEDhKHZrbcntIEntE3ZTSHmxBxSBDy6qacaaS7/gxuTNdo5cG9lkEi+
lswmjJ5tu0m3FRax8jfw0x2I7bFI54zuSIn2ci2IVJ1OZ7/YBaUDBS2xDMBrTM/P
6p1mVc6qFNRMBMXAjEkedv8FXG+IExKMnq/RPvdupwovyAhb8HgAYZOQVIYZzMlo
KXfYlVic9LYBgwzWjAi1dGwC4xR7DskB7u770TP2LeCiDPDmZYgUTON4rnqvaAji
QD1dDzV02+OQaUVqPLJdpZdaF4tAhkVxw9cOxeuAU3TbbOTNLxhWy6fddh5aO4aX
5VYiDEyWwPbLhKXE7PilTWb1UfldaOdL8NjBpgV/ayS02MOpJ6FUMgK+Ws0mSiNl
rfrz0ltMyWgdvbHsQ81FZwLcbdSPeBdjXNS6uRGBmso8hcSAoHCuyWmqiXlymO01
QlxDvUwze79jK7FarWJ9NOnfx7oto36W9qzl+FnOo3JM0tSDKiAWP3oOKs4biLfs
iZPIkeeGP6uouuZ0nSMnHaQDDZuee3ET3DAgOa48kj8z0QtvgcxDenKN2TOh+0Gd
K3gYAsowQjzJshTlITQjEPx/gkpjn0qbQfKa47RMjDTryFWFuJP7cjWfr1gDwblT
BF2JQDF4frJY/FJW6cDkczPGj7+yHNNMj51aTTztznScMUhvfrtr2mKqyOhI0Dqx
yLgqFfyBi6fdsngziBJliDMb4pzBsjIyIiLL6/Dn58pNhqQg0TEjhKaYoYzGuLVr
mBREsRiz7h3xwKx5BZmR58Gpe9ij5U0qzm1VIPleVk/yLdaM22++1wkvkJa2Swny
22NlzFO4Kz38+VEOE0R52g49EupmHdFsNWLREKeK8384nKU92kJZW30nerWXWkSR
nhe8akBCw9+8JdLn2BReYAJp8FnUEm2KzJ9sn3k/OlsannHD52QPeYt85UWnxD8q
wbAieG8sGnyZvBjT7+nWs72PTMr8tzRbS+Utb2IMtXr8uqqI5z2sZb5bWqQjyYsU
EpxkwNAZLBfC0RfgCGR0O2z0tOT5kjA5Kr+EBy8KLv7AG9656jeZBlT+BRcZgA8X
pi3ASofj9IOQ4LUN8Tnyo28iXINtRNiFskV5/NbqiKs6s5s10FvcbjfGsvfpWc6m
Rmw2nrQ6jK5UlVp7r0cypnk1s/rck9WSLLWUUSrvt/WKfMlbP+VuSM5eid0EWOj5
2A0CDIhdj3DTjdlYCLyZiWac06nw6AhVsInAk2Esh3luoskA5FVu5udx4wCGC2JK
ZMPVD5JPV8yAJEke/V20GqJ+ztYalekt4SEHh6B0Z+iuWEbsV6soSQDEjQ4FbQRm
eb5qkqZ+NIvDpM1zu2ZEZd1fBEjcipzu1mXB0SgmKY7vi3R/8Kirvj/r82NnJZZT
50FzirgeSbv9iKj2grP4qfZfpPyjTim7SpYXj4Ti13vr9y/Ev0FoGtxXCkiE2ar0
nS2TeIiUdpv3fffgmuOwyXH+XOaF/RQ4Pf2t+7E4Nf39Nq06VSxWirGqJmvSGyCA
4y85m+jCxO0pcubXS77je6APQDTj1M+3WATuZ5RfoAUIUlXyfbuaUIKy9A1bjaVl
XbgD5LFum/dPXjyeOSKGnKW2maC6u920cYyC+v7jkPWcd41tcbmRjcWvOAcIWW0e
fTFrxEBpT884jXH4GvfIjkcm6wouOCkGtb6VWBToK5Ngod3lpjdaTKa/S2KOlRz1
13s62sM88pXIV20RIl0tAgBCZ/GAAZcGZmw1FXn9iWK7iTlBml4ccqaw1K/hJB//
SMnDjhWI2ocNt4fKmEv+RFEvtVd82We8y/Nh4i32mde9xcKyaPI8EgqpMyD7qr21
GTHAbEKjShJHPLelpb1/yh8TuF6AtZrpRar0Hs5TbJDpQEDvAF5eXvL/TJ6oF/2U
SFnWMUqD1O41Js3V6tBmzNUd0jzZ5/QTUTPoweJ07vjPHP+G5VjTftMccLf8jDDO
006lNA3STj6ccFzqU/q/GHtQOuHbwObMPzKOeTofKk0ATVUA07vBBcdiaO1HOMmx
m4OXbGMEnZzdIVYhX1yr3QAdk0gOT8h1JVD/AO55l+Yk2uEJXtXNV+AtZGU6vYQX
b3xIuANrT1LY163VMrF4CK7r+FtnMfwjWTahU3TFileajWF5VRLtkVgjhJMyBosr
cT6dvCNlPCuqoH8WBjlFH15uzEek1MWKqwE5JLrBxRp27cwLU7ULeBGV91LM0BLz
WLjnG2xcpZCX/SfcEBA0yuZ7wbtUgYy2h6UsY0C6pE+MHubNZA+DXp3yVQNEj+un
R16J0Mrxx3E6FHipDmWn9DCo7TvWEKka5Zecws0GbI5Zl+SNWK8szf2y21XOl2mb
tunAlV+LrmReMaUIkgekJlbn8SahHzOfd5M60zeAXYsREbTrBjmAGmm8Z4HFafKf
GAAgZiV6396aeapnNfTDkZxNaYVJZWmE7gEclGvnlZb1YtGBiz6XhJOO3vz9+vSs
sqMIFCU098GU3J1ymIzwDlYzLs07J6d+WHnM6whyqpATPMBO9xeo+zGRZq2UpsF8
qZEgoKRdweGBYode76Dpi+EGkJ4IiO3kXqn1sbTBMd3kj7j3+fvayPRghTOjVd0r
dbvlyOcjcljlogmqN47/Dx2o4jS16NEC3srr4fbY3wpn1ISVlU2gbqxDOSeEn+Dt
ItHOVF95cCXT+329XorZC3MFnDK/ghUIhChjZsj9RJdR+rJ5IGpZubggmByyWMiV
JxNuhHcwEsgYjh+WlFw4T/p2hspDIua+vsCrbNrlCdVR9ZuGlAVpJE6h8k+sepfq
5A6EaBiFiVU/ye14gNoIJmLEU+526R//rcNpf4+/lIeWkgWwY4klAlcTPYSv5+XB
kCG0m6A5uM3uZDDhy/LYUUYW8fHT3ioFmDNu29FhP+tj0HZFBWC6I5cT3JyaxecU
8wdXIr6dRo7IwkPygQl/MBeaMdURdfdafNK8yA2cXJ5ihlAXHGULwuojip7g92pf
RBYUJBR7ZsOjnBRIfDx4gOU6xUpnndxJyVJpJYINfOn5jtrIXqjtToh+zYDiN7dj
eH+6kBNb3IQNQUex39rE7Z2nFD5H5YEJiViMf2edTle6EO6QpSRc7qOT+xu4TYh0
NfcOEgVbfTttXWwOnyJEmdeON6MM69Nf10K9AjgOUmuWoSI14rqJdn1n3B6oVbOO
T+g3JVOfioNpHj1zLVPjoA69vxE0u8TI17Hb0b10dzS0X/0apvUde0nyz/tpke09
wCxHlFuf9D8Y7/rKPjVVLfyXGioCKL5X45xXEi1hjh5LDJRwW8iS0N5gAwxnhrUq
z7ZJEsM8JLLHxpjmCV6cfoHn/5KTcXM7+V7dU1OPG/8tUDY0qKLHiuZfdFO9vcol
pZs4ktm6EsR2q6AgTYBiHHTkyXoQ1C7vYXV4oQ6vLJgnUYj41GEKwR/IfXJvggCX
xtqQnH+DujSkWt5gkLh7Ps/XQLbey66PygmQRUyhBoGBdopE2pMgIz7oakKq/NEz
NFfB3K5IpwfV6vgdpTnMh6Nz2KVIT2NyRascv+SuuaC60aNnYu7Vkba2IWdzmp8w
8wa1GizjmXihNnW7SC2+ktmog0unIv5KheQM5Y/hCK3LYACvR3BnO+3qExpppHbA
bdZChduS1U/nP8T82tBa2bJi6wk5AR+vhDYXme7+17weE6WRwwkF4sO/MkWAlOUd
gugmlZHCNtkxSrq+DyGnNXBAZmUL+Un4ISLmUm+V+J9MeL3/46Rwsf1X+f6DKoW+
knC+WQvo1nvvtXiT0ESkDScLB+pX0SFbzXPnKcmMCuzYEpYK+pEOm3IHKZ/Y7E3V
j2bmdZLuj+sVg6FzAeqBTC7q5rj+Sw+vjln+bOQR0aDYA6psLjw9S/qACVrnrkyE
AZu0R8ulPkmJ+BGmIzC/toqtBzpAsUfCwGZeFptXdxPf722WvhUVXRlm1nXiqApw
tzpoSE0d2TsytwGdQ8pALY1eyI71tg8Cx9/P3edXL80Xce6McXbL+0NgjUWgfoyX
1q6VrLYC3BvvQqAbtNnth2caeMcgNlkRhhaI4zpUl90UhDekOcceJ/udSI2Jr2S0
adgzCixzd8lzewRTqeB5dIdqncQFu4z8gEbFGav2VT1Ymq9tZ+d+px7hlr/P+veK
BGmAc+V8txHa9cZ32V9MEcFrAOhaiOufkhBdLVFkiAabitdMzJ8MAvivMQjscxRn
ExciHGkk4pQjeTTLo4M8GW1nAxxnms3LrYWAfi7bZBaeini4sxvlm/4lQCiaDcCJ
+okRyOtFXqVawZ28ERbwqbV70QtkvSReWO063sky4wgFMdSCoZ0R0omFcE/3ZA8h
/JFgTn1PwGMQMIlCMbn65PTHeIVSFNb9Bauo157kxzSjK1iPvxIAM/4ZcFEgC/Bz
SuU9LPjB6I+rYodRNh4N4yIgZbC+lykFMRH9v+mvPvoaFkNelhAzBjPV37+LmxfE
DTz6dinKvhEKZPuN4VAcBKwNXSApHOWYCGMtBjiUAmhkc/5Ir0OxGnUHqfFuQzXj
D1EdmH/R9nBxmNp2e+V/aQrF4swXLclN0Ym0FhHZ8B+t6O2du26O+aXwlm28UNg0
Opc/webBX8Vr/0wAwwvGYEL2640p8lOMzE/eyMcAMAwPeTwh56oGAHCrm2grjnvc
Rue2CIlQkT9sGg7aihz1WIWEk9R47aH9iquzHFZxmdHpCtos4ioFQ7AvkIvyv8rR
EDJHlygD+klsellkrGDjDg7gvp2EqaF0NvpT0hIwuSDazcJBSsOdKPgxh+FS5xKD
VHTWUpI3dYzco0LBnJwOAsKg0jvyZKYb9J4KEVoSvycd6GZueSF5B6szPyCpWWld
VbrgRybCjGcjjktHMBKEgxguGAsuUrxls92h09eHR1xjHRXJasX1fjgpBngZp8Zc
SFAzV1lFKJ5ln1VkLFBPWyQS6eTivi/VwQctnDo74L9O/t9jtT9HcrlOd1BqBjSM
6NxO34mRHaClkAn4K8PrnrlRt39KraiLl/1dybZTgqXw7LJYoyrsGIhwER66zvCn
VwWNzSA7z7gDAX/UbetlTkMDEW7cmrOiR4iLbYKj0R8k5auNRLRlzWsS1LXSRQ8S
XdHEXHpE5pxm/8ki/0nW+72sCEK0k8ABVKbQyJA8EuN9gVhqlUGKWl49q/QVItga
iUx0HAZit0KSlgkiJXyxJAfgnFFfCrRMbhOaLaLzrilu1xgSnOumORq7OA3QjpIG
3FWynTDMYLMsAJXffi5A+XygZR6Bez1OefofKgZoN0tq4XrzvrXMbqCGKAyiXuDV
9NqNK5WvCptAG3abKYgqMNJ6FKYZGAH19li+W7uSVoaVbARrJcCgnrnoOmj+lhxB
bfosrQswLS0h75+5OTCGgIHQgVnZNBc6cpM50zXOid6+FjJFuHoVp8bP2N2bzg95
VbVxVrW78fgmxjTRYQQLLRsxj8KK2Gjb4Kwm9VIOgkBfeMadgwEbgDivvH61Ie0p
1lmERecEKrgFRAZxASZqqvaNyY7kzv7T0Ag7DWN4ET+WHniEwzSYi7Atii3uIHws
tL1Sg9HKtDXed8+Pinw+ehFpcqPdulBgKfOvV2VzCADIh10sFgnLjyFn4w4U/4VD
SZD8S/wC/yFaEpBHeijw9iEHeIGYA5G884blwKpu3D6xtAdSSXJzu8Yd8oruiyvA
dESuPi4p1z7S76ZggZmcHsj9DxFOYf1abBluCe35MfJ7Xjq7uNdjuY79ZzzYf4vj
XLAu5oNVzC+ShaF+Es2zalH/XauFPt7R/q2os2CG4ygp7OJ5tjw/9P92dmEMJuC4
kbzMHB1veaxPeodMYUgqrvFhGC6sxFArihpcj6/4f3ecZ+y0krctQufHJFbx2nD+
l/IaYHZ32lqA/j0g0SQqUulYZyHN2xHaJwxPDkT4d0/acAhJuFL1U6L9n5dyrqAm
+PzgMIM/q5G/TCNcY95Da3Zj104Cyzoe+T80q7gFI8Fo9vWUvDRO+S5nGfTojN+I
9LSNf48ARy5zkbnSl+uAAnVYsKl7XePRZQuWVNsuYoQ3Uuba42PBnWdNt0uNFD8c
T+L0gOnSJzAr5MbmIHHDtZp9oqbd+EpNRqaGektWTGTH3CDiLIVC3clD3LoxBa5I
Q+FlimmTHcONglxfevb18Lmo1rtiZKFUkiABY/cWsbtXVWjPRsWz+uyLc1Y5/tdn
81B3oVHiHakBAaKbX28stbMBngIplgzlfkQZzJjdbNj/NikxKdFae35JBx1RXCQz
MQrtMZ01/dguoO83MB3oxUC92gp52VXt9czU73D2oMp6/Jxc63ZunhP8M+1pd7bq
lU+2CrcHFkPkMgC+moidZUeSCW3cXHYV5OBr/qU1wnI2GUuOAVDW/K88IGERJ1vU
AfN5kOrVehpicKbK/CjcjLj8IQW875vfcvJeMduP0kmhktTd9cLBSAB8MpLViuh0
AEK5IDcNDims276mzoD3eu+LYVbQhD2yJDQZd9Z6g+mGLIqMC6FJ4YBh86b/84ZE
82oBCyDxh+j2pzHut/lJF0kcITia5pl8k3jQwXe1V0pjHmiq+ZJlGUfDG0p5b+0f
L8rXyYOE0ifVIlvEGy9ct3iFvUuFS9sEIaaJC0pdpruKZVAGghfjnCPQgmb2vhFQ
OrTBLERODw17bvaF2NLw/mFI2+ICC7BsEAUxJbX25nsh3RNMo66wseTxGo88kSP/
ZGevz/Bnq69hBhgvU3wbduk2Tzkw1Ge+cqz6tkUZ2O+FiUOOt9tD9lPR87NCxtbj
BG8bNSUwWqW3GW0AUGbRDyeb3bLTjYRsrPAvT/XfwQ26gg9680jjTClRVaM7t9zb
UuJtHrPwgpe9oQbqtn1xjnbyg7Ir/DJ09NLGp2aaraM48ntPbSjXqukc8LdYf5K2
ReV41tx6xAQ11a89Xf3BTfdo2QlIDZqB1vMn0Jj1NmRNwc3PQJltTkOSTFC05WkD
gH0xAqcpvuJDc8qUT4JgEHSNvjoH1GgVKLMG4pJlOffhFVYNyuEyMcgxrS/790z9
iDDPd68UZUX5R+iSVbsGnh/8HzeG+YNY2CWlWMKPF34TgGtBS1uDQCHG/Koz9YLH
lXuCeegRl0CREiq/H8JhpgeuVpawkNgxheaGHQUlRjqzWz91OagPx9IpKjqRcBk2
UMfMe9ASyB76M0+Jna2uvxHo+n73qgYeNkQYcmWqL/IA6JtvEDWhIWXLjNdUdrIF
6XLUepzk2E89u8axQK9G2G0SA2cxSgcMF0W5Xet6In+oy5qFwstaUFmT9yzhaOlO
GBo9mD7s6Tr+KSgQCwZYsqgoy89p9ZVpVfCkqp6ftERvxGi4m49QK4IjT0V0Viw5
/CM04sPYfb38wmgaUHM4QeyXi0BN+9bDHcejGgHAclo5q1GTAF0G383oGYz8mzyG
SXTuB2IxqxAwA/4gjcMOdCwJZy5tXGahQqRZX5MCOzp23x10OScVs+m2g3GGvMDy
hVuiQzL85Dj0Xy9O/tBgAg53TWxwatMSvb49+MbIX4tr8sS+0MrnktrWCbbPROlD
MgyiyixNRwBZUPgNntE0xDi2iW33hXFJspyJiiS8pb/x7gfMdTf7inTIz857Okt4
ROsB6vb2yjrAeBNnhWY9m0bv1ewPKpvQrjrJBQeQu+vor5oXLKplmwjZw5YvhGMm
mMyfBAlpJzD/y0nUnpJ4trgakMrA7ov7G2jzsr3CxS6JtI+remoaMNpXws7AMS1s
Am/Yi0tsLB8jPU+tPYDYvc/hWg37+ratrKE8xhaLJEdTYeXBfm93det0V4qYWoRs
WDgmbSW0B56nt8qIQPYuJqnCUIvspSo35fVydbtARzD6TtEzxTJAJ1gxSMgdaEd0
Wx2HibN5ApZi8CMusLln7VbIG7MZfGtlHlAXdOpAi63K16hrpODUIz6rD139eAUx
dueFOetId09FI50yvceAqcduwgTuGS/T+ZekFddqeCblFh7JqVX6TuIgY9YnoLnX
FalieDLI8RbZD2AbiXTEekcIDe9tvZCmTNiXYsCA+LwYR5xvbcr7gKacF36gRosg
Jf54gQMN/OK21A29GDsgkQ4BDLpZM5ztp8xknJZuyvjxVjQ+4GOr3eKKI+hVm7yz
cnmAQb+Eh3/CKt8YjmpmHeAkghPA3Ag31Udz3ef7PHi7GxqtUu8tiNrZpa15eWKt
lnPE/hKncX2hAqkqap+68pwaEmZF9bCwQoYg6HRPU0PEjfLwDrKXIFkOzgOXWRPu
DskWCdHwv6NtCg2Ji32y8TwQUNXiToscj+ykkfe1dYYtkGLozQrlncqauYf/Sf6E
dImS0Ft4dxLgcqWDLBk02Cs+iCGASFPYLriTU/1/RMZoxoRzWO9pknIT3gYrDQ2Q
Bz6CGQ3SstnwNncHNt2NVXxKHGeoLQ2pcHz+L3jMP0VCfmAKJxfiNRSTtjLNK50H
ZbnjwjiGyPD+0FAeKZMM1wsFYEoOrOYvcGvqWYVsJAENPdURugaldgQ5YMVfgVkP
AiXDHxkM8GkjS1i7O8Cy4fqcu3uxZPQalCCqyXQLwMigYQwSYji4PWfooKt7n6vH
e/FYvCGGkhQ5HokwVOq7+MYTbL8NeBFWF3NI8g98cPVNUAZhcIPooGQSDqMqDb2u
qtHl06izDxin/AsnF/JXqBZD2rWi2U2e7igKoaUpg4/5Tf8umj25FkCgrzNgSxjl
mqnbhp1Jpbrh0afDMhKjwHcIdMp8k13OQbTqxGNkdgz0fd5SViEv3X6s3DimPqhG
B4qPGdlKcEkoYAvkKZvcjPosdwAgsDbnPUc/TxWTrKEybJaTbnAW2z//Ay6qsUIx
WE8+lpUOCNTQiik2RSQjJxjZ7NuHUvB5WJLpKZxQWYe3Vb4iQ4OdTDNcqEft9/sm
cvA0pHnf4unc+eC5ogyzgslt62mgqK4fU1e6K31lTgQwtGVpmlRzEuo+SiVdFc2b
FclokDkxYB2JDqrFeik7lbJccFZTtdbeP4EUJNDITJ2MgVEMwAxDP0pa9HQEXcrt
E58XhmU2DAsJmQirDELI0HYFRcTxeEvZaFvsmT5PqXKH/dyGPlu4815WkwcYt9u+
OxYx4X3P6TW/u5LmUkntBYF8y8xqENtCT0f98HFS7GFHQ/y6Bn+jtgiR62qRn8Yw
HQ/3nzYpgDor/JIgFQB3U6av4xQ39/JqscWYKqtLhb3H/NSq0IuQAEM70h8oHCav
SJTERbWJxQabHKZOOnwtpqvDqaatlUY5awzOxaCf2iLdprEiYKXatfAZbgctnDMP
CWJIOF1/zXhgGKoAVrxQk3+qGrwdyG5Poa0X8+EW/lODWyJYee5vMaul5tqy1G32
v30B77T+NRMqPq9xmwLZs4oIqfTOqi49+yTmRUc95abQA3d2eh8/qVlAlRuiNpIn
I7miOROkhYLKBvPh/g5I2SZrzfNONl2+EVxVUGx+PoEnawZBvZp7F8JF2waF6rZk
1uFyurRD0k7xEu/kdBHjCe48q+IGHKdty5/OgfePjIa0m95zangINbZ3Fq5hxehw
ah80RYVDzOlg875SdnIGyghukJe16nR5IQzOskMv+LffwaiQm3fFJ372/XTuNldA
RPp+ohtxDPEEqsycNBRmkbviFzt+1EvVFeev0UYb/8RqQ63AzrlmMUIoIjh1qD8I
xde3RelqRXA1k6XU2cIEtsK+NjtElphwvmsrtA++mgBpeptBPmHMXkhe0/l4o3f1
Orln0aqOz36VSjJXzamRST6NmdG4pL3HrKVGmEbKwfO0lJhs27c9o2YbTcEl3IUd
L3EHRqpkDdC0flPN61bxtRHfRy5zP9w5YAVBDvlV6XDDSOu+ohl+GgGtV/m4xwRm
dTfMS9P0s+Y8oLuuwDMSYsg+4ORiQ4TV80n+eU9x5cvv6GVmcqYgSdxwYG0Cpfyb
EwzORjZoGJPnA8vQR+l0gZFdMsCBSYRK11LWZyhBWNp8LWfyp0VTSi6XHOPBRfBW
Il2tUDqqeStBXKX++hQ7dGcuKlPSfognT77rSR+IEcukhGCNDJYfUl0iXb4lUJGC
KGZsn5s+CnrPRdw6AyIGvu3x+2+CSsw/BdiB+b8hTz1Hb0e90b84/5ON4V8ijdTY
OIL3loqiBtxLw3FusWZDs76/KkbXWRORI2psmTgrmnYpwAyfm3SsZpFta6hV8POp
F0GFZUdpYAi6dE4buVivJpkTQBBObZMY7ZYW4NH2KjkwyQhqsH4cafKkwNefBZHf
ZJFIbNUvbAtpzWUvt+qJburzZJwuviTvumdu7vAHItbXST+PID0vbfTWc2IDhdIw
ZvUKRughcISmmQuLRSBNjM3nd9T0b+IEEoStGTwlYqf82h+sBMyf0+KXmvuCPx2b
IWCrgrYpWjW3KPZOTR2YgkiOg0fIJvYOuAdbdEZAyYbSOGMa0d66xGYLdrge9yim
0WeDkpHhQspYmGP3HWXue+0Y8va3Qgyphb2NDwaPKDvZuDQgBajvkuahcx0jvWhL
qkbwVqHFqnS858sd20DzBYIxNagd56XoPXvZ9ArLQe/lkxBeHwEN4zDfFoKSdaYS
C8k0ArA68fUGDXbEKzWs/UZ1c2Bpgo50bCzkWb33f8g50d57UsP723wwKXoEsDf4
2aBOh+f0bMDFS1CZy+xY+aaDzKEm2qVHrR4Vr5c7nEdU9qUMIgxHssg2XpnBPSJg
JtivXtQr/5RMUPrGmJ2lssYLz9e8fGE5M4eizb4GsBnQDiQrFDxChw/pHEaFM/oZ
pTB9g9vlxjKxjIp+7IoO4nTvV5qaQpEcJi2t7lrs5PYoPFC6Nnt/Yx7i7kPoRKO4
CccOPNko5ys5Y+iTHOxlPQNcL4zpzgw+fF5SvRZadpv6UXI7r+rVYKXS7zQMcHhn
8ZgWLabij88cTRNfoFjPPCBliBCFUnLJn8Yq6Dv1uEx7QvtTZgmRASNdPmR0hOHQ
kKbaJJ7oZJsXecxVHhbuv0PkuldWd39f9WekAv67eDYexeyHuJwmQ2b1ySjplVpx
qj2EkbnYMMtJFnDSV9VtLxIF89/wh5pa5AyjFgPCAbIb+UUZ0NU5p1QCBPKsV3QR
EHcHNflBdHUbuX70UUgXJUqrAsaE5ZJ8ZR/dn6cZ1mjbrIQYxnmAIh2H9lXJncsa
Gs3nwjXczd0APM6yClRlDCuPAF0iXsnTePTnqHOboiG6ZOZJAYf8XqUyxCrkVS6a
lzqDLiiflUFyTygbwg1guXmWsXNIugSZ+KK2SN+KCl5VLE8yFalybInIQBCRXeKu
w5cU1iebYOUret/tQSTyUtCVGA+jSbSU+8USqXTW2hLziNChM+m924UTYZ/plWVv
DWrqJk9xbvBCnJer++E40zxVXnEASBKZCzJqIRMEx4DVnKsjbkp6raza2UGT9F5J
urG4AMUQw5SGEIyDO+iXkUPqcstEp6sAuYqWITqtBHwHAYhXcSLyaeZl51FWTnjC
ZucggjMGiRje04nZvak0lLGU43c8F1O6C/WB1J9VIU2tPLXTV0TEoR1ZfB/wsQyL
iPKTmBvAC6u/AicacE2a+rTIqDXReGMKMITjevQ2w9sSYlMLGS4P7COmLqwLtIhV
3QRkyHHfY7vjZR4JEwTTQS8EtUmN0WWVQfna7SgDrbqy/YpPXoajc53yKiAxptfQ
8sgbnJXLa59MLnQsut8YnZ/dSJ1WJkSP2zx2kD2RTrzleW8vdJH1To56BHfmZeqA
fLtE0GVq7ZPHqUq0H39HyUAYnUlIq/AU3UkkmTldFQIiN1dP4l5YA0PgBA0M2zGR
YVUlux5jfh9WCp7ErCPpWXoVDmaEUKMPlU5t8BPMObzUgFySvubHYwLDRnNqj70a
wMkaRBGz8oMhslp9rs11zukxkjTXAUA8l5BYFSnfsvuPOQNHYc3Fy1roB1eTqjyC
kOWasbptP2lWmKhXq4CRTiSk6iOmF0qGXLZesLXBUsaWh1dAPAxECJkqAs8jMPQh
doRhrXDuHu83ln2/zFPtviAcmNG3w+K6InLBxOEDWLFHoq6+Jgp1nCdp9cbPtEGq
lO3dbuZX/3CxGCHjk1eJNzl87Ma9hnYSvoGwQ/wDQ+gy+QHKWEVNY/admqjw9iqr
u1d36D1GtvzmtPyYsVqBylnvk6KLBLI0Hf0TsmDlB/I4O7i8tKJcIHA7ZUwy5J0U
WAxSI+I/yLrcjhwUFpUy8VXF9Jsg00mzl0ZPtiPyCXeb0WbLZg21n8QeuIbXtYnY
eKxjWiiwu0ymadSNnjPUescjxFEMM0dLuVcxkXINmYKbE3ed1AufG2GFiN5ICNWz
1Ag3wM3/pPTOwOCqEP/RkWrxSV2kVn97ZDtm3suxdltWYKqRiv4i0OHrg6R3nc9e
154hsepm0zN4MXFVFQWbXea8Gc86g0an2MZvjAl+QLdAEEB4LxHYFee6NGViO/ot
9/2pbQEMUNbkAXTq+nLajWZY5Dp63JBiOVinwGE9/ljcUgaJScQStn7lTwL4ggWZ
PQMcagF+AIw7zsYr1vNIkMBrlCiFA9a6+BSjejd7mct9X/VmR9rjBEF0woxNbYrX
7qAeRzNCv7Uokfs9kmobv1LzmN400Wf2vYMkBNgICSV/ybOZET2eVRwDfSKyjtlJ
zaBSu9ag+uG8OkEmAWlR8Y+uROdDX6QRcHaBvujRo7kauSFSde4PkqNH09j31c7B
8uq6atBt4ZEVD4eCCNgGEzPmDDhnZg6jJVGvabPI1q0Xk2tGGuuSElrkGtrUwOv+
wPfq3J7i7Se65wV8wT6tmgSgtC6ZvdJ6HX0+YhCnCS1BkkdLYGuudv25wPZtAKiA
rB3hgrIAneOlSzA4tEHdV+RZA0P3Jxad0XAoKLQcQIdUCzQ8iRHZd+fDhMrXaj5f
gLUTnZVV7nuBOuV+JZ+ClZOYGVj/YH4qKXhUVfIp0Mpa9zYlzV8WGz1Tb2WwJ64A
wr38hvciI7lXw30VhhIquDlZaBaW390bGDc2qS+AxMUsvAjMB9i2/PO3sBilc6gs
A/LwrOILRif16RNupu+yuiJKMvYUCSpoX6LnxXo1P0MDd4XzFWXKuuobIIML1WWx
8vJdKvOkalIZ/rrUNJDDZKEpFy562lfRf6WYx/vcTpjnyr1P6yha61ZDlTeOxAxx
8fD26UC+wHItCRTmsvyUe+48mnoZnv/UlLU1sbI84V/51wLbxukI7flqKKcc8iLu
xnchzT3Tn23TWSfKzL5493bBnhd++iE1/4TcvIODKtt+dYRhVfYXQpxJW+D9f4t3
xQK7Iw48Igr+oRnY2zw7SOdvwl2+ZYj7+NMF9XSM+xSXEfY3An+XL2Qlq0xI6drc
QGUwFoZggUiGc7jKLbAYkiqQaa8bVUHv0RDKAkva85nClRN8v8AWzvFfV3nNFc/B
8WxBKqB9+ItI6GoQNSGXaeZBaPP4FipW9zAqiTp6YtPtAK2MG0mLb850oaecz2sP
sNtnkWR0R6zuC9iQ35cnW7+S50nhiuQsEab3DTGd8DXes5pfejuQeEkimzUXJbvF
wpAYJLZd7fOuZySfT9FYoOe/0AeG4acRcH/Wc/mj01eRxhy/ZLAgPE+o4vwwA/9M
z0h/0t9urkcwVU14qvk4V6BsOXijpI31swVWXjHomme+UZ3Xiz23o3jxrnXA1Pcj
NQ8VjkqcU9USHT9u4uWMUDM2Wc3qAUvH2jDor8hU+gumBn8LBWLYnMwNbAGODlXS
qowTtNVwgY+OTNJg3gb8Qd4wunJdynhqQXnZwhtCkrlGe08n6PmnGld5BIkLbIwZ
l0VoXpmWk72beo0cgrV1FTLH/pQO/DrW8cywgcwPVdRBgtXm8evbzO+ponJCWdJK
8MLb2FbK6EqoMc2PkZY2ROxubIPUfS0XvBdFi9b09utLWgb2PIV9qZaySkKRAiM2
OBIx9x+2Y/nSBticm0l1mddYTYrZIWes3iQS8NOzqp+cCroHKbV+g9DpllTQFUUe
ImLsDqyfl2Vc6Ud+JViQSKbh4ti7zyaeIup4PSK+Y9Id7/NS80BF5AXHvd/7kRlL
U8ZIAa6Y35DmXclxr/bTkc1TOOPi0eKhzU5Y34Ug4HfvdnHrDVsFDQzNRsvORXM/
ZyLCKqU7arlSF46VE4kRD9NtErNeVOFeA2isBzdlCCpKDDzPr4Y5qa/nTU3dPhxF
so6rPhT11kehGm8eBZMH9cwUDPxsHyEP1mc+IgSmKjzrRDCNvmcXCWwixouG9k42
kQFb+LdlfdEWpJttt9cZj7dMVSSFRPVwYasaGk1dTgxtjeofia82fZ94i8Ewta33
v4BNdAXMCw8kCE8UVAGC+PsTHXLK4qKKrnhY9ZgXGIFlHtnEyRGppfPIaeyaBV8m
61GxWN/PArmpOJNTiqop1CSV87qEfLwazwnx2WU1aBp+pIsSi4DvoW+HaKk+XBo7
mdtHNmB3q3XSCBSTtKwsiktsKRfs7SHQJx3a89aGeoQAYYhS5A7PU+Zap9Zq6uJk
80amKKWag0YIpc1JRF/P4+JFtedTT9iJ6oQ5Cjkt9P4B1pEzA/fE3QODFWuxq5Px
9srjo435K80ewf+bP/syL4VUJiTOEZoDDEqYbm2I6kNxCTme8FPR3CyJDbZvPsZF
7WrrL02ks01zmDwAZ/ejVBfFxG3wzhmPd/l2MQkUcdQnnOB4W6yph5guqFi0QKpx
6pabjGUHMy3lujhBgLU5IVhc5OiAEpdTgUOtHpLhYJp90sE4iGMgkuItcCHgF2Hp
XblFZf9Hqgen4YTqHVYLKpGLtFSXROK5EYvxmAFQoOKjNWcYBtRCWJ0UsiMSpk6B
pknaS9g9k/o4WjQX9TDs8Yse1w/aUjoHR8SIeb9L3ooe/D27evkQV2Rl2PC493qN
jeyXklxJvOIfox5dFPEDpyBZwMFBW8bPuM1YLbXfziyiz87S3AZfQ8n3ACRbfHzd
Qi+yGNhGPCWcLC27NL8xSw8HhfcZLgzlGE++rA6SNRb3jACUSxDdrAnzp9DGZfCy
3TByYVpe/+28bo/K/HtOjFC9mHACA9F4Hj4pS96qFuTc4gBRTmHQtASGVlO+lr88
GDztOOZc6hA53vM+W4RaP4dBWprhFXtixVQo0XKBEYdtQU8AAydP+kAJyKo1wZPa
DcTt3h5lveZN01wpDZFyMQXtsmF/UAjSexLqWHwMxPhvTUjU8wccNGhG5qDEH/ne
AOTECEeqvVumW6cpGLqi3mFuPkmr9fGwZ5/Zzon/jfRJBjDXkP7i99FlKjc2+4aV
drP7MZVvn4z8zZDxIRA4kXEuy03ceguLzvzJfy4K1Ya71z3EBqp3HM5zi58j4kE6
jHSlwKGcXhi8DQyvaLk/WoBJlpGV4IUMcaVKc/+rQ0E/WIaMpUd3fEETY3kTRyEd
BkiFEC8xrIs/xURlyY60Ksr8azV3GrIkbi5pCtFAU2hFTXekBrIjTMS6wI9xH9qh
0icQNqVI1VTpPzxg9ZNSGFzqRb3GfnAd+JOqD6hT9kzFO+iizMozQ8K8Wq2h4cJI
GTdVrpdrCqhoMhX2hwhtQcTm0L9icqqLptCU8S4NsnZx1ycZAMJ7rTgFAdk4x4zb
LZSkYBoubzOQqM+UH3DC8MKxmXQd2mo8GD4z3yF7kWU9U+61pClIwCzE7IgLdF5M
yqXLhqxmI0R4d8caOSsQ9QAx+/VmwLM/MW+YUqoFa73OGHTt5vgRiDTCu06B+0VS
SAL3O/o3QXRLJIX+I4qstbrVDYGDZOfA2mcKUPncTaH3b3lzTa4QqvI9bHdAuLZn
ADat5Tavlxse13j96xvWa8s0hMI2NhQeA6WsgbeYvXiZQgKFguO5kATvvvfjq9q1
DNyBOZz30IXrrqG7okkUfX38DuoXeC3Zdak9mlVWPzxvAij9TMgA126mNH/UnSMz
oyoD8mFL/x4cO9/pqYGxBco0hiicLucAR5O+j2rcAr48/d+yM1/uDK3uWvN+/N2u
HQMIaKWE7ca+kXfxatXqYGHaYtwNd//sGDRR2xsHTIY7pbhm9K3Adh5nhHljo9sP
A66Lp0yZisl5XVYa98rRrDNxD6Piv6Osvfzz1GkFkzNMYOYZagWZ/PsV0+EcafxI
sZtoc5dFnr/ltUmF+QZxy9D1io8lpiaBCXeUikzjnrEuh49jAbH5Z/HyKKmqen06
orTTX6UhLXnsaSmoticvk19J7eU+RSoDbdc5tTPzsFhV66NLtA5mSqpT8iD4mTmz
KnCOPRDYm0kJmbL6ex0mBf4BcRiZbq2+Cn+uxohLLv1WXFV7lbTbpPSM7YGF+nr4
4NvjOkB/p2qsa2hNpoAm05EiAH7Pm61JVlF8B7lEgV8KZnzh1QPodYR32WUsIhdu
AHyE3Dc0smAxhOcN5z7Vc7d4fOzPyFpLpT5+Zy2FVBVRqgExddHdqCpsd4H0nR1Z
jFJe7TPyU3lTqvIJJxBFcUIkqcq0tctRFJ3GQ0s5zW2NjNK8fLHNzN7KwEUB4Zdz
R2+aFjJHXVd2tnQAfhYYEFTag6s6cZ0x6jZxBJcKfc/v3j2xycnxpPYX8XHg94x3
MfJfO+knMynYRjuByCWDny3tCbzuJba/kDBkez87lrhTl9xK5eladuLw+BqisFoH
mC1xgDKT3zjQjakDFgXYf8zo5SNjgG7kANw9bwGAs48ykF0Q2E9bG+ZpvSh0KJrb
RJZqBUpc0Pwlqu+xftFPoJoREkEeIvrU6E9H5k41f9VwaLabtQmB909TiOfteAMY
3duXULfSVb+/NXh4404shslXtD01Hvf26GMrSnEOU4JhljNWc4Iwngj9nloKzs7T
a49kUuynI7ME0qKOIDJGd611zwbprJyH/Xci0eo/9vOvTYugultqCwgFD9ln+FvW
yZej8d3ZALrtzB41e/BXbN7TcWIKHdzO2EjvRtW5H9b6gRn6V0PeQsi9/Y9wruOJ
Rx8OGqba+Rzwi7NPSmMjnH22UTSSPgfWvIk2luOo05ikcuHgs9pirvtetewh9YS7
Hhc31vL3LtGuNs3YvjApZu++0aIiTcrTxT+40fSQRKMjURuiONjCHqeKNxiIz5JF
hbZQM963mhPpfR1ClwamcK6cwhG66bGVECtX50SXBqFPmHISjYKlBOcHkrW0Uhvx
5oLNyEzgMTrZOAbLvBoc7Qmc1bGl8D9fo+1ybGPyIdT5raIKmajYg9XgyYRdh/aP
AJdFJ45Q/3XRwPXjrD49c4XJS1M8F83PJN0dw3n3l4K1izVntU3oxQoAGLF8JImy
Uun8nrQJ/+jQQKLPZ/xf00SqVhE6vCRy6bRHDAbjG9egNMsWiDkCwzyi19IoXCQs
azbAasMP3cEtr/17ue6N3SQVT32ZA6550ibVEUsslFMYfTGqjy06xxMrefgcpiUI
nm1WTyPrGGmvDOJqU8zKfcfsLe8jdl87E2NbwjQdNusKa5hXHu96kPKU6qVWX6Vz
HTXFZesS6zWHgMjylkuvS7hIUtqzLyRmwKxVCTDO5JcpB4jrQ8A2bQJekvsfY8eW
WlI2u8ACNeCxtk097vvu77CeMmhVDYUue5o8E/iiZOVEvIbgYdbDfH13CIqXHGRO
gQnmxFYsNC5gkPP2EdLnnhwjWCxMLmejSaDQaEDJIUrnhLUfyeEIHFbmAk4L+HJi
sq/DgynT652wIvSLxrT4ivKDXbNOkvzS6eS7guWkSFNoYhC7BuvQHLvqWdciiejX
l0HlpfuQoScXXzxmODm3eUQHVcMYZ2y+pvfyrf12h55vTlC+bCchQ9QqY9Ze8o/o
v0YO6XhRLBXwg0+S8ZXg/r4hcPT2v0m+2oRqJSE1vHjK5Ckpp4FxML1KNpv5Xbhp
0y4a0XynLsUZ9bJs5L+Yi+gPVvdgmnXOeNgvzEKFMbK3T8AtbriuuWkBsx14isau
RQt47q0DKlKEXtSqtoclb5vwZrD2Bw/ns2lfeL70t8OhEJnY3WNU8Aypxxvq447w
9QVfsBuhXqck+WG+d/ZIXDx/uYqI6g0VizP8RbbZuwD19imEoiYpcgg4OGfdb5ze
AAnKvNszgJtz5pTtRaQ+bYrZuByxTzgd/ZE3HntpadBNnfMoRTmQGmtj4XKrYvMV
zlDmlHvwSyh+sagAf0HqWIvIxQeS4ltsyE/+/mgS2UYEQDpycdYOkMjzfWvBKtTP
zB6UC0kxktaNvrekBSjYtZ+eJOT67QtTOBClvs5y2TVTTvPLLiGwivpao/mtuXwD
D0vWWEB3p7zbYsXFR71ileNxFNwtUZDBFUzhoWse+QIkSYuHqcW6ZfxynUvvKjLX
Cjl/q0ozryoGOGlFYMPwOMqDuZ2/64dLFapMi/L1TLPRCE/WwaiLuK/GWLVRlPUA
2VY7ySCKp03SPsHLmUAHWyhw9TDqnQuwpLLKGZlJq3fxJxGFmAe78ztXCrwpWHZt
I6U3Cn/tzzFd94XM/XSggR2mZf8dOtTkv0J4vUKVrPDxdngJNeZW2xscOpOGA3IJ
Ws9HPVdGPMeA+oquG/x2xjvBzhMq1kywDpUAe5LcwPlhx2Qh4cuywnDsoQkkJs6m
4xBTgylPzp9y8QEDXgqwfHP4tyTIXpd1fot9CF9PlflIAFdeubDUIZVEO2Qxp/RD
Qlr6gFsKlAt3zl4FhW0RpB0554HrAu+xkm+jrlabbRrkTA6LdorKwd2FxC4LTB4t
9TvfhuQIGfW2oqsBrS6J8py8kF1GR+RsaPG7ClBAYSoL1uby/8iS5QFnRW3y1O9f
scvrvEnR0PybG1N5XFxrwBljFDuRtlUUIlkBTBCkYBQzV61gWk+ve5F0S4tPiyd6
kczEX1iHlzvEk6X0FKYzcA3E9d6+DvBVWHMO9CR+pH4VWzUfbo6p0HZHpEU79ZKD
dsxijrfPBWg3jbTv8WORDL7Z/iNkCF9H5IDjFhZjFEp+WLtKY2aM+FS+dyjgpmpS
f7plpQ8auX/6OC5Fa5ahU+o73gMZyCOkq4x8zFYcz6EYExqZdTdTmskYcyg2RDjC
QUIv/EUPjYbRa6Huc2HXDoAKxSY1pSJ4WsPHgBpeBEh11kmjsxc7vFomzfzb2pFB
C+27fGa2BszI2cjzNuyGE74jfU5aORU7FC70l0XfgS7ZM146UFTkCHAIO3cIFHfA
pDvKgtkKqX/V50XwkM5CRNRkH9RugXnIi40QBTz5MLCyRc5xMcgzTRpBh75r6iOn
MWvAxf6Ws/Q+qebsekGLcmt0DKHx7zSH1a1T9gjSQEnEKxRFfyruRQ8YQaf6upmS
zD5uBZud6TI17YLvnZ/JbhmgWeEv6vDQafwtP/xyjiRbrsy23yWX+X+5LaPyTXTk
DriqqdwQhSsxcdXp6trNuEj7fpSf8F30SzFiBy1ywqFjmZp70foLZ7RrqFebiWeI
EYqWVGgiw5F1d78sZwei9tigof1zcaO+jtYgon7kDGPmog0whOyyTckvYr6wdoby
13HygV6tL9/bP60Y3zHu6EekCtH/cH5tBDLQb5NNC3o4yTZFPBk/ymZ7HRf5A1d1
Td6NjwI8l71xzY2V379NuW9kaanSHhtnZmtTGUKgJG89mAl78xdnxEymKhAqqvhJ
ooLwAAApl1YD54GYc90uWmj+5pNhSzwwKz2+SMaS73OOVbDA7xyGsJ40iGKUF4xe
TXaXSmITqKJIn+L8j2zZ5SRXu6sHXDS7olhYM+Rca7I2iG3mjU58m9wTvX+IUEfA
U8glm+CZyHjhf12Ay4WLPTDQWi9YWxPUGrTGI1gMmb/7vjkbjk4bE0axdT3OwDGh
eZs2C269k8NuqwhdzDV6tBeLfpYi0f0NfJG9lAWz266CXt9hQ3R2Cy/IcT3+TReS
hOSlIyQ/4+chSPnf+gFlamp1QEnQyUXb2LKyB1yWneFF0sMzqcY4xcW5jn9QLr/b
cZ4YEqa3TfXd8SFNisLcBep78rNye5nhjEpLOsOGuWOIbI8CsPhUEFOtBTGTHZnl
/mfJJ8edk6DpmFL2NF4+Klwyxucau0rC8hpoUgJ/bhUaWyHJwETv1GVXTHAjZreM
UG4uwKBmjIM8UdSd//1szeiVFO/pbJuOeB2whtdBhLtzrEwY5NQQ9wNuy3GFjLyt
y7leU5SEAn373fyVbH/fXXwe52bdzyCLhYXdoCapUz87aa2nCFlF+T1DSx0ggPMZ
7unbe+Jloj+S3UbP1GpXjd6AfDiPbJmfH48FBi+4NhZf2Gh9YA5EnlqBJFKRhz+P
ye5KuZQiKYG/oOCm6KBwliswjRCZHG1nUfpmuJLcxJHjBOXHGRi9aAltnJnkbhRS
1AVFdFuA73mFq/bZT9WSOoYdky+9Nwg1CYSc54bqgpnwI6a+T8r1hLlwNj7hh0Lp
TMohhKQnBojiCihbMWL+ReocbHLPmtu1YTvCMw57nms77l3ybBw/GAwL2xHXdfm2
TyIePqopKHqC03b+Q+97zcdGKXrCcfMcs3RBkr0blTldBgodqASrwr8F6+7n9GcT
qgj3WiIFHIy0ghYjxbT8fugUMMYZ4luun+02OIdV790g1ynx2tsXhbnGz/SKD8xZ
4jKT0C2l4K2tGh1Y6XBeT/TehrVI8PaDQj2iVCh26z+jvYjXLndsmapzICrhV+2T
Vtf1HGH0Ylr7mu/9J8RG9e1Wbi3dBHK8gMc4ZCfB1AVAVdF3qXl0wIzcphSNN0DL
4h6QXWrZPfXZ9His/m975d2Ir3chiu9D8wmQHVkeM1WDRjV/+hr78tFUuSNjRYAc
IHa+OriuQqmyEg+BSptOUD+8HV8EXqu18IajKAiL+CL5DHosdCx7d3WpurH+w/Db
3ftxAS05uqTOEbPM7hKGVDPB/PjeIHq2s8vVucK4GuEO8kGBDUuGNZOKUAWIlRd3
QNHO24wYGS8MVov9EmujwZnuGREHpjDWkiFkDObN7UbRCjZSbQIx6O8U3PkP6XPm
Gxlhyv/wU04XwzeyPujek64Bf/vYhl9vO/ncOVM7lUtE0P8GLZlUBf/69rQKInfd
TRNSNqhH/yFb5S3OnaIMbrBzZ4i2nKBjXLD+LBfAMtR09gr/3PjaMy02I/DSBk5u
LrQcpCVWbx6l7ImZuPXC+PuME7wSOBwyYQaPxdClnC86hM/JR3Ta4ooOb5hGTM0m
HbVNvhIkECXWprOUhMzGPF+AfyvUDV9ty2xwk5RjkyZqAUhPf9l3fuxNHN0AsLyU
ByG8rjo6UEZ4vJ9c1PcfX+nJ3DOhpvfSWd1D76WBjXXaQdGom855j0cx8ocm9U5i
JukFWbF+VFEXSlv7N3dEop+qhOdOUdslAFb8nr3ZxZroIaMEYfMXX+1KNinOepiL
MlHDcz4tprYuMxVO1Vyz7mpWDKNS6ew+6IxYzKJYoZdEaBxr2f15QGRjoqxhxyfY
w6LuwY4QFFuY9X0vfcS9gLkrlxejqWrFZKD2E3zc+855M3/5eCfmAu+trCmjoXEr
ZdJllXzelR0Dnpmlg9hZWhuGcxnNzsGv1ShYpVKIJ3kSIPgFCt5BHoH1yQ3qaxf1
WGnpvGZU/ePNA9ShsKGiIH6Brs5K/2TIjbrxK1MPjAeZlsNPSijaUjrt9/PWEL6e
IhKo9Ho6BqU7IvAC/zUTPG1P2iOaSjHTNqYATaKBgvICFXkdP5DD/MwJ2o1q/yQj
RFz+01V2e4TOU/0Wt8c286RrZQgPMZxZHNZZ0D95/akj3Bt1QEtI+DwJl9hDR4tY
1B2MvUqvlmzKrTgisS85yPd5LttoTzPse+yAkFOYm+Ene6KmirObj3++YZaVJvJp
UcD4LTV0gp1tK0K1S9s+nwdZchO0/WoZ8PZzd2pKSNeRoDmLY5ZS+7K3jQXhM5Bt
ydlLJLYY9azaQiyu6tutXc9Z37I0580X5XR2HkVuRj5bxXbnxT21eLabwCz+Jrvw
/MvBxS4V39fXV7Vrya6fV8eeBckMHnn3TY+Xmh0ZWOUPjdm6A5R8vw0EtfqwqxKj
vLV3gRxmx0nhu3qD65vknKi42wOsns6zOjus1M8OjHMZeWWFMYgRC6CPFIqOTPNO
5YdIMmDMh5duri+l2i4hmk5akps9xfR6XVEXPyZ7JrPqe8b/KqQL3kQ19USaCrFv
/4vU8s4f1y20NmAlJkzmlEZCZViqu+AGAWyPM0EMciF3cWK40+E2SWKSCgcIAsUH
54WPSdMvUAi6YM7KGQlYHqEQkTAoVze1/X5Ubqon/gt92RB2zCokf4adGfRm00Y+
uL7VhS3PZtRotoGuyZu/DeDDXqq3cOgdrM0NnkwE8JAUF5oH14PfMpPeD/XH+amy
0xwgWe4ObSVm3zTvR99iCbo0vBWeXn8MJI0orcQ9ihKlcsUIfklotgQXZ2O8Sb1t
c67Jjd7AdgRDUhU6je3spPy4pJPQXSNUSDH5x+RIQ5UqWHF70dUTTPEAryOz7qFF
a8q4FbVBUhgIIzc6KEJ5ZublQxgIjmfo+f/xVXTdTToCMir8+DZd7HMbefLrkDoD
j1SxJlzvcozwes2eu3QpzyRttFD36urhXlWVmwBnS9scT72kIhCp1MX1bYDq6N1j
y8DETH7L/DFXLNYho3X39PTe5Ls2J363kyQ7V+I4HgT4vluwdJD2Vp8tzMCISxuL
BKITB5uWmRIaY/fkFij/WAzsKpou+bsro23eTRqTsQ1qW3q73FSYaaft6UX6WsNa
Dui8isvOwDhdiL1C7fHMOjbedSSiVvnWosXwIEjwv0tG24XuvXMwScfXgrLcyALT
aSkG+YoC165lIHsTMTS/4DauqllBP1Y+KUmtzF6c0Ixyj0WOUwFvljdGTY9Joi1C
5Hyo2XDKw0xT/U3B3vB4Tc1xOqw4a4XXdd+fgVwKbNdyiFB1ftJrH/hrrwg4/a7O
E8iaC8Qt8dD48n1hJQjGdFUcVoa8d/TlD+yVx9OK4QGFUqQ1Qc+C1Hbjl4Hx0W34
BqbL1L8WR/TMQNctXALIvsHOEI+SD3901/AMqI7ugv+k6EgXtVf8cL6Gir3Zmppj
xOtm8kB7JSOvtRVEqkUVxYYoCPASzQbxhWuRzuBwOlWxxfqPc6jFg/xc6+nFTQK4
3IoDQQc5iG9G181Tr8db2doBWtbfDAJU9s8TuhHXMpsdVYt4OBYnCdhAQOTaBIfv
v6H9vmoZrQ2070QdmQUS7MamR2B6TqFaXRiSBZJ7ngm60z+dn8wkEO9H0uIBAi4q
UKi/CVr6ltVWEXcmuZX4pOxbADw2DenEVGaPwuitMUht07OD1iWaGYloN5b1Qi/6
FifS4yZHi9bq9kmVoUSBGDSDVikMf+VxAmSTktV+wVDWsNHSVCzdjfWjLrKpVaIr
/QHdhw12baX1jP1ZDX23lMMqs/rAjjbCVfZONj/lMWqloaG21iGMv6vj/6xMGeOn
cddgjbj+2Fr3GGBJKgmeRKWoGtv1ZysaEoeLsx33/cQWAG9Ay9aBPC1qjpl229qu
nJP3yiWQoClsVbqf1K+1bjOwaV3TfO38dWHRm+OOVhJITHraJ0TwXza9871mICMx
enRMX76Ez7tPXYUmckSvT9H74yDktoIzMwRP+r2PVWdNslL0mxZs1/kIUmi0Fv/X
Xr+KNm+F41iPEKRDMhNgOHqEjbgNtHQGFY/puafOi740E7Qj4huviyc6x0fR+mMN
4oJ1+r+cj4jWYfRSFJwWOo/jK7m/+fMlvirZjOCZnlXuULZo8hSDpUIsV/xM8shb
VnGGtZzeSwo7gRxMQRqvniuRAo61qBM885Ep4XhzVNir2BQWWX98f+c322euAJKJ
VjeH90ZCs3fdYUPoBisE0A0w/AdQHu4rrRitISs5lE9B2duypmCFg8MbWVZklTA+
wtYq3LMlZNtvu7EyYAqeMh9qoFyXerahhp1lfJ5oHQeDaEL1MQJdD+dCo0Rky/0H
2mbsc32pNVzTV3a+tDPBp94tWI/LWcQl8LZ5oXvXHJxNdfmqyh5W+/G8CaFMWqfF
wdvIfoU1WMEPnN8n6bN7wdLJzADBq88cgGupeGq8k0nmK2/mbLbqREvXJm365Z3R
bRExFRBW3BxuONvBiDT9K0K9Kifm0aGXtD9PwRsVSP5DL8xNOrFIR9qPi90iVFLO
giKc9Qv3fW9i5atWnWi7W24haGleUsO4VHWFBrhiVmPtlSgNpP8x2bm1DiTp7kvx
SWCJpG3b6RnR8HWR4LFhpzPhz/xLZ2Fut2W7jl+Ii0mJ9TeH3B1i18bDcaOQ+2Ts
+dHQuO/aGneB8w++ItvxvM1GZybOgU+WDhpQs98TXZcsVMhqafwbOgDIUVquW5yz
A7tPy8Ib9Y/e/sIirzBEhQHmq9iqpe9AXWPTLKukow8mw/kpii9ha3RCLBrTRNm4
1B8v2KDBasUHxD789u/mS6KHk6KvlAWfvz6+V/rX6mq2OSZ8ExUNB/XAedJNgOLO
rvQyrE17zLDzLYCSq8w2pVQKH1AiArewYdcfahIiZwlXLfNw3EhWpHYe3VKjIx/K
1YPSGdvmUn7/s3i6pcMNrVq8q/YfVIWIM3oNRJMQ2tlDIe3OyrHfug06GzxaCmq8
OW09IpEH1GwYnDusb8ANLHLutLbkxiwlx45MrZi68B3nik+01Tho+oxg0/eXBZmh
0BnLQOezCPwgEUIdo/kFO/a8gJpcUYa4bbcNlN2Knx8R8JiFAjVTKstbxsvmkmmd
5izurzoDCyzQEq/ZdFg3D5t6fQtbwWbKD4WdE9ajk7vqf4GUGUJfX+8e26+2sD79
Q/i9VzEekD8Fy4662dn9CFflNXUDQtcH2eAWhzBtryYZznQqM2dNzb96RE1L5rHu
vl9sJJil3zYfv3Kr2oc3vWIEYZfbYkn7sdWa03vhC30XymheYLS+ncsIR9SEf+8g
rdztdulNZfRCbCCnc3V4OwJ+dQ8+ItNwKIi1xEaNJfyHNyGA88PwJ1Oir8WlHRa1
XV0Km2hUgdC4/Kcqky21AtfTaqSbENfbTZOFQWsBBGuMZ6fQiwwLmWaGUq6BGljn
fbk0uVbEVARMUBY2n00smqXh0rq6MGnYSh3q534Kzf0vFGI3r67y76F74qtM4V0J
6tPMQDqRTWWRzDejCt6Y0DXFshJPAmKSeDaI2pejrNrFKe8zjHT0/MA7KlsIwBiV
UwKjrIjDKKYjyrzDZ4E5377KZb1/JRkHos8zDupHg6voidTZq3YbpXK3hmIqlwnH
y5j/ZBSunVAj2ffWWZmtX+uR6KDv1t8L6/4QJYNUBpDWmCOj5sSGCDs4fvD9K2Ao
kT0OOcXGbdmLcnc5t23h7C0PD0UM2d+UqR7AyQ8OR6OnGzWRPOQmTPEHL7/9qV1y
wfw+XGx5zOeb427BHf6GNV9bFEK/Mc0XkSQLcwNcz+vf1T9oJKt5VG6d6fonfLES
yVITifE17y0/NHGagY7GAvGvf1GwIu72Xnbh59gW1PAI6BRy4DcEgT1vOv8Na40m
nT9GasDSR+vlcANg02vSqM0aQHLrL76bzmIYpHmwlmNZ9Ya6T/yPB97SKil/RNMP
T4C0MCLr90+Q9GRVWrceMbQS9YlTtuwxn/PA9lnLETWqDQgT3QJx/M6WtB+7rO45
L/anLEjT0jkeO0GnqsYdJ2WbJROCuD+uOiB8KgQGJv9bYjS3S5wnEWPrldtCpkvM
8o/epH7Aqy64GuC9f9/0jTVtnvxao7INRE2Zqx4rhkJxiymwj4XN96xt21fiPuVA
fxvqZvt4km5XBSqAvp9G2bmb/cjB+OY/oexosRcn6UlOQ9nDl658fuEqs1O9PNWa
FKITVeqZAi0wSFftQd8ib4MpaqbNbNglGpfwTsUW82vdJ2WY6oPpQXj7AWUNmELP
+jqssuY4hyjfE2KqIV7d3o2qGxZYmsA3RhSSPfKr80x59PclIVqdY/zk7rkhgISx
+/6OnF0Do0F6imyRS34nC2gy2o6aT0GmIH35vbgcVZ42j/rtJQL5c2oGIpz5WJE6
So2N8TT60M13XVVHsaET6FYYdE9wgl4wkhsVenxHnEnoLSlU30nw/YeYTKNRj57R
lQa9UnvibD3jiq44IrVVQYNLIplwcqi6heakGx6fNH2FGyHL069xK8RHSBvWFp72
VVjoQvRRrrCi3cYdyEcZw66oMfdJdbzAl2cxcFf65839iN6V6Ih7nMwES9GXEGcq
i7qUjYOS7GVdTugToBax2pcvSf7iGuimhw3duNgIYTyl0eUlFFl//LD1H+/Zh2xf
yi4vH3JpI79qOKnnFG/xADEuwIpiRIebgcBP5cntUWTpiGXyPYv17CiohSR6Hvma
wJPyqg7h+y+7TVzLXiVmiI9qB4OGRSWDlnKRAdjIodHRrXW91u7+vCGA1f5zqDJD
jZaxPpjgwBGW4Zx5TfOombDQl7C3b4DFNwgNJzNCrVNpEiM+BUrbSwzpQT/qBAa1
GthkZEEaY0hdZgWzaH9EuBNeF2L5Byg+LEB/0Q6tJy4YhSaaAUOu1x9tBo2SDyCc
Nk34k5H9JKv8SRD7p3ztUvwC0H8MoVt3RtLTLyMguPzVOrnEyqwXj/c8Vn/yjoQP
0NU7zJm9A69pr+MBoRG2bi2i9mzvIyix5ajNr5CM7T49AUTrD6yVrHb9TnQuhE4k
vfJQG+VQNr0QpT4heWapYfsdxbK4kcQQnebmA79Mfs2xD9P1ETZV8gpH5R6E9UIg
8TZYRsjsvBkzohvOz3CNYGeSM84oQ3VeWPFu/D/hdmrfNxYLNtoxLkFOFKE/YPul
Fx1To5q6U8k861q0MAdJ3oOwlPo45GnbDyUCKQCWZpnJ4TAp4ACwOeA7DsNNG2Iq
tdybQXtd7usFAC36nmGGXcoPYxuBJXPocg0TTBJIM2M4e1MHGZ2unenIruihu/M4
TcXWGLE/pskQ3LcaQEyGf36Ks8GDayIOBtRbfxA8PeCb0oefo7+WuViCnQWx4WQJ
rbpofGUINvRUQomRPf6JwKSKqZ20mEFxNZ1WtdNzZyVBdcl+2rodUJ3MUXNVBklI
9pf5SOfOLkPhH89xHPqxOhYOIZynF19+WEN9uiXZtV2fgVD5Xjbk9aYQsMyQ+UOD
EswLxieegKYgcTgP7+Yq85yk8lQ/HiaCDTecTRjfGvIHXz+y2mDKpGH54XHMm9U2
ss6lCZjl4CSXSYnDc079aKZnoXAyyqKn6XnhFAyENS0QJJnY7zvYOL+rr03mgzaB
DnPm8ag7FpGRtP44V1Gr0ZPqib7PzUQikscLGNhzlG2cUyH43+1hKGS4y5xP1E/J
WRLoy1CkNyn4reW5jy/mfVyo5Isdy8LXHZ2kJDBHAiQI126F0E6F+Vg1NUJm59So
LPxeA3yFHWrbxY9VPHHj2o5MVKLcC+SaTKbR9gyzhaGIlmRd+shiFXrvhSlvZalV
nW7mJuBtihymArPzD7/f+I3gh/6jPQmUbmk2OZ2/LKwSBm5OHZbT6V8tMq7tGH36
IQ986rr85YbIzq8ucGD+IlVWZB5LBxbHJcGGZDg8lssoaKkGJ3xehRizP2ln3O46
RR1avgX+DPcT84BmS5sjCRaFo1sL783G1URz1U4eEhO+DiAZsci6YVcHzi9Y89p2
N4c/7jaO77e8p1EPWtIP6tzOHZtLMjrcjkPA13xFAOjrVgcrgCwvI33a9EooM16d
F20zKDg91q07xcqDNPbC1hz8Afwzs8hKZ2nFbCjAcGgg4aTHIRqcHAc2i99VluYa
/dNB9GhzVV69irLusfQxvwa2tUCA+3r/9dq0BqCV4HIYOfvZ2ZRuxL4LBTQeuqPI
xlrJWCOyrPEjXxzy57qIWoB3Yzwv/CDetMwQaxe8s/jLLc37Ij676VKKTJmHEFLJ
mLSTZshdqVUb8UoB5NzxuKkJkngWNt9jBmkqtLJcqXfoJLo4A2T5rVeCFCxyaKcB
aM0ksMOgZOJP/ZKTBmmBVypYOHUmQoM3O5Xbb66QOIICJ8aOv8VU6l7PFx2XGYQj
eZ2hDY2XFEVeQCxskkPHpBJdKqTpePiu77YuQ7kjhHeAHCGSFXB+JZVYCx+UzGa/
Cbq+PagKpZ4quFXWLJIBnw98hXe5fWW+9AtcZ8vegZbsh6r3mnH7i5v5Lkao3eCf
3326795VuXKz32J9NiEilOgZwyEQjLlHENYQViQFUnMOlyxWWlMG7Rj0197eSB54
RorlitwtXTgkVx4eywS9q8An01a2xovGsJv5vygLymRlbOr0noVQiJ+wKQGLSRSh
8kemVAURrZ7H8k2hBhTY5nLhH6zP+4sqyu4aeHMUUzSwxzf9EKXE0RL9TKrkTQlK
XWj/8UKWa50/tL1UD/UTWLMgDoQ2umhnKxd0PXr5d9ixbQRvE698ROuKdJJYe98+
mnL/76RJTm46YrhPE55I4XDIchk1GQ9nOz5ux9Zx+gHfGpRnseX1yIR3RfUYGCdD
R2tBBJafMtSPXU+8qDwIoRC8hHYREcBHKE3oX6J28o+iW/9utZhTUrNSw90nPrm0
pen75euBu1CnRQcPHAvX18x7csYcMSQSdbG3CSZicqxQvOOF4doLPMI3TvGSSEHE
Zlj14QlxohKYs826V/6Pt7yufhFqI5s/GDfL1IHeCDuTidPs7RzuOsZQei74D3Tf
7SNJt9B2fATEiPznb9ECHP2yLhgBo2vRrHisYuYFPomafmk3+0Ix1X3s2Xbsug1o
SlNrpLI9nYBIlBw9oAOtd0BKtZ2h1MIFEUP8Gbq6tJvK1P2IoXinVS4mRLrpis4/
H6VkEbBTiIGbY4fi/xNZjGsy/gsr15D1n505hJOhmf5x93NGvIRX5qzF+FxMo0Px
hj9BRdwaK0O+UPq3Z9XDjX2SV+SyBsfcAQcJ34oENxkFz4jR+N8MyfoymK8xCmXY
oYxa+fbfy9YTd1ogIviNVsmCc2C0EDIO6+ZZJQ2U4+Dr3j4avWuMGsWUBnh4IT6s
fZhiipiH3ekN+vZVTOP8JpQii3TCNDCv+1AYgPFIO2U6lO+6yfzC9t+RD78E7Wad
ufgd6tX7c4bnpn0q3zOiI6PF3LIQViEkWSqmJBbErMRBN82c7wMH1CDBHtP0Oo1/
jLuMp5/c26hFDRjdrYrGatSs0Ovi4MYmCAVvs8ISxRNv+g/n1C7fUG6tkVMfcWyy
kXzkEJA3HXR3Zs/WPBMrEVTGx2qdEWhlDbCzn/UGWQ7m9+sovrxvoQJsbIfNBDmq
h0ASpx0NdObdAEr7/QrFEMTLtSmO71l0yT8N43i1ATCV9NxEdFmmw34f0aIPHA1h
khNLiX50vfxUNCQ5F0kkHxjWM/7QUkwO9/iA6AFLstfW2K3unuNqpG+0s4jvv6e7
f+PNccufVwH1YsI61iEQ95fdJvcJDugBGpTQ9mZNBNbs2hm/SwGC3qs1fKFbGGDD
Rc8qc6dJ/DSNzcCtybO+xwpwiEbFBIHQT/KiPBPk/zvswUpfZniFKTWldIonw3hN
E1cH50rpK3p2XB4/swzpdhTidP4VvHU6myDFx25vqimbmduERXb25paus2h0ARwS
F21+FFrS3cOu9hgchK/aWUdByERFt84nF8Kb/iYmUBFQLOjKzsrQw/o1aEK1qHjV
TIYjjH47EYYfoHFHLPSC9zwNyb/SbrVwvqK0gf5yGFu76xf6QqYGb57s+XKNae3w
5f2/EtCXjSABsBeJ5y3m0TTycg2W55AYS0u+M1r0jk7AmM9TnGhe9s4lK7xximRp
SF/C9/Qg33DxP4fUCrNYyj5K/5EXdKgcWoLu4oBkiu2OsKAJC9HH6T5Ta+OM4TQZ
Peu6xbiJnb63evLhzMvLkTcf/iiSOzpApygzcSHNozSlyXS8P9efpSgiOKqRslpm
VbTh+Nc9H1LvUQMjJDqbF07m99Fm0NYna/RZ5EkGCo1G3C9Q3vjGcZqkbH27GfrL
DsSkDcH+wUCq5HXE3eYU0i3CJw1T6eFrY3FlHuI808PRUERr6mQuAWy1K4FcJcpp
YfPfgVvcwaFphQAnGy9oS8CjIvv+zFNtB3a+0QFf9iLnM+PfJ703X8Ugit6U67cy
gIHrju0Mj2D5puBj4D5t25z/29KfGyFBcNud2/b1P5b2njrKIIZRplRAfqG283yv
tB5emPj1rTH2tXRnwg/WsH7PlZqMIPqFdnqXyvery3ESxsDsvnFBrrAXLQU+mjUi
JQgsA1+LnY14zvuji6tJDN5itUIKSd/69VLUy5AItPEtZUTtcxJya6fNG9RMR7Wy
jEzUUmrilxg9eCJG2lakk81UI733LfOwGdiFobYL6kJWmcdn5G6Tizfn4V4ECQa2
mDr80UFVSVzX4TWbqBIuI1w78Xk9ixXC34VOcLmdQjSLbI8wDLLl4TBNQdGa9dUb
4d8I9yy+wMUOBC6f18KvKaTDoPeDmrSjvBiT+KiDUO6PjvYOY4BbOeXSE2S2qnpp
rpxBUzS9Ba6xtyNVihqwXK5bCP6deOMcbnG3n3Iy6S0za8K/25QSAYiGOnb0I3aw
Z6H8xnPqnE1HtGG+E5/COrqKXXfG9VJB1bpVFV6WC1dFKSf7UHngZ2QxD1m3KpnG
2ZpUSdkenueU65lB0StjTZl0TaqgeqNBqBoUoAj5Q+OrHYQ6nVo6idniqvio7DMZ
65dvHW95wLNq7dcDSjQQ0OgjttfIFLfguDba7SjVvAox9sugOrcHn1Pz5NyGXNFU
EitMhhcqFqJYYRQRAF0qdTO9ET6R3fLnkWKBHMaXBaOk8FE5cxAi3mNMl7fnybcR
qHZ9vVtm1iODPG+k5kTIiNCSS+2MI+xANHboHN7b2hVTCp4JNmsqsK32wJazYR2j
s+opVSaUeJCrsEtstE09A4QLznz1FIPW3/LhI0HoeRM3cG0T8ivwups5Ejc/GTh5
PHaXabLQcrsvVWedCKJW+8BvDeDjY55EiEvL4Faojns9AX4kRmGLT1dt94L5D7tZ
krWFmtxPfDh1p9Xno0MDe6MIV25Zfg0yoxZOb3tXm3CvtmiYVCX9CDljaBFzhulB
SrsG32einex7OrVIJZt2Lv6lcojd2drfBcRfyxPl0irP6FTLz2cLQknOH2vGbLRx
0muhsQl/regpC4oW4ctVazOQJ5qpG/XAQDYQAqw+63wBQeU91Rd65dcsKgAjwYaq
Fh8D9Cv52MoHY5dmaBoOAcnH7rLFntl8ekPakbKTqRX9McOmHQiLiJ5Nlvq4br6t
tcv8e1EbMNd9DNUnhB5gsVtR5kC7T09DVr6qlKDDmRrzHuwm22EUFL91D6NnKQ0N
U+m/Abc+4/5dvupTwNgaTv7ZonW52rhVl4yidjxRnK4fkVgEje90BmUDB4wjD2Wb
trzn/yuMnY9FnGpv/Qg7HApzqdhUrR4xzX6RgG6mA14XR3biEv2L07S4QKixkBsg
dddQS6bsLZUTwhpxbp2wUKzYBvNfcug4UTw+/YnkHDYUkI8YfHBN7Aa3SIwPLkRi
cSoH62QnPNSjn0E/QINvqKdK2bEmzlnKrZ0UtqWLaflM3xeu+bzpVMYTkHJk4v56
Jy25DKFZvIcFpe0deH10rFPyGCqVM9dyqbIE+NrY6yzSC5ZAa4Mv94dgP2Yztcv0
+xYlXxlBOjU/bLB7YZ/EWMy9RdIwRMGtUCcaQQyZuUmtUSxX9nUl+5yHDnyOa8Ew
AgIf+kaAIqjggCAjW7uWJ7FGNrc9DR2diPnEuTLkxNfgUBAflTa6B8oUoQNPayNK
yKQzT35NhhSQTfR898odh4+tpYpp0lDqP/PpFnVhBOuKfgByzFAPKRKjEyp1AZPe
SIr1e5XmuzMjrlwnvWt5Ubvqolbu7N8cdcMGPFJTf/CzfJoG1D2n7Wk8yG7vdT54
BPi7Xh0FgBeyTao/TZG2TrJGZtp0QDxMH05tixiQyrqgHhXp2akZMoAtfUGZW3B6
WABA9zFfqvY81P9y0VHLAR1rVqC9ViuUpSCQCgX2dQoMe2Ex0Kl2V3gFkVs9E2mQ
i1p7Hn4Sg1ls/aWo594oy7rxsjNQIB2e1D/17Uzs6C6xbbMfPZwXCMgZKnWYiobQ
eKUovjz2FGHYB89dVDMMpMV5z1Buh9eJq6kBf0Ko8hYEWGDe670XhWR4vu2VxkcL
+XK9jId9gUZ1IbZaLxHOSqUb23t+2XW6k0wSSuzKVR1Td5Qf+X/yUZe7s+OQZEbx
w/qnZ2a7tiSuay9rGjH+eet2FlejdGihCwf5RX8TfY0Q2G1loC8iMMJF65gDaTGn
ngf8QBG2+6VTzN6acAeuDzyxUIqWJ/iBwl5wuu5jmMjscQcrJtqQQ2+kVyKFPEtr
ai1U3O/LZ6ommTGqnAlARVwp0MHMo88NcFNYdFg9ECJ/5LIfEi8HrAmuFIR5qlNR
8ympg0q4pgEeiAj2WLLm/Iul5Xu2+613vpwvm28ytdHcUCn6cTjlQkGtzCWDqCt3
ayEPp6DqWVTciz9FUEmXDzgGpqdPPCts4VxWPTl4Z/1h4rThiRjFdDOoIltb+tX0
mybaY1a18Sc90aCKr7vTdKunNnfJc4QghP1bzGFjgXjd8lnehcokphwlpQqSA6Dr
aHQfMkLWJg3UbWD8vMcmZiCZvJv9JUngAtKXEeay/YHn8xt/mIt29A1cZemIJ84h
bfrsAsgW1GDeZH9Lj75ydlyIp/zR1VhgKDrGh71ij86cdxPX4y+oO187fEyfkRrw
Bnb6xoHhjwZy6M0QrF2vtd9CAWPwNPpYgsOwv16K96f7FHOK2957Us41YJj+iv2M
fR/uPN7C0fXuVpgRXxHGtUjg+oFq4BF08YfIpxjId1xlhzW+7KZZH+SY6wJs5F6o
v4302TH/bUkbfAYM7/Myegg6FjS56mwFene4vIooiczY3v8R9ec6fV+5v286SjiW
llkKvqiKM9N1fZVbVCK82z8LdkCZ5ExEAD3UDyqWiCGoFzKsUiGrAUEBCHEGvFIA
jy0TBZtu8TP7uPw8QA9E3lDo+sJXwu0fNiekLHvxFgNf8jPfkX2sJHj1WLZAmTse
EfF9kQM00PQl5PdPpRqEPlgDhPh3fdiN3lg9prNtX6cLGHOSX4k2iSgxatP18uTY
ObfsT24RZzBobh0/mCvmeByqovuDTDCgsKvKr7H8WzvCBktduOEYuAtZiOqdXqDe
gxQ+Es2kzqzhZAJHNDV0vgnJY/SYpwkU1vDppbmaijlRi6m/sRuR+hXlY/FWrUSv
2BrZDw61hNNtHQv9TYP2loFI89482bBm+kmtgTXgvZEWDagURLjJN1//B573xbfH
81OAO4p0MRCt4BcsdxRAXYDXuar53S0ZqcgcscmhJOWW8oAHF4TfIFzw0UZM0Uwm
w1LhSJRIVBSg5BrpG0rXeOvcU11NdvGqCS1TayGMoTbZbFGiOC2ZjStpKxJrOZIY
FOBgjx7qzvGqWmUv8BrbL/2LPIse9UNMv7TTXw/LR566pU0w3LZojyFZK5/de7tX
zdTzsiyi727UdJ+l93GkGiL/CATcZ91BTcwjwf8F5J1JOWGHKDDtJ+KBWQuKTmRp
SSFZw9sOz1DEGUDimIgceo+lrD7CnYkL8Po9bSRTN31tjZyklFfl96xhC6Jim5W6
PjoVNEO28X+otU8OaDlI1qZmarxoQQ/+xODKS0G0pIL6KVbdsNHycxar810oNOpZ
JHTK4D9Y0DnwBWxIX9+3r9BqKfYqzW34Cynjzh7OJrfjR5UWchiq56ErotQd4Vd8
/TkqFZokNYylRSln8ok5yOZkX7/4Wv8RiXaLix+hFT8DIcOdiUxEi8+KVuM5mZ5m
/YhPOzSL8ZSxs5g/K8S0IzgIVUPt6uF49pKyTGXVaHejc2bePHMS/tGO/1+DFsd5
bQwPNbiPBqERCnPS+5BPyyjLTClYi+8zxBkCC60ZNsED8ZT2YZpfyOcdRn24vY16
JH3He4P3uQsyFyFBOWHccsLopcJUeTwUOlGxTHA3H6xeZfnXDapiAuRdjS/ynHRf
1ZHL11t1xvVQz/tRkdLzlT/mC+KO2+KxKDHoCMseawVNyiSE/vNeSlJyOKEM6vZD
SxQhNEdahk4iUkLsH4e+X0vIFB63AcbCj68eL7bNd/o1O5+HQ9FWHE3iGI9SVuYA
mqiOSyVwdn1CsYYNAibpcV72Y4VAFfmd/nbgBhtd1X5mc0JrmP1FqfYx/5yKuMRq
J4MRvMHeooSjvmTZeCOOvpGGD7k36lMDRJvlJFEJAU8FQjRob39BtcXQttqm9bLE
7J4I1BUkY6FDXe83POc6TEtk+Tc8+LY8DqvNE4j05mUEcc7N/DdxYG4tO2OtCVoh
SyG/3GWFaf5C4M3moM0q/cSK4idCkXn8VrGLd6g91eA3QzVr2sj2bGRgNQj4ecKP
cxeOLpkX6BBY4PIV1ePaz+YsGaxmIhwdfHvLaCFSj16PZF4zscj3Umv0TOcuqM+f
I1KxBcV699TwPN8xRDlUzlK+ZO03EDYqu11d0m8vY2QrXcBOQataWkNXavlk/HoH
C6709JdldfJ/x9mbkDZaqn9UoZagr/BmuzxV7BrcMrjr0dbq5DQByI8sMMCHeJZf
EkXwUL/hyUimbUA4K9APyz7X7pmMpQu/QLPYf0xQO4DJFXc6rPFi5VmgfKn/eC3u
BRZmKEWfCk1Bo2eyf5RKjMjqj/kGwFOSrgI6n7JlgjPOhKLIryM3y3+QY4zPBqXp
mx3Flk9e9vdQFMUQEC3SBuVMbQweWMGT1rQ8BVjcfPUD3GUCSmYN2N7XNO3OQB/t
8gDBOsjimB5eXbJiyHxN3aSkVHNLtQGw5bzLMpcvujdgb3R/1Mfp6VKRqU1IN2YX
XUMws5FyWMWiFxGVXcOHTT4wIT59WRvKXw5TzhMALV5GUf3qGdin3hbm8e1rFiIs
WxwHp9rB8mUsDST03/C/scRY4GQg7gknfDTC0Wcxy1ZuGQPm5ltqPywAd9xUGM3p
tCR3cXwAkG8wmsvKTSlAIa26KAbIBBaABRHAThQruou7CAeUpc6g2Itgu0iA3F5D
rcgRgylHu7cN+IcynIimj1X7QVBui/wtgYqoAVItdEZLYVVxY4EQa+EzOK9jBtBJ
93UyGVkLBdnwY88ILy3yAjkWs1W3HKaFEI2sLkpB5aQzmv97kG/aFuo754IkkDIS
06ZY6o1cj7mx/nbx6Fig70mFkqdaSJ+c/KcUg0pmGeT6u0GPfYVap80Ly9UQ536w
MS+2vtEZ4hmMy6N5G5Xr3PnBrkknWwRUbi6xcRPh0yHxIZJs8Cjfv3cpr+S9E2tO
tJcocNEmmhjlQ1MduqiRNxDwDLKYBNimQzqeiHpChJ3Pnb8+7qqB775FwKaPCfuB
1JVQapJW4mo8BbwKOMQPM5oV7cUOQB2hYzSuyaMt9iBxnITMmuN1CKj+Sx0G5ZcI
udhA69lxmAHZb5wzIiSSWg3cQTHQSPV5p26tw3pUuP0tCVuiJn8BH9MQRwnOE0jb
NY9rUZdvrEmHCVDR/Y04ewjMhAHTrX75ptEJFX9SBf21DJ/a419QA9QcZE3DXJEn
mP1Gn9gHubKQ+QBqyeLiy7zW5NWff+Occj10Iu1pSyhA7DUGs+i6DgkJroQAilhk
qNiEUfJKPjXnTcPeTdGnR220MuTZUna07ees/aZtDU2Dl2V7kGh/Gqd/Q/CY0gjG
uk8brDb+TWWVDtubkeS7k7ad6HP47wSgys3kj4avJl5pIp1i1N0ESUyLT4knnJYR
BBSrgG9b1wI0as5neVoAgZpzuv+f1KGAHEc1Sbh+Y9s1FRk0VPo+2Y5M+ts0OU/5
cxTq6yQEGnKLxX5JqARyaWUMTXAmabk0+JpAUkn8vCnTE1cSxS1ETCewlI6BmXCv
fe5iPbsF6oW+TK1wVNu+uEbCoOmI09Cg58REhkJtkH8meQ0USE7eKtYc94eg8w1I
bRW/3PXhGmQl2OlVIRlmQprfIdZw8HaX6rsyalp2k+bcPSs0Gqdoa2Vt8w5wEcW7
M0EzMBwXExgmc7LRzHT+VSS0pjT7JZOgsY+BKJGxRO3/kumxn06nhu2LiUcJw0gS
EdE5o4VOLZpvhlyE82GImmaTL/cB2htf/TMn8MGRE01QRCCEMvagQBu5dPBUXu8D
gw89AMxmKMdU34G6tHaZ+tOaxFByDNwAub7hnI6aogX+ZPOaa4ilzER/Ofo9WvJF
magntkwtMsQuP3C4vMcZe9/DvMy1gGLLn6gsKc4uXT0p1fSv0HJ56lMUCM5MMzph
YBUkB7hAr3giwwsQmH1J7264syKiBgHFiODUm9sDMpLdsnL3qGd5a8gQO1bJR1Xp
5NmWbLlOW594YFDjLJFRXY/WR/8KCZE88gXy0eWqXpqehjAYtlfgy4kUC6fPtbZT
7inlPD48e47dMbfmCfmRTDXfi5bhKeQ0OzFTT+A/v8wDHnVfd6EWvnz+xSabNteU
DGHp1C2t85RPNyVvldc2nO6xFLRfaUHF4Ba0EK5G5Ja9uXX9VMim1txvG7hwbEM/
7x3p/M96k+weGfXYFKfTqcp3ly77jGmRkA7/ICwx7OKpFKYRUidTNwHJoMUzJY0g
8z5I0r2ZP/64FfcFz4I8AVMsvBzgUiyRkFeon8q069PoQjRX53rnCCSUfaoNJdd7
+Mzq98Cz+taJ6g0T3LvGo6UM8uhytShFte4hitvp2B8IN4briPiFOTBv6KHq2gGL
WQLOsrvnuTEVs8ZNN1/qgul+hlEk5dz6ARq39hrle0sKc6OVhOMofxcALPffKO24
DW+Z1JqMctru6Ia0kmwCcxTDsCUNVjD2eBCaBBXgk8swKJO5YvYtp+54TOE15Umm
t02ZJ5SMupOj5yo4M0oitGM9aP2yNCnw4NvwA3wdTqv/QuHQjFO10Aep3SbmXWhw
3cssXvrs3kWkImNBifAJ025rrlCg4jToQXwMFyr8mPBltNHHGDLRjHQI4sbHCQTp
ZXSM17NNRZx+j/NPPq36/MKgCoieyIPAZA6FOgbavPKqMUgpEuZlAkOvBkFf43ue
4yybYQI2qKk+Q6QygyDX5NpRlSmtQBv/iFyswJMKkkKFcPDqjKMY+ZdXycOqvmsZ
TNsJcxOJl2/xLVejmquOhq7UaTnWj9eeN2UMk74VhTGdJGI2qttGhycQ0Tdh54IS
5rK0CJMUFMQpb7I7h/KaeszKNLrdbYbA9+FG+nnn8GPtgdZ1YCxp9n1gW66nYq/5
Wfh+f3FiN/d+XiR720nUQpiWqfxI1DgMR23ALz9zp10h+Vy+a0O1cGh4rroC6ePZ
2dC6Bca1KgS7so6zkwEZVfrOG0N+TwLpgPo/Dxjv7aPdA/1hscWK+7P7eb/8Q4fj
clW3oMMZrouRDKenIjzVDBCYzl4oTAeuGNdpne1+j2CABT9a2P51iz4JonjbSEqc
7GwrDMkp4uj/KucTVk2HO7Rzn1PXWPGB3YIEArWhwV2IqIZ5aPvCzsMV7R3Hqwje
wNN9tYcDV3PC7MzF1ZEnGbwJddSKluUaW7HluqxCDDksswVUjXSnz6TCC7LYYyDM
Y2QpmyeRO0QkD5x76bR/C2eM14M9YjKEi04HsZqQo1vg+7JBB41wGSTYRjgqLkyz
d2hbEUQ58b5wRimm7bw4q4Mm0xZHiI4Gaf9C+2V4mtSkJj6RhntkXuPfUB5Pp3cO
k0oFff2BDcOQJ57+3MtIJ8DteYq7+NfhdGFWhoCRAENnllDYc4kNmnIM4NtDxeso
Ke/MtSTGG6VCnWogPt5d3ENzhi9dPBWVojKJVn0WSZxtbi8UiwbJbKFVJwRqmGdt
xFGfQVmLQ+PyG0AsSd118TtN9NaXa0E7c1HX4/r27jKTygruhe5pe/xBQDcQDM5Y
laY6in54MLXznR5cvn7rU9zRERQfYSxGAdWUKAL6oVUBMW2MspAAgh6+BElpQB3v
XVgJ3wccQHH9HiPWK27/TebkoaW8g+9drmJPIMotv5xzWd9jmj1WV+b5DGXYGjPf
yj83+NDcFKS+pyxd4KR56mAELtcKJZ2/eMaHxZbT+uow19Prn4zAcA3wIC+x4z8u
G93QLPml0Y1M0kqm9plIP+jKAsd/1XqV8wJvZx3oAYgNUJeVPkkmyzaOQ2hXvgKY
XyirhHXxwfz+UxGbdJeOZWNaJI2FVrZYLp0ZJ7xzSYXGyqJ7uVYkXJsi2m12p2KZ
BI9AZR6P9RCCa1FnAyBAjydiSEfkfo3i587aRTmDnFnnZKCi/ros2hhowZqj6kqB
AHI7ICCeJZK8ewyiDKc0FxGE2BkS+ak+KnLLG7v/CebGTE4Bv1VWpx5IrFAvHWnJ
iRoRxjfIze1aHKI/YFIhIAoQHfzfXuIvi6dzrvkWSIXc2aphTroncJpkPVF5divL
R4OodziOJmq/7qax9jlQ5pjABKgZhOQB42R5mi2M5dqncMy5I2GZFg7dvSXaI208
vzqQIHodxX+ZcBA6eh47E9Xy8U5nlzqXmSQ4cadV0pz9RV8w6HnqJavi2D0D9mqu
Sy0aT7ebQh6ATr2ix8YDDnT1EsQcm1BBY6tntBWD2YWb/XPwav6JEP3pQ3YLQJZD
ZH+sxCH8y4eCu1oRKAjH9WPMW5wBk/YJCiANXmX0P6e7I66uauP68EtMc2xJH3r3
thcpRjjtc7cFlo+oz/CEoAHo6ginMB3tiqVOUx1WC48DXAvaJPVvGjRjslfCT0TM
ZTjGUEDVt/wpsaECAQJe7UsoAuQhaid5zS87dAb/PVO78PqEXeun9K+vc5WZrYzF
078ws8Mq3Csc2fHDqZresRPgiM6I/ZXj8HMFPPf/jIUoyqGK9ub/grD5TWNWnqYd
4rHQp7tqocBKfUOtgnHJDP3hBfXGTb438uGrsHBZwetqiy+jfFhEYYhifTScgelC
oedfRREON6uX3DrHGrL9EbPmvfgdhGyNRq2rX+4hRa3jeQZnQWlzIhN9YoO1CtJO
fVuJC4iXVQDtYC0IrSMlBwZllGWksRrDkS2UlxPzf7EvO0bvsuCVjo0IyjwXJa3j
lf9zeXggEQ0qGia7H19CB5AXSX0BqTTvrh7M+Yc9dSSb6p8RjD4Sj8mppkGIzo+L
/L/FPArZWkDG58izMkj0vIAqAAEcXV9bi3xA6mK4BurNKt+mKwK0Bahc/dFaEHqB
wr2M/RPwMj/L4KQcicxdqwW0jbiyGyvjxXVnosItx4ZJpC/npqh81uSUYvHAdh14
24Qn1uBV0DhBIGm4Bf4ziNBi5tWTPyqtyKfuXiQMZPW8bJxBeN0HF/8oZ868DKoX
3NNRCqf4dMNc1UsYo+WD/RZ8ou2+HBcHvZxCydtTP9H9GkUXXULPV9OpmB9dGnvi
b2aoUr24Ku4IocHEYJqdwtpYDX1UW0DSWxj8csDqFlak0zsKxCcv/i6lThTCSDxH
Dxa1hFVTzYppqOR6iD23IPowsNqJRnYW7/PPhogq7bo1FG1z9Guj8+3rLKQ2Tugm
UufK9J7aEF/HJwNH22Hh1pb4Vm6j9y6I5oZK+SYhuIe5lf8lOAYXgI4adzmDuTM0
re7fmtqVYcZIpv7gAZUsBLwiFuNnKvOV1L2yN6SQVsxeSWOFM3nNsWFq4LSSMXLY
49pWfiMmQtEFC1aTW/A8pPubygc++Q/QxFoZYYXQkLlHRPDJCQOD4Og4piThZ7f8
OCTGs2FUcurOA0eBnkrKgotHutiLOvjVecOC32SGXXNVoWWJWq4qDmTiGiAbIHHu
P4IUFhvWe4xPH2KZ65v1mWoRXv6+tQHmEWnn/5+vGCkcQno6HfApmeH6/sQiaW4l
/LbD3fdfIp6fDEAXdx6lL7W8CuSuGY5DVWfzhmp9ByoRcgr/DR2xvAbec+A1Ua2o
3ba8R11/AuatjS7b+Mt40qp/A2jHUk60hZ2uzmJQ/BbNVTxdWtARmncn/xnJmf2B
GvBXZXf5zMg1hRFZtnB1cB9tWDbkyTUyl8r87c8xBnW8lZuRuLcJMCdPKHeXXgKS
ajE13fARO8WKyojJ8R8657Ra6IZ3zA+cvLWqxzck0Uq7QzJ/GGV9CWVtU9SZCRz+
FxaZmlRyicXJw8B2iQ81mIbz1cB7JbU4mPlz8I1eeha+EfcWkWjZlp02Hgci79hC
WIF8Nq75nKK0Ii7YvcEaf2M0Ew9osLKdi1a1wpN9CeCXZ7RNFqDosi8vtzM3HPqw
GbHKPIUCUcsopl82ymf0a9PHCmoCP6znubrVYspdbc3TFrpJbu+vVyKmlNdm2ZeF
yX3ghTU4f7VhZaVC9R6NpTGao6oOUk8ufUzPm/s+OC8ieu6NF8rCl8BbsjBg7rJj
8FTy3aNqE4ePqKds6G28/XPrd9JkzMCY+pHLpYV8j37HHu/cjtydXcbfOo88b9Hf
VsWY5qEc4VYQq9VPktl6ubSEBHvPVxAas+JXTnsImkcMsW4zixu8QwniRFFCc6sr
0AxY06zDNqZNFhA/34RCd4E4ogvUU0BObDJPKFWQSOLpfZFRGcLdL9iQLDZsiWmi
oWvbB6WNIMZ7uEZA8+Kkq308tRkr3/qxeTmu38vx68O9ubc583gY32doCZ6EDp6Y
EEhMNbqMW8X0hbTNFvf5+13x0q9ANhTjUBkybZthVciYhVK6VRnd2kjEWS51mKJ4
hG40BYTfbVJuPbst4UxUVo6J+JMrbAxipR3k7a70viTbmJ/zvqOJ8lZ7TTgk4QcI
bQ0sBD2wsLkjFuFSvOY5q3z0W2r/8ltPpALTHxU/8g+etiFgnhOyaicMlLqeaumL
pN74Hd5BhhkSKiPcR1+eefMga+vN0F3d0VBuEoUvK6+f1mxDmirgcURsWwN2s1FS
szYQLigotfBluLgWFkDKz+jJQAMJ2u4DFd7ovA3S8WekU3DdwF+wCCOIOSHVnLRl
hs9a0LP6SE19b75OBkO1bH+kQN1wrmANNJ4XMBlmYnSs1i71rhyVi63VHRyrA/zl
+DEf1iMj/n8C/IyoGzGd+ZeDbpEWh5Mv2Rx6NCMH96IR2vZ0Mw1tRZbE4Di6buui
2aEpowXwqv/PDGW8r0mD2Eq4y5a45G7wua+E7yI0EOo+vwMV+QDu/Y8pqMGdT/dQ
o8PGoVNQ87shIQdrZ7X90GyuX8T9NEzdcUUjT8bQnSN8LNm0erOww8DWVLgJc4Xe
FF0+elz+wuw0JO+Yvpa1LcIGfFqB7vDoDme25L6gEPNOIV/Awxqmvrz03O58GZJD
xMeQ3jL5WriJNIHk6vglHbEGVfZeQ9oS7mLfZVaUmYlXy8oBIS5FnihGQvh0io9E
1jWFrmzDZ76oXLyyZiImu/6R73DbtgMPJk1Kbwbsg1Djjyf7PYg1+UqlH96m4xj7
dysvRCMoVsemwi6ECEbJKpZqB9jPij4O4RKJvrVLm/s7E7j6NY3ZxvvBCj/FrFCi
r1i45qH25SndTH1oVEoeYpR23UECgXOKK3kaY8+fGpfM0ho+PPG1XkNH3DHAkSSh
+TolAfgC4R+A/+csLfaC+sHTsMNgoSISF1gHqL8M2VBOgwkSE6X1zRLNa+zd2sv+
LTteKx6mCXdQzkIM5PMc61Fd91KQjsN9jx7Ome6kOofU9/tlQaJQYKXFVgTofv0E
0Dv0VLFrusR00gZ53flaResh9lq7xWxTo4xErsyYy7UqZdJdL6zNH+8M1/sYI9kf
Hqe9v04ObLrn7paWm3LxIjSkkx/s2otRbrP4SgX0NmJgrXoZzKaxzcLxQhMEZy+e
pS8riRTPzVL/Y1PNcVW38VEoxAT2mM+tGzoFEfNmkbgpJVCKk6RsE46VhuLEB8Rx
W1JzOXTocMCljM/dgH5j+LoEfiGT4SLLeHorOpVw4Aoru5bywv6tyg4PZk2B1yY2
OaS5p1jKAv2O09Y/C4jEnaW67dNklQWErp2OTd61/NuIxzd80X6GOBs/d/p+R53N
T5h0dtazcLVhEWGV5HLcRvf+YdafQpEd4P1qszdHadXGoSvsBjAhoVemQttJwyu/
d1JdrUD4J+ihcODU+bDiG/im4n7/QVL8He9OXJdmw2g0BQTbKHDl5I4NXDuiIEpD
EW2i3E0qGjzdqN0kCTYJ9GzsWexWg1AkaNkXA7t2SXxLEOQ71DWWZ0m+uVAQ/Y48
2gR/uCR+VpnBmm3bgHrarZV8IisoEyA6M9tTffwJYmtp29r6Ii+JDRIPSW0JNCiV
eAxExa7HHUv7VI2TQ38affMpaORGrTjOI5Z2UePbK53u/nzgx/9PTxL4pmzieQSc
3lVd+bwgfMsVWnpEl/5Q0PJS0F24WSkUMGTlKhaqcGeq8czae9OFmWU9HBk0nLDi
kRjMxnct5SYFQOJnupdFUVBLRy+39iI3RtYLGbStOOjyT6wSaMa0y115bYdSV+1e
jVTciUbDp/nhslil/a4mz3N9YDxSiBlkgr7alxdpT3/3gtTbvBBS0aGXlc5zKHzZ
RomrlVAuBqh7IyHb2vpqvR8NLtIKuq99hdSlUQZPAxqz65B/atmwnXCwHG44OdNK
5a9xkIz1FFyNN9RumWHzjDOW/f1CdrbEovsAh0LktwPVk9PaEXyNdGiZle/Ynl19
++iXr8a0Jim3HfOmQbGzxfyTSyZjU5Es+V0P/yarmNAEl8BmUy04Ld7jxQZn1lHS
U3Ddo8EU3h9WxKlmzkICj4wkB4Sl5uCUuJd1c6SmO0mTXO00c07Kgw+Re6hQi17c
sw2M/s2Rrbk4QqvtabSvsTSC65dqB3+mebw4f+DV7NK5quLcgZDuIeSguxC929gb
A4V20jas75DyX6du3OCiITQRDW2oFUCAM+WNi/oOD3qk4wjYliIb0IO1a641uzsd
PXe0nosOKKoyIdcjuR6z56cVW1yzw5AUNQtaKOBywEjq4ofBOhvgq+T9XP+MSfmA
hseRS9hLvyIPQOcpZZAGrFfaBGOOhu+xql0oTKFR1rPLt16MyVwcd5smnA6S5b84
S0Dat635E+z+tIMNsewPW2/3UVbrMBd9X/01MgfB9R8Q9DAPhKtPufh9MENYdAcp
/o44j272WrPrZbjxbF2UI2+aLHQJPWV1CVilqlQUIuG6zVZcOEfSoFDodNm31y04
mDfKG+ZzIwtqjvWCvvUjwuONqLZnzwDAMFilUligkHnP9kkK6DmOJ31Wd2ppWElQ
lpUvX3JwQvYXXpSaHcHAanW0pi0L0Gb49pK+nnlRNmzHSYcewsMKyrFBHHxeV6hm
P5yRUErnfXCjtVf+A2MLXuQj9kwcm8O43ypW1SKbj/hZ64182WAoyDkDX8fqpr5x
auTcRWkP35TUERso2NnxCDvX+0HMDdL7ecHqZcEuG3DkZGko57r3F7B6nVgZlQ85
ptkN77ZlReXyHEoAAFTb1sKXIya39FVjqaWUHUMtv3mZsTNLCCRDEomX9UCW8f0E
49M7Z42j7Q7073Nns3Tt/l2u0JdaaCl87mV6A2eUejk6+2i9QuzvwkqRjBo7df0H
KjSuhk1xpKuYSm7czoRC6ufP7e6aTeFvBGVetvzff4OReHxuiwUdFmNyjWq1r9Tj
/C68ig+l0D1ZmjoChyI5Srs49GNwa4AxbBigPQ8pqlQLcQd563WWWobWalS1g/ig
Ekp+N8PzV+O6LNeB2GqDvgYDIB4RODqdSvH2E2b4uk9Qki+DAK0AXuIT+Z9rhsL9
ebUgf7ms074UXT2iqUS1kalyg/s8epXhMdvaOPOlYYTlJMYN+OxhKs4LbDR/bDal
oQwJETDJdcUW2NN8aMEqDXpkHtvras7br0s4YoXNGQ9tQxTwwlWVZMqlwvqZASqE
3lv9vcA/XxbtAkeSYgo6JAk8LAP8bJCQsdmX2qHmBoQAT6S39O5KFCxzt2BikqOo
aPhRDSH1Vb1Pl0lLboi6w9UPhHVK+NnOk/K7qmZ26kvOJI2Cze+1XkPVGUlzDejA
D/7v9Pxh0A5dHku+TJWCrVVzWdKo+TA/bhtaEml1TFvEVUPQSBUcBmKH6pub6vhD
8+ogZ9jFhFnyPLmc3I787XfSPny9RKkNbJ72feo0S6FHBp0Jc34iEBOi85ctqCh+
cf/M0QnOO8bZt0DhHvthsAdLXxVhk3gRtTcPnEU37uvRSnd2JEhsgKhg4dOF4Eym
n3RyqBCCARZb+x93AwFHvbwIOxVv9wTb0/+6W4d5U8jJGF2wd3e5ZBU/QfS1teWB
u51426jDx+OBM9KOvn/Uje/x0CvkcRB4gJWxck6FCaYHNnZq6ppjK5y2xph3ui+t
beS+f1l6ZhKDMvhm3Nru6d/CHDeNzrF1SaQdf9q08U4J9KcasnASCBh0rF/CMPQi
vDMV27l1Zb45Rag8tPHOQSrB5eOZpEUdopTmNOq7hmSaV/WJI/Mt5FHkNS5Gy7HH
G3RtT9raj5nSelXpjkeMDpSfltITUYeN6H4RMrO+a1C9m71CIz8ZT9PJoL2vpVKJ
CZI11ZerDl/M55AMJPD8pDtJGLbZfUNvhjZ5SuTS+ky2cNhvUu/0cr6jBOIgaA1l
3Xrv8fRDgjxWmi/vjRitRZRgGqd8MiRqpTclXRe5jG4Nx32Lo9uTbqHFkg5OhvEa
mlSixpczX5L+LqIbeCLjkwpR5+Fov7QleY8QFxsH+sd6EkN7tfghFx9l3Px8Xy1t
k2ti37YEKYvu0RgmlGcOGfWNYkLJuMmSKCJQMKha8cqZtAhghX2bPKexYVUEoiBR
Jg22xrOm8MtxDdbUUS54Y9s4YcutrThw7izLkbJPywGXw/B5RtnFO75fZRGNvpCJ
KYqmTwaICqy2vvb0Vt9TZ40RXit7fIP/QzlAtsFd+qg8u1sHW0JafrApbHmSU5dW
0mqh30z/q96cXRwAxV+RUSMXh3FLG+a6Yt3Qyx3E9HUr/FyboNFnUlM/vbMuN4G8
LrHJvJnZYaMSS9jIpN3kLNKxd5yMOose7ClzjALOa5gG/pClmj1W8cA6Y75ILMDO
W2APQHb+Vpbhm5FGf8bXCxgx3i/EPBWiHCKRlUO1gw73JC1py3+RW7IJfktwpKCZ
OhVe4aEf9rFofhKWREBhDRkmyWXXuOS+WEhnUF+2cHMsxtCG2ZlvvRXCTVs7ppEg
2nNrJ7gypbYZ2Ka0V8+01iM5wdYUv/isUjs4EDxLKzLJJ5Hhml6V/Qemny00Dqw/
JNiTPxpjiTQQZkJwB71jFDK/VosMEmpT2mTRND48WMQq4fz5ht8UzjgWCtmvLmiT
u2b6rYjfu9t5/vAkNFJuGIRYQICBgz6IuQP2i86PejiXoVVZrsqMYY1M+4lGhcD9
RZTLnnGda9XqxhQKbx6I/Pn890V/FCZRSKWRBFRdLqEA5ofaMZfOm1braRTUXbjW
dNhaZd6QH3bf3LLi3nuG0o6voxc0XH+7VjhfOZutHJPHrlVIj2uBDIKo+AEdl/uh
sfVVfTl+UL0gTOA2IgfuwqlUpLMpmIcH3bD3Z4sV+zfKbtoDoVc9oNiYKKA4jUyy
zsjvle6VSvq7NCrFhO/JkCqvF1eFroqOoOSHJi7U6tsYPUUNQSW16edOWUH+8YvP
EEZk2mhDt/AIuOWpeLyMAWq7111s1Y1O+sZtso0dwiofKuUfscl1LaZ2OxuIE3V1
lw/cFllO/3jocf/G9DZDxv8RjPfLCeL/RpST5ZPfSO1O+oGKOkdvcO8vC93YADlG
axI/mXLlSWXn8GFcF2BpDf53PkiINZftSjV2r4F8MtRr6u4k0hRuMrN8HgsxC0sO
Zhfrf83YTRKTPlO1+pC6c9UPt7uFvE33gulOMnIroG9kQce4zKEu7u6cx3vPlGKr
4/l6H9oQ+67TZ9PigTp+oOK5ip2b6IPp3/3TBKRS03fLnKUlGlG3vhYIpPeSDJmx
GMaF/7OaXVWbLV82lZRgKjbT/UeimfIOOWtAwCLxSSflbr4Kcb1abcMnNlUjEneP
UnkiLZN37A2UtxTbAXWXecR4l0XgmPpsYMSIXg56VKUFUsAqgmkcedfwgRYCArZn
SX5h10XPiA7L9IIB8h9itqW2rzp/GjKzxO3esx8O8PxBOJYB3PnhxKUyRHDiEsDR
p3m3nT8zKSso0GEzA4kwfGVj5jT8aY+3NCg5OIJErhIQotVn7uat/jYQpMs+sUOq
tm4NPWPHq/7vEQ14AmQEhLKUtGE0CQ8FEBpbJ806vlY4Q4xUcuG/zJmr/0xR9BwX
/7JI59mY7QiFQh3LIdUk4EzogumiayOBkz0+7rjCNxvfeX4vBVSH7Mp3eqwtL2uP
GjDLq+QkMc19gP+TOEVNp2foZSnZEmUfye7hpEpGSf/Ua1Isxtq3c/NdZ+V/7c+7
BdLE6jVqpN9F32q0BCp2nmLsBv12lZfbbx4yEXKSxlrD/igPvCMW4HBMUlLmAQlT
Ytw2s8dWlq0kRSmE3prU0Mwfa49urr2MK3P8h+anRePncGR9W7J0q9s4ax82IWv9
wo4aDLWkHF3MRcIsDtRKdfi5E8yBizYFK77P+nhOMXJiJqqEKEoRKGNB086kUCuI
vZWvi4BMqm6Sa1dxDXqsazW2sBScGpkojz1QPd39xlwyH4IvRrNo8e+AbHWdG6Rq
1iRi2mEai4ZH7uZ80sYhl/XQbMz7AdiQGYb5C7BTHzgaGXBwYHcovd2HeFioz2WH
GVeL355Syz/Ygq0/vChazQTKL1gXSLPDtdEJXgKAmfGwSRm+hqIDrpybx2AMKZGv
ckfzhTZCdrz4x4aOyJsdaHhriE221C1H3WyMBwuWjrmPXEvyiZCp90jWTJAGJbFp
OgZk3oZWIfq76uDV19+3t69xoO+v8h0BmURfm6GvTIcj3/voV2ks7hyWHWTWyKOy
pkVwIX6wZ5u0BpfKxue7xLKarCXOJzRrONynEUwzj1T0VBKg22bAbDc8awOi9HpU
1J43C0nDGRyVRTP/jfebHLqNB8AdX7/eR/ZGZCYzTbpZdTlbf0A86OlzcH6Dwdq9
kZ+iXjanuTzQftfk3IwFV/yZ397a4MFDBmMHU14Sp4wUcrrO/NKwT3fElb/+PkVa
/YlcZqbbyOSwfsWRNn00mhj+0co5QZvtyUsGi2zKKsrdp6bPW5roC+tVMCoxe4sV
vEN5Qb4nhNT3IUsM54+K3eXepQSkuVZHSlApcpSespuQPDqupwYVjkM5HJKY5xV+
RJWEsXk1v0exBXEuj3vDrRpOEd3jUQa3B6yhe5aICK0IGB93teEBuisi0vfoSp5p
MUlU+5VFQSYMYI4/xvzSHxzbKIijf+zzUs9sax2YvUeZi0GJWmy5oXNhKrlGurQd
eXdQBdCRYOX5zVwwHZuwQyHCyRy/5euN7Jacw/Z35F7sQCryysUrpaEHDYKC7MbW
brxzCUix5NrVBtHP1cmTXEvRTRbMuCoIZpIwHDFH7UpmaeAte51EDCKNFWBcRVNX
t4LcY7Omt4Lclttvyz6vHW8zHIdekaK8pvpPPVA3jtu0aeJ7vbW8WYJ3oQAjzkUV
KwZaWsIClaW/s9uNlfGIQbWIcebV1t2dIBx0MVJ+BCmDHP5LJeBzLrsaxBrG7pPt
DGYYhuYE7U7GcYpdy5RcgqNwrk7ChV9uVfnCOpuVG7/Mht/VG3K4UBmyM35aOVw3
QhZAzQTxE8Hk4Yz4MCxGC0crny0gDwbwo/s8DkcGK9WQQaar7CWjipFsa+aUSunk
mgOsd6tKAkXOyOXYRCVCzV1Pj3HwIqME0AkTcDYpCFh9kl/R/ilyLXjgkHeoldj3
Qf/qz1pJ5S3EVU01+EXGrOc7qDCL9domr4+JlLhirLHnBbXZS38IVxukleuftjvT
3nqj9UkZM/g9PxMFuolGhRaJkfoF2fUviTXz5UCZ0EZ8wJn1cabn72jXl/EOUF7B
d9+YR7GyI4xlh0UbQjVO8FmdMesXtcYYovQP/8uTJ75VBDVfJh9/pPv+ujwb6fm3
LBzdjZgoUCQRaTwNiDtGhCt7HaWtUc9HmX8AZsDUWycTWlOFxHNbLZ9pnFvGcFrJ
hFQVcBsnkWP0YEv1O6fQJ3IKfSlmH8atkGT/EHoGH9gB4ME3QWI/jzoRquU/G8Ir
pWhewF5FT/7ce+ferPRZk/iUNNM1QabM4VnLcilMB31iTd8kD+GkKSPQzP3F0QnM
vGkHT440SPppf1pqoBv4jmDU1bci2vTbG6iLdypExEIw82VCB1Cf8jE+wKrHgcx9
EJgI84d9Og6HSidAXk0OjxpGUfLFWUztHytQnMDE5hhQH0NzIAGOKB1v573A9w4Q
71PJRqbdFJGgW4+X6tSYCQw6XFrhD/MzSdJJaAEbnVVzIf98MmWaUPgSnPllmKMM
sX3D4c1qunBCnwGgwmbsEaFQhEHZJ4Fov8gsHkaZg3fFR7LJqR4MFD5u+S5y5xqd
ec0OcyWf5wDNe3gD2zSS8LPC8Ydy21CwbQ19N2IqwzXO10J/5Uqkfn3gAAox55So
y8JssMEKIdFJwc5QnIKo/kPyyRSZXZ2zDb6fRjTfOszOXoONQyZcILk2EKazC531
5s2Y7NZMJWNeOITXktGcITOg9w6dpeV+Bau2sMYAHKKSJmTMouIOoC3G/gWKvCNr
togBz8N/goraO6ugOb/BQdOVvz093kyVW8S0PY/LVTRyemmF/cnDqSsh6rRGv0i0
vHf6IlOb61q9mdmxBbiV2MmOJnUMs8qMReeVf0Y8GmveXQh4nFXbQbpK5yfvmdI+
NzZJUie0h84mKYBUtG1OT3RzadQfNqilPRvLcifzopbPGklXSzolFCK8dBm5j22j
gGLgPIrVyZHwCSc+U1Xy+Z3ovu0OX5AgrKdVuNurZvH+jZEIZpZN+M/6ipWfPj4d
+Hk9GdX3dU2DgStObdJrd36Blp2XgGjCmPebMCIsp/WaEHB+CB5em2qY9vgsHAzV
BWJoKFAoyuVZ2erHR0/zZBwQbKthOW66eEBxvulDkU7cdSALlNr4FvompPyekCTG
JaOiDb1xvvvTbsxXKc3q5554MgeMQdDX85jTgw9tgKpVudVV4YWdTJcqbrYk4/JO
/Qt1bVx1hDSjyS4IZYEElLq8CzBcEEjbd4F9TLEjZJ7NwCVsArcdCqR+9s0PYXJb
yU/7vHhcR6cT8xWAVXdltRBcMqn+TEvhjvzZ/JhsgdEJVSF03beDp5+cEWj5TIBv
x3GY2dBbPLpVYFfrhVecfYKSc7BgjIEdF9Dt/x/VKvzNADHWC0Tpdin2ipr8jazg
iaAX603SLSoRtgOBY9WS3S14zwTrljJ3Fwj7tYwCzxBF2gZuv8e02VsDtTUEg8Fn
u1Qv4VNZFQbjXLan8CzeUTrHewFif2UjfLPRY3lF5juK39jRK6dOpCq3LQZPVywL
pslETPpgZTHqYXKF25HdVwL5Trc7x4Mr0bL5SWJF3yzc+en+QEGU8RdmDU+fownG
WhdkCPEUO0eRO34FMw7XJhV6rb/YfTFuNNbjdQYgSNCPP7Jdc7hvzz8ogNJYqmYr
XVVCPLt/bqaAfGBTwa5rtZvhBFQkfRkruXoQ/NVDeq4aCQWnqu7d1AxI5cvoTUQb
efK/WNzwju8ba68bgLMnD0lZPYIZ3iNjjAoejuMO8jOO5QP90qVAzMveU5jIYxG0
wcPLgKcian8mVHMUS1v69VEY5RReSLPtnvea6rC3iCHXrq4NQIgN5pze/xki0gAj
tC4bmW4CQtFFunrkjjaFG0ziQoqItq0qBPVBSuM1CcHoqlvm7hSNVJZd3GNNRMwq
hmD+zprQ3xjWKK2+nK9ENOtCli61RVdEpHLj1j7QOLTqwpm06U00y4EYdIgdXhL3
WI3uk0mecdd5p5sH1NWYoYTqJlyoORyHaXICtC4/b36PZ/ij3mKIUKgVmEWqxAzp
N1QfyIDBDjbnSqybyGlmISLp0A5rOBXImMMfTWVgj3Uxd+N1VsNtzWwJn5dcmBkk
aOEOWeG8UkL3Bfa0JvnDPZqgwj7rUoHcNiPJw6aZRJg8oO12YjYmCEGFyIfyaDeU
qJosV7kXzH1h60P94+E2XC01gaooSlWHqxVpARlIoPvBsmJrIHjXWb2O4Nd3BiPd
S2qOylO4/3rEnYojGB5eEddRnEyPb+nCn6PPg+8WDUoMMWYTlfWN3yp9lTC8q4d7
P3Y6f3KOiFNvYQAOT79F2YhPuob02c8jD6q+vgRxubb+FJyPZrSL3szdWoUXGqcl
lZXiGAFI8end1/IT7nT+M501k+qjV/aUosguL9HS+gnc5Y1g+IJcfyj0weTHhxeR
DfUjD+BHTQc9Dt4PZkbGpztiowlb3OxqwXZBDmhlOA9b7nAUQyL3540u0W+sn9F6
MOCuFCqqlgutKNToZlkNiGGGzpTYQrgM9AuhmeaWWoKdg+HA806FKDjanPygvisO
CCRXxCg1xEN6QsbBah5shsWkK38YcG3ghrIawk2ZRLrdbhrlF/JiwDt6pb14pJEG
G/llREGEz9Xf9wTjRse/4MaJkoYuFu49dXRRTVg6g9nge9qpBA85WaZuxqCX6U2k
koaEXVVsigyBFIdv5ATxWUAopYfUfbpYwRgf+rzzuSEqeRflhEno9pQya1MKfScV
i9d0/5BirBFecIbYv+F8FFeKMbwjxD6fMyWN11SkajETMt+PNY3E4Rz8PhfcsEJ/
q5fc7GkYI8tE+LajeBZD5pwilJ2m87JbjInhzXQPA+ph9PD2BJYL+ts+7BHRiyCp
z919Z/nMsTk7wSlv7agsNgwC/Gg2ZqZGX3ra26QTOftEjCa9Gfuq8v5gKlblULH1
7E9LIJf5BFzQ6tFaKTCkV043x+V31zms+tYJuOhmgKop4FttkrwfVl2amDkbwu31
8nbIu9eoO2sEbPnpcFQK5kD8hNeS5OfODXe/mkt3kdDhemhZiUNOKMcEr6amdchG
VWHAq7P2PPF83ZJsidb0AdFcLwpkXEi4bYrRlLhm4LbMoP0C5j9raIkV4fWEiR85
7snaLUPGs16ODQZVB+63yfkr1gUxFYCRdEXl/eGB7lziJa3+wNxr7fA5W/GxcjBn
3rCU3SeHjEaSrdUzomugdSoyLZf8IMkWCwfWHZ2VB5lHWTp3BPJlyXOCCuGZUNr9
n/zKCFCwk6ElA331tp7fRIZrVLptxZuuQFwbXcCbsi0c4oMIB6DoPGcp+js1cT7i
mFYJjGIyPcQyHua3Gz9hSmzr/BAUapW6vr3vW3RYHW8SRJLqz1FlJ0X+w0gk4Sk5
O/q2hlpFmANyZapK2FPPamgM2rten0uYaEg1hubHX1jgzXRQwyWrJ3OIdUopoXtj
sr9tLyuCCqge5OJFx7QVs1qah+zHQgFg/d0DW4z+7M8u+5qeDSCUDnW3ZUCRyQt1
OdO5yH76leaIxFhTZqFTuMtfmaNgkvALwHqVK7QuOKURpGOYHp6GIjaDJs2ZEm34
Jgz8HPbuQsad/9zZDlST6F0RK1yrAgex1vKB3Uj23oicsXQ6P0EcvwKJ3X/dwzbO
Hb1/EkE8EeNqaArIl5b7LgzPEQ1JZzC2TYy38amzMJWWCc7ZYFanUL3RZL4o63gD
ofLwW1xqKlxuhIRdaAfHqZKUOTYihcyvoaUsopiJbGxoQOXrWtjHeYlw1EgY0odw
KKPwakba/h89yIWeji8jlMo2aMMaKCe8ljP0d952gifHmdOZRM6QgN1o9YMvbq3a
wLebdsB17QUjkoiLwwAU79QLRupF1QXVxUpwynvmZ6lba6x5JW96kmSHq3t9oGye
K849IMB/vWnGNg8PWi18ubCYoyBy2wATRVGE4PS9gBmpuc9Jw8VIDRH1ycxjWNHb
px+a72axwTRFWgjrweYqELxx66CmpbYwT/J7Km6To40N/H5RynACJiK/9ipEzJkV
p8d7vVQ6m0wb3o6LWugaCgIClU9ygs4hXKA3nwlzieUZbgV9XTcxBmitlgDCRdBR
shfFcFwTIkkri0YINl4lgQp8iRSgYJwpnYq9fK15Vh7nq69u2+YTUOruQX2a8FoA
sFqXafdz9HEaIl3Rq9hiVdW3uM1IInsHRb6qlaGosxZn+scBwRi1DjFxzceKkpE2
JV1PrLHI0GZx0rpon4Xmwpyw2ojGKDDtboAF/XcvBfwV3PggPxVbdY2zFTkJaIKT
1uoWy6HgRHJEfwU+DVMTiVz/hyqIIUU1V/hWiuYHV2bSA0ODb7Vpzx6xHOUSLho5
+Y3TnKg1b9fN6Zs/k2T0omVrQSzhLNvlT7j/DmBrKDvtE4bpGCw/leJ/O3jXlg4g
DnDoqwCd7oO2FX2p3/DtxlL2FqG7Oc6tfNtFnft6PYJZJIwajMPu8Njg+fzvTY6I
oyLsqMmj6pECWYVaWGeTHb/iUhiDbQ9WvP4Sw1+BB9eHljjoiYrqYKauE3p1+Cxi
JLd91/iHpueA8RpDikIQEI5gdRmwiqvoqImT9HBYpMOebLWPmscxPJ9LIAeZZ4vJ
4lqhmopvDqQp/i8SCVW0dd1mYi/eex4vnaNsWb366v7LgE2i6BEYmL9q4nUcYjnX
HjCQLWMv1e+ZfFrnaa6nUS64PqqcbP2SEdtbQdElZbapHPfVjmvrrz/Oz2Buu2rn
WbkWqhGz3VcFYVOWn0+iaWEDdB+IA4iBq+wLEgOPNrkLJkmAg5nROR40AxeBixSl
pC5s4MTmMT/pYRFBlMAGxdLG+ePOeq2hu45n2mvmg7NxAwKvJjrRDGcmuvE7qhyL
4GZuSYeYViYxxvvEGTRrOGEFvaotmtpe08yAkWzeTdO0p5H7Z46wu0At1l3miJL+
CmFyMeXRBDYA5u0WPMT55vBY2/GirLQ+aHbpKQ9WoxeuFojl+vL6J1rEhW6X8r9Z
T/5EKKtsAzfhWUHGcZkSIBNr2+v31bKARGgqPB3GGkYAAC1mYCKEmPIBca4fs6aG
qpuUYpvA+djsvX/lXA4X9LXuXqJt4ZnCReFMYxVkXRfDiDAXoRtOPtmi7m8tpyN1
NaapWl/+XmmXHqvNlmyellcd9juf178C0UAHNZOX0xscd3WDp4FlCdEZXDde7Jnj
0I9ofd+EAyFo41akUwJ5fZd4udtJn+pLjnVWKZxpwE6J622sC/Vbf7mGaCAj2qYG
KL9jXntpR6H3wEO+m00fi9hvFMJPk8OeYrVNGCO8M4ISm08esUlSXCOOBts4cbST
Y3Rodly4DuS0DQvOWiQaRb3yaQ5lphrX1Hkp5yhmV3T5JXokM6fABnZQc7mTOGTY
2aYU/WHrNx1lEbOnnLuvaB0kbG/d3DUUVYJbKa8pVCIpntFd5U5eUfE7gTxHvIo4
Y3TaSWfVja1veY+gha0SB2sQBlpz4W6QyIwo0EtWFi2Ym61KVGQvHO139+BG4j2c
Gcm9yGyFPvCuTGqNw2YqdtZP4XgJedlRyAfCA0vB8J/Atq6chVW2gGUCm/L3Glrz
0u5t0sEyO7F0TK7ZD9zwZgfkE84Mxe/dDYMiBaQIFkWdLA8UZjGobEcvbgVfYWe1
O+J9nijcQyFlpfQZmrpTSdE6Ji8H3cmSzqqmz1ATqCz1dNkuPXURbKnhcZYkC3pA
OHW4Haz8nkcw7QCx2ZP861QuLr8PSNRwEkWXVfk34KTJUU19z4oGmiezZoDlacg0
rgCeHznXpPCStd/aCxGk1hZ4Hx1Lii7VK206//hx9nzcYf9slwPGoIzo1NMk46h9
Sb4JseZXYSaYmLvClfLCnunWKfZ+JztktTeiUxn2c6Lp+jgJEUeTPVjYTGUAo4gK
6LQmZGjq1Nb0yD5E5fyt2exrFgdb/oLTmi9WvwGpEHiFwQlYG/pnEFssCOAnpxXO
kCKMqeEUaLDmZ4lhUeB5GKDPhq+kbl24yNBHtynpsG2nwqwpnch0iA2lj4egAaAO
JLmbovKuq/gs3y9t3LPIgsrH4usfweyjRJi5lYuHPNZtGf8+au1srJUKadbrfBmR
qndMdWAH8MgTdbuUnAUBU/5FuiNZwtjriLbnGkri6qIwEHUBikSS8AbWhhX3+ivl
Qk81RzISDzqyrijOv4jXIhHLeBbFCqAtDlNEwoMlV+kgOsI99YL6vYaRCe6KOhB9
9e6h+5a6d/PLCKfcpenxLfAW4Fpd0rJ2FpOpkJH+vAv3V911dmAFTxg744W3Jn6u
eKIsdLTUrRK5PIeTL0zlNYtKMl5aY84PmVNzvN7KQHS9Wq2n38T+lcrdshM1XxXC
OgznZsCSYiGxNizo2M9hHBsfYUOdAnz1rdeY4Odh+AV5+Pir7p8C18YsXF7QMSlM
l8K66KMpOzMtNQee9vjRvgEt60KgsElCdlaJi6xz9isTyXuVXY1pQ4yn4BZv/jDU
PyEMZXIhJEl11DDgmgqGHZw65hAQmVRtwWS+/0g9TAyZi0ttbnilgoglTn13I/qb
NVqVhJiyySdOecvZXNj5D3k9j6vJL+PWVIMHct94D7oR6b0Vbme2Skv91XROkpEc
hUkNODHX/MLpCYZMcr2oyKJtk5c8fp4raAv8FBAw5kHz35N5Wf1EUqt3uJ6JPnDH
hLGFjae6SIzEZcicoAPNtbZx+zCNmseT5mf0kRwiB+IZcjaxwadUK+JjO0OHuHCp
6+zjepyqZ7dDSYF3wbk5ITjl2xI9uXPUcnC5r5DkkuIOff89NT926VGrX/8iPVIP
FvT3RHTxE8+JFTNR2pfTKT0wqVq6TYTA9izP4fAI2YlSfqg5TEuW4UXb5OCRbZ/1
ETQaEhzS4DoW92QjI/n6SvOSofVOs7UrhjmOu3hHIhvRVUSAw2fGZkcQvXK+s/IC
4yl+sGEsnnam/shsv2OoYCjMVbphaWa5WQmvIL8inFpqrUG1hDxpbzvMgTcyx1if
5ZH91AIp5sbkquYZdNXlkAPXQLQ5/4sHNM8G5SEy1CvqpL/M+L1lfzfhZe7+Xr61
FStB/KRmY0kqhaAaeuqOusQhfmBQFR7cXxu31aU0agfaN8s0X2TfCA5NUIFAS7pZ
EV930X/b+RP3lKSazhSP/IRwIc7kcvHoE+5dMRPsO0HcIDTmi0gKsNHMjpmSmJuX
yx+77nyYkmn0mkPU6HtiO2Sa7pMAdSPlgCe8+Ozlah4ImeW16sJRHq3J61dZyZMT
OlfLP5s0Hm6xDSPsgZ/iD9apD+ZLJHEMqkK1xRZ0OX+sLmfkK1+FteH2nT9WJFfU
2OtmD0anbmxmcmK0gW1klxVU32BukuTeMVG8me7syWiKoJEhj1k2A9PP6FdodbfW
TCBVbBnmT2JJL9wDQljt1xteRcyCWmEriOU9n4xJ4fqjTgSq6HXcJDo0//ToTVqk
gQu/pT6nYpDHjTPozxrpIZ7ruT0HlgKWK4J0+QgBA/hVyxl66mPwZ34Jb+yCfID1
2t4WW+bNZEcc4Zo9sZW5SuSIHkF+4wNJtTnFC/cTKeftuIMvlqgO+pmiJJEqnusM
jisTGTI9BU4rJSiccB8rw+skQNMcRHu8W9kkaBOgkHsKZS0aQLPUUOrneIGUm2MV
Btl52gIQYY45FBHZGgFtqrESPVZmonAwhAMCaPfpXuok9vUUoRzQ4gcDWp9JafWY
R1ay3juoJyA8MJIbvssgVOnQPFNqUvoXCMsGsuMari+dkraKEnxKa1SkVwIO7jc1
HkytwvUKD3qZVX+CLQAIdM4d26R2QGvzziqKKw58mss0EQ2T9fk0NFAJ2SlgGTQ9
xLsP2SLiJOJzpjW+BUz86Z7doAAwnmBb4cpx8FcpvgULy+iVZ9A8IpMZLzHef9fu
yakcNrtiPQpe8k5PVYHn9fcWpqrNPaiExHRNgfotQm+obsqRvF13WPXAUpWun6Yi
8YHY8ZcfUhbH8juCdJ0c5b887mdgAbtja7CR8HnXcYR/TzaabKhYdtnrOlLq9PZg
sBXliK+LtKybv3BJp22e/BwE/GQ584iJr3inVvFimTQOnudSe8yQO1ABiyGb69UF
0T4HiHOZhS9T9zhanJRSdMoSOy8qiEJeTqdpoRr3c88pO2uM5Tej/04h6LkRYn9p
J2qmeCryDadyhjDIZcuojMK6kudwJ9cQedyF4WF9KYh/nmRtjvDqWBOwmG33eXwV
nXN8LeN3d2ryiYCRE9CFgHoV1wCW8o/tAYgrTL/heGJBcatvRAdIZZEuv3XdJn+v
f7ySBLPUbRnjjfVOf8OvyODTthl8EEQlJXsY4shm/JQNhE8Wlw4G/jvV25AxY1J1
GAxkh5OK/hmAtHXBwklTnPcyDcfqhfHLDFrMbLw3Xh7vAc6si12PXsbOcdfIc7Ep
PraGnUGYSVJfLh+JfsDPdJwwnVtfK1lFWLWY1FJDarEirHFePtHcYxNvVj0I1Nv9
PwGRemqZTsOaVuxw869SHpAN6gbdluc/sSjOxkCYk6QUR9qTAELXF5pMNPaVha6s
ApWmlSeDFAhTgAPu4niHcdMwtFsMdY+j+Uoeqz0FX1GC0hBNsBtUAOZQQtkDgNXZ
s/vi0IYcOQW0QKHtI4dCYxukZNhrrkHOFp8ejyAg7ujMqGxnRSldrDTZaQKhEiCO
1UQOQXXI5I5rtkMTlg3rHWss6Q4mTvXF1LpyLww7ha9/X8iUIl9E3xYEQinQfFw/
aiyxDgFt8BxcnGKbca3hIVK85uDbAWaxOmihBZgJ/XFgDZ1ckO+FMCYpaizx3Xt6
gpFZX1zXF6KsoxRPJFthk1SfXBZTueJTF1LxY7s49/hv4BuyXzfiTvB3PP77j6W/
vlHJbBa6EB+igYQmq0/znznNNsV4atCY82++pzxmxhZlHlWEfTdoM5qu0LBGMkgT
eiRdeyxq9uIXZQKT04JlQk/5PH2n3SEA/sXYduGtQ43UjPoVFsz82CKy/vlsLFAj
AP11WdZRZQrrSkL61yIYi9QJd6M6HVied1rBq3aSiBmDqOhM/HduqhQ9tgOAEhaj
huYkq2AH9MYpcdzJZ8Rbme7oowgQdNNH6okJ0eX6ww1xe2l4I12PAmKRyWoL2u8e
+e2/mneWdLEpf+DeYTH4VwV/tt1MBa9qA5eoORyNQ0b7eTDGI0mxojNvyo9oLkCG
G1st2jTUNmiPtKPSYVPbqLuftn6zNSRB/jU/1H0SBNJPjjKp+HfiyQbIrKQcv7Y1
04ZyTP356vGTN+XFl2N/KP/6XPDTzaiwuzOixbFB/psEYsrV5sO+54gs1ITBvm/r
ZnwAvq4aBaLvQsgtV+FwSJKxKAleIX9vPtt8Fobav3R0ckAGU5CXCkh9Iq/gGkgG
9l7dvjIpJasHYaJGohnyf83mRDfxeOayZSs0+ZMoGW6T5MkVIThVUL0Vwope716S
bbWHyKHI8Y3aayPC4GTJipbhXRvWdYQqyxxLHc8p5R4r9FwXQ+ntuJXOVnCDuvDL
txmw+J7MbK6nFm2jIcmawhaXwdsZN9xVaA+GTfM4sDa2QljuxJJ/GBTW5SpvmOvk
3J4Inj+Rb89def/LVFpEmaOtgUHcKzVqK152W51udjzDjPBlkYCHpY43hZ8EKbDE
3LzICkfUEQ42J7YKrMAoulk/DugUbzZAPOGPi7ZQxm0+G+AOJy7cq4vr6j26DhQw
R7qmTU7mKRJGcBVEcC6dwy9OYIMsjs9PIpvq0vLeAhsohLrCnFHOJqOAZ6V5VCUm
MBHLeCCQ5yQuaVpdl2BWUa/zGgGRNeTIiNnpxndzzo5CQr6+mMlxSUWeeBs/MQME
kFsey8ecquYFVFNEoUwia3ja4YNPTAUW/Hre5SKmt7GHgIhRrNg4Cv9F0TuKHCJz
OpDMX2P8lbZPi9eY1vSGuN/+E4R2nBhQ+dXqZSDZPsA8k49MLH1BoXEjO3gZKvOb
Nv5K6V11bQg2kD2KcSpmtgkhuQZrkoyr84SWpGNLJQof/CdrYZ4foGHDvWGqzbJ9
cR7XTFDQhQ4XFCB+4iYPOQKg0fHltrzfZ5U48T5id7RV9mB9L64bfRW2g4Ang9Ql
D5EvzKHYPY/Wwcm3hReRIjzQRUz0NfYzpA6RARkw1kqot1+DbMX3kPtp1zzb0erJ
CouP6EzHlebekbdWWEu6lZT+CEh5MEZPD1pLK8+O+JW6nlUetCVJKw/XYrxNX1Ew
kL7B6ejJuYrREay4l2QCyISIJsVzNcl0QAqr0Loj/hYB9ni4VTefNXchhNmo+O1C
0OMAoGZHiYkdgwgz7RPrW4T/CQymoS+oafur8+Vq9p20Pzii5Dk0kqdaNwF/g1GD
Cx5cJG8JcwADrimCZaQPNycWvDTDyA7SepswaYIBQWHFR4r09d2L5YoaCUaP7CCc
GTBjYEGqoXlK9teqsSyWYHTklSMsbv0ibOD2UM3UvuYjITPkTEfov1jOzt0BMfL/
yQiTgbIo/fqwbzjmOD1nN/tkGRo8kTdI6a40vR4ePkD2Zj12BHMAplgglnYjWxez
UswudDAOv/3k83HBC/57h7ahjWKj/N6vt2EeoTwA2ALDlAkocSTb3F8zq5oXl7B5
sYlrDnBQO3hsadw7MPYpJUpDlgskeyedvv5m1nWU8zG4fYeDEfHdQhTid4AMJtX+
oXvC5WO8SPBIPd2tfdzsPYGMJh+kWx+n4r9Mb8CsPf3Tn1fyhDRjj5LrEy3O3X5q
J/fa0QO/VAq7d3AY+iqcnSDAwrnZgc3redegRvERhwFwJjS+EO4LCp5/Wnjx4YpP
x6yAir+tMnwf0AxjL4g7EB32XYQGsaxdGpqdQX36wB57I4OYUes1rLoC9On/0bXb
2LVmt69tgANS1+XOz6dr7FeCYkdiaLcqXy83ZE+ekcO0jCsDieNWc2mOZtndx3d+
0LjvjBaYO6gIJe1ghhmgI3sNjIywjkQhtx9I29lmxCQY4zXqHlvQTYFqYsz7GzWm
94hYYd1U9UToaz1ChnlP7dHBu/wp2L+Otf8wtSvmdG38s58y9HhhVfYdHY+eA1v/
DZJ3BmzSeMysnSmbbxtJebh+lNMjiyITseCWXNkG5lWlzPBAscsjsTX7NdDGOkMo
ku9eaKlJpra+qiTz1qDZBRCMZ6ppU67fN/GYQMBW2U3i7Rk0IfwKx3g/LCOWytlC
HoXTLtTQB8LXsn6IEli5TOjnWYu8auLolxL82KZKFOi7xwRgvwThJzo7tmKgIxie
gY+Qi6XpAOq6IN7FO7Y0hC7pjtNMRieQh7WSJYaEDX9E+joPWxL48gPsgwi6Pl0A
Bzvik7JmuJrKkY8ZNXdJpM6JiGqlyv4KHlyqQru3gh2RWRjDoEUV1x6fefJiPLyZ
7dNQuldzdiZf5lNKqLRMHHqN0z8/8iB2ECyE93fZJFxISuyxXmLJNduyx8w+ovER
TF+J6npmjpNsjmMFxxUSJJcNNNvBNObgBdIzMPXLjtSF6u5GAv8Hky4xQyB8KRf4
xEAV8R4LJD/t/LwJqsnb8PPVxNyvuH+nJPtfQmGZ83mhQEaoRdpKJuWIJOy5zNwE
uMG1inXQJ/qDgn9NZlq7uvfVCO1DxBbYtUkW79ONurxWRZY/9lrhSB21bNk2azdV
Qnb7vqmDYQKMdywIjPlEH4CYYuo0f+mpPLiKdc8uafwNFL253OZ3K4dpzrtcp+EX
2acyErqO5ufz7IWkh93JDyJaO+8pRUyC/kw8IeRdKGSAiNDLqefwF80vyUnSOnlU
UJf/sqJZX385CLdmxCWZov6W3Qc1P9+j1IWmwpJnw8DJXMYxNi1PxYj1NYDlLImg
ybYPfga2hspcz/TpfmbKNMTlB480umqxhylYs2TpUhrAmJPq5Mekh2rFXCHlq2ia
29glnnXGxsPJjtLG6todGIpam9UaqAaA+KofadLoFFOiSOhNA145E/yV605V13LH
NFPwaiKPv52TCzv4ZNqGbxLkxHvqkwpH/t26hHITdkrJwrigeOmVxVgE/fzTo3lt
Nqb7zp3qq6W9nXuP1NaDxRyeAl2D2huaWG81vghhCiofsFxCq6jPtscgtHVDview
7NpoFZE2tqP8yhTT8farr1vOILfI2NNj/a9xI2VKbQBtzQuIWQACzEJeWL3tZSIB
cRsf7UGwqPPBu6WPbyOpLYMomAhKCg24n78qBvm3cA52cB9fuKs/iob2fl9WC6KN
26abHFXCFv78x2sWIldd4QWVEy99IDPXjiwXYHeZYl3lP8ZziaAKppFjBqLJ7fGf
k7rOnyKz/LsSlwe2ViRzFP5UmcFWs8CzxIph8YTC4NnjsSN3ubC0qf28Jt4LTjPR
Ll+gm+T8wzTR2aij5eftbvZOcHdUG3gSdZCRqQ/cVh/MpOfS6WgwRiWS1cjp3TXl
jyzC4bZdwEb8CFO6fEkOnG8/TPV3kyO42Awp1YRcA42riKE5+/54YlcBoyxEglO+
jGr5VcN2oCW46PRo322kwK4tYAxgNTSCrZ5zzCxg3FlQBRDR8VzMlqYNKj7lEihT
ubZo2TxTZjtwFRUE0pjyRSCfHzmgkLGW7JKospOlLLrneN8T0WzrWfstjcNflNX7
tqfNjRbri+HlsWnbiBLlwd9A5c9k0x01HjTlXjTjxrHXoPI2H3SNAYzR6xrOp+5G
JSd3Fi0LpHR2SWmCP6pxIqjYMNJVNNxmfXS6TXZPZdfGza1q/dtisBlIoBVQ2mRq
EE1tHMyAn9h4Gb3gl6ydqiErzvQesyf0KoU03fBYppr0Wc77VsSRd7FRFOnB0Ora
nxE8ckOKakkoaaWhv2BPH1yoWBCXkuxNojHCpJNRmTans/FUXlK9D2v38N0HxLAL
9J4VGsI4qIPFgE7t3Cpuygsriv4nQuL4V88DhCKNn2AytH67YvRTdaYtYbat4bTy
HXUdsWm9NcUhyLkpBrCP/T/12xRROaAJApts6DBQMWz1oemvpkvhYZcoXPx/EzVJ
vygyG3mCcvtWpPi0Yu4v+CjZ75ox5/y3lyxO+AvEv07Iw4CF6OsWv4axgPkWrG9v
SFPpn6QZaem0k6VoadCvgyZagvRfYS1zn/4eXr7RzyYvc4gQJx1dzqcItnX+8MCx
Jw/pXyQZRh+WGQd2I4+mfZJyBvhLSo+C6tC2dB2sxFGTGigK8DAoA38C8gi3W368
abaSa8FRThDRstncESwfF2rwD36uhbAYhOs/76HMs/zHE+rWu9t1xDkAahP5Kloe
CRgUQ1aZeBwGiVCK6HG2zJXEzjplYS7F1Pz22AJjMabQ1pPlvsg33eCf0wzXniHB
IMorXlCYoodlrxlYNEBkMooB/aHssnpYKQYpGaHaQSX6nnVZu/FKXxfrtpH+g+6w
w8SvqMi0BQVlRuLrsQitEIHxovpk8/n/QN6PTG1go1oC0YRKyoA+p74Az5exssU3
6YUcK8lpc9ija5B69HdUBE73sUjfVwSiE1o1uUZXSlv1bjkLSnl4LvDPjhwe2ws8
6hFKswOMexiPHgNvToaTKPzQKiyA40ZfI/lGPB4VrMqDv0ktmn8W28HRcR8SC54/
RoIe74LrlvTZWNi/2TxclP0F4dd240ryLsQjlUnMgB6MAvX69NyAbUINYlEQCiqE
jBIHACRPUv5shv7UxGRbKF0PpMoDBKEt68fm5vzG7+gLR3EEL1zoUIgvxQxZSOaU
dFRvHXuR0tgOSab98sJ72xSmn8IGV47B73aAvncwQUnd7QG27+Gzj2aDHq+ou5mj
I7XfWZ+/QJFDfKwTSXSe+2Eoyy5B9JK/HkdQ6cOF2KyiTENHVNB+L1Ji0960dQ34
skh/A4YlD7jt4SdVyy0Hzyb4M7B+CM2wVpkUCLWbxDBXAj9sVduPZxPDuYO4lCEV
8HvMMkYMHXce/JWg6N9NcTbvKDqD7ehuZgDWcWKS0dlOcejVwoKImmNULVkilgPp
SMHrS0uRCxQVOi/CQNcpqD3pPW6qvRufXJRJzURZFcMF3/sT7p/sYY28jNPoif8C
IPBAu1Q0p3gD1QiIz/yOBhLI+F1OgstH/B6ySuLlmaT1z0pzX8RC3NOIMT6g9+jX
gpM2LmUWx6RKzaU/RwMZNn7B0fNh8+BR6tNB4UuGqlUuO0yUcD3xQLH+oC/MnWZt
MdWtCxI1FKHZuquY2qwcvg7MDkcByG+HfFGDpmNURxJMr/wGXhGv33/FS8ujJVx6
kR1F2d9Z5HkyNf3DmYORdTVChIYx27nfZQ+wnVYNKXY8w+IugvLHFbE2SgGFKl2Y
YL0JisglMCW1HAuOLNUyIwej1++k/srdZjJdR/7K+5ljIo5Vjb944vZtvAJgHHhp
FCJN28MNLivYj9BQyx5fN/zm1F7BrIzlv0gwoOR03eeBbYqSe4GKImacDe1C84AR
l4quViBc7yxf+RY2OhWhfSBztkTMFPS4JxQ8LOoIEJuAubyh6RO47heOmXhbIB4K
LqFKIalyg6I4aJR3LdUaJvBHogh3sPMExotpR+oSIdiUxK7cjaSRruEbu+u5Kucx
g96GLWbLOvLJCQGYdNOWqEj+ok5+sovAVEzsbwIZmRzt9YhPSxRGuFHKGgzUcZwa
7Zw3bRknTKrQ2/itqYz32OkpCRSBV/9AOarKieJIxxFcNY6Vy3o0IecIpjqKvFFw
DWWF/NIbPFH8pauCz1VDzjdPgOfDpMjlPlvN/sQvQApkakXsiAYNEzVH6wkuAYDb
1VluESR3ylaYoGOxo8qmR6ZJ8Q8fvXAcAhUThNKYTPnnl8lcOL1AtKArAaoaccvO
EIpgiqFwCJNe+t910jcX0V89Gjm/0S6MG8SjFEP5dbYGfFL/pTGYNKLRUl9O6Ukm
JLWqrLQ40jJnmp94+/CjZg6rzVEX4W3DTN+ZHI/tLjos5Wzwq/ZYN0QTmGpBB7Ot
HUpXSvsRzge99KC5BjYAr7RgHR2nDWBLK6vy38dkKYhq66t8KBDxWyDLXoy5u4Js
LFRu9eGWahKfZABkyiARShZzUYSZRV8MxKcc7u4YlT14qLpHRqP+Ma8/kayinDMO
LAOSaDMaE4RoHYXcA/BtcmoIKTDDpP1V8vVfC7oJM+ZUpg8TCbgile35PuxPTMS6
aK881UWx13Gc5BX0TMMktYjJNDkYUWmnTV70drxMd9fJ3hEAN7/QjU5/bg6cpwC4
uU0KY+g5EeiQkUmNQX7slHskuUrZXmrITxAXTtkPkja92qGE6hyOmzZ4Pt1a4yhT
9MlSihmIL23SL3jl21akHZT8NHhweYdkVr+5lxz2MedIk2FTHARppM5KCb2FEIkN
Jo1K9cXXPm2Uyl6g377/RpEt0XgYPWEz3hezENeylgXkdbWRW78R1M7bau1yjbbj
PUl2PiOrez1XIOT/2Gdg5pdbX+YE668Sy7DhRxN7coUcZMFmyvVCW5odUMWZRZJ1
CvQf1Bb+Qf3sY6cMxs1/f2MBc1xYxaHzykeM34wnQFMnXPCwW49R223oRqggMPKW
DQSh6fjC/NJMNkW82a0Pq7W8eAcM2pj0WnL4asdnTKeGLZ9x36Def6W1LwX79gyf
4uYRhnZngJmDf3UZM4B7G6wr2lQ27pq4Anxjjy3VTihC/PYVN2SIpbh7YOKWlDgv
+tGyrZ5xtaRn6PyQOlz7B0HzeldkzEh6/hxauCa24GCgYIMRtSNSCdaJpmyVabC5
LsiYL5HQqo3PJldDMOOFdZ9JgC6lyAGO7oIZeU+UXEPIdFqtuSu0eAdrpnPkL12q
UwWq/YrCO49j1lh7PGkZodO2i7501CKm6U85DO8aRrlRJh9Re8Hi1sS/T5MCp3sY
8FqRBfsiLIzYSF88vbWRL9JBWqxhgal3LGlk26FpE/plI4B7lZIMIZ6dgUxxYSzU
LtdLUT1PlGwHKK62zUL4rGk0xDgBD8Looah2Am+Ern2YyeFEa24Wwi/Wh4TlVeB1
Yq6jigy/ZkzGOPu+ISa8OSuS8ab6DI/cLsB85MGP+w4r34rl9FhFtSzaV/79cO01
d6C6D+4+x6lD7w0XPwuL72aydVRk3NxSSTRIpTSt1KLje3M7Ed7ysg/nS2CsOD9D
3oaQQdbwSYM8VSXpQycaA/UtG6nJshfFkjeVKlMwmtz7sJyLINksD5PJ3bKnuthk
ej4k8EcfH+BE1tcfTmgjj5GBz+PvBa0uyrpCxW8JUw/fdV/jMX5JCBsGjVTsnnKt
5TSIRo01LY0vDF6//ymBKL6Uy/IooQ7norkaXxZ/DACZWaXAwC9KmHf73HbzIfqi
JywX0eint9L+tmmPTYoVmoNjnPLCGvS8/OKkg1H0HDVzTXK9p6yOnBgz5JLVTMPD
bGn2lJJDB4ASC56eXlZKoLdCVqjSNWSLRc6AYGVDvL10RF2svgDt3TABXogWKnio
YVbRaTX08yUfLG0F5oWdR00Z8ZihobYnhH8n58ZFch1PSPv9vwTQvfHHJErrPTo2
u3R8mnYXJWcmbaPkHLFE8JVHAXB8plSMiyLOzFFLB+zPx52xNeZl7ysLOQv/RroA
AWLdyZ2cZHSM+nTV/Kt1VrzM/Ez1L+LLo8WhP7FhNorbhdVngTaEau3v5AyIGQEy
RgxpQfVSAj7AEJJNSjLXWqUArl0ixq1epoo0QetbNn0HMjZdN+3lIkgUDkEoxTWS
ZIWIrDorzg9A0FZaQMY6KEePDjFYquf36PXPFSm0MtXwXHtc+F0BXBIQv7o+0EWs
Suo+FHHyduofjQZNeeM1alIKgu82WM+H7UGnwYPTGkkkvP4581WDyNmKVGObsjEt
tO4FpFMR+A/7913XfRxDRk4ngFmg6keVxVBW5AQWizstp5SRtDaYv84/ISHtWrCr
DFBJ12E8IiV6WoHuxAzDK3NULiw67VXy0vLHi5SeuUyXFqQuvyU2K0z0go9KHnCP
cxQwlKB1/2kFCFHo61q4qlRy9ThTIM+VXJlz34wvqtlWmhwdgOVfhmfbh8TCoqzh
SuiqVCn4BdbNdYaVcFiFGE6/wWVM97vUNAbavnRh5g3MwrSzwHAEaSdf2fto/B5K
0nV2bUqbHRcPCXI5XmiB9vuPSGd6+r5Q+CWE6wIU4odl2plK+wLdyB+nSdHqsFXN
Uu3LQHXkFx8c5DGkuLiYyHLhQC4qf7Npq2PfwzFoTVR5YxIGkpybXS8kk6YoGPeZ
bFSa4Vno3TUGsDqH89OEdP/tw+Y9nqsuZ+/lnMfZYwhd9Ku2+T0QTQXV0bnn1sUW
AgSSURwIAKbQB74UM3ExhF+VkA+DlIZ7E3PoTxdBZuuShFp9fABVqUwtM080ygWI
p2ho5Ciy8XWnLg6pPTUH0N+kzRShwYwzBo5TfFvHT6tenzYYvzZSLHOlF2tpiY6A
HFrUid/EQjQ4vcxuDhaUlsAEXEoPDJjzD1jHzzRBqbUAmjwZXsooLwNp1qQDxukI
fcgHFklpoBtWaNzMFdn3hm6a1rUzDIrOniMBtFuH5eoO7QY7djHFbDwXFqLCvJgc
9lzl14NLkV7UpeKeYSrATrfStVReIqVDIdDy5bkSFQaJz+X4gdie7548SrllHzme
222pxRsYBNkjJn64N1z1VJE6Ec68dAbdybynuJFBv124PZzYFk1gWh43Fal6D3W+
RWcTsR8Bj/l+omWPslu6kwLrBkmb5cR6VEQnfMLKPxjZ3lcuaHbMwPYFvI8sb2wl
3EseylyWbD/nLBOQKN/kYHdpNQtN63FVxXyCkspDyrL4ENW548OvYfbVUNJzHKXF
9EmQGX9JwGdYJFlH+I9WQkuA4SAFWV6tprTYwT9guBBq3C7BwwTducp5QuMOvAMg
z3RWIbuPWLHg+C5NieTootVgom/F4uZe95PMJCIv9qcdJtFk9lpuAsVINY78XqHi
8zgNqWEax7kBr3WkpbjDslEQyOZNgUl0xnW68ThnVQ424gLNIkzIVBa7arSC+eeD
S466hYs8wVpfJc6r4UliSiQwBe9s/BOsx5n/lQ8UQMbcwQlEE5QJQ9nlTifbsK75
N2njOijd/aVRvVWNorws4Zj8ojBF4ZVnSd/MxjUWuhSBhnwdJRxVvkyBR4lXzaQU
2iByIG7WmvjBVy6nD73dGEcC0F4c65yvgEgjIMz+SI1tc1Vfue0boJSFvC0RVwWx
ORam7F/9Tup5qiOF9TTsEVoNBGxvgpC0zzRTciSRmQQIp56H0v84t8wOgGKMYKtq
12BpsHGs9DUJquMK+ngIgXCh3wlF8RMwTYnGwUPbzXV3k+IdCcmsOR/eIWz7Irwg
ql5+jDRTBgwyT15W9rzb2MVwJheNFk0XtAr1umZFbsoDUExT3K7h2bmjyvjQz1Sp
cEVIWLhbffXitoVve3vghpwYjTSlEbOzdVUk+qEAt1vCfnO7AwKsfKxk3xExDFKO
LVB5dI6CiZo+D1nbLoE7Jg4DOOCDd51XjQEHm/a1zTu+udKCenL2k1W9Y+kHjI0h
MKDWKrfz9TplkxbrFYaLOb4a8vqPXoummOMl2CKPrqCqYtKJRgfKNrr6m7fYNy2K
Sc/bINm1PS685+eipSiT+NvZg1vUoclPhT6DjLXP992d/fU5U8Bgtwr5ZsMH4x/6
63tyRPVyxUxOksfD9OY7NrahLos/0iymLw4BYdtzp8UTlrp8QPX534xOBsZbUAlT
joBe5HJMYrfVxFZx0/XAIaV6pQcg0nGy0/OOlDlwEH5yeUSz2ro0t4b/6wsdaRub
bkPlO9xD0MtHpX0SlGRG+FMqlwBd6gCwKpp3IQ3M73QI9LGOSUD/E8TZOa1YFKqd
5IFBpqtsSYTfpgDkiZW2KeLFUSurC/yzI1e9dAw4p/bRs77doS6ZqK9AeZg0RZbT
ndLjO+sYiqzovAN+cnsqLJnkG+twPPonE9ambW0mvNghbTYkw1hlJGiLSvdczUYS
mA1K7CUF++mBoCgFEeaZemRoEsmbh8hp+YGvsMLTs1CU/Z38+028qtuMegMyAFza
eF4erzxLdVbtiXFxztXuNaanVHWvWT2A49Ls0BrTc168kgweoZrMNuH7wT2mhWtP
pMfqleXA2n5xrFBitc3cfIa+vmsCaFOS2u/EdSnjdy0mkrQRI0oTY25TjLupfKkc
dZrmuvdYoJdx9viOV++6l5X5g+HWTNxs8Vx4+OBJPIt+6cokxN1FC/29mf2kHVLK
SvMkq6apjKeW7pgUATbniTQXn3FzU8jSzJO4azK1StrTCnBuTcK2g2KlkU3B26w+
cuQw/MjblGRkUkMBH7kHDO3nDpsG2ylQcWIk8FsFiGuJZR0ROybfOEA4LtDQswfM
6vUZCDzQeFDlgQqoi8CsTb/txp41NdXOF8rVADL2SPwph/Jw5svji7zJdqjRXQqi
HKduqc/H20968rPQe+nd/kWuKFUu+DtNpvcXKUuSdqlFDvalbUUdGJKbvJfwRvH5
RPg2HiJgsl4vRyv7pLn0X5/GCsSl/VOw1ZLaal3brMpZ4Siu6r7l5pQSiFlowtHp
KNqPgbIe/lYxV1WSMJt9mX+Lt6ypIYaG+mzDHHQP5IjJAP96eUa+ezVSQ01nGHfd
VyRtppQ8Q5ny+cbWVGh9+1vHuOcPhHzWBixSdPAOpz+DOyZj8epPwAYQUsiVUetW
FrwabGS9S9uUJNdcvapMR/VB/K6Gk+WuKeDqoYVUrqIl5qt46ycRaBYlWWhpzmkR
nKnaAb/aYQUaxI0jkoenaCRRXDyWQhR7ksuy0AFLMVILbgMbxUPreuu++axXBaJ/
RYjvq50r1ifiksCD5ls4urzpbqee94Ui8jyxGRjAaWyn0Kyu04SiBxfjv6+l0dJE
EIq3KoO+95MkTMtxjtqXh8Bi1sg9orsDkFTEqWdcYlxC0M7RKuGl5NhbbyRheasF
RVGsOsCzT4sfdAiq3lGffw3HH7TEQ1bladSPIwPwLjrRai5SkEayr++QlSW56QAa
GLVSFPF1YdRF4w04cMFCImv0ThPOqaW0JMwajE7U4QJhqdbeNDngXAn4+Hy7HhX6
QAT15CLZDY9h7G+/KM2AOP2ZkcfTAy3Mx+fugxMQ68xWladdiZhPxN4asOVCQ2IW
pNehLiUq55ODmavspL9xldMYQgsTHSmOV646XgjFAA3yGsQmkcSP2rFerWB8A4dh
X4E2TyHv2lfmd0UUAH4UsckKDEAZL4LbtxprkCw2C7aspXhIM6AKsFxqWb17x/+z
mJfkHUOSwWCUQhUCk9s4U8eBr+nLCZZbxV3GfBnYXGX5Ubc8Xq5fpf/PA4q19zZY
/lhPuF5WonI5SFc/xfDvHRvcsFQCM9DH3sXO7bJOzRT9EnJ3zufcYU9a6RjpYFlG
Lex0/j0OykNRzHIo1DwfB74tT31H5+ReqY6Dc4xiLlII7tNlGydZZjgUH0dT98lv
CGlKRbmDdKI89F9VFn7bB39MhUwlYdHJyUOVL6UnRj9B9c2XGIW+v825Vd9w9a71
lMxUpbt+OByhde46PL6CQIDq9SojTwDS8n/UbXd0Tbt0U6REcGHWg7ykfVVhvtD0
bpfZZ8nyZ8tQI7aGW+3PJWxq4zjRr9tn5adh9GofikrmXz3ISU/7768WXcRqV6eF
QlAKrS5e3S6mkRFDTCRmVS+EN9P5hBlgMJj/kBkDmijWxH0jbSiGRaPzhhQEm77a
KR9nDunbn7nGdKvkKy1e4CIdhw5l2qLC7zCbJO0luZi8cboWUvD5c5/SPsbPEIck
kuSuM7MBLD9AEIIZQrOjvPetpEYW/HgeLjemDsV9GIqxsf0ATOR+Y9bqiugaRW0E
0nVFCuhpc3hk62vkVqOOsY2wjHPHuSth+NCgbMksVJYeTkzh1pZUohOA/GTfGfbE
mewf2X9CiVmy9UW1gd88asXRcfnNwUjeLOI1xSsUoN6tYI1TOWmD15x3bqCWahBu
AxtbtuV1o6azLrplv8ITs/fD31twn9X5gTlHnY0F5sT5uvMT+GScEEAQJir47m8s
evi+KY/CiuS+f+fqUv5OcDkG3c39MR5KVlYEKZObddXEuo//f9MdsO4fuhCzcV+S
xyvuskz6yWerrwBLmZ/N1/7sgEn2YZgix8PU3z8C+hDZQuxLx5P7ExMiEo1SmoWu
hgOnjPb9oQvB8/dBbZq+a6JhyOy2jXrX6kSfg7hO8uH4U576LO2Bw6jvqh64jsGC
3ztG1FIyILVFGoiNm8F0ZIN+FIE8+trzkW5LVxL5xM70DQD0W7wJFdfFRlhoJelK
4AAnalEc2oPgNB097JtCpcxSa1LPBf1yy0xhS2WX3q884z581SyTkUx0XzetFqiX
/hH/ryr6tZZHZU6kwEraDjh2WLWm1fg2T3YFWvzVU5SxmHc+FF0yhE3DYkb9GYnA
TqQA0uNmRNlvGAvHGPjxd1woZ87y2pTZQjZ4+XnFj+1wcgEYURjufEOkMJr53sO4
PhgybT1jXtW5rq3hzoxKd28MOS59HeUFKwehXADDu74a3icM12C7L1fgCR1lCpTO
T/d65/lvO+ct0wPjCW6bZ5Pc3SKvB8HVpz+aus5jrGP/zKj0JhcmzGBYYwrS7IAK
t1DSvA1RznBB/9S/pvFoJ6Hc/V6ssO2+e4UZ++tfGKz8SuQby2qlyQeAch6EWde3
ITq6eDMpmRPDJb8yIt9PVnedpUKJsHyc3X2kHiAU6UW1kHQCiGykU88Tg8Y6RplW
U9llb+dNO5C3C3/zZyxhcz/4F2NqQOiGgQuO0ejuzc9DQhC5BIF74pau8HRvQyGN
+0nPOi62VN7SOlQfAH+nyQNicWUXUbnhsaM4rlIKMPLNXQd06pA3G8PifwtyirTY
is2TyVzk597CDsFpRRFMNF7iYvRU8YLOVU2KHya3QleUq7ZyaF+PQxcq9qwwZQtl
XfS/iy8nHZwpa1WkEATlxzqWNoqnLi3CDqPD/f4l1goZ4VMMz2G1RMixf3bbw7CO
b9hW4B3AVsndxcaWZFx8zmnwOLg28lVDAVnuJh7QBlBP3P310xR+Oy+n88swSS6l
8KJi+pe0sGQJrYvW3AiyI69yRuYk8KryE51ToH1CQnWcsGUV4POeUelUsThPOYk6
c6oTge67zU04Dczg/5wPmq2xonhRlfJUMmwW/QuDVsPLkeWiwsJ5IQx+zCYkfqVI
3tBV3biphFM83LOlwQClcU/57zOJZC46V67aMSGXEQF0iG2MeUVdDzwXMYKv0Gwc
PObqCeMz9+j/v1EwpNeSUdEtYLpdjNjy9Fxz3F+sacTMD1V6fDnGnyOnfN1tcx2V
mkcU6o+Qa/kU2zlYB/vUpg7Xqgk7gJYREuQe2bHL85fwZDVzJLyojZGo68Tty7pH
7fxxOxLy2HUYdw5qgRUeMK2wA6uRWFuLlQ0dmcBmkUyIRpb8fMfWL/5v2A91TfLV
lHR4xYGLbJyrmPDzex+0eFvNokD7WoQR44aVRB3CS8r9vX2LAhW8w+xVsLPYpIdi
o84DkSHOWgYnbz7nX7XLNBpNUTp0Ui3+lvgMF52GseLAb//YRxDRICnBtQlR3i07
cAhYBr2JWqMcfgQCZThKrqT0b6TNFyNx9K7RQ9o10ptKzrNGCbwTcumpVOKIQ3do
XQnNfSooplvgcnvtnfhHaC1UPFbvEKDXYGeRqrJkiC2MR9xAvcx6NqQC9mSCvMxw
0KbfcIk6wKi0Gujbe2cqrW46kDjdJgb8c2Ycmeg1NUnNYlYekFzNJ2xnMcwsMjnC
6xHVBI65T1IIhx6WTvqtjk6LbyKDfL+TOL/PzancgHgv7NW3uhMPwt1H/6Efu2Km
j3eC+GeFKIsOjYGlBKaqlQXAA+6QK7ILUeKOmgVTFQk9STqurU9bbPg0DTkvJh3k
kZQaARDpGR0EzBNttp5zCwTMcSX7JxPVmmdvFZ4DgAmSiFuRSGO3WCWZUxcFf2cO
rD2vim6wfkVlYXU9TY9CZXq/szZaFAMcjcY3bH732eM9RTX2fa44ZkecaUut6aaS
YUVpqfXYC7zpJqLWxbAqhdAvUEnYKkWE0kLvAEN/hr911V5PvwyAMPCnJcSzYckh
lJ5GXI5/iydFyITHqZam31JxA/NI12YjGukHiB4PMPSDtJktLyM8qLfp6hVLC9KK
okqxJgQm9tL3G4JqNMdd5fOGdKVrePg7Q2S6GOZ0I77ulMAd2AnqZzPb1j/CDhLR
3xxax0A1hteYTEWdfuwTfWxYXbFhuSm+wSvHXaJWkwXyLbJJ/Utj6QT5gEzOQ0A3
bfo3yV7uSV4+C9vdvnbd5db+S3h4Q8yUkwwJvrFI+qOcw8QbNPemhhmDUO320533
BAuPpJ+7asZR54Vi+vAB1l6L5dMzRIeRgnzRbpoYCBGMgOzmcwCiwKh/cKXrVkzV
bm5x/ZGCqYbSetRw+DTNb3NSBm9Ki/tPVXBm6haKPXeHMJaO2zIvluPEzXws2h6R
/1j206r2tg/xia1Tb0xXzT5MDfUT+Id+vOwuPNFxFlgH/YN3LpG6ziKnv17747hH
lwUki7S3o6ZLnqrRsNpwSjAqlXAbJWL87hCEitKzPXdLQVHZYjleEcA3+ypTHRnf
E+Jq1xT5SnUt60wim4EXqzl6HzMFmOF6gMYepgObvlaTeO1LqQIAmmEcCNxy3BB8
x0K0Iuan7vWja+NDovjjQOraAvfcU39P2isVDTbc+/rCdm/r64zrBWySeS9i6qq6
6z+lwQ4ntGrc/e4v2QfyBK1sB5zrJfwy1Vs6d8OI90MBsg6V4UBxLAb5gLw2ni9F
0jWFkeK4imPOFCjgBvBQe6D82ItR0v8f/nbSzN7IYknlt/lpA/yRDlPn9WNJ91By
Fi3CHphpD0LZHGrtt4MUT2gH0KQ3aIaw7Ob1s03/xhuKwCVw5JKIsYBXegg63GcN
4CBxwvm+9afMUhA6L1FxegTzEXHuoMx47T6Gs2iQUW8P/D/J+SoDqZE1q2cKJ5wj
cJBRh1tA1n8iMeHPYVC9Eu7lxZpBrG1AO7QVyyXXprHIesJK929+LNbU3wpdzHcE
6olIQTe73qtzxAEC8tyaXB1Z9cAf77dxy/tMvh9lB2GvUJ5RDOPqUjQKsABR7Xw8
H6SJps7qfN3UwZXo5GHN84+LbdxBZHQ8M4zkah92ypHIHP3e607WcDEG8eVbR2df
ym7FuJ3CqDm6jx19V9YSMk095JPblScS/ko8dvacMlL73itTvqbI13oBC3gk3QbV
B3CMTZ/fDTY9SdipV5mCmCZjjWgkWkGN1RUzVLu4v2V2P38D+kg1XEg4MwhZNlr0
o5E6OoX7rhnCfcbCN/pTNZB8X9R+ms2WZvMENlN+fW3KuXbzalvxCrsNw9buo+4P
klxv37+cOvYSXVWLVHupA0DSk/ivHJOghubGE5GlQtZ1XxF4ZEY75P0JkflykeJi
bF6K205enJ4Ic35nPyRr6VL1ADykl/AH+lm42id0OqwXQ9nyR+q05JNfvQzU745y
/xDAxfpJE+EFVUHsCgch3JKkWt732JqK0yobD60i96cqgZ3eH3hhTkGg89iwgRPm
Yr9Qa/i7cA2cqHLeB2hr7TcYQEjoIAhmsTvgsGgmJEP6zzCldDfmP9ckEZtjxWEg
0AarZmlY9uW3cl1MSVktCDvVr3pb99TaXGkoiNCQxSRp7RybA+s86sV5dxGD8+j1
U4/mo2vVuOs5Q7j2YOXnv6cOb+9Ic7dadSnrpmuCX1QZiXpyGz5bYQ1JT2Bl1+71
3gzsEP3nKybO/EFEF+fZnqNLXmMedLr5Hw1hX9f25y55tLbLrsuFwnCO88aGBVVF
ISvRO7NF8Ltmf/xhBvIyuAJJFOAAWXDCf/WmszeQVFk4OfYiwnshLiXSPJ05RJvX
h6p/vbMS0KwYpXs6n5n0IRpKIUueBgGUZvksAZpaKuELdurXDyIwlYZLoNrwmZfD
GxE3PUw0awpduKRanRKjZ20IfP8bbCDY6teM+w/R31hpilqbyGfjpoD9uVxEK8TE
XgGzqxNqV9BFoiDylKwbd+cbufB8rwUc6ApoZ1EXMOSG42SXV2qboNlC5x9HYAs/
qGMLgS7MQt8Oq8HENfCA47UJChCFRFQffkPjgr/yiRWdTg7zKU+YtJTKyQGLLRGj
tWfLoaUwEPs0wEDdRKGsAJFAIGh21nnzSgPJCgTUCF6ldtIm3NeErMhLsN+k6Rfp
37sO3YugZEyPQVwEMBIRBwY0F7KtUoUuha6WNhc/zQSL1k8+wGHA3ubHyKx2dHxl
DNby+OHEp9MOMlZUS8e7wSKwy+UyDLTlFUW5xk694O/oAUB7IYnt2jvif2+ezxO3
ihVfFwQ6a8sFIA63Md0NMiaw0wj9Bu+LkOyeNyAEtyRTBV2Bn3c1+oNj7LFa5ILa
1BVTIO6vg6HRFIjsLHYvW/89SvEfa8P2Q5GYETUnQy+TBcRptuHMpH1tTJ1o8N3i
v7Q5/9JC3dNCIWp9JufPywys/vSE4zQIkwjm1WbSHuMRljUbh9SI5Odv2NpT20HX
gguDTt3nb0Xelfx9DgZs2zlWasEsNCN2Z5NQK3Eip3rzoXxATK0/fm9Sz2YbOTbd
e4/ZJB7LBikv+b9XSL+GqMyJ6r5igysZMLqaFzcUvUk+SKFiGEsdXmkv5PvaQdzj
AM2ha7T+Z+vTZHRb4bGSRMHP5wfVQzB3lMxBr7kIxkKPy5wpxT/BxoXhYCPf4dyB
8wfsAcNQQ6SlZBaZIR0HEQ1wp+gFV2jVlmUlcZ9jZaInJ5wfXjYa2VpZ1RnFIBey
l0envo5BV10XuQdfioSwej1DwcTbMwExEb5Z9QjrHYv3ONQQ2erp5hCphw/Pgkev
XA9SD7xrV6k/6mqhyT/5FI3kM0ZxzZ3SJJIShIuiYF/LZWk/cxR3CAKa/peuRItD
18JKsV2nrU8uI+iVwgH2iHY1943yf+lrQd78YSZ71sBMcMbGQgZEmhkP7D/NEK/O
mijfNE1jbRkxppv5zckalE1mnbViTO4pxSIoLYXZNAvS6KNx+xlB2vh5VQ1jVEGw
xzRVr8rdJYFKOiQQP+KjNBB+81VlTEPYH/BREnKcd1YIN5uiL+kYRkAYw4U7kMdx
h+2hSyDLldrvDyego8D7jkovUzfsSOkt1mYSCuyo48HNF1GZi2KgyvYsQWFi5fkq
sIFf3ieCfSMouJPtTRCsbHkn5DJ+8E/znwdXl/lCzWLHavVWvLkn9WIIlzfnT6XG
gH6j6Dg0BZJfmPM3yw7qpCp+/8+CdMxBpdw1IP8LSIDf7vaniAyfpTs7meaiEbZ3
73EO9zx4BhBnzA1UQwL8sNHOKXaM7VYkEviJyf/O2+N+PEIMf386wDtxpkdbiEs2
I4eduerzPo/AiCw+nNnFgGG7FH5WoQmRDYqdIzfDFcz4dV3+x7XvAiawKBofn1aO
LAiy4ehDLidhBJhZqnU3InG1W3bIOyrAvJ5KykAbwCgN6rDYPVYeCpx/vjZwNhdp
LuPMEt3CKe9ti4wXpryO7ZEZwtAgWX0LoEmR+eOBGbFfN+momqBlaZT4ZNXx3eco
1cAGCctNvI9Mx2vtbeBgiq/eYt0Sbv0sFjo0Zh8Yb3XragrYL30/kbJz3E/Csb2g
/HBUSVt+qOw5YnM1cUx0ND4WXejzBA1w1xq7jSzQE4T6sLlGllaaTtusI9ZocyDH
+ucSyn5qQhL/9BR5Q1Rir1D7buzxMe4zklhvmepJy/WQXbOopHOTA+jN28wb8+4x
WxqCtGy+zDhjf7no5AjEuTalLMd62IMaBR+tKb1XLZaftGWkeVGHq19pkLvYv8lr
rHLJAh+1f47Gi+qnqsm7roKFpYpDPuKs2SimB7cCZoHQSR7fl1tik4TdvGzygqeT
eZ0xXgdV+ebcO/7JJkpX/y2A1nqrG4SwCEPN5RYTg1ofIEXHPvzw90tGw9o0INgx
mAP8sb47cJJOHgQDUobpiJp+ngGTOgEin7GapfZ3ZeTUD0fiwdXjJNM2zfvdpDrO
4Lhcg6rFXFIM9djcGxjjHOAS+92Drb9IqBIVQ8O7xEe7plzw9BVr2B6NAGwuCI3V
+PIUTxWjZ3EsgzTNu8CamLmHyINM8iJ2mLjai/Oj2PS2hH2hQUa2/ng5W5mxHSkI
j4Yca/GV+yqHGeWuBkdbOZJTBkP/WekD8zsPbIGMljPoF6pcYyZnpf4kADlAkkts
Q9ZrqVD1LCYzT0wYPlM1WjeoCXjGPZhviMMe/fIy6n1p6mzeCZJ8uMlAlfgd+Bjw
gwVwr8ug6TEjWnIZDTB0ovWkmhgwKrcTimNXKZzrDaygAU5XHEEeggcmQesnj0Vj
KFMZAJ8Qn6Bsx2O5LKC1BElwlGmF3aAwBiJO7Ffmz9jwLGonoTRt5WS4Phv+Q2uK
TkL0OSen+IPAq/fjkoKbxhF+9H7RRUXCz9k2EEbHrFTWQLFQejPQaIxL37I7VVyo
vYLSNJqM3apBbfgjAvWK5HvuT9bE255tVbjbBavW8NqTb46LQh3+XX15AnrCwWg2
zFR8lXVYqCzCCtL8G9HrDMx12Yz3VYmpRvdGhwQn6nCWWGzqCOewwZPnJwa4mGrt
HxNYTXEVqtN4GOE81D5UJQnyha1aZSUJyhJuZxuM4KHLmb03oMGnzsgN33gVXKxa
J53CGYar0LM6tbUtzX+o4Wbc2jG5O8GOVkLuvztdrwE08DZ38C5m8MVx/WgQdH7N
uQ5qF/Q7GNsHHqI9NN1U4NtvWxcHe9QXXd7EwkTmq4dl4GfM8k7SCt3sTRX5U9Kl
dKyI6BtEkPD5m3sSsPyox1KFUE5ArH+vv0d4yhz8PibR3HlDJL1vhwTfh5qAeCWT
M/0L4/6lHQzTBYRUcqySDwkhpn3JJUCIYC5UdO7zjWKkah2Ic854iNSqOnFkrfd8
byoLsI+u0ChkvVTv3Zn44282FCyIivo4/9C0kSph91QJ1PF126iSBv2K10buKZfC
k/OXAyWqhogQAXiYNYym1m71cxRm3MyyHYZltRv5uVAnnN6//iDSr+T5+1tKFSBC
oxPAIXO9eAyT71GFso0CR5br8ppWcqdwYWQ1BaKfHRRHrJuPkzRNAQZbURK1+Vt+
Pd0JJoUw15B1/nhaMkiA4fX5caOKyGetO8/wc40GRo6hkgeu0YQroMY5JyDfqrJ/
zmV0tXkZu9YX7k2loVvMrs9/fELAox1fu/hUoVujTOo3SGcFgs1jv+T+AlODvlVk
JpvXiqFGIj4jvPMHOeQGEKstyZtH78by8gYM4T92vvoCMqhmTWfaE7XTbrHbV92K
xc0rvwHNgbjKLoMN8mhj3J2BThgiyVbhKpvh8mkAPJu2PAELG5wioTYsXFu6/aLu
uDLnWP9lDpOxoRDGOWW92lxy3GexvTkSfkZiFH2jHDJCZoZ5me97/n69DAvxEnSN
1R9nt0Qy8kpd/bK4CKeQyo94KmenJGqEoGNQB33YIav3N3+ANNYQCC9x77rs3Iav
uUbHro+IPsC499PLXJUjDPSBmWfRmQIlkQIlfT35pZC8t/soL9gEg59bbTezkrN1
QAYrgUuobjd4N5ZRe92LuCBbPp7RtU1k/BbmKkcyEZUAEpvvlkeHxDLhdXkbFdGJ
Ygk6ZS7NWQSffQFJoYjZ+XssCu3i5IU5Tdq6RTBvVJMwO84Exbm/KDTzSv1TS6ot
4BchOBJk8g3waDBDOgA4YO0LYxlObyR97At+aRtMr+RSgxQXeQPqH5/hXdlNqZfq
9gk24emV6dUjEK7WBg+ggbWApj5FhI3i7HF81cyNExgrQPKrbEHv0gK6r41SSUW7
kxH9fkEaSlsINus33dYVXPxoJxCmUeNiwchv73w+Y/U39xq93D+jGwgwtMfZGzmY
IN8PuVlLxRHTKWvWx2QFjE0kFqi8H/2GAmArHCx6YBv70L2TPI+AMzSKDcAXQJAp
DbL1RcJkk7pK0umPFh+TQyRthuLQ4s1fmRZXvHZPPLy0klhRry0+ckLOhBvRjXJZ
f5XAvyFpAeTiaFhU7sTIwssqAMEd4fDU+CMzWUvJ5bK+zvv3ieAPXFudL9CxEAjk
cV8rpfiFvLj5fd/xwQO9m+4cyHkrAduEw1Qs8Pf1pA3eDCR0iH6IKnV/5wvmpRs0
rQWdgxQ1u5RTuh03MrENtu0wTb24tL7TOQq5OUsn0eVBTKIElwESSIbnLaklHegT
7q3eyd9H+AiAJ+ytrzNbIaNBb0KA3VFKI3NThH9r000gtgg/pqf20pCNP+AwsEXV
yynaegduPRBlrnrFHVVuDHlCjMWLp8oiCInxhnWKbJZz0vuH90fNmBhI3d/6XBWu
ncvwWvbFNgAcXlNFlXgWsanyt3A5udzXtGKkHEUImoHGziZUKCMwZVs/LhsuX7KF
o8ld8yoE9vs8P9klI9HAAvBChOjhv/SjWn7GI0GpESZhNz33/JTx2PDD8QbTZdjN
4LKTS+vjZm6PAIBtXIqxLk1fdxAmTXHStIR0M4lL6EPtrchDe3By5sCaEw/7HxoK
MFzhOdSt+PYgqqu6LlO52bpmviT6JHKIRD3o8dEjqa6GJ9FSumsOD4wl8PZtateX
7+1p6qPsDzT/QKqqMqC7UzcLRhDT+B1eQLB0074HM+w9gMAt73n2lW4FvzP79J5X
uKfMlgeMcmzUA60BErLsmBCqKPCNVO8wG3eVUhGbbQB2zFIqYG6LWKUahxQ2aluL
g7GDfRY2IzRtcQPsXpBzeRCuLl5GTqR93Z07JXdB406A42lPJEUj7D9XzeaZOpps
La772OFtRSVkZtyG0BYMpNoIHJkHtb+rREGCiLRYTO76RvBR3ulVgOuQVmhTBmQ2
JLrr4BUNvx1SozrqHEg0B/sEF9PM8YwUtoaP4EuUbVRsEpLElXnZX2gbXHeepKGc
x0dq0wAM6aDu1+pFSZhGER8BRMqpr83s36AHX8cdT67+J19ABTLK2N8P3QpgHHZd
MnsScFpJdOTO9dMJfRiIUzqr+ItRXr3SQoMe3aJhrK6xNigyXoJqD+0J+AATZ3m1
uhxAdCR485/W0a+YXSmbcHUczgxQR7p5KVyIdA+V3u/CclFAUf4YHlj9EIxbXnsl
pnxjWzpJX/DauP3T1PXyDuEGb3ZVqW6xGhq6KyWyh+d5+VqRzYb3pUEvKgL8gP9N
28htxa882TOpUy4AfJgxDrq6CXlzP4rn7QgMfX/zHBZjAZ8x7SRTl6vAlWeUlLBN
bWjpiwxiwc9u7f+YsfYzXqLu9CBx+l/kiEvXqPUu6/xS1mykB4+NzLfzmc0gWVE+
xXg9TScdYy/NBlDEBGxHhLgxHK/dgt80lNqD9NsleJXSjm9tHPM8QBIest5rtxSL
Gznqq3fJTrXAdaFtWL/jquI1KiCxiF7kslpBbJOEoqyYAdlnmI7eYNIvEs/Jc5XH
s5yXKIEop9ltxxtegiT5fvAHG9/qwbemtMrFsd16aUXL6hQ/4HqVGEPAEqqRmNMq
zjA9aNnvr/LSLGyGpWwcE1B1KtHVYE3POaQoHBCNdYz1l/+gG3kMGTun0YcI/vXd
X+sdzqZh2PJ4qwDOLFlTbsg7y0WvND/1OdyeEKmw+qQjLZUsPdhFzIINdJPWr+4A
f+IEYHOahpIeDUNvCxhas8KFa9PWrDcLaq+jvRsNzzGh4oAQoKm0SywvSK1/gC6C
S6t9FUWM5bYr/JWldQNz+FSnCVkUMRFCCJI81btUlVeFom1wRJod/mREz/t0dnZ8
Wc2jS+8ru7bCNWG0QZD5yRIsREZqja0ze3MaMKnZp+ZpODaq0py3O3ldSZsGd4A4
0A8+5G749W7bBQREaWh7H7whXp+Fugw4zGeyGJG/6qjxShMhHK+SpalcH2NaF7Ec
YnXrjPdY93/oK0v+Mcz3H28lkG9dyYprw5ZEmq/WBBG/pCBFBE2NgwHuqss0mwql
vunkmyJR8dGUm1Xqf1YuqcASp72k+q93fYjUF1oKTy3aU+Huu3lrzq+hqA15w+Qq
1xQgsV8zQw1Oij+lVhBjB8/A2c0EPQaYzWWNYx7wB/+mriRh6s6P76sCAz+aRe4D
GHBmqC6BF/3jy8uBEkkWhm/8M3dXdcMv/wZ60wiFwYRmgzHfBtV95yGyTXZpbN4D
pkPJUJ7M8NMkmpAk8riBbKeF7qxsu/AdDX0tl99mINbCx9BGAcmPcjOGxF6A/yv3
yOtGmimAjNIzeynE1Xdx/6V2A0EMENSyyUoGktIThh8+N2VuBCCoYyIZXgKUoV4P
W4Q2cgcCVQburgxbESu3TPa+i2LqR0tO1DfgMiYCFmTHnfkogJqqty0BFTJD5amN
jayND3cURYGJ+39N7Bo3N33bcrBvTT04rCjaJO1bCQjbtf+FNXVie8JKgNdbbpzO
NWe6MJscTE1McxWjfFeU36+hCIfGy0zo9G/ld+BctVRwDX7MtsEBgY0QfiNMQRhe
wBn1D+1VXhXKouK/SsRu/9EyZ20G1/eZKJrH/YiMOW2WYg9M9trIlhfkKecq2lzU
ui2Jru12TRnNBShdcw0o9NfiiOzw0FFF5WUv/ksCBb7yrmfp74w4IrkH6Y9Xxi6T
FVfImodZiOONpwd1nIGiE63VFF8ySHNcDhT4QpPYE8fYzldS5/J5cnnx9NSoZRBH
L8Z0CdOjM8j37sczX1rgAWMCnZKHWQiM3nVbmsxPwSt9ccyQzJaiC6BQ30IYeAVK
9OtUM9GqjySRsngfSB808dCkzBwv3NMP9wXvnUemu9scbnGIAdfoaDolUhrr3JFW
I+IGFSJv7P4gyc0PEcXvgZV+kwY7u0+qooeBK0wnq4iKSNh3bL496PWrHeyBCTkD
d2dJULDgXEqfYzYA/AOt3RgqF5x6KgeisuuQgy50qwihYUl8V9WoSDqdjfh57L4j
El09yuQlF6u268l36Ibj5+5b241chAqxnD5ZU5vU8dvQfc7GFmGKrpPj2/4AU+zo
XCzlR6YYk2+RP9gTD4veeknCw2dSzW9qXO3Fx1BTDuwu0Gp5hLx8CwZfU46HXXw6
ho3bTpS9eb7OzMD0anSMbjH+bl5MgCyvPkybsaL8mjtui+AxZDgVdNelhyDVIDj/
5wESat+IwBG+C9Ts4haHywHlwqk2cZPiVXwrKwko9G271j3DVvh71y+sG07jbdDb
CHhftwYPAARoOPcbGgw01QUnexMSqWjci8ncRn3/+Ov+iYQCcYJs4mDbithFGJFh
wL4eeZG95NFcX3DLMJBJlMZHQ42ERU7tR31S5oIOmAJfTmhSLuF2whjxDH4P9+x4
avlpyG8CnmiF2J/4Imgr2+pZ/3Cpmfd/JlDqNISPUeryYN1t/D0Qw/LI9SlxaDBt
hmu6kWfwXm4A9q89SlnxBgZJHp9gsDxqpJU+ySQneB701ieIZN2ObXHHnhIjb2u/
baPc6pAAD8ms0YBurATQGjHrFr0JUEWWsR767aNboadFH7cSqi2jgx5/9BgPFlzt
76elANPgP6We04M74+9xy35Kfj1YnXeBcl/8kcCxFncrEplrngfJpwu8gT9i0EQ3
E1QWA3rQKFQ2wJ8lNtPenvVqvsTh84M0lDVYSvvW64uVN7PR3Rx8Fa0kEJJcZjC1
+JQWNeSsipaw9VKKRSN7mIJDrBufaZ3CzSB32RNxVOiGRMHgeGbwPaO6LMkdhQkZ
0j7hAYU2/Ivp3z+NWrcl4NAXLN3iAcHQSk6OvzjhP8B5NmLAnRrRTDBbanKx0e45
Psdu/lg5/EOzt1aaOvUi9tzrti9cNiWcFQa1pzHIBZDQzcGD/BQX82CCN0efa9mO
zJNh3ewc8Gc4ErKQm14nGr8muxF21zwjoin9Yr9SH8C1cxwwBQ8z/3RZ69VHnsSM
triDIdJJUWCr/bv+4VG4QNEbE9rMzDQiEoGyk2NKe7U14Z+VqG3iOAGeLepASWDf
cSS0oD0XFtlRNITTX2UWn6jw+yH/byQgJC3Q7M0XHnn7bm210tAsQrzW60TbXkAl
E6JxvH+qUqrdcgx4dVyF1Lu/HGFCv6NR4GRko5mQGSDhPyDCnDv7i7NCVhAxkloU
BsY1zFdr4tj8fjhda4iSI8kzdTUruFsWcUd5FJud1zoma3emi0D750OmKrUueCGk
KcgmalXGH1kjfCAA3ZiGYlKlZEEYMLavuKMR42TYyFyR8ZTqeEsu3FYol4vjUPcb
jfog/emF+bPFHDQvCG3R9H30xvzwGqw8LWJlcW/UuRTDVbZsOvivv30SQgDG40aT
LLoT/pAwjX0A2RmV+3VIWDVwKgpBAFImQKMUZa9N70hImEvHSY9GYC2LhAgl2af3
fjSYyjofH32N+HAip6uGrBaMbgA+59CrDWUhx8P4Fmu56SS+JhRh28ZFRjwqddgh
rFtSe3/LnOUZvjvHETvEW7fhq058X2xnTQ4TS2hawfGWzd4ElJujncp9BFP8jhAB
LPiSxx7PqV4fsDDRVeDvj45H/UsHf9Kp7/vzQ/jdWu9nwnbn8npw5rpKqEnl5ntk
QfCbZEYmAJIhCEEilpRdvbN2FfsTM4nRxFNZTtAN1kCbHDtjmBLaTj077KXLB9vA
E4L5yoaBcTYLOtpIFyEk2AQmvDF6n1uiJQIDSeVDT1zY2pa/42D2dzpUxFY1RoRs
6fUALtdP925TyzqmZ+CGKhX7Dl966PGOvKv4laHdprdYtio8nUZ0vCR7NkGbn1TS
pjg2+47zyZEQT8rCJUWNA2JwjF4+gpt6S+9jmYM69d2GQvSWW2xUtQFQfY9YDzf0
DNQJ6swajKDo7M4iwOg5enEuyxB0sU5Azk5A5o0oMcypwPP6ot8jVdz+4hf54tT4
sxGiQgYPHSh2t5KuYz3gZNqluANVgKlp/kM4l1AKH+1yyxk/iI4YCAudcqmqRlZk
xRAXkbxmt9OyyPll0+KVh7pc7De1mfN06B2o4bXr31q4gPOXdheXYPCXwdjjXJOw
/WmzzO7/Ft0if4MohPg3PEvTdDmtpoo0cXHBOa927Ykngc2Yif0jSBUc+l7kuvmo
YyhDSkHEUzBJ9XgS7+ZOEuAVmiDjjc5F8r6iNq1c0B5oGGNZCDtUS0hih2Z4AGTh
wkF0bAS6jorbzLj49vc/WaNrL7EIA+MYrGTKdKwJxYutnXJToXWPplqJj1odei5c
PmMt94hKbSZeZLENGBGsWTjrCP2vC9okTNA5a/NUGXmC6zSkhL43hgKMwhwQzRl1
0MnmByhOeP/PSk6qz4KZRwjQt4rAL9sXZptm/4qYN+EnP6iuykJbz+hmqBLVXmyM
ILwxnc+rKdz6Vx+QVIT/zmy0NCIP4M9SwwP3P6erNMYFbFxMggPNOc5QjuYJqOoq
Xhn80mokUbpwfj+hay7d589R8wnSV+VmwoYWgtN/VdTuW3LjVuzJQWjbHJ2yZzcq
X63FaLQcDVSkPLwnv72700LiEzoXjD7956GSk5WvMhONFRtBW1y8WYN2rs94EG4i
LYSnKccjDLgXPUp6k2nKvOqW4NrBw60QkAtLgw3/aVm/+F/DSvJseP2fmYo5/BxE
/n2Aktt4B3v313nwCCPVcZnrM0IojUhjsOWuc65mFfLKSD2+D/GYE/wRXSGIhjcS
uudQ7/SblH9SgmvfyFmkAOAgdm9kgj7b1nHuZcqKAeWAO1L7zxXmHg4yyRt8CwH0
QSxPzgPiAGikCec5JtSGYsrap/DHFuwMRqtCbZpG6CSyiyll0HFMAGWeCpxWdYEf
ps/kz63J4jS2GygHyz9D0AjNIDGZZ3bkKUHqFS8Kpd4UxLONs5WVubtS58xKLudu
pDJTlmMZLUzajj3AmFqjanR7i33xKX+wtKlxY5eGQJtRALWi8lWMLwAus4/QR9vG
pR9vboEI6c/hpGZHacOsmBvjPVnaZRfLoIiu0TBTDLB6n4eI/w5stPkINUWdg+93
GXFT6DlvwreH8e661kZBMATkYvu5sEOBCeNJd0vAVyDuyYOIFukR3cmA9wzRr0kF
x2MY2D7wXmt51EXlHKkMZTvN5NmrEZq6qSplBjMe/hRIIkg8n0l48xCrrPWlWc7J
JwWctw2YAO7MrTSnAqW0SfwXtOB2WLsBTH8+BpgqPCk8cIXIhWInPmkpijslzM/7
iEUvB+WSRW2NAaot6D5X/7i/tplHg58L06Zx9MTs/QUVGM9IDvj4SbYSsqDnhS02
lcent9O6js8midrUHXnTCLm2OUULBYv6xabESPgfc03mjed8ltAlvES4zPMISmdg
BCs7oWy2SIj/tyyEkSU3POsaxOnR8k437ZSN0mIh+bv10+k0Jr21uCJat7TiH8Xa
0MnK8cm6rL8PVNQMV6JqJM1KgE6wXWiI9U+CLxpRQ3HVHrWKkIS4crJYyZSf7Gz/
XUTG//DDL0HJyxB5I3lIN5ZWFgydxhCBx9Jo7y5V2byQoKKXcx52SXKzLKVptisz
qKzx3wcSed2Dn9bQAbp7fpsff2YJDna5oPPGYd2XHtUr7QA4EEvPKeCUa0mNTNAx
/0CntQeVI25YRbzmNUudle5M3Q0cW4jahkU7RayYD4mEVNkTDugl7HIOUxPaqyTR
AvUk/T2BO+Ey1KBnXzlbKYd2WOI/WnnUSj1cilWMH39g8B+MPelqHTn5FkIzVlod
eM4boStUr9WKOxRaddku8kLIZbKBQKb/Nu8jByEcgb/Jlw8TCwl5AeWRG7vwMUx3
5MEJA22ESQww3u1X7uc4eZJeIaZXkugUj+4gS73W1AgIvPchcBkJyEOTvkrVc2dG
oUthZo+R0vD3HKRjey+MSeqTleUpVTzNj2WVodtTPjgfBc04Mob76Ln4JPm+Zzft
s4SRkQwt+3d/JDiumTXYjZIkua3t8/CrA0hzmaYLhgOM76s/0J+t7LVDbMkJ5h+m
uLOybgk1udV0L/wgZ6mjY8U1YyTfH4quioRDe+leBYEQd5o06Vjz1828NSv1I4Ra
wF9EJgGVeOZ9WF3izBvg/qSGUuqVIaWWhXiNY4UbunkaAwO1fMTQEfivNHqhZZoO
4+DWy1wQPXtoNAFReQUJr6p5buLNwkZ9xVW4RXpdrS796gcTNpELHc+A7AgvibCI
HGJn9LI9DYMoLR8oGIggGbwLfxEJgsMYy5/yAU+QdZHm2oc+v3FUFIWYRnUaSZ4k
eqaLsjYLbnFxsCtr8MfGJdyOCNbUk2PASvoLNrpO3B8hf+kSVZAKx57mHAsgJssD
PeeuLsLwQCpK6YUjaak4PR7zLN6t2EVxMHFqRslHwpnSNBcqrowXHvjqbIPdV3hP
Q4xHU7RnXL+fpVcJhapO9kg8ibS80bVC9841VW91OEw1UnCIAPCNH+UcOyf5hxmj
vhn8UiW3eTOdTRqQmtiUHguGjMmLKlTNwXXpqojHdCWZ4WBdnkPqGiSSIs5CjFNq
2O9yaIfv6gIOTPbuR2UShPgfFpGVvUyO2O/hUPa4R1qC8k0dtiAeoyOZxeIqLhK7
NqDnX58iWJkGmIJtRb1Vpthzt79pbOQWnsy/9ZiccgnOW7Th2OLdR+tFPOIDS9kj
HaOhLfKORQFVdN9fephMDELecLw5c11XsnqJfV5yyRLgWlSgAKLFWvJ0xUbZr0UL
5eTJ30C+LpItk2bLIW8wpG/2NH03lXD7zdtNVdu7Ydn1hrRJhFYY5oz6TjZdoqJ6
mz0hI6rD3VX1zTcyQ4hGjkqdtxxyoAovbkPyujzrTlXKCiTe2r7MOYrwNiYctwJb
31q90ukNN4Gz9RVGaFx7VtMy8MehEV7pYnTRW2SdiDmrAWLM0M1bsJ5n0xDUEFyB
3YasKbvWZO6oXa1Zi7hQTvW905ap2uLDXPUT5nFGQTDhFcLuh+shJJ7wISH6289Z
k3ThlowT4VMH0x42/JLJa3P8HFN3JCGoCoNHnZ0hGwp6tJWcPYjRCbW8gwpdoBVn
ltnnTZD8TrnXfrZU4aAi7ScEk+kFrfCV0E8dtfborPjAhHeKMkiejrZJd/6v1yWF
Wxjugf3NWJvqHoUFV+2kFiNi8/h0cTXSHcQRGZW05GXY2nmgPLYS7jJ3gcp/GsrH
qJdgF9cIWKpXakuoA4Bw4VKvyVa9M0p/SJLQFw3G67CfYf/I5FDWaslmJnenEjkU
CZTYYwbMZZEx0yGaH9K8yoXIdeYwWdNF2hF9DgxY7/iAH2r8IjSWN3U2x8Q3q435
5CCLpsBGxrTjSSxds6PrbRn2JnwcVIhJgvr6qH+0ylNcHuQNL9MT8OMrFznDiPPm
gP/11QsGJMVNLpRnKGyRgo4V1N3xPFNXD/gae8N3VgpP+MEyxgCrftaS3Mlgy9NH
Wkj04wgbnajudX9NBjg9SRa3/gE1By9Mn920v1Jks/OjLO7CH1nHKufiF84jVqsn
g1XxHEciLQ34qf76s96Uw1wv0kgzMHPkGQHO2/d0Xs64bZC23FwL7VSQ8sCyzRQM
smxJ2NtbPoXuXxoCmlkQ96Qph1sp8FSxTd0BQHr4SFgHvZIrzc6WDRWBAlEFzrPJ
Jpf+mu4v0c/Rz/TYMZA5YOYdh1qevA5LrFmqGJfRQL9/Tw9R4L77xJPVilQXsNbC
9Ob9B5OKhs79awl430VvIyHnAVqEX7P+NVNLxnWO6hP/tLEb4eDEWmYEzpUJ0Xxr
MIWe350iZSqzWn92T+1W1Lgy/pPWiPhQ7uVkvY/ffbbk8WGB0n9DAWEIELBiYgaH
YYeVlMUCxHpVU4HSbsbEKCJupmAJ3ERxywokQXbgQIm759gY8P/Pixisa/1Mf/s7
saeMbhS8HMG1/4thVrD3WF/gVocakuj1QXaU36UKxQDhktwb5yJj9N80V1wUW3AB
b1EjwI8BDagmXkKCYpAtA8EQFRD1S+GU36N15Qgh8xIX1ZiPS4o0Yvfcc/NMX5Vu
MHTYbqwaO2ux3UVpt+X0ZUxNUjTdAqVovDQanA/yYxaH2Qga19oJcOSogdBei1gz
RKBQQ73auAphWD+NW0hrfYqu0KJXyAUufS6YmJjUtwxWHRY7DI1iuKBxWWk7E6In
OEuqurrxU9qx37AtRNAZFHvQzfzPM2cfZhxK6foiztE+9ZSVC+aXFCRh0f71lIlq
SHUJo2l3RdDWQfPS2O4s9+n8qa/mq37B8cldrO+skz5QlqPC6ae6zbCFLomM7bxQ
lNd6WWBgaWMR8tsD47sIYFdy0gZAq+2RdXFw+3Xg8gngFgUVAFJB8UlUP8vmDMNK
0GeS1qSVIbBbsSiGhoNwOPmOLkpBDlOwjclD2uj7/a1SySI2ZxQFE2B5+PtJooAT
MMaIALN6atee40Y2ZZmJuji1pNj62NEBMpXgc9caMetSzHH00Ms4rePu478ZhB4O
qDIobri3jLOFCSGt8rKlPx41aAOXb1ohM+L9iiYh3QvTRG0uNZo8Gv+yo5ePEhx2
izbQ1zbjlUZNC94+22YwjOngIES4jVjhftJhLeWJE8vXYgIz7Di+RMXicDua+I1a
YTtPmHB8iSe2H23IR45totbtv8stwPtRtlfPICpSPJLmPGvb9Zwuk/WrDSZYseCf
ye8BXwPNwPdwy1KgB1OFnEfDUtuuZLPkD6hR0UehQrC8PiD9azxIf0u2miRdJgtF
gzJWULI+X64WOzrzZJ/gVcsTtJSWe/zC5PQUaqfheJ25V8EgaFTK5eb3NCMxioFR
lXdPFo6hsimhRP8WUhBJPWv4rBo3901ZuMPb3A29bw3cseFkikxHo3gFyCzVJAtX
Exmxr8QGf1Ia+4kbc92DxQqf/NcIgtCY8gfeWTRSPhDVKj+ONYTwPejhDOl3BhZ1
9oL0P0xgSLBfu+ots+I+dsYxmnAmaqNHAQF6etYbchncd1JgxUUgl4sfRXkg6ogi
QQACnbvVQUNOpTUY9j1YjplrEwGiuSal5OBndJEaZlQMOPzjYkXZJuYtf+rfnVXT
AMeshvz9SYPIpKZyVNR/Wrvd6V+KLSbsiUV4Dy1KP5NK5biRiufctWCAaTbRe4Vn
7zMpbUK9qzSWLL9cizRf8XvePN6lkCljeGzDbTD++XqVjyIoSG2mPnNjW/Vy3J6u
Gm2nAwm5/LAue0am5XhLcuu69ikzNSEznAEky87qHQ1LOkeipfnQmNwlpKHRVq08
z1W0V7497t6zzEG/OYvDZcQkqWoAOPrugmzeD8gynaRRLjKna8+q5zlShFhtwVWk
qL0ph2sKvCpLmLJ4fkdZKfpsKsUY1PkiNpMTIRqlr6HWUCg7QVoXGR/srSdmonMT
DmKvV5+T0qC4gBggkUW0O+S423Y9XVTByF7/EvSzin59gxbKxDBcjfcKdG8SjLTc
WYvc9vzrJ2JE/0vt1DWZCBGyma2XElxiM4P+SDffpxCgrTpJ92l3ctCfQaQuIPSp
3oJU05h5X2UdpecSCO1IEzXfc5oM0AFN5z25kuQ4Fak7u5qKiVe1RbpYlDXHgkjl
b7TjJiij/xaKpQw8mLdAJZCtwtLlTh3wn6SA8w9Fnhn0YtKXRLNi3n9w2s11axGn
+VpBbuGh8shS0/zbzyVCddrXpxCo1JxnRfIsu0LaA/WTmHgMrv1LPHH8EHGvzfpX
+2zj0BuqbBdBCCFvwr2tesCZuq/keyFNucJfmCap8PeMrt+dcgKJBLwbOWsRK6ml
r4Itt6CbIW92DaEDrJ0ykjVK+nleMwPwYA/zR7OT1zcgnBpIZyKDpMfGuk388Oqy
nuGtuE5ErTM43qwQH20jyCnWeK1mY0ZjeZTkvWpbRV9fdeDjOasLZTnLTsSK01H4
VnwCGFxLKmVTFcMTgjDY+YMlxAp4NsOH1PvFG0E+vQy3wKLfD1fUvhfPQXCnkTLR
KE7JoMMiKKDC08lQ5GS5Idf0lhRGi1BKTnr4p03k9C8dJ2epDXEteMYBCtaWTZlt
v2kSWqJi53JRA5NVxDcwRLsR7OdUsa2Ob0GSh37vhIlYzqfQllFsqhUujbi62ZyK
ixuo2LtB0f/y+Q29RbAWoXWjtDilfvsVYRog4MN8a6EkVV54Fw7ToOvse9LoA8k/
Pv0e+H6uhn//UcsbhlBqZ9t2qqRTytqdydOAkCgqTy2FVCDMhJztIHdt61772Dwz
ECdyKQUo1xykHrVkvi36m2gL98StqGE1Za9NrRnKGI8rqQQrTcOLI74JiSJtd+1/
8MXNkR0GmjmHotYqbwHIxmv7SVTTYAcffl/bZ/NV0Y0xJ1HELNeJ/mgCXxZqTUct
Nf95/E6ES4Ms9il/BJ3Ax0y6ZlKXBD/XGDycFjhJwykV6d65bg1z3G1dw+IESqVy
Z6TGkafudFzg7XG3fkZTROB7hnEkJyVcJjBfBns8tVAgXcetI53U+fce8kkQ0EwA
WJdwJ/bF+bu2KuMRh3Mtwc9bsNQ+Ev1Fd0BENhdpRe+hKm+hKg6CL0o3QctT+hmq
mr1O+5zh+XAo7rkC25TkFEF4GUfV6O976Ho9wSjDEZfjXD7lzcOa/511Zfj65LBD
wGgtU/g4xPgRRRci8BTcz4lHy0DrB6/gdK029UZ4dd7H7FVqe0XVgADntVXa9/pp
M0SDFXXo00U8yCWjpBXbuJGl3kC1xphRKocE+zu/YUK1giQNTlU1gd7USTNdZUry
ZRmrhijgqwpKeBCzkdqkrQJSWDiyeu1Sl+SnT5hRgDmmF/GUi663qSIsBJ0urFeh
uo35xAyfaRkwHG1ioYatjLH0vqaqm3Go95oeEfn1Eaj9CWwQMUrrWiRdjoKYa043
vR2JTOcvL+liGSPLBPUDXpiuXuFmmOsgxZzP9x4Xtcc0+tccw2xpSHFs44g0E3Iu
qYoTJgiDmKrYgSjCKwyQtFQwKiWnBJ6n5TP4DfFEtl7g0GrQAuYZEVDvsMuZyk2G
WtFy/OjQlyoo7UhFXTNPxC/fG+LbiQIMgfnFCAeQWz+zt23n8pY2DjCixaE/hzTs
LwPWm3MyOnnr5ouA2Q/xiRZClf2H4wRwq9wEkBLeHIrdMJlkPoEcX7bo2vq1pE2K
b5gFDvKuisioY1a1Zi1sKDX4jK35ldrPxBwfYBmaOVKe1jM6J+r+VwroJHDGWZ6I
POBFhrVz1Go+Kkm88+muxBlL/GCAQgWhEt2se7zwoL05hfExkvHpCThx2ypidDMV
LePhROkUqSAgpK/FadjjDS1LS7EDJ9fLgIMdTj0owhA9qu3GFUI4SrjQKnkeN+X8
CLZxvQyMe274kg+qJntui0jBucKJelQ1jS9jb7R1NI4ghMk/pU+wcx5NreQM2ddC
zNIDBnNwwAmJgrs6aEE81l8tqRHhpsXjhdwi8dJBupigsoGnTkSbmhYfL3ymSFzr
b3+l6qvEtCdnEu1YWOcDWLgUnamo847DaPayjaSlLyFgwXJhYAX4BYibieLDTRpp
Lbcqf+dukoq0leNy9XgAdUuW3tSMEczYKAnDpAxxeheVxU9iykOD4sZJE2CRRvD/
DGjS6M40wZV795/cIoIXrMK70rS5eWLyfM+02eT27F6hvgCXDopAbSM4HNi/7IWy
QGSCKvEPvjpu17QBZGQkLux1xjDJx3efxtgayt2R66KgXFDoHqHo0FpQoNhILob4
eS0FEgnsOLiIzvjucW6RVU/GTrXnvXtJbcbyX+CiQmG3DkpH9d7iPZs3mQSxWYQB
6OuaFlBF/3IkV/obCSV8KtsRU/Bh6HWbR1WnCxB3kQb/td8Gz0ElzDdLo5LW5a2a
Ik4sc/y7Varf3uOSoG0dgCl03MsJmNIC7+dReQ6PA/zYyZy0sHRNbVOuxpW97TqJ
PMQuQCCOBx57RWZBStOZmCId+pAEI8s1dxI52SV0pbn8oUiZkMUuQiJRltdjsCCD
fkHawQ94G5PRy6e7wK9K9Gcid+2TgeNL2LMqQ5i8jJ1vWLojywuMLJF7Ts5lgsct
x2yEb/00abFvstxSLF0t/E1V/VcenyBbarMMX1wHulgVSUVShUU9yV+b6mnTlrWp
Dl8xDjMHeo9TnVKh8DerJbNQR+g0HmxUjekansBZCpggoDhT9IoYp6PLUXmqyDR5
CB8gK/Hi8huJH+U9OqaGClCqe1in9VfDy+Eud7HvoorxE6zhuGmEZhO3uEY89loe
xEFtw+nrTUN/WIdwHcd6NbRHp8z8JBKEZHL27LgESP9DJ7MglONB6T/pqnwWz1UK
ORpkocJMFJt9GAVFu24Us/mNuuh4BBrypobWCPIlm04ybvCYgk4637FJnwCcapM/
ksyngLa24aGsNAMF1GhQei5ErvZiRGUnE2Q5Gt2PSIu9R1ZXwgvr/EBpQ5YqIAud
0es8lo35NblxLImNdPL4TE3LVEMxdpCJqGHao9YbFfKWpsQ2OEqceQrfJ9PCKBes
GsTrwehXMjxp7Kwz5OP1WZdSonAo+eeUDaMIw73mhXo5/wGSdlGgmmU9sOJ8S/O2
DOe/vKKB9jI5Mcxhs+DtV9DI3c/XoIabbTvpM6BD4BkCMBhd/He6uhgfewzd32C3
EhoE8lTAw6WXXt7+5bONlxKhwTVvcqPnFRxw9GpojImDLc6kvcI09Nm5ELZUaaYs
1yfQ57sCDZUaEilKVvfvpSTqQZkmhDzEQ30I5DsdHOWjzSIb0463lAX2cD6YQ6KX
bShZUICgvwjTo2Zy+5KmYEtO5/ENeDYmjHaAJOdqHAghaZCW6B32yX5/nQvQ3Ar8
5McKhI7mpkulD1HOsF2wTt8MQcXB9eA6lgxsMdsth49c/Z0mBoGyZ+9RKWlcER5t
Osz4RibVEiqysDVla3icDUfhcihxQC+4mgPzoolaae+dQLT/LReM3WFmYN6LAEAv
OgibQe4C4c07qc/Mj6Yhl1AjY5j13tMJ3ZBxrklwb6k9e5vsw54v8ipNaDdYAWys
HD8Q+LM83kKiZQRkkeO78BO4UT3+glmziBASv2p8vTf3+HBxSKwo1LaScCHa5XrP
gAPTVIlsSLZetDMI5Gi5TCohnULgmviebOhUy9FH/4LdiHVW03WoXkyJb+HBnDtG
xWmodjZLENNhlbKdqzEhrS7vl10Zk2WZHBZrwuuLAJ7YaSgaUySCMYq7cjS9CC58
SvZrK2hh107B9kPizGBYMgjzQ8CiF1k+tKGgzkM4PzTBzudNUxDdH5kY0X2nRIqz
PxS+thMXX6Gg05gjNtpKhQ6Mk/jby55VFB5xylxFITUZZhELmQfuCWwe8HYf6DQu
TOctTvFRBuMeRCG/CSBAUW/e+znyof7s9q/zNY6zsUkPa3m2bLzGz/LFfcqqV1Ar
nH8G9YHVTtmsnhBozC28LYq+cdPQs9FKDNeLui9JHJrfpQBTGgpMbNY0Fb88mDLq
DwE3RoHUf598GWoFFotx73qBKeW4tNyj+R3OGMr/tB91dMYqnbINHKAL4mUHw1ZP
67GwmND1pHLYHQ46Fp89AvJcdxRfjJ0pvXJuzRzJrbvR/mfOs5ZUC4Q6jf0k77nk
twyTxVGm5qRaSkBVtFmyu9BtfdXN5B24lOcdvzPaiV9455J2xWlmM/3w2PZmaNgW
5mMXGgiygjIJCgZ09/UdzHlh+ObJUjEwNIcmtieSnCgU7KF1kMBQNaGAkkD2PDTU
JJaeXtqnpViqziP7EE+i1XOJh/FLa9Cnbl0nnQEbGcI9g98bNhS+woMpcn4f5qQT
OF2zbi0AasVZPS1zGDNOL9aShfRWee8qCMS3nYZA4vuCPCTAEyfxOsAjj7ni2vka
HCQdW/rM+iDbf1z/cOEV3e9RmuxPQdiNk+mog9Q89CmvSLpF6nm6uBfe87iLTi2P
d86/0+SmJVF3lxNVtUjX0TOiMvUNGaqgrcGdQLOA1W8QT0AVQCWTjo2gqbxjSK3v
+PWBGwsoH/I2gP7Y7J7R3hwJUIpiTLUuGOQi4EFaXrBiHGuARar2V3+/Bn0ClITh
48I88mP/31lU9oUefvi9Wfr9xx+ENqKxMQarEbl6j/gn0fLW2W/TIxEe8GVU1oEF
tzESBiUlnncvPNWNRllLtspHvSpv+Nae0X13v/fQY8J8r/8XIP/GAQVd21yvCi6d
594LQlb/RxEeQ7SMfGp22VYvbx/vmK9aXpPlgZA27jTl9sMp0H4xoP/D/TiWdye9
LpL2jNH/YxSxFdFkP7lIe4FOM9csuG0A8n/01Tzcg+PKSl32kuEojzW9fE3jKNZJ
5SyqAdyG3wCwEykVL2TbzC30PwIJOxa3g1hv4f2HPip9lUw9cPpDdmRDtn94Rk7S
J3c0HUnuqBOQG80Mu+q4LmwIHgG8qMoMGtjKB9WYoLydwm3ai0KxY24lOgJ/EwvU
QH2/wrl/wXumrwaurBzBZ7sLyAOFXf4wXVtqtZte4lzdU5i6IEkvltFBh+swKxV9
HlNjjHSMHc8UB19IHGT8E+CpF+EaD/YVTLSqm9zjSM10wKYpr1veBKCBrBMQ52ct
Pr2MLJyiEKf+SDr3RSjWyA7F9K1w2oAkS55hJI+X63kJCrgYaz/54l6Fs+LO26wd
QvNDB+ngpwXz5rKsgLerbUN0LvL6DmiY16ztN4PTNafj2lVAsX/dhRBHbXI3elff
WgZAWONdqlfj6LeBvtcrBDLrmZANzMi9TEJ3Mw/OGm0ZHWJvfCFIPPGJa5XoZgcz
xU68FH+Q8RoSANKAEUSqgw1m1SZHp8LmXGmN7vIGjwNMObUl32m0ONMSpvristdO
7Q5p93HFyLr6km85WQYnmb0MPa+XlhI5nKfb/+5gWYRGOdnHOyMKEaRTB8Vju6yd
vLZr30uAJBSZ3GPYihsYYFwcuYGFxsCudAj85zfcWWAcJWn0cT5PulUGoVhzRi6k
i+GrzAYamcMp1ofqKdaAdV3OInv42WD1oOO2HLUGX2GE5p43XHL5bu3itrRLNzJ8
we+NWaTR0LHP5+Kj0glm1pzFKdoz/CLNsClSgZFXmzSh6vRrYvn95OFlKqKIZ+iP
HcW7VVTaj6zTHeKv1tJByNPUe1udv6OZQi/23JGLu2GSsByUxwAee74dH33HGFuh
/sP11AozxwhT1H6jGK6Vh28WdRLPlOGz8VK7wK5VgHgiYs2FmvFuG69tmQVxLCDc
V+pkRLdR4cpibHTd8Xr6EruQyqbGzc5ZU9uEZnUFyVb8prD+gxuCabb/ZByhA+vT
x/CWhmGM38exxMKdb9h36hrtS0gP++632F1fbzKIu+3wX3VkuSm6KXhQiIdoclKK
tPyjnWr9Oi2utLQ+uXWF34C9KO5PMPitEtu2T3CS/hs7OE6Wff+C3HOv/3Bjzn8O
GGggEXa/+dS1w5SdhBIcVzqCrn2CGylz89vMY6CuoqFbATrcCuXDuM5WLN4/pK2c
t1+WQXWh53S8gvOEM/AqVIsaCVObWa4AcMSTFQN7hGsMMftrpeL8CHrIXZdRqFs7
JmZYM4fz5q+3l80FC8Cu4KLj2p7mhcGEttdyAZNsEQxE/YGOFIW2utWgCPa4zEIV
7eDk1eeyFTRR7/NXSGNB4hcAf4gE1MATXQouRDUrx75uGzOejHUaUBDI4YmmSPdB
4wImWIcnC1UfHfagB3+yWCWu+nNJssaufWcPm/rBSA5Qw0pZujVN3XBEir2dc6OY
GsDL9RBTPAl2Frqdh485nlYHTFWzHBB15qUOz7nKITGzbEwfCgmeQZkialnjwLtG
PqbvUx5MYv2DBjL2WvINee2d3Ix8P/TyE5Urx9K0YU8QcCBZuZ1ZzDiv2q5CwxEH
1R6LO1I3xBgLJQKRwxz3UXxP6q/r1Jgslo3zgL5iqREGq/MgLy8F7y3HIAl/gn1f
z7VcmCUO+/Rexm1KDneOrWu7H8AeCYo9E9tDf2JlrjF1UlrmL3y1vfxQYAKlnlOS
0N7EyZmPOW7+KxRwjtNgXLIoJaX7pGD2woxOdwPz9SLKOFHrYOKdHD7BIIpAkAlV
GaXpQjmyX1usmzlnDDysM0OEA2J21opehEsiyFPIkv/rYFxOnU3AeatTmG8Lpbzh
RUOP69DT1XQ6rmy7NE3j7bL45ZzDnq4zI0uJzo4ytM1OMI+aXDVKN5SZLmgqSIJf
3uBDA5vdLItFnqtCo0b/AjI8gnJxow7wzZTfKkfZJ1NBlD5q2jtu9snQkBKDEtha
RF+dDeWP3jj0g7R6f6oOq3Y1AuC/H24oc/6Pq2kQTgzHYB0m/AOso36wu7UO+i2O
Q5Bsfj8pnGQMQA78VKDjemt9Cdw2WiHEJ7lc+17tCG6+oYozkL+/+Q/FBPa5tayZ
O4XDsjwnGjw8mjyizI7EYKhuCN++KPfJ3Q8A1x7bl8htF3vWVSd3P2zh2qLwiTNh
R9ufAX00EfAChM2uOnPned5UV0RKxuW76xNOTAfwsq4leijxtEg/FG1wu/pzVu+7
r24vE6ovw0eWxe7aqzsPqCDX/s8vbehs525oLAO+p2PnV+U5Ge3GTQirpn9aeOUX
rN3rv1PEkh3ju1wtECllmmv/KaC1yaEd1GNwuoObMzzHbDDcusMSpAiP0vIlWLyH
DSZ3auMjw3PAT6L9iLsem1aM4rrILiM/wQxwi7+WoQX2b8fe9nama1K8xBEZx1/v
1twqUoCXUwglAEoRe4dJf0lWPPHJZ6/FtWDCHL8wfK1QFxy4QF2jr4k/Y4vP3Vx8
NqVQlEIHbp51ceXQrPUWGb8mLLpkcJLoGMh4mKU+H/d+t++bAWCFVV+MNFBDmDcX
4DXLPfTwRQwWbEFO5AZWFMHSxXxbaQj/7wl3qHKt7Sz7DO0b5xSULz0hq8gT1oPY
wQO4oextaq3uY43ZfnjFPQLLIk5kgXJZAC2H/PIHycxdQcf6+QciyoKO6MZ7yq3N
5hQNC8VsR6xMpVUZf9hAD4eLdKfbGHvp2UVzO+CJFL9f1j3YBm9w47KUy4OAw9Os
0WRj6Y8rs7+W2BwK7Ww43mnonndFMEr4hWNmvL5eU520I3Ck1mDDm8pZAw+uONEb
0veJoGX3FjSYuNosodfoiy8BVUxAIv6s9KMWLx4ezICQ+SArPR8y1zJtoFw/LSgD
2HUm3VcjYeDYdaU0wE/5doeZGp33rjmwe20uADys/IGUZvUy56ZhV4GIBjeEjKm9
K3vmP4twmp7aMT+U7DJmGdUpRboPzy9yURg9qgxmb3H1h5bY+2E1+ozi8iSq7lYZ
PyYbBY5nIPwfuVHkEki1+gS8XVjlClmwXaLM6AKYWUMVfrswfy8dgpdHzoVQTtU3
M2Qsflf8Q1MJT2/4z1ZVdO21SPt3WXLzXTSE0542FuLo4rbcl+qAmGj2EEmA1L9n
8Zo2G/awzljZi08dGy2GZGDOy/XwZRtIEGyQeeSI6QsCa00dDlA5gxsI8Xa04WLI
/MRlWoNZdfK/GCfWJ4DfqzIqAUx9PRzEACtV4hkNDNVOZ+U7LUh8gnckhw0L9yRw
M9SCxfyZqB6pPpieZrzmety/kmOlNInoV+llxcnjE5gV0QtR5JsG4zmNjNVSStlW
MTfE/lBoMqadGg8kRHWFA++3Y+a+9LkDuJHa/oG4KR1ma1NE+jyx/Dxaq3T1qJsO
mRMlmAdPuPY5Ch3WqqH1A31z1tCd/h9AT+tjVtZLBHMxsJA2kHmwjQJb0b48pFRf
4MrLImgh7KmMaTBGRsEvX1kYEXUOm6Q4488b+LUHITKY0+ZkSYVe+3BVD2L7ESz8
icYIxkLwbkKarkRG35N7Ru+MPaeDv8Ci4IHKn5/5Ag51egIBTGc9fHIwngJ6Dtws
Nc20+0NPfMlfD2f8LNx54CrJMTfcATmMyaV/UtCQWlUNMsy86O4fl4jsM++EZh26
1Se+CvhTarcavdw13QI9T0Pfyr8u8CKktTOGmkzj7Ewv28A1OPDS/nVoYzi2tzjK
LaaSHfW0V0xmqJK86wPt9V152cwGf/7ghzMA8pu/4MeucUyPNFRKsYhU9fGvmpO2
c42xe0GWTPKsA1PLFYpQpy4+yJvG17O0YjuxRX3+lTxDLnY9rV9aXvpOrUlm3Xr1
u9iC847KncdkOVjgTR4njVQs3RhjZH3MtarC1xwaiQUy52mRcBOOXEqoOwryz8bP
9Y2TWWPyYCDBQYWePJa2AqzDw3YJeBn8jrf6eJ2DJLorfxRsk9ahm1r6E0/J/0wO
Tu0ZSWLgJOE8IXC0DaWCpFAp8W557Ui+QRpl1NaA/R0xpTezUF7DCK7TQnFu+vUg
EB4SbqJ9LbyclhlHXj7pQ5mR2tko2WR+cMjEEutFdv1nXYZ9kp5SL2kU/0zqbd45
Gt922F6XQ/a273cfqYg2Lw2nK7J4Q9Fh1BG9/qL28sWeD9jK/ZhaW4SyETxfjDg2
Mfx+su00cX+5O0XKRylTijHlkuDYEOY4SAH/V7x5ly9vMLuCQWLrHm8ruBfZIKY1
PJrZ3mA3P3pzKm9k9I7HzXEtUbteRC9MzNyIGQKe8+Ayg3dVOmpAwQfwEsi+C43h
oHDHXuO7ZvE1FBXvBRfrCvg6th/8X7o3e9c5iXpVBdt4/vZSzxJrVaADjvQbTnlO
00aXRNONOuoNPxOs7VywhGpwMuZTGjI0MjYzeHpN0VKTD+1HDQwlbJTl3CQ/qrL/
imHzm1NUMOGbC6nrlyLeQTgQCM5oOCNzK7s4k23HJOpaoL2i/GjP/Xsfc9WanIcK
lnNSXz7zKKSlDbKReaCt6qUJMdp5aN3YEtQ+mxVQE9a8zO6/Brrb/JifWm7uelrp
TS82EbjU+4kdF+rbAAHzVAp4opuG8KYDYtnn8C48HsIwB2b+r18y8S/qsZ0YsBeg
BU4c8qxKnuK/uFP/UzHFynvF/FX6ZG7ELck5ehIHUEiCy9J5gU9uzThhgIYgglkt
EBdUJS/xla9GvrZec+ri0c9kXN3EI5aV0Oivu7WNG5Fxzf0m8N2XeUEuz8wyemVS
FKvywSWVQBEH0NbwUHd0VsRn7trQhUO4XMgfY+S+0BRcpjlMte0nltO64l8EvlFT
8g83B0DtgTgHb52CbM6sQRW2SW2I1PRD/nubGvhWr1YAfCVA7KX5q+1Mr1EUyWhb
iIkilQrLi8AidU7JzrWAxbfK+f2dZgi+lexMj1wvmo/2k33CMuKQsHDOCUpmoi9t
rPlHbopyNbJM6ITexlB2pJjGLASqViRouiG8uZjyUDLFUhNV/wyG5qfjjNX39gVo
ynIOOG83stoD/98z/og+LtC4IVOGr0mde5IDUWqNR1rcsL3TxP5mJuiLsjLa8VF3
5biUJWzBsiHOMIVsLcgLUiPNW1su4RoD099iU93M/7t+ocvpWA5/1pP42/GmXuW2
H5P0anW8nXtOxdvQgXFPTuRpnhJqwCzpOlfNotfRGIjSm/IaLND4+JNwALKp32+e
OITz5DIYlKuJcDBLUvF+7dbx5AQhiNoX1LeskoUo6ABq0cI7eHT0CqIGRu3bDVaT
e08b5VPltTCWeFnc1IWdhpQH9kH5X+gyJvsbo8n0KHBCi58fymsQkwU2sGoxlhx8
hEtaYt7M4gevOekpf2fZreBBcZBpumIwbBwjukLXGxBpgTnP0RK3KIQ4ggoZVP+0
wo9jMXpdx0nn4o+zlJlzrGXy7bm5bddD60xCUCATZWXNCKgjJPuWcXIQEwlIqsq3
pkDWxxJL1ekc+2NRm7QE4kmpKOEuu8JeuMncvXusSPVQjHKc9AEdxukbHErhBgCA
cQa2A65ji9JelAW508q2x48hmF7KVxDYLz35LY4LVSULBe+JpE9XHv+1d0CfJK4+
s9fIotmmJ34NJVNkKMDd7+iC1Mya8zBF5GXA1iXhc7WGZsqdv1j/kZI90YkDlWjr
rK2oiT4dlYHWAa3S3Zyw21pJYIjwp4lv3Vhqd0NXZzpRBe9Nnq5z5/4v8FCMlzGn
6vIbRztp3jRCizE9O7gYTMdstZGDneqIUyooFCNHfF79dwhuMOepTAzytaUeY7dy
oOMLkp50RdohQKr+j3IKcTjlbh6NC/JM4HcxNRMAjQZNFXuoYjWkT0T4uH4FJJw7
LMlg9g4w/X3IkL5WTaMQSES9wwKJkvC5NKgyaXKSrsD1kHTkBah1fapibN5dTJlc
T/dgR14Z8XbmKXQLYL5LSo4qe7hGVn3uOC1WxaIjgPNXsrCHEdJ8uAVOZOdH3Zwj
4rZ4qdk0H3hqL+7Eods/+Yji63YXaiV1dWnTpbtMnIEc3nImMBdhVgjrcw+tarF4
7CnMdQaDu/iEvhGs14ajhZzwJCRwjdjW602+4/EEWWbhC+yC+lkw06oEICoFTjbF
QwP69ZbO4wnb10GiuwA7zWvHchory1JpGq/Mhmm6F2ElY1rBY+Od3ejzO4Rmgx+z
rk4S4kt91B4AeEA6RfnWTcYRLHekRH3daMA+O4nCkpcHoy2bY2LpTccmU+WXIT6q
P7agymqowHBf7guQqlRc8Y0vc2tGr+SoW3847xf+Ih1MD1Seljrfq6AcPWSEeVKq
2tx5xmLKj1gaLDistymWlpvlJlsaKoDkT2ZcVYqKkwC9eKZGrQkB0LX9N4W5YcuC
wqW90n4izFuly8fqTq4icxeVolzFWRlMhV0oCkF1mZJFTIX8U7k3FLIMbW7MCcKg
Yw78nIElwnCkOa6tAzED9Fx8kRAiXXHVaqq2zORPmR9o78a82mYMflETeRnKqldC
18AGx9VMl67/xkq77+EKNmMuRg1+yc8SYonRcCmNa+xYh/RL1u+SvIZOJW3+vR1T
OZ1NH5cD1ncHhRIa1n3dsqXN+uHVzBuDKKunuYD8JIRv7hFmhpy5hltjmkDOcYUe
9ldOLeJTLSow4UQ0ZkvxwZ7gCeCto/LE+MaNYk/873DEG7Lh9TX5TXeOOQ5H2jk2
H9ris4YpsSczIMbo/vDx78wb+VR98/NaXFvmDHb0dVpZefQe/4aueBKTpfclEXRw
pO8ZTBEzDdPOnn7BgCEv8GE6Uabt6GoJWlAiDNKWDxZadfclnmem6lTCa1fZHVXb
yp+gRWTai2U4wkBMLdr1Z2N+eNKk0w9waAc9RC8nFjABNvGKTz6pUONE0rZs02fH
WoiFymyZ0Y5Jb7qjzF85olDqvZ2APxgXDW9o40fJAa8sMMHnCoGHTMIdQ5XOi5Uu
pdaPgk4Z96DksGS2zJU7EAeE1n5Blo9DIyX4ypem/W/ronJhdCF51y1HHYpkkn7H
NT/y/HjUGFNV6Bcawh9hHTuRJMyUKzzIRkovo+fAf6FhmqrwxT9R32D2B2apl61Q
xQOO9OLV9o1WOx7XR8maFs4EZ9X/kuR8qkTM57i/b0pIz9dFNxxCR7AMeUSgVh3t
24AY7wcJBGWMERhFYQrkohF4joZdjN6i1C+tk+GFGampgJKskUSISyrwI6+aTAC6
3P0G3HalA9UBSVjYAuaEIjovWWip187ytNAsaJ8voD7PiZprbyuUxMJynETs8dZT
vlKzFIezl8loo/5/7ZNBFzDUUUIpi4yXNppFS5VqZX2FFseH7iZNf3qIcZ1uvpPQ
OoLTfELWmF0/ckM8qUklvdJd0lca2yKRAsNgDc6SOcfpU8Evu7FhM6LoeW9oRkqv
FHoqF2cF2srWmNJieD4Otgzk70UvNmfFfkqYKTOtmBSLJo5Vtl256Wwp0GlsSuht
WkwDx2JIKkRsYGCyUKTgIi3n42Rg5TUlgeC9BRoOvyatdTVpVupbTxWrNz2YgHKy
Q9yCc9+klX6er71SR7Lc3fuDoh0NfLijEmI41oV8GxhZnYs67tm+K2f0kvNcWPhy
4sL/kE40A6ouqAkI/RwvZIcmOZaaDSp9qv5A2W5q5KtG3Epg2BgGdUZPzm+E3IRe
01YFWMy0f2TknBBZfRx9y+uq74slogYSb7j8hLUR6mnEl1tZgZTcrwfAnSjQh6eo
pgUY0ygdn8nKM9HDc7KkV2dX79P3EOnRrAGpqF58b6BxZABs99MvuC++b3yfW/kT
BaGjDX8qOR8uwgN8t6A0xXijr3lKz3anvWAxH/rt65iJpNcvze20oOFanOr80SrY
0lFXZz0UfiuuQHrnJuNBKLshmPmjMbbJc6828PoqhS+8xYkQg8JW1tSwbhKcGa7r
mrTOmL9INtpfDaOmDG/8pa6JS5gZWEomF2lh15q8R0028tz8sWelBl+A7ZIZ1yXL
Hu/G4DGLEfa2rOJm5JkDPRBPjtpPnB68/zhLRveS1GLhiFEPm65hmIgKzw72QsUU
IW3AVmVoiK8UfOZZcUp4Kx3sH+06gmMVfidbvU8z73R0zrOogBaGUbOrJ7EWLJY8
FWOXwkkW6tolPL7U0X88DLzUed2kWIJQ7tKZDmmEFXudh6rKnjCbQmsn/rJI/h7b
2wgYEp2+nn2+FX+lqlHDGGLa9pn8+MDclvtAXg0I0H5GbR2GC5J/HoOrDoo2W9wZ
h7NVc7pe7YFuRnLY6llWug7PRkxrHivUIJ5Oc75Rlr19u7+MgM4/tsnxkFgf1kAz
Vb7klAhTzkbBnWE0Ue6e4dD3czWkkhceUUEh5/S1d4zxwRJyzlUAdPQhfNyxo7yv
e/OktSRfQhZYfHzEF32iZnCkdu4WawjruE9twN0/nxmQMkSW6xti6drAi23M/ZWD
/8GqDAU8HpJxszFlXuzkGkmSE3LdcFq3yBW5XtPm2qhBY+xnxCLayffbqj+kpA1H
vA36zmwdXqrxJ7r5h/NIVJ0WnwbpjJ636av1v1mWaw4D+6rZD99t/KbH1y1WxTBd
+Ind9csBJ5zcStB5wHds9QlESFAYuNXfWiCuEeSqdA/+wYS+pb15b85iYtyfqnvx
hq3BporVe314IgKtgF336GaMPWTfKeNru4U4v4ZMUCnXb0lq9HJlfl+qg8NLvfx5
ApinTayh1cGsZUXPZumB4kMTzduDFSznRTJSNJ5kjxVdI0zRY8pNbqBR6qtRTa9J
QkKn21o91/Y5nFwLNjQv/4LboU2SHzC5RRJ9oZzN26M7fdpCEVX9Vhw/zL7I3xRz
v/myMNKRtljqvgrX8fLsQs3j6XlM1daRhMOhf0I5R6LAszOZEdF+9CzvQ8DgG8yH
1/AMF2CAOsa1C0GEK+5lLDFTT9z1VrTMOnf9bULgjQ6Lwq83DdlAHvCTg4HbFXiH
ftPiEPaoTtRK6IVGR102IxGYCxM3JjxWh/WIK7PuhDcQWFytFFrExUjx3cv6y0RW
V1wW88yXOsm3ih4f+XvMMsp9fyk5+laYRin7pDdbmbNtIiPpaQZ3QBVhIsTmKUGT
078Z78grW2A/lYpEYfx5b8RCU45qeQ0p1r+OL2MZimGLUrnztuF2p7SKWJHwf6+9
yAjCONdGSj0btNAysztHOPfG+2E+Wpk5dQM03nHl7JH5HF9tL8SkNCfN1qNA2uSJ
OEpFZb7vkA+UebguJfGmU1xsfTmbN3RTsBi4/BMN0LQrjiq/4l4Zagp2H0sh0bfu
rLvhICoQ1w8Ax4FFUf64lBQ/Oqzd4vRZn59lByUn1771ntDzvEz2ZDtJ6P2XpW7A
KCKR/mRQKXRTch9ldIK/xWHNWySXIugMqvq3g5Sryb9c83XSRnzhA/HRIgKZkuiY
Tav9C2no/LfY9g82D+csvxxTkW2qQIbNxrs4jSQvfDQVeVZPa1fv51wWFIHzC5ex
K3bWDaItxatgI1D+CnZ6XJ/gjcOoUvnjqOlwQ67sQHn719cwc+X6ZurIUKqSoA0K
Ag/MfMLM5mh+qB2GVVArWCpQ+44BnfOUf/R7S3zf7snwVzkIxForjlkAez4HyrI6
NM0il1DElG5jaVcHd52wkT3CqwhbcuYDWsIoVc1eHOZaWX8p0jPKNrPuA4taGg+J
AvSLnQlKpxkxY4Gyflip1+wCmun16GpUifNkfgsOuI8OaeCPb4Z6RJ2D3Sj5WXq5
FX0/9IpxI3YFK1l579OKPCPIIiKJNCM8SyQ9eLg53HmR+04mmcfnv9t8XwL+5Hky
XpcllqmXIlOaEijVTaPPAm0lQf+4+Z76pEqHXt+OCArgiSp9V5vqwzvafabFhYOH
1yoNxDZZSxnXadguP1cEae6Nhe2SGynDnmVcbp23An057Lu0xsTgiWKNK/S0D6Ur
GOQO1zVpDn23Bq4dQDyq/np1dKxJq9SpleTfmXKDHSNO5be410Jdo7GbUccqilor
37h0ZcYDZRvwqYsSDtaS2k0gijIPQSr+2clyNrKILdnldhrQ1Yh58WlRsaCjnnKV
WFAoInLRgcKWXCiP3pqr3KhVQJYnG/yscNY1wThsF3BTixcpgb+1veSMUpOjyS/d
AnwGKrRbZRplRSivmo9ZI5Ba7bsjTpP3vP5IsU0UQCmLasm4jLM1+0acB/OvktA+
qqZwPllFgF7nyhTP6aOC+TlYoMHhaLrg9vftCsBIeXVnENOXJOeJzd8ca+1xup9S
9qBpchY9A7wa49NkG0WcP8122RsOh0fPwGKdUmpJSsNSqxXiEPZLQUvIW0pydkvP
XL0L0XYq414en3IjVqsGPkQPPRhCEli4FBxh7tdJCjJ20BFC/AnaTS2dnZUp+29z
8vsqxp93aC4f4RqTOhTIGMYk+14llgbxmkS9yXVOJbIb+XEaIQWmoQvpqyQt63o1
q7Nx+sNfAc4RQDraGZeFwj4iviE0HYfVMQabOp9mLAr2Tyr9T5zQ+N07Qw27UMBR
rznVcAM8rVw2LGYP0aUodSZF2jc2JKJEvHp1p9HihBiCP5GsLxF5UJy8SeGtJVH1
6OI3fyliHJkO0PtTWbrePoxo4qW8E2cDTO7P+BN/Ff1Vj8beiXOTLuyXo6jkLRNs
p9V9i/aT7KFpZd6i9zdo1QqnusWZmsmFu7f4lXix36JU+k2YzxKhRkoQq2qbu+Y4
53AVBUCoijCs6pOxYI30fW5217yjgqf5bgoP3A0BrOHRKjgGeX8+c7r7UWcRmy7+
OCf7qf3w2hOifdtPW6VfnITq+s9a5TB+ju8RivZtC7wZam3exwcySkmhpp5Ap6UY
man98SD/43V6XcaPeHM6eHSIfbIRJmlnkgSLxDHXUFF5fk9BUkSuvfZmGD9eBSeI
s/DKk48xMKtbYxdpPEh/VXumX3lsWpl/9Qw7AypEqU4zHr2efKgpSvQMPGbOM1vW
on4Sw54MCIuSQAzemqR+9m7g+QTy10FA6l3saJ5uQ+F7RMGwCiCPE/8h2MOgUEuM
sV7PkcJxc5XglNdd9R4sbX/XLNOCdCIHM8KiZxT0bR4PAxl0/38hku0OiB0scXDi
hdxQK3+hQiFGeKLXi2hysPS0Zr063soaJkSVxNL3oi8RpzNe4Hu1ifgWWB7f4SGL
/lXNziYAbtVCtY0YRJZHckutfnfVNuu64lrnVQmA6QE5Aqukx9ZQWm0djnPj4zIv
8gkiBxK9XkStbXUnquq39mbNtob/POzVUyKYmRxD2c8BGrN64nHPGNbatql9BKp1
i6i5IXxkTFjp7P2ys/NZTYCs7xqq611DWd5Wv2v6fOtQ7+dz+61TJFcN4IBStSt1
iqcyVsReFt/YOtXHRN2uJ2HLIyAxGYnNp2qxBXrdkayspOl8/oVHtrWidI6s1dyT
x9jHrTWD/qwyNj1DneO0HYDIMQOXoyaykrSpisC8KcwizZiw5t6WBqHcdyYo2HSL
hkaT3jvuVgLiELmDAsWNy7fxI9C5gHX+PeXwq0YkGrlXkztZhCaM5oVscl/n7qKl
6ZPI0sfgGWiAsUIeN3T8B0fVVMG+S0b7BxF4PhIUBJc1/7J3UBCLXt7S91AWHYPg
ll20MR8yTCswGk16UpoxIuPYu+v+MpmVPX1DL3ck8namQYXes/4xlHT1OknZVclr
pyiKmYaf5EwvaoMtXH0+nml5QkYQFknQAxeBTXlQvOWOx5CpU8NLC46cFZubTcQh
hXsK5ZM1FbVA1MXKo18p65qXcL6VkUcP+QI5zDlyZNU9gxpacSF5/K6OEC/yGaki
uWskjHJsPpNdJHUZuQkaqezsiS31BX85FV535fYnw0ktZK4JmI/kjY/YMVEpKUZx
qUUQrnNHlna8x09sDrXDkIrVAEW/TJG+FxXPFz8FU2R+G11QQmxYwK82+wm4+8J+
fje/SI04w6n6lGv7FsZkwfZc3xGagNf8FGNbH7XAowHEblBCUJDzzQUJv5/HoR7q
7PEFOoKFTgYTN/0KYDELkw/WrRSQHb6GaVskUOmj2tZRGO1ZPDynooRla5K2vKp3
Xs4l2GI+V+tFRje6U/dkIYgGuSIN0VkwG4N/6G8JBXEHn9VlOQaS2GHXs94g4O+M
+Xvnfj993HmTDn46n2Lhu+Obhtdsi4+TQr1pGQ8XbbI8p5IAYUfRnoJbrY7/ZLGR
8MhCX3KTTDl27Mcw39H9EcT8SApRBbksw6pHARHlcTECKye3CyvuMXUVrzRZscWd
o0V+5i81PezBCIUd8QYAbXvOzQBqGo944Zbw/BeUwVRvC4QMiWkfVEHeo2Fozpj1
gRpERnvm4JSzkVN7xsS80m9tOvFHaa6ZSrn/O5rs2+6qLZa0hnIwS4JiClGQ3SIs
sL6CeIcJCUVLC1Ie5dPqLR5W28saJV7qw/2ASjEBXgekQ/3M10L5W9//9rAI78po
iJtgcyXzS1Pj+W7+BtcNd/75XYZjcpfdjaT7tc9XqP1QNnMkLLPBL26wjwu1t+Tc
1HFZG0RPDLfQ95nu7CUBRoHIai3WeC4LjYUCNhF6tguTU9qKP6NExtJLCdqf2oby
wYU0Y2fLnbbbEwi0KGqoDr19VAnHjp3e7uXhWWF08kEjl6/R0i+N2gevXJV/nIzH
//t+ZQJ3MRA0PoKacIcPeh5yhc2gyjgUMFSNtFohKSSWt99C5eb+6cb5mfAlhK7C
08IIIkCl8VKPjjJjuNoHQ1g2etBKHbnzHPCbQiNCyQ43vEnbUjxUfGzKxU2SzjjS
P+EPfkwRWu5iw+CUWYvvfDK6qa3VfBIb2lmXp8cS7VwV9A7ZYIs+23OxdpVQlGnX
EMFp2Pwa3JqCImlDJiLley3NFJ99TmnnyDqTtdkqIxGkt9z4oTM0SkXUXMYvONWV
f1NIOjB6RIiylSZ6ijVNYFIvGh75DCjwGOxNL/8Xj97L2cfzbJDu6b5wh5OR0I6H
U5hYNG9dON0flXrrMldo8c60ZtHUl7azv6N8TA1nSEHpdUmJWniS8/tp/Y85QK3k
aq0AATLCdomvplDYwgpQaLVrplrZKCuZvriUWBOkTqN0QuBZGIG3rYlCsIMbg6L3
qKeD0xr0dCd72G9EQmsjDUMj2sMgL+3fYa9O1xF72GHYuEN0zYZFxVg0r0/hO18A
0hO5kuRC6h+8C4lbjy2uk9B+2IPaDhN1jNoFY/RvRYOKWhMyAhIIpvJi1U6Zlcjz
yDezKiHPPD6qwFbb8ZV9BUkwlmFZae2wrN8otn1eKqM9DP68M8IhY+rH+URsDRpO
nYJG46slkUugAY6J+NJDxc8A6Rkg7EeL5WjlF8q40N09i4uv5rjf0qNa1DmiSvvo
k+lODHgcd81Ko6SQroyzDeTcpI2xwF3Vf7CuucX0eQURWngpW6WaNC0TTWl9mw1c
+IVPP4AYR3lEb+Mh+j4YoFdAY3m1b/tSUysNOysnibQefpOHsnxfbwfgHn8Hudeb
uQOf82p6Uz8Hp7Kt03VTIc2L2xxnSM5G9AstH/HSjnnrLCkTEUhwSEtbyHpZ6png
jkrw8yg00pibv/RsXbYqiHAlWo8vCMBQuCa7ZltUhU6YEAYEGlfucF8rH0Lz2YYQ
wGmNj4FzN+Gr6hhU4mfchm8JzG8/Fjnc0U7pAAoHmAXYaKOU0x1d4Ox1X6kPxRDt
9InQod6UahCrMt4+pFyuzGIjthSlyU+b/dOvFWH8Ybv4F1r1xMwUZyoSpnydcXH/
RqTUJzLMK2kIccKAy8K61S827LUYWwwAMGZFn8NFAfwVFHd18SEGgUqPJieO2LwI
9KryEEOXWZDm8hITBB07x7yRVxwMuNBw2syUhOz9ecRivvCbkz9e+C83RX2cFnpD
9KHKuzyqcPjT7ookCuTYQdCgAD7TEDfPPmqZ0GKyAcmWX2C1yfvJ3HYnlKlnjDxA
I7801jgk961nfPDslzJzKVxHzMnp1nPEqGKOpRpe942VuYK7OkROFLFHLuFbrJH0
WsDXYPkPecYIT7xEAJVuIAHnvvq3JdF3SSZ2xgrqQKuy4KIwE+a2qW+3miuUee1U
vAIwrFOYr7IrZPfFvYqU8nAuLfkvNau1rOsx5Z5rodAhKsCpINZYbIR/6CNU772c
KCA3G6BsU5afKtL4KjNiQKSO9j/BK77O4HIGGUHEihB7K/aPXwMa/4gj4BBMNEr7
8TkL9kEnQok2WSBWlq62UkzP9skayXOPixMwq4Zuh3c6qoCTA+Gam4rf4qzgyGX4
tqcWzp9UdhpZNt9iGmZsx1A20M5cm6cG/CsuEcDTN5qZ1qojXX+yQ6GIdFA9/qBq
SKsDxbPer2fjvxs+k9L/eDYCp3M0bfm42TqlHwJFgNGWNwMxhf77RPHJKiwb4ykt
ne4Nj+JtgbFBLzw0imVcd9zfr42cagM+Oz8lAOzJ/6bJ+/fYJwuxqqBO0i/L9aZp
TFOho2laq7FdpmctoHqsXbKvpvKEfT9rAC51PwBepGJgAZjXekOpJrr5J5HD/fUK
NIBL8LjlRppl3uJ6/S/83iNriKTSn2Fao6FE/5SgquSkpZj1e59JuCxPfdu2bSGN
iIfJHAWGKp4Rs+SnzqFSpuhXs192/cUOOl70jATNdGwKnFZv4qOttecRWuxo+Ecg
eXMKQNkaYqXnLKGFP2GqTwo8E3Pptw8YTxaDEZDvyzVeD2J+ggyAeC53qzkHFH7V
aaU1iV99UyMHDZSQSENXzesUHKutdrzu9ZQvpfpP+6r+gmxiYmH7lH2W1xAJ3vdI
0vKZQl/J9jNBpY+P++9n0i2U0mt0GdmAOrHyhnYGH8tCkxCCEXVyN7cGlEp72NLo
irPVBy03VjPv3w0esWqeNJg1Xtx0ou3FiX68W4i5MiKqP8Wobn1K1CjsIJwoB36v
k6JXb1mh8a/o+tGzNWCklMvF5ouELDJzTkvzG/DXQQqUqPbqYe8xZer155mvwogg
QvQp6wrqLFnWUvmn6Ep+AjQa4a/XXEpY9x8M5pVMbQxkffiUEXPtgCY9qZpob3rG
8WS4t+mV5rZxVUICeRBQyczBPR+lwvDVjUjvdzhav2CB6N1IcR1VHJqMAqi3s4Fv
1QNrg7QLDLQf6jEG821FPVKaLEH3a3Nl4V6rOW78TcVlluMFFii42mXUROZ0Zn9D
QhlWTnaJseCgAGHmeKpWSewMlEgxtN2pJ2ClN7Ib61bvrPJLD/lnZvVGc5+tSMiK
nqqpP2poPR/G5F3SMhNvKXaid3M0HrG2e1e/qpuuIwIEUQh6ZXexGaeuJMe5PXQ/
7WdefsFFaOjdr8kwB0zqRjvyKTalaifszIbBN0XFKf2kROiOY/FzG8V2hszTpb5h
kQohj6HlEVHlocwQ+BT2zCP65k4PGBVvdRdrEF31Iyid46QnqzTddBnH6egMHuua
4IFhi3wBlfNvFS382aHkLW1Cl1YOGd7OoUXijMp9+DBprfMalCCyU17Vw7+CQfI9
G4oDJ6KeaBvo5vj6/mIsZuZZVqH1viYborvmpGCa7oCEJ2YJ9DAQ2dpaDh22oNmZ
ZZwoj5HP7wbFBZPNhKMdWJhGqm6xh9NCaUsejJUbOwylza2OX/XhgU9wV2XCknnv
F//VQVViPCmx6Uzb7eb/0o+h/0gSq68oX2CnlFQYWjFlEaTLxv/gxpchcHXvJBQz
yRfFpprQv+L1sxcozaSHuIXiw3oQcViDMz0EMBejB6f9vgOX3Z8zFRn0WwmOJdc5
gdBn7FXlQ8v7j1KVF6mLJ3bHCUy2izwourHGf/i3ncvu8z5v37Exief0cxZteQ/d
uYe0YDPUrSF+Ht2GiHXBnBx1jOJ3v8+dI0LbG1n72q8rJjqb/mKlkc5FQn4FkvkH
5ptv6Ccg3QL5kYepKBP5eIykI+FEhI8e+807N9aN5JxmWy2KptU+g2gyqFOOi4tk
Wffc9lS5phYwUIEYc+fLicXkD0zFoHqLNIEP0TiIiuZDzxyyw92gEzlSsG7lb97s
n/mJbW+mHCHgE5UX2WRQbdCkjR4OJTUQnkAJq0Gimi73QzrLYpZmQrydrjBBYnKA
S8GXUZ4bUwVQZoEqoXwscRVfoFvYA/+lF93szs9Vb0ejo6L57DoNaHqxkLVO6HER
KyI1fsiYoN+lSZ2E94CsrKMumF5dS6nPF/WIeL2KzAg5s1bXllum6HBZbmD5Ys3r
xCIE/ISHvnFMG2BIwuOLjxzjMD1NmiOrayFhrbyOBQSYCLuTNUbBplHMiJ3oszXw
+8C1dHckdtDF3qiSfjcNl7qG3KjX2z0OzDCOwALjiINa5I+cEB+dnX+ejYc0Ew16
hkVr7eMWVXfrEFJoXD74ASr7ISWNM3e1FtJHqSa17j2AezlH8ebF3z8mnAZRo4ag
4vHCAzQ2OuS9hEy+wM/zg/F34O2zbN9pdXM0Qh8BHYQ4IlSx65PaNdm6l48ua46L
NnmaEAiBvvb3suy8N6hmgloLwUNoQqA1Fz4tkEignhuuLaRxuW0KzvfgdvP87h00
n6bveBSr+0w8ypmavSxGxGAoi5uh9uNwtOpPiO7/vfyju29gXFsw+p/Jd070eGva
HaN+e6Z3bt+9ErShUG/SFMWYisDdu4uq2Vx/vjwUl6tVmy2sUIZA7ud84wtXgfa5
zSFjkb2SgQSCzeNrPF5/DzXKLl5HA6fmDUqoXxzbyirk+XL0Ap6qAGAE2zrcZpZW
v6ES/rlm6jK8FTtgSzBdzDTvWojs/EFBQICOrp8XpfYpC1XAPAQuG+1xyyiu9FV/
TzSlvIiJfL78nTx8yeBYITUCfZUMulnZAOoeE/U4EKlIkGXRsXCG+gqJMqthqMMv
cF1ZIUkb9UeJBePcsRwF3M8ZW/IkMNEsRArnUzaIHg9yd8JbtTTbAwAvulX+IZuh
SISiXpQ1l3uJJsNKOYBazJYCWRLAmGzsAsOZwE1TcF7YF0723BVbIttei296Bys7
AtVvR/ENF+OmtkWWO+nc7xms2JYTq1qpKKI69fWjVnhNYYNrbQ8Ni8frVR10eh3m
hPX5AGLI/sP5Qb1ul0BPtYDI6RaAXtjJUUTv8ML56k3YYh8YP7o3ak73SIjkiw1D
MkxBrsp0evtO8kRkdK/M+RPxyHtireF2dm5i9USyjW1wguJZ0RtRAUTP0B5rR8Wq
AOOdFIE7Ii5N5jQA+xA3nTomDeF7ZSf+R8VOSii9J5GcYFoaxgym0/IYZ9r9HOL4
FN2qTBHBZfPZ9IEyD6CetGGpSBKIby53KenAX7HTFxO+scWvU/pRyR2kNj/BJ5RA
JlJk8uUD0fbP4ZpJMl9f3T/CiEc5vWgTpVdJobHf9dx4WNgFcidZ0E84aN6txyC5
1mPDVj1oUvE8wizOi7lAhouujVguHflwT9O3B24JfAl4JPqBhVWM0cmcYYdqa3/h
AX8ny9mmy7Ewayl/KRvYMKJwD63duRCOZF50OX2Jk5gN3fvsgi/QMogBGFBEVULF
T2aV4DvyJGms0A++9OE/h1XiN7DU5VQudbBUvbjwpga432YEXHaf47X0L4ic/zjq
KXz0FleH3VBhTs1I/NTwAKlVWoNVtHINTZMWN7eJE43Jde0phXdJwOu+UR7coqA8
bD4Ubzj9eyYiBrf0C0cQIr6jDPz+BCaCHLJ1TnuO7RsBfR6mtHWRrVbbqsOlWozU
zn2YT8GVyHnNiyWRA9Te5Y2Kwn77/lQZNV+J1gbdxWf7TwbM9D4JBTdieP3eMGev
QCdg1bIZVwxDaXVE9KjWqElVzIKqjvkotPW7D6MtULvel0y/Z0WX/RoADOHeb9Ij
TsL+r029BZNigxcKn+nq5yFpb31ShDo9DCtCa/kqzVe2elqWMZ5FR1qyyNsnTNrm
XACUY+BcS9TCrVJvhmgTl/1DtqiYehNAMcwIfZV2agHclHBrbjG9xuw3kJMx5M2H
nam5nzzVKThoiaELXxQNH3Z54MpsLZaJoztIT7jd/yw0pvBkl1DG94YQWrPt+8iq
U9GvctYXxmGACOYTsOk9ikbxLrfj/gc1jL+9W21DIGkQAVTYXU5jv0XAXvw6DT9O
xSSE8AbDQyFbNhrlHeMhPqi517Sd/5rKCua3gLnXJw3F1PVO48/bhIrNh4stH0lD
yY/+PZdCznNxxYfgEDWdNQGjP/9XWrKhbazthelHYDacK8+m96Pvw2S4AREYzl5s
VY9Z0UmnnNOiih5gXMhzLiDmuAb4rUyqVxzcjqEHXR+aPkx47MjLnwLmcIxV2qt2
ZRHX4nnBTmZ06r3mr/yJMZq3Q8VnYTkafMjmIx2obPY7J4aZzuggLocpW1cCOyoF
6DV2MAGcOqCeHdn8i/7btwUp87DznDvO6JxXQX1QurtM3yK1uO+IGZET0+sbA6lD
nnooFQE9xp+ruZu7bAM8WQZBd7MszAt15RF4qpdPtWuIpp1QrRFkZxqlUGhRA8Pf
TQL12ks6lt78B7A53Z7H9N8rHjy9vrQuEQ/+NGe98H7PVLPk6DZoOl1p35ILTZl0
sGXShAskEThrVe2sddBiB1+0IAA0WwCcnUBi37BndukF3RBflluGJUOgtCy/+3bi
ZPqMZCaA0vhuAQDoEMRKzCu9vuV2GjxXq9CecHsP5FhzEQPXI4RGTpHnSVr4mJdd
henq93OIQ5HXLqFHeeLweYibuSP1W7dgkpi8V1GFcOHuJniolfUgj2q9ne50/Ynf
lmU72xe/8e2xpeLDYuNyCwYAX05VEChYl4wTB7+KEd2j4Q8TzM1qoH+l//bMHbZ/
cEoBb7bkDOlusWWa2tI89iPrpKN+3q5U9CIpGfniU/ilzxWhRoTOGFnCwpdc3XKj
zOFc1PQoKBvbnwgLOXX3Iqos7dcb0wd1OpfPzrZ7l96UIqhOsYOiM87mpHuzx+d2
xG/Ev9LX0YydkY6gu9UyajvDhsaLOyCaCAKylV/FHkWNeQICEKGd/mvf/vTbhlms
lW7rSk6RSRmfPvHs437U9ifHXEl0Bf5oytXWBgONlgRj5n906XIOYVULRuvGKB6h
rn3d50X1YeY9SjXH56eRLCAtyPrTX56Cmlupv36oVeV07pupmRDTyUmFXUKQKgzE
gy3tEXlqgQFrorFV0/rjD1W2dizJEkkEATVqZEf5CZbhZWDVx6PB5H1RvCQUHv7d
HzzT79M2sBOfR/jJXeRGvzA4On3j0LRie2zY0/AUwLuzJaT7GjjK4xsD1on5HvAP
uEdFEQCGAWVU/SQRZUTMvzxlGGCrWTHyTFwf8NcnjbS9uJblx/GbIGennF5dRmG7
zKsPRzw7WydWtw3Sas9DeKGe2URzLqswXVqWJWY/gQpqkaLLvXoRCbP5k3Myutok
fn5xh7Q+WWJ7vtF9MAPcxbF75T9s/4S6QB2H6SWRQsA2LBFhDC7LY5wxeTnIYs2p
lWoSFY+JEgS0RnThAW9mcdiJykeKyehL4ZbNC1hfrtGZpYWe/5LIh/XtO+jA3YBZ
9aVpbVA/up8ev3zTFdTNxWqpDfAgSdn5A4JxNKNXIUHYfkNskMma7UvnMIovb8tu
4PsPFyx4+p6HDw1woHxpyqyEitBhXCeJz1rP4nGoKYmPr6wobHzQipgWlzPCrg63
Avrd2jkT1ZAPBdixg68OSeEF6vIITFMZshejZiUsHsb8lb907tyHgIOK63jIUgQU
gUnI1KmyPufHTSfz6caHhM0baacyPCiOjRrlu2kaL9rt+eipJPeKulNsC8ilOxFT
4+S+a7zhxqUcHlFNIXR8mUnIEcWhoJRkqHlxlxVLHMsg4bPXuB2/67XzR89X4jSF
YoM6I21I2gazTh1zx+Ww6/gS07J0o5OWFMq933ccKDhH/lNeEXN+ZfzBRgL7do0F
GCJaac+t59TpE6Ct18qrtn42cjqS8EBRvKJ5gIRJyUvuPoBoag4QYENKCrV5Giqy
Oq3BMwZcdyi3b6nz/8vIT/VaK/9OlMZnRxrfaSTjGIMUA1vjSCMvczpo49c9xiyR
z0jyPj/bPDXrnxMRgdXFdLQVN9RCxssGwgASlKiUtqTZ6Ezb/rZ6yMHIOEF2L3B0
RGElq56twTauD82ItSjsFnZqFKw4/K1S0iYt1BMImR+UusAzQ8BPppX6JhLTRxTw
qyDYx5FBe9A0f8DiRNKq0nbEVtyAKY5KuC7cUV5D93SA0lsUQpbMMX5YlruDlpS9
6puTnmEA/BU66uju7s478XvQhJhjy40CIL4rXOno+O/IkBKlzxDgrWcKRA7F1Lg7
dxinGlhs/dmSFqR9TAgr3SetS2500GB3258BL+on07+cpvTX3HAKzMVK4ZzqWNyV
ljGcMVs/GyZTmIxM8fdkpPE0K45wssNXW1/IjJnjEGgWrWiXIyRA8srzCfKtFpIA
umc40r3LlkLzWr+ExDkPCEl3mFod8FHdKGqdfObyk8JlaOhOg5XRgvTkGkuNTTrN
86l51K4GqYieDp5LToQYd1EP17SfaftSFhiyFe79IS3KicLsvoSzy4Gvy7frbykL
+vxz/KBp18FXg9wsEazm4G9fJHSinfsUnh488AIv9wbpHwvfq2NfvSzRUOVbD7u6
F3Dhl3b5d7rWix4KwAwvfe3r0k0u1AQkROYLcBmf85U7bx4AScmi8W7OVIbmB0LD
//awD8jrD8ewLtbqu0doOxYyBRttg6/E8FO0kuukQn6F98c4NNfT5qJ+X2VTFDwf
552Sf5lx7tneJWjMo29CIpIie1sq0CSYZM7XzsuF5sns8wtgPsLOt16gFel4hGLR
Xikt+DWeRjfksYJlD4KGi21t4tSbHLWLVgs/m5KTST4Sxk7dkl2lgvFOai+/EbCL
LTh5CjanwxyZnqFtsWxBXHGb7fi5qrBCfD/PRe38uOPgguf769RPo9OSgCYrFyEC
i0NKj3EG4w1hz1UlGtfTv4yIgDd+pJYUChsV/Nra/kOCoMaHA7kz2o1kJW6X86ZE
Bh6nMC177zIvXZImYdcgrk39+/V9MmjR1flFDzfIdsNyf2YI6ILxngIxcPEwrmPa
DYufSuxb4+wFgeSV2ziGHxoywtXv2SoMh94euQ6ym/HmxvLLfpXVnCpvtEjUetUi
PvDN3jGPm9PlgQ6z2KdbKuHWIXCgHqJ7bd5bb6yRLE64Rj4GotTCJKDDVe0Uh6Ep
Mb5sxcH0+bnnjVyd5HVGz+Rr+ywFqOvtJDeX5IeaF7N/MnUrQVm8iQESEdJbFwln
JDK4Z7FkROMiKhlOAKrs2l5JDRElMH0G4GpGaC9KYQjdzaG0qKERQPYMQ+ELI/db
DBqkEoNLwFKs5CEJh5Gxv2Za8e+JeOu1COZ2M64gM8BfiS0CdQm9ODxCvKY72iK9
FJV1kG8eQyk8y930z0bGKF3B658+VPsykUZWYbDvKAcNYx7JQ1QF8tDG5wgqBiad
NRkwDzIB8jXe/cRm6+y6c0s4BEDXxXa23XZNjU9TcA+vSH1SNdA3o3dIZ1QTjPrC
UkASA4DA1/VKthTStMx0KUjxrjWmMZEJDAp8ra3E7iO0X3rWzenKpUFvK+ODoRYN
ELD6M45//ZROJYpR1b9Qk6NmNegnrbVKMada+2KonpbaAWMZD5MMTmB23tkfHGku
wgST63v5Oi6ddugbi6jFNavgT8NzYebzLAhJs2tJ0KmwIBWD+dinZcyoaGw4nKDa
vp+yRygdn7OSaJceJJrm5EkyWpo69MyH0qAwMgydDiuvn/j1uQIs+fnEEnWz+f23
IcGD2nbIDknFMs9EanCyQIBNRuY7mZbYCh4A+e/zeEhEMFAkyQvU4jl3yPTldM0q
UCiqtGpuUzJf6PNjlRaD68sYZBufhre56nj0I5llCw/odETrDg95Qd2EWKuJ5BqO
0AWy7w2svavjxoJQ4krQKQwzf5VZU91uVeVEVbemeWQLgj56c1mQ5EjD9MClZuIv
oqWJggRodkLQpo5OKHsPrID6mX85/MfaJbMBPe7kzfK/R9eY19muquPM/KYVsMDr
gXGebAxtQ7RMsKzh2JbRgbeSj2PnXhiGEcCggFmlFZQzcIStvRc6s36xq095Iz1H
lfK/18uRcgGRwkHx9UduOtA2nIOLxkCCQ2aEcPIKDJVnk29kjO/65iCw0YSzzKqk
jNPbdIdaeBeQU9Y9179reWlII1wtnZqUA30fjfl29vlvoBHFEudy196edExsgSfA
cwjAeh0PrQIP9VVFYREIbNAmTE9LK0Pc8Yprw1mhuhXcO/nQiPBRwnW5H5Plrwag
l5moIdYSp/HGJPFc7cGGtm7ixoVJl51mLjDECU+DtCM+NopJK3qIJqlwOOUXmBeo
J47xMwLHTvSJwW8Lto2mRKfQPexRB/CV6HV0R2yAW4cWvWJqDB7miPnYw6zvG+F4
gI15TkPiwZDR9qI6vnCkivWQxmXI+4ILhYnpMXIffxTIce7VQuWYIK4dWf9Y84UT
XJqozi3BAn+fzXSz3YZRS9zZuJCB4D4tVBI2J/wsqCKiT/0DM2yTHYHfv6IeVL0p
ovUGHmFyn7z7sX1oBpLdpE4nTQbg7/awoKe7aP579k4UokNND9W0qszM6IThUsBm
hkgArjEBkwl9iEjuUYm5AfS5/oFnv8TZ+D3ncwYRKjm4gdxgYwLqfwcK+nBUm19V
IIXnD91HomdGHmGcbpcEwacM9P1JFklu92CnC2OteXvH1OfoDTtCTBETVECAQj8q
ehHoOFYmJCBW0KHwLFBED0ibcCY/Zu5xtAJ/vmxXZr8DWBKyV4Ri9yEJdACJg4h2
4/cfUKmjh7NupPWS2qqranMPuc0iiB0lN99AOe5D15fc3hl7HEJvpEJhhUAmcNiX
OZ4Zn3PdvNxWieezAoOCq4GHgPlvVnde8ggE3cVnAOvltvQKA8vdDItspKQWhiMH
EuzNWjuNCdDza3/ja5BZDPOzqhh+6aUeYp4afcS9VzzJaMj8MUZfHgyPc2fmdBjq
gl47q+0bJqWyLny/yXLTPLDfWAyWWguOeQbo0pMNhdVdkG9HhHX+WsK5aCXWB2YY
y3yf9i6YvBkwYaYDmHMNkwBK1bkHkBPbCqyeVz3jO0rnSIczbyanhoSOK4XBqezJ
iT2OiUk5OCKyNS35V3SPb/EMyDpJjwGXVpEewAYgJRNIZ6QIKX9Ye8JT6Bn+MKTv
Y1XUs4ue9/a69sx6Uv1P4oRDo/WPitGr9azQjycBRngWmEVyS49w6gdOvNdRCBFT
MgzndY5gysBXAyyM/IMqIkUHQ1ziKaIlCs2UHl10FC202oR1+W9filHG7hbT5MZ0
d6luxZRSwFNTMpadtWBTU9HWnNKGWxyqfYBw3/NbJddgFNPfEaGeeObD19zw7AKL
HQxIMDX1Q65wuKMNABFqyGSCwp6lPEMCbhMHblMc9yFwgpR6ihSYikHRBuYchj6D
vx8kMjMOGEdbGL4CEcOWW/6yiaxfPzMxGt9sk/QqZF4rNNlkyiTWp9YpdOS5RAV9
fH+y4wQU2DWzY+/QudoiDZkOVi92FF+7XIb5TQW5iOu6zjxuZEKm3S5cnvBgNs9p
H5odj9QjUDbQjlDPdsuasnDkn8f+P/RLpSNX6quAUpCCxhoYVSQoDYf9hWw9Cw9v
Z63PYgwTr//AAFzAk/0Kd0bAmurCc/G3EQw+79NrdfcBbG59ZlTuJe0rSVJ6rMbT
Cg6CqoEFaGxSFWhPYNDwZV+LkTktJ1Uh/SXbQDaRlHZcMRRid0xeZZQRamRI8vEW
/3xs9wRnnjpbN8oAHDulZcmMhl/xSJwEgz+UVtHPiZ9TC5advPYV71mOknzKFOyN
y1Y1uYqx7sPGEyB07LrsXfyyT+2INgy7rmN2RBCDoVRzjTokxPzpxcj8qbFoaROZ
tM6aKbhG6Qd1OW1Iqi9W4cgGh04F1gg0bI7UOdKjxCvorYXGeAbyP0jPVMn7/vHS
7iIqAuCDuRZYmHG9GS9zOCDHNq0s5jKNg7L973mLXAstv8b3SKTmFB84JUv7maEg
pkZzIzgc3fFeuE35/5ueo9QHQWhvuhpZ+9t1KiTxLNSBrE/O3QohzBifUWL9fWtd
h/funOzW39SrOmL2jp4MlXBrPhQQayO7eLMcQQ00FVbTeHHTMjLFxpFLqZ7dE0iH
H0FRebY6w6zOkrl9HpJneUr99me5rmusUbVgOOkgkN8Xl93umEDy4b8AU6CRk3TB
NhbflHwRp1UpT4+4VWN+VmelVIUkpdS1YjDfhGcF28NKZC00P+TBNEfU/p50HsSB
bXc7dd81qGw16TXoLuxDAMlfF21vjJybnSxbbbFredOfC9n93sIl7KlTFzVjeNfb
6ydHO0v0JpLdsGMiH/djVVjvhhcNx0YlrHDwhNO/zSXXw/03+Hlw9GKSFzcQiORy
fR+pIYp607TuMNCSvKruEmXd4VeFyfongnIwucnoGZTQiQv5eqLzHr/C99LNbq6V
UINkYuYH1XsY/G5W+Ylt3/WfVChjvwT0Eagii1pu34mS+qlqcD5A+LPMdg7iAAws
h6CLVl15rtmEgkvgtQKmQrJiYnlh6P1q9nceHLpu+C+Ur60NfudNT5GPVFcLsHls
JxB0VVJh/nkWDFh9qLyPiquglghsRakYZVI92z9YMel7v0Mk6nBUS1mL62MhWbny
Ey+iHolboYg8WAWMeeURnBsEFT89cObeXbQMsLaBXYEgypPKRrWe0wt+8BTzW+d/
pI3M3PCJHcvnayNntZ5M84AA9n9fFu0enjYt55FUBnBggjCZyo63ckVvoqdh6wtg
F6XnLupWmsa9dMzzW1409yGGfW3FZJToLmtfAUMapUbfy0kaImak2vjpiPKaXOxT
r4TdjWs+5NuTnECJnt35P6DBZ8DiSFm93AYDu8xYc8BeBqesx4sgUUCmHcuJZ09l
1vbtMmLhyeMlAetnuaSpwG6/sFH+aNaHl65YU9P7B8xPcgiFaNrfIlAzKBQXxtRj
efOQ9pYOlDyndobWY5aQ0lkp6bco3T4r9GrFuC3ans7U/przaxqRZDn4vy7lwqDW
VeyawfFr2DG426KP6SZzZD+dWEPEEPOpkVwFYpkqGvBM7QXUF0p7n95lzlpTI+Jw
7/e8tb0uVMG97FfBBRpxMYWRxmKGCKVgLpu2f41QYchY+LL0hsrWwPN0Y/gcRknM
oMaCdBuEk90M2B4Govy8nrg4UEYd3xd+zq0UqGBpZNLso0o+CidjQ93WJxn/Zp24
rP45oX2MrmhFrQPz5fxQ/rR2GYmQePfHIvB0dnkLiQRuyShwkGsLGC82WdhInFO2
1Aejb3HNTAe2F2bLBXo5Xi0BNEIV7x94xNL1swDgAJcHh32294mcshM2MmNm7LAC
BXceUIchESYeE9PTKGN1kqtlnE5eK84SBvqbbBMNzVo2exEwTTLZtOsok9Msmanl
hMENnqlX5K6CUBdktxOXeyX5ZZcKLCyxL/DuPzinf25HI1F5U0In/VV4Uca2MXSW
NhMnuIuY7zMAKo/cqjOO9A44n4ffHEWCPpkO+RXvWsZCQSs05+zt8JsIygv25XE7
j5fCFGyz1pOelW833482dkWSwQylBWUgEhbTrkLmS0HO7kc519soNlsdZLlEGeYD
acSer6DuoMNtLeBCsPtKVVHLbE8jDpi+F60f4Xv00ru+Z+w+9WoT5Q8pELSK2KGD
1YWNUGm8SxvIooDNL3WM8UNpQap1c7+d97bpLyhrEpjhH8abESFYPQym1e0C7IEZ
mymQkA70DxZhnZQryyFrHb8FVf6Raq/cwsrFpLMefoHWYbcHD3xDmB+LuHBMyRWQ
YVDD7S2dW4m7d+f8LhL1lc3UrSrEwX07i+4twkxDXhbnoYlYbmpbTfIwIBXwU8oV
gm/wxeXp0n/IZKdT29o7Jz1Q0oHjrTbKVn/cnE1SXh5t61G5IfFb5hfFjya2O6O5
ybW4jK6+M5j/lpqO5F68rwk8/HblaG+sPLEPtOaizGoBpbLD7BgXxKtMRVgI2mIj
zDvKwXr3l9Bnr1n92SvqGEupnZVyjIGPn6Lu5e0Bgq1LyIlH7nMj6z3NEjCxFp2a
SyPAvddk0uV4Sb/ELQsXU0abc4m1ESZj43cgOqHc2xsVquWmk/x96mSXBUUo6hrr
NF/4bVnRuIRx6fNAbzPuZ3O1yP4snuHmGU34WsrwE47Qe1Xm3jM07hX3XpnSQywA
5iVraMFvGN1pSVIteWW66o/H5A7UQbfxuhNQ9AwutA31yLdS8olDVEEw2KqeqoBm
NmaD86uKrv3mlcds8WFXuUwzhhJnBi2Cpvmfwr5/El/LEw6d1L6Uh6JrzNtkcPll
916gBwRxxIX+znGXtw0Z2fD4aeWKQ1HQJUC/ZPGeUN6WeckBh3QdxH6ZxCk9Y6g0
UlFUDZnKn8F+4g/y3Au6jJE/0F/5R7RoS2DkM0emIYSapSHKv7fy+K57QLZynkDB
k3hHLpil8J/IDq/cxpHf8/rGzjfn3CFsSGzMBoX1F49dHQQ/wCYljEVkiaVkeF5X
WyDGmt+a3w+nwk9u0QLCUc147XLBegXepLRCEXUSbDq0xzOUJ52bCtAW2Q+tFtv0
F36Wq578pMWrrv1R1qvcmytZt010cz7ZAXfYDMY0JzHVla0DLvNea8v+ikce6906
LWeEtNV4b9KpMViNLn7dLo6CsGgfaBWx474LsEocwVnHeDLgHJ4zU4iS6P/sHgq0
Sqiu2mwV0yZC92y/bvpVweZRcjeibs2vi0hf+Qt1R0cloSk7Ua2eNeqQ5gTNYEX0
jITlgEPfEaGeaSP44HAktxM23B7HKn+hPL3kLSr0vTssOAEkMatyTDImd1gfGnZa
30ij/4Igxehgi5mF70DxKbXI/B4Shy01L6Kyj0DIUaVvsQEgrDexigniQ23AfDUU
+F66yi8Xy7xJTb5q4s6vYOMQ6NOqJwz/u1Qy4G/ME9dGtdM0hVMiWLytpALOYLAd
zpjzcOA5PdhARJM1i0TU5lj8wBsuWkFE7GEMhvOKmBRFp9h03/eDpqONquHaC8Fp
tGMiPKN1wST2B9EGCwjzq08ByKMiap8eeHZAUXtkuiyXer4WUh9N1MANyLVpQbBP
uk8xc19DwUryu/UUsuN9p/AvmcbFPOlcNNOc97r89dfwCUwSpfccyBcpXyGVL1uZ
PqKuGIMcRoe8ThUjU8uAUHqXw8p3N4S9hlGfwdS9kShkZslHHMGgjaVTunnFfstx
p84MRFilkhSsJDFjRFaK7J4X1CZKXu4jMbWzxckFgSudSxBS+rDF42w3WvyYmroy
fQ9a96NGyz8tC+kp54iKhpbT2fGAiWROeXeA15kmwvm9+w3qETABGIUD67ES+wlD
XAyGhqRUSwlMmRmyAdaIbQqk1vUdheaf8DtnUsA0gz/h+SmAjrct2+CAddtV8a7x
wrHjxkw0dVn0FwshiIai59p+8idkV17ao/DD02PueY/l8j8YwJUS0Iw4XsQUECud
p3lmA7+JI5CbT7516nNLsGyFHw24HUUxsexxhC0tKhHl+Dl1FdfiHAne2a2WGw7u
h5nbeyChHDgpjbJwtE7z0dRwLru3FKSaQfQ5r+dreIksPDaMr5k+U0X3zXDLPhSk
tWQbG7VEICJ7Uc1Cim/qugwHRtLW/u39YmfSn8caCet7lnDLaBQ3hvaQxOiR7W3K
+V9X9hr3hqpp3XISibfmVvWyFy6AIe1dvEbH4yJw+Bc0pK1DniATUXNZXQuvXbu2
fDgOsNqqQSm1HgO21TeBTWxe2bLglVOflV/DT/PttLqJgqrI6+4bO9rPX7tSQaEr
eAiOrz+Q0m6toh4J9HGB0rUMNTupuSw2vliaHa8RZqQmrprYHGO9R/VkshitS3vV
shanhC/6bS/xCijqV6ht8FU+Z0d4rUV5JM0Kz1ngELRnB2adn7gimiyIAiw+qPkr
/1Dypo7T2U92/mlDOcwyrkq6KlrFPaewQYnMKUP84kAlvNxf3K4qnX9UiMIVhBCD
CBfbL8D4rcjFOWKLZC6nH3p6mq3IeQmO2BW9FWoHhofNlhfye3Msv0PP79jKHHYD
gBM9iMF2TrkMeUDSR0WfdTsU+8PMupT6fSsgg8+idCwDqj2Ctpbu8W1jmQGfqM/4
eNewjxBZT8UxYp5Rn8mzFWTFk9lZrrAHD8izfLOgDKuHkeiSyq7Pq4uBR9vAysHT
ktHoe8iKX0NjPuiNujUN4d/QcUGGgWkYKPoRNxngZzSROh4CTl50CiJcs50usA6I
C3yf9Ag0bap7kyRn7t2peA7VjrEYzBvE/lZGCjF1vVXJFGq2ej2ohHKIYn9xMi8x
F5ZXz+QbwbjNk/YjJYk/1Aj9Rs/VZO2qgumYCxyYaHKWmHw2PcUEWea9HmeLLgFC
+HA7i8ju6NC5PRyHdNUfHeqf5ok+B65QCTIUPfd27OkV2L2VQGb7PDdhdKz3vsgS
DwzK1Q1EUY5iGfpW1uOPLgeACKKPIPmrfki77Y1tdNvNHldbGiSRwblk81xfdXkm
Iel3acLJA9F0899OApV2f0FdsMmOBKVfwX4vgfsvG23tc1BmAefOUeU2GjwKPLOo
dMKJwAYjKsQQR5czznlHYx/JlliWe2osX95TJt05FMG9upbZWUrGYIdjNI6tweHd
o8fD8MnSYjIXsNXicL6Pg26hyHt0HMlBtippYZCfDc8hbFL6WJq+0VOHhs39ro7G
R896XrYJPqTgGLERWBnRjpYO+zYaKdqE+l3RzRQ0vtsJJjz6QVNhkk6+XWQA54aj
2R5SJeOx8jdalTJFkugiKsoGKE4s5cnp6mjrdIwhqqkKINAeZmKMRhJl+m5gSxJZ
U77j/+NfoInNsW5tAGz3xe4E10ejE7nRrqnIf7Zl4Ybz0iHVRLMAQftH82KNvKTd
UHP7INNoFKY+my0FCOl9aJ2Cqz9+I7eAH1ZGl8eVAIkO6UGhwrg2ZiVUXPqBFQo6
WeW2eKiSBCFmBE4EndjFK7Z2KxPQ6okpRsxV4aZng/NJoIaOWt9+1GI66DN71w1I
nq2YTDM3i7jMFKEMxFxw0jU/VrdwhrdNVlpSqipXZcLR9MGu2h59LdfHqykXFTeL
YqK6jElLlcNwfaey11cSvkqVGaEFbuZnNXtval6lSqFrtqd6wB73hRcorc3cJ2Cm
U+2NKx9oiU6/JFpz02ycvgh63QxEXX2cTZq2rSTZit7SmdCar+sv5uNpwEUsTu8f
wG0QNkT6XJIJ+jm5kDasaPCvh4EaCVUH6+xTDfhLPKTpQEe3Hbo4Grf/qs2jfWgK
gFFQh7CG4/UaCfTjtfBGssyIV9NErWgdhzgpC8Ft4DLvMTx51z6Bx1zCBlbvXtfD
uAQacYuhyPGpsmepXnMT1P2lualHodyMEU2YCFZirS8QlvO0LZcvYj38RtsrzSXT
g+5cJ8TQW41X2stL2u9Zv79W6eu3MMD6qYqKhoI7h/VO8+2dukuLS++V03WNUBXL
tndrW6x/3eP6gsZ3Cs7wMXnIHq6KNwb/EgpYySYzmACXZ46iVceqIwaJD+hYaTch
p4fYe7D217jW7aNqO+kLIYKfVS1tntI5b9AWr9kt+m7H+fv4/uJGla+lKv30Qiad
UY3KF0UFTUg/HHW2WFMOmX67rKtzoyZfpTVk7IJJwOPq3D/nQicQzIe+b1eJNw7t
v7Y6RCMN96vVq6uWbjhTFpCyKD9XI7HtqqBCUKSk57zEknc93rXsYQivVdISGr7I
gGUNoKzDmRhNgq5HZjLV/yV+GuhVyKIJVdw07XV9Y/aspmisURytSeJIojdz7nZS
uBX9f4G0Fb0ycsNKzODO5E3a4ZWBg2SgXJsW4nA1JNPGWrydPRoSoG8txAKw+Lka
V1r+mGOKQx5+DJ+S0huU/XshkABFBB+gjl+nWDYY/wHR3uM4VucC0PKx4Q77h4uM
q0qkYygxHjej199DaNNCQ8oYHFuu110hCMNlX+qesOxul0ew9XgeytgQ58r//xQT
AOjlzFDXqc4gI2K81eqnrbkWH8nVmFEV2TfD+7OaoHEv5ckQzT1azCQZ3OE5/AMJ
IRlLJpXix6Vi5W/q3lvypq2oxn1ONxjpXTJMSQGdyuPw3iBR40zjOQ38X5v8wB1n
b2TQxiokHjlmKAdvLmbEvPiXpbIG9CmnIYw+z37hsmpKfUMxRChsorTG5wtj7a9t
n9P/vDJpEvwRQzdY9nuAFckG6cFdHH5oUPzy/xLw5C3jkGCKei/j2AWm0rdsg0wk
5RNDAn6mcJ52L2l6q44mTc0Zjw7u8aejCVDVeX6FcpGqrriohluqH4X0Lk1G/0Rl
wx8c3PLVnXtKUNCpG2GpYFHRoE7KJrmqaOElmQn73eaKXNCegRv/zRHvQL/A4C3a
SIQPa5hcTChgWYR7F174ko47SFgBUIFg41a/3ytgQd0tCD5pk/pWAcFnlJWpCfh3
sYBI6b79YWxYG/toVyF85gh9MrUzvgrRu3vJqVdqctac0BouPixvonIdhGdnLB+H
vfNvpql7i+xDI4AkWYJyDPK4u7YjX/Vx24qq21jWjCb7PV9Bn7lWRyyr9WpilDfo
egZY8UCrdnwNg7+KuHcx42xV9S+DU/V0Ws66d6FiWxQDNWZGVw1E6YATeJx0I2Aj
YwPbUctZV0f29YyycPqZ3hacT1F05ZCEIB5hhxDGKZorm6D32deacWVBrrexcDN/
gzd1FyoI2efv1ldHKMuoKPDIcvi9Ke1MP8XRag3aJzSyHCwI3nYcCtdGgbWXMgpu
bz22pASqG/uzMs+FYErWB+BcjtVWKuaNEcBagJijTaKrXFpeHN/ziCSIBzZ84IBM
veX5RteuOFOYh8uUoi2lPT7rFhc1W7NtWyMGF3JEstKS646diTchXJdjwKfrhksR
n3AyLcNl1GsmkuX85cTglINHie3m4VpBSoOJt9xI7RDL6ql3RgrOWxYtCETZLvDu
cHQV46mDWH9+kXaUZ5l/CnMTyVGvw6fKnZstznhwix8PXqoQCXfukRYyy3CRfjy/
licdG/0GRqOBCVFEiQgXJqfRph5UdJXYBNDA3Dc/CLrMrbITu7ebCWFBgo/Ke+mI
tmB55z6S4j7gc+JEnqoE5g7+p4HovPLvSf4PNQ79hZvCEN8sQbEiYtMbYUShTlHA
VWO5GLUEgL56hVJGbG0OJGGGIeK2vTVgkMBDmsY5y91jpC48wyPK/zzMGF28RUnE
VeubzIvUYCrqitEQ8b6miDc3Icgmx5UX5qOy1S/IU15bY3mcASuhCT5/Rmyh5kZP
NJLgDwtQ2vjiyauBAZde942QmZm0lIfOu8PmxIOW7sr/tKdt3C/w4cplyaY1DaIO
H1UQoZEtcERBrVuwSBJjFq5XN0ZmnqhFWVkKu944X6UVQCz1ynvmdKcOGjjCCgaK
EGbZmx47ql7c815XT6vHPZ4DdiSVwInDZN2FRwG5KngCG6T6rBZ9w080QXJB2cIx
E2APYYSAxDPa1T0kTzvGs3gQMXvrAvZec9POH1PsJiIDAEsihy8EyPIbHLb9xYCd
/Vghh0VxGjo6ByLujGd5NRxnJl78nSXBJMtL0jEmQq7aU4vu+iToEz20rW6CjTuz
ZRJVDiNIbNXUGN8i9u1X9KNFX96RQNuzy024G9tcnIeI9T5sSdnpLlK3dJGqXGRt
j6aC3gPKZeDe2Ts5vCooKceoJLFqgB5jFrqzkr9nkZjCRU0RJGvR+v7HPzWVOobp
KA3FprEMyAgLNKE3Rw3NAYPFwYgBGgSyvBoJIxSyNp6u9UNi4gbo9JHfu3UzdJwC
4yK9Df3zaQLF4RNy3/iGaiR6cx52jrC7bA20OJEat4oGwN8qDfI32o864fRVoZTO
WoQzQriFpsDNIP1t3xwpesYOXBALnAX3AHxMYshtU8oa1CFIH4yXvw9DuwEz18wz
w8KgKknCJUQcfY8/+zfgOyt7gX6YZkw66i8pA1M3xy+ynnn2gAvCYSR0YOsd5Al0
zk+VFKwgopvaW4A60+bYCI/RtqBN7HSropoy9WAlVjDKgaD9vLrJEmCrkq1Xt/64
EA6vdYbAkfjO/TMzvLBrDL2jaVJs8TKhfZdL4cE+6j4a7R6wnHzNwOyJY/H8ggSj
h3I2CVvYuwU6WIfly7MeF7mP3AFxOyP1Qgc43ZRYR/Hpm+bAZHp/Q7om8hs0nIxV
AflrskCWD4c0HmtOyhdGckTCCZw598Mq1Nneiht7VrW5GUYEuRtXbx1H9P8YhqSy
HwOv+OI6BsaWOJmqo0HE/0wjU3P/TMIAcaD5Jf6kvGym/F913BjU2kdj94B6BPg+
w2N68o+xMx5f2fEbuvY7mTPJVaHF+S0GDl5l1YDGlwPyB+fDjs0geBmjl79yeAc8
A3UmY2GbznGAsNjU132OHqGINj45fhg56+J+iFD1MDClXO6g630IGGFbUeQ+ICA1
Bk6+h1HAqLQLMf5bA9bv7jY541ICye/SAi1aK1SW/oRx3XLmyVfgo28C5LV/ivzC
bXoNhuuwDRSLtULgxIE/sRzfQqDBPtSekt2bVeQc5Mdey3pCMZa3dbAeURPX8Lgj
iZt6vB4kn3OFEvGvpYGvSpva0+uRzlNBO2yGA/CyajaoMucXBiaNpYc5ZqGuZ8Fn
Fh2bMrlpTzmKsREWYFoVrP2Btq/NiaCfeE7oRvreA4RL+rLqRb1w4jODw/BAU7zw
n1rv6GtolkDqYsufwxcPKWGQIgjgpB370kwGINIsgDVzOqHiQZh3ZeJ1WoOhq/mr
4RbVn7W+smAFVQnFykZtYrHH0UAwHxvBCgdyZCICCxOmL9+a1PRejVhUbcrUObPA
9xR1yNwkK05O3TIr7CwNMGYFxqJSWYPR3jGVm6YB25/40xPom6GU3agUX6JywVMM
mAEWp2/xzXpJDMPuRVa5VgM0/gf60CmqtuNSTtAn+8IGXdEKaVcrZGrYl/zPG+wm
bvql4Aeb7bQ1vOrVs4rGKDfssOYf3vXjC+4WROrqbXYs1JpOqsKkyb46zoCdrGiZ
W9wR9y/M0pdhyI3ePOtc4B4RJ9ZmgGQ6Kl9ETG8Z+lbjvR3W4OYTYlCVGaDtt/C+
PBy+khVFOZy6vzXfKj8AHPw+SqRiVxdNcZ6rgjDlK56WK22mcbhwyoftN3cBCgKF
FtTBgnH0DInBO9sAbRnfyqRCpND7ow53P3uBZNJiFm15lbh3fl47ehYHKrFUblze
TYtuXaeVz+Xsd3Tg3/0j71Bs1TteqbvteQI5s6tTsJiKyLFhs0g3dgtGtC0f/Hlm
1eShsIWMazmvAGiPhejXJbs0qBN/7n8avnu/7+qrI/5uPLmhp/zQxkttKp3qdBDi
2TiKIQ3ocXoDqsGLMGsDeoT+zwkZU/32dlSFg0EmuK3zVDMxFmSH3ztGPqKNjQ33
wOxJ7YAI2ZSaXn3gkubb+46UYdO3x0UV1DiCTWKpXgl6lHNor3eRn8PXSsnJYZTf
upZ+wW9TrAg8MAxnMsGWOgtJ+6At88G2yAc1v0fosOGQo52ZWy6ufNm3VKWy3OMC
K2M+jmI1CggpPLJq9r4TXAy4keS2bMBIy6dpupkUbZATAu1srRdm6mLBVHBbhwlf
VOZr8eMa8JajSEaVrjKf1aJ8xUfHTAlTgTIJ+tZUJpJM+PgvKIWjB5KpOToodn66
IMVDFIWCl5ehz6tDsSwPjac/9+uomIPD7cZU2jGc016o8fv0UpUWy4Che/g2idCb
NpxX8nlZ8JEtM8JuuXVXy6s6aXq0cd0L1viBTQfOn3G997y3eGRQB+abWLmsmU5W
eR9fhOwlPHAh1qtPa8NYStNZyt5N9pHmibYYWfkXFf0K6smGNcQEE7MV/JzVpQC0
5WRLQEi76U4IklHMoa1Xa+Dru8nhTvhGygJniVYyNJniyAXCmk206uwj7W54gltA
MtD/+9kG/9/WM2hdFZvJzLfJQJx1zna2tlOC74GPfHYM2HCTw2elp5p4UcQVHR2+
HjwZi3zwtf4BjT/f2MxcyGAs530a3AwoS2j+k2mXjhYxf/R610S4sPTAemq2r4CB
7YqBtwvC1eYIoi/iHS/IJrmDm+dKK8+WhK8r/jUt6GimbqT98P28/rVD9pE3vs7I
tQjkxYBSYHAeFcikuoyPM58SU/CSPsGH0tr3SRllk6mlaBekk9jOHztrXGGfDbRu
Rx88fkt3RLXoUOfZuEQamgyRQ1Ro5UlG4wknRdIhMOIztENOKGBSyKnZBYDn0IEd
AkbC8sp9m/sQdezzi745WyjD3gG7T00AzLqLFHRPGogYHramt5lurs6GbqbMOqxZ
gwVs1h6RDT6AEUicg1LiGROltkoJLNE5Zwgz3XGMIKj5jJbR4PSewmzwDZ2VbPUM
ssIJrf5ZaIh1KkiqR9yzOE2KR8eVNuS78iKuHVdZ6ej7BA5wi8fsvvd2Q8UTf9p7
FDnOUIMzi5BFjozsZKECUVTxIbhCr6PqGP1fWuRN+mspNTlFgXcsZPo8TSMdumz+
DNbkyj2g1c1NQYs4olNqHnuf5n5CypgV2hH2t1CjwLUra4xD0OogK0lZE3SricpR
64XIwGEt3VxfErE89JRX1MeB/anA7KHV7RDUUu08JxIAvbEjui2RWlHwA6ecXPKR
NDa5AdOgl3bvzeFpOo5jztrKb35PuiubxCUT85wnf0ZAOJFR0+OkzNYedSgVi8Sa
1KxiXWvU0Xo39mQLBo4hRpItuPON2PPuX+v9Mqn2zKc8ga8M08hEd9NlDK39Ff+e
cpfspIq4uOQGTA7HWbY3nCLobcSY7w9apQ/20nD+iFLJCG/3UgyStbV6wA8AKkg7
GScVZZCf3J2euO3SUZ4kOU6MmtVhkY4rM7obR3DzcQCfJR5HiBr1Wi+Fk7Ysa4Qh
8s1xjMS6mBEJlrsVp/0pm5bnVrmVTeH82upWUHPyrHEZodf9tifA/dBynIJeFZpq
j49zwRfKjdZYYzOkZcOa/JDWHHphXF1TdxkY/zAcxOF6Z8DKHbuqg226yktz2Jf8
G71S558Raimc89WETBvGLK5afGkLMoJKf0uHUg6sQ//O82wF6mcNP2lOKPmfNDhW
LjZT5xRAPHpcdTPXLRlzkhf/zA6jOuO8z9FC/rz0GdvqdlVoOPYnIb8/ruza68mL
qps/zldpGODuUPKOnC2egfCcOEhDgr5NNtQMoHn4tkkkJVRgBgM6zcpF6iU+7CZb
XOnTzPvOF8V0ex3RRCvfjMdfWMLPFRBEZxjRj8fdINASW1N1sN96vFJPUTbNnDVN
in6b8KPIJkud31zGRuYlekOsdtPvN8D1s3G3WD4RAa/thedNQOshVhcbS6sHzqYT
TyyUU3tHdE0HIx+CvNL9Bi+7cmv00NxZ547vtySUg3cja5kYSOEuTjkhW0cBIodB
i8P3KoqNB7kKevCx1ZKzwztgqMmk6eyVecvR9EBgmHg84XXeg2We1YohNIJiF2ub
1KYL4zDtacvb8ZzbR+/wli4dpSa/JAYPKQE/mXxB+Jq8M/c/Bu4nwzAzF72wzXEW
gpFhcMlUQW17aGO3eULftlv3yOamlu1hkj2iyjSp1MHNHvD6Y7PrpXXKOLbnQqMX
qkskcwWFi8hgidsg2VGb0J3YSM+C1j//Dj/zTuVEI7wALPfEp/BXIWiGwvhv+CEP
vlCh+OQtL8R7gTtSy6xhHD+UpE9ZZrsSy9Zngz0FHctKekPBgd/+jnNRwpcd764Q
GAXOJVwUQJYg1cukBBsCFvJ5FMemcUP97cr16qe5LrKRyZeE0oqqs6K9wSpWQMGp
1wl3HcIww/W4fpVjPS4exYv3D/pgxbda0JFieZJUGq+lnuKa1BgosA3n5i7tZ+wE
zDMfpVB83S0kY9Bi81LJkbzZJ2oVKamEyB7J0HYQvm1kfkEILfpm5wu2aOgGq2KW
+4Ud2MyKvof/YSH5JtRhv7F2ZLybRnHB+11ct5Sf8Jp4U+hmUumh8OczlaQ8hpAD
akJTIWPsV5A/OrdMMJ3voESFMnniJ5WizeQ980zNdTAPKfRt53FltFr1rbELYzaw
XK8jwDO3UhxXOejb/x56F7qxSKOSZpGpXM4mnuPWOHalROSTeO4PKJSGzWPek2Ks
Un3GPSd6vyrROgF85VdrZTG4fc4EI6IVQxm6H57ppkIkewBfPpoqEy7xmHjgyvSa
dI7TEypVz9X0TmM97LLiX4T9nCJY2G8++JGuA1yo0n7z3tlzWWo96QYnQ4FNqUTN
isKpRdxtJiQEvDjW+Urjd2EsPfx6HzcyBRWsxO3jtnDzI8pVq2JwY1V713l/wwqz
hxJaltEOCnvUJcTMUqEw2P/j8x1FpbhUMnWpvQNyRsB3tMt2ebC3RKyi0LMLMVRa
ZSbmMOUDRt9j0I7vLVhRF4NGxfgaLGT/AzHnat8yvlLokrYq1joWndN3y8BNFTNW
HIFph2WntK9WgqpO2Cv8fpqxpQFUAWqVfaxpml1JoCNmnLnIgpZDMfBKIuE0GVND
TMFXQNAD3ghlzmUFMAz1FxyzFxf0wFOTY3io2gjQKB0sOcQQvRVlasLX9H1rNvOa
UhpUt9upMi6Tq1TkYRnoOWH3WRGTM4+NG2mIjAy9qiQJPrUjr+Tydy8u+w+r6/CO
utLNY03Qx4ksXNr920MYlEnXJRcKblAFDXDCXx7i14Me8PXtLf+tpylyWHe81JDg
UAgnWpeITSLQsNFwQCZ8UYzTSjFLShg4/1yLt9fZEeya4TztAspP95dtIgzXtr2L
QtH7Tzz96wyXAXUEfB0R49q8ntBQyZk12yMK2AH2j5DhyrVSQFWZJSkOvkz9sn49
K2hlgqhF0iNbdo21ItrJMbPSCR/8BsFTSk2J6i0W9AqAqc9+07EJXfLVWQjnVgUG
D1ZTzPatf9EmQg8aTmeLohOYiO+gKyHNzH7Q1qKzyaPCf08M7wMIXZGybDiB/QvL
lhZ16iFMendUNbnlFbMfM30k0vtzr9Xqqk6Asdz8vMKAWqMwsFEV01TSczgH/NM4
YFOeGUWgt5oVCA7C/rYfPOcoh9nXSq4Dy2SbtjPXNFobIZRLRXPVqA9Ch/5Xgknu
JI9+ffk5kCZm5527phx6KQDjJhVbzK//3KHllTbFzJKQL1b0mANopPnuh5mxTOzv
7LP2qBIrN2FtrsStTd1m42ewgWhCWaAYUnSuMsCQENe6RKCiV25RMk8xJHm8rwdW
y33TjR69mA4P7rm+NAP+PWqoMGysTcu5c/3XRJUlbXz73d6K6xCZDL+8l5e7Ioaa
p2fvP+0VWB+v9vOmGVW/NhMHfmn5jyPCseMzRL9HBKbbbt+F2d4OPE+gpiaATwt/
CWh6uDQzu0uQSV1oPiUSNVseOeirDhd8UROjnRRHtAX8MxpSgmn93Ntuq43Uq3aN
YAnTfq9XG/aGFbRLS3D3wYmXwvi3BEIEh8hHVjB06hkbzUCe8KzlU0ubkqiQoPRm
AxiNagWTLIbNfZugbWkKYtIIIhHF46UIYBlPIYLnFId4Ew+8BxqI2VSp3gaxTJ+1
kStyJ//rRu1pmMy7uF7QedAshYb9Lk1Mp72kBk9CHKSStV1zpLYyidnX1o3wTsJy
sW96PqLVdvSnIPEZ+bBo8xLwu05w8Y2+AJgCnlou9gmGYxGeCf82quzeov9z/Oer
9qZ8DqsFmxFlmxo1d4MixU1Ij2eqKxMWBnfDWkdknRfGN5sOUHyLKI7cjgBa4Dt+
vSRYbOji/0riNqOTxWtzcPhVo46DFM+Llptg2eKRBQ6YuVGJryPz0UyjX8vMJmNY
SYhm/+PmxwBX+OXazZi99nWbd86DJTY82TlK0BlrVlFz6CQIWADPceDficKQ54Y/
k60SSBB/ttLNS9yOVCPodCs/m9CQPCRY2NjCQWoVJ0RyuhqNBFzeroRUZfokeG6/
DI5SrkT2NxWKN7sOFur6ZNWbSltwHYp6REulSlvfP0nIWaFwnXiybDGxmYzdBpm/
mxwEWuBVyzT/mvVpA7XVxi33DNJbFUCYNELPV/jFbRSHRwA0OcNvcVBoRKDYaw2Y
tp3FBNywR0x64HiU1DkTiC8ttE/SZz6v8p+bOwI4NhO7FkuxTFQrKbYLerIiJEKo
PKj5MuEhRpwwHHV8JbY60JGeP1ula3Vda+K4izrfqC/elc9NOojhJzyv+nCnmNnV
gMbkYT092NzJ4Mh97pe9WRUWJgXF8OqQMo2QTNHB9Dg/nE9LVXTn9Cql5ABSTeWz
2gbD5Iphi0+tUlFguY28UZnpLqV6gIXndsymHCaQ3Idi3bCeybIIvf7BIvlGA7nL
3kadwUInIxu4sH5PxtHdvIh1m5lYmEQONBxnLznhY+dXH74yOHCJq3QJRVtgIIY+
92FIVemK7OubFIofyOKyTh5/IBNXe5NZ/EqWazdkURBsGPkl7cSm9WoZK5KpEr0Y
WmAWLh2Nq0m8H1WV4PDmhWPbI2shCnzZytlvpLbWUWb3HpuDZTJbX9jRV3GBLeBH
6zi5I0c5NV9T/DgN0vc1h4iKQG6PJIzu6N9h0zxje69rhe6lKrJ7RtWyMVBEji5w
qWem6AWwDXLXdSePkxkV1lMJ468tFLHouQRR9jyM5M73vgrdRPn8TarqXWTr6Kyp
aU9z4vZ8d94b+O990fYpOsvY7az27tkuw6PSOc3qhH6HiF6959DNQBYNQ67lpIIe
vKOSHNSpFuN51ENqMdxMzlWHwWI6sfbwbQ3MStDqVdKq441cF5DeXDjiOSl5cE9L
gQdT0dN2Wn7fHg9H0K3AiJYc7TsSl8wA/DbtDVuzsBvphGtY/UDL5l0AJ3E6Uivx
/ArLDHn75WBQNZFxxjO31yFkacxOgKZKk3/QpbtgrOeo7OWUbWs7qfqTs8Sg7hmO
c2NfepsnqLIji9gjFKPe7SSD5TMUEAAwrFWU0QY+e3/tR8U5UPSa1o6LD9vmAPfs
4pv65aoVy+MSa2RePO0Zo13C9wVhsJEa2NKnjkncQ3IKkHeq1txzXX9bTeS599Tb
QxkbV6eI0W4pKvyDMNN1OyFwfYlASHYQkkQXM+t/gVvXxIa2KaV7uPKdJ0Jx8pws
QCTlKUuywRC7gx18s2Ufza46w81WwyshJbHASqbT0ySRo1lV9K7MiUGqv2QZIBaA
dSJB/FJ2OtLqt7pYuT4KDbY9sjxLdCda+0AnMfWjeTmx31P1sbtA8bmqSLcGvrBf
+jtLHLlVtzheh7DJfDGu2ddUTzpbcYtvEAVZSNM2Vgiu0/ocOvLGemucXEs5g//G
WSBsFwoO9DR0nk8k7mOJB9bJH+NW9SCCkXoXX+b0DqtMQqrG6ZOAQMWriYEhc2RQ
Pm3MtK+2z3qwKfVMPTwbl1+RAbrD+3fsD7NGNHbLUa6hs17mHC7o9G/Avh+f6bJt
PZKoINXsbbz66K/zeyBz+OAp2qGimnJv5py6SJZOmGpP5o28iEhczOsEE8O4FZc7
ubsxVTGsrWH3F5dh/y5Ec7w5BdhrJB5Zujfz0dzpjQTfMAuorXATZgKWOgwWu4qQ
+FpB57/W9ZKsGFZE2lvQsBTACJ6S8D2BPU7dQxdIsqhyjCRTvpgaAZxACR577P7S
ekuvt13zfxDQvmAT6QkJi2gi6Uas3BI71yXI+QAgdC/pLCGVz3DrSDzd2pUpyTSu
xOugL8xAhVgMBVV7XZPEn5PnVPExufw0Ay2ZIIRPNFhTKBcj0S5Dg++otFK7FlJ3
cogeTU/rlG6uU0ZmDwKnT23O6KDoLp3zZ+3mZBOH4Lu9W0PnNeROkkUvMSO1aW1Z
euBbBnCT7eM89Xy/ucqm5nmcr1Oqg/sHZpzw+bbWKQeH3/AjzsEJVPIknYDzDDpY
i3pGZ/Ecc3Q3QJ0w0IYb8nQ5XFz0K1quJCDmm8E/cE6b2O1xbHZKDgHOsOihZl8p
pXFVddjdKr0SktLeDHl4KT0uuogIcK0l5sEk/AeMC7A6LlJO5csWls8S/VT36+qj
RVaezDwq3ExoqJM1oP+uizdYFzJPSzVyZ1b133LJMeE+yg++QMgxDEHOOMBKqBcC
+MtVh5myYahz6yXbEFgJdOcd43ELKgyWN6fLdUh1kLdcq7xHhpYGqwTS4cwJlA2s
UFYNz/0BoR5i5vgrKgx63ePCeUfxsI0F2qwnduidPGxcjG7JE6UCXIWPJUuvwYqr
X1CSXoCkEgCkO/kOgceLUvMBDeo6+msye0eLD9qCx7jVRQnHsS910oxyinIZz4F3
jQn68Mbg2rv+ksWooH/4VXuGKTfE85YE1WCByRaFogG7pwKF+bOYNhdA0maEzSUl
jZxvzg3MolX/dOCCaohcQywJBHfOYGEBecQKcumsVXACoC0oZX61KnGDjvuTS0ys
FQuPFQdb5jKBKwUHYVqpxkNt2zXnbBpBDxnJ+4+2kjtgwHWv2WByIAoNEGZHQfV6
2EHQtQ13Zt7jWjk9JzsJuNbpuaFNwS/wo2dZeMv9XxJ7onjGWPSHLup9nWqUUS37
rVCZtxmtpqyZPmPTb899mhFgD6EMW1M3665MElvTbzq6Y3RARLxOQXBnlZ551W94
lfWX/4t6l9g9SssOciONvTZoLSRMqcOUvwVRp/wWSqPryQ0WlTOYVX7S+ce5kbyM
6T6VDmdm6S9UFrH2z6bSN71+Y77wx6CpnqMVwLI8cG1hVX7rMBZlsjRk2FyTDY89
nM9/4X5p40ISltrAuQa573Ad91bOANgQhR7/XUo2VYCleci+OQUhmTJtWJd8vxon
QE2zxB9c1W5QYTLzkFKsoxiRLKK7aZWoj5+8cLFRlYBF2mchqseBya6xDdUrBjbp
KlAceD71ysUYotmIPW/KRvlGEnQU7zXIBmjGOgfC/HO9j5siavUFbJdaIUCjWJjg
S2wB8BFuMDIe2GFXUF8h1kDiEW6DXwBTZ7AD7iF/k3NaAvedFzOZ3iq8Beeqpjcw
fbf7uFl0NjhQh1JtCbnEH5MLhStQPuT9vM4rXWHj0mwVJdBc65pcuB8qc9d9zMYF
Zjvo9OClQ/hzr2YKw2RHzmkypV0VdqRtkpDZZTA+vmR8Vjm5n7XGbyzSYUC2NT/h
osDw5Ufd4Mee5C8yt14S1Kui0bcHL1fNHE3gY2jf4F47J7BKy518neuiANI3JmPk
5NMB6105Bb9mmozYZonlT5WahYq9vn3e8HYoR5cps6smpP9A3N5tS8mm4oLlCotg
r19dNdl6Ext3XjqRLSxykX5x/qHYWVjRNiEekSb+SUdWFSJeZG6MQRlMOGEB7YbG
kLbnxVnqUV39ZE9PuMWVBuMLP79RS+mLaUOycA12qNNjhFEyHfdFbDRDhEljjTNK
FwPh8vED47Ix0tGRUlno2y90SEZJV/AopgUNRaoIgNWNFSQsb8yEngvT/G4weuZl
Vbhd9jaVANhKrSPMwQ8DhZnaPeERH5y8WKk5lBM2v1vOROnf24W4aRKUS+1DnLNX
sFJLHbGXl/IOQz/Ob30eCzu2GWf2ZtG7BE5+vcFc47blCtLgp9+r1yDCuIfEghzM
pyPJGPH5xGs2DvKekt9RMbXVklFUAGpI2g8QBhkTS6CfS6O1XCh+PQNJoVLIspgE
FxZUL5Dnc0hcclaZfEZ2utBE4/r+0SYLBk0m90M/+a1d5nwPGHPg9vXh/khMWvI1
x3hIHpu5irMcueBKfBNl6E7yD1cwb5rqmMO2cKKSdTZ9TYwxwPCFF30nSzaG0PAw
kg+jElmyv694KMzYCpHHZIVonqaaJBLxGX1AF9OX/wNhlpilX7bR5N/9ng8SY34K
IOkrTFPez/lBM54koK1cPGXwkVrspgrwZK9ZMvSx6uypBQAtH9q8zTxUQbq9SHex
nNm2sD1aIxlSPZe7x4IXICfeHanmK9z2KE2T7wURNa8nveYO0j5QfkmcR4ZKtZOi
FAKAbjuaJIZE63epneLGCwwhf8Dv+eGHPxdnhXGgza7FXxm0QzrMwZXwZ3W6ax+a
aIoxtv93Fdmmhmw8FQRJ+ZbgXHned9XlLFVIfA3jXw5sy562k81YxqrfRaoVQOko
6np88GnSxQl2WI4XQGIzK6mOfY/XDrkCWHzXyppEVgQ/hHAoUYVINQdThzytWWFS
e8hMikJBLDlX20hRcRroKR+LblYc2ClFNYjkSMfArwxPuVGSkPLHw1KMUjGbR6t/
iATIULoct+hwTsMy15/s8yI54TTx8FEGNV6gfW57Nopk9OrUBMxzI0hGVjhUwNjJ
aSs4jUPfZOhfoYse0WgDcLJ9gqJQeqmpoTe7/zD9pzNaX0SawVGyt9fQxAxSri+P
6ukXndNT5k1URkQyYm06zUs8QNxBSYpX0nqb2xKqJ/C7V0EBBcZ/pBqJj0DxqHgx
9h0vulPqfRkDKoxrOdkw1JJ8WAiGk9q0Vnkh0vhppIpIsRoUR+BpwAei4UoiS+Yx
b5vQ4PaaetlmDON29HLnvLVpNteqtBf8aPB09XJ2jgHAb1naeBYAcK/nO1ZgcVBa
YhTImrkJH9Sc/5q5vntENzd170IbbyNwtJyKcknixl1gkCHaRl55AEUNEVwOKXJt
CfuVVNp+9VuhYyeCGWv9JZrETrVE/vS7fanRbDqVR0uWqDawJNXRIAMz/kiIxWmH
yN5vJ/+lkdTylYVNGx9iWOo7gDyjpJt8EkaOu0rCN/rbDFgkypYaQi7V9vcoLNeH
ELwMgT0abVIewyag97sE/kugIYBB09ZIisv4MFKYXBkVYTkL+Ys2xLA+5+JrJFyo
awQzefHyz74NnXfXVsPv8omALlOYmT/UA/TAjTfwQANuZtJZIKqet9z0pAw6+EAI
oXib7BBHXVTtLaeVClLlKLCcXbIevbpQt1DaAr+SFLQctlPcMiXx3ZFeohwhZWN/
wwGcQexT3UpIzSy4MaXJKYkcuxrMWr4ONeJbxArXL3McCh3WjSe7t9g01IxR57CX
HZ37e4M6t7MuZJW8Y0rNCLQbJxgRhVwfk53pkMA7xnSZzwvflDGVrWjKP5vXUFiX
HNz+9a00jV0ud4Z/N3DGhq2c+uNH30NXPlWO7FSRoFXY79RFn/QJ9Wper4sO/Z2Y
OXuZulu84N2RJee2yeigw3oU1/IAQCHIAm8gpcAir3+Qz+Mn1eF5kfbB2+delocX
trJHniU8JZSpQ6/zHzVKSwfz27iAaP6yov9rB8/WkDNRMElIkTy0Lwd+I/sLckeD
fCuEv4ktNsvjGOMEeoILCkJCoJG4nARH2N0DktVS4fT7Z2e4XwxlFEqCPMVyjVev
bRjBIfWOP5Q5o1aE6wKuUZJmZmwMH620XDPV1RBKeLUksi/LJN0vCf0TZoQcswWh
/CrUCJCFDbkW8zEiU6/030IuB7/HsfvdHXuRUdXRZ5Q20rSW9lx8EYbeKaHy7BsU
Tzcs9A2HvpaN5dJ+pCCvjowA9xeoDLDkSFa9Cx4qhpcedw3H2aLr/ej66vkqKcqt
WFaJBoOXg+p0gHp96Ppz+DPt6STl3Q94dQI8XCb01CihEKanj/H8ef8DSHFvfCl4
TkghA0UjxaIEa8gilahmVxGtoNa3fApv+URx3+5h5j17+CRqyuR4hWsMBGobCEWh
YY29H58Fu3yrhfkWJRDvSxGiLU+ZJ7g0t5qix+5Flqhvkt7hweNDKyizETJ3C1YL
8aPPXP+v6tawKki1jOlB8SRZrfwk5GK0HYBdLe2IQCujCk78Zoam88XNzcR+tyzB
mvva2/eS1cpQOvlX7mYYaf1qDbsvGKP3HQqRyzXVoBIa322M1ck1gB0COj8hSM4U
OHS3mEQmxywJwIKypMErY+jc2/5k85VqcfkhUHO1Wq3hxmnT8aj2CFPtLrYBWdEd
WnMmzDIALkvp1QNt+y4DAJARqmUCQ8x5/UI3XIB1B646T2vvbuFv30Ajli8HsUXH
c52aPSAoiu83wvhzm7b+TDQU/AUBRYWgRTNvFg/6TM5TDktrG1xu6t9A85Q8lK2e
TOmCucHe/NvI3cPuSSgexK/lKrJjnb5YZKrVON7amqQjHPp2H+X6FsJDv9SRaWjN
NRIUpiLCOYeOdZWrF1dQfugTXL7HyU8VLhu5PF+S7vQQJ6BkwoipNyMRXQ3VrW7q
pAEuLVSgYzPm+A7AMc90Y8KXVtgcITPljxz/JyxltwiT8W4IXLwsLBtUhda3FFVY
9m9ZvAJ15iLB/baN533MLEc1G7+UqWfmlMlRUVIJ/c0frbj7JoUp2noYMkOVPg/1
vlqsqQ1BzWzgsA0Bfgbf64TGV166ZWKkbcThAen6zlKc4AQ3bnsXpxptH115QvuH
DTjRrFAjE43wMhsOGxyEpvIdK7UJu+SvhvP7STYnPOo81oWUEHrCKajpsdgaT/zI
sMtrOy2vjd4DKiaBAtcRiT2KKw8tLUeFoKVONRDMxrNwkUWnaIDPvxqVSuSrPERD
glx1/FvXaAPzRhD6hohd5HHsa6wkiLs7GCvMpEBi/NYvAEB/10Va4VTbYETxU/TL
72pFsa2y3jeDmoQsr0dGqMtF9AvcucNU+mF6bkMZ2tDx1GbZ51/wKeLKVLlPGHmS
ZtZ1KJj2IJ6THCRnPMqvlsPUA7ygItp3ssrIJ4kV95u68ywFgJVd3Htf1jMvoQ1X
AqhDopMQLCMMpFPwOV84fGIwYoF5g9ob1gEm27UYP1J+n01ecBisXJABr+s0vJKC
Y7RottlTdRGBuD+ZilUh1xBeiMlGXG0n0uZcrTnkthRVp8zUHST6rFzGdhnUoq90
3ypQkWLvmC+petXchXKe3av2x3CNi5uit9/IKYYxee8s44nK8uDpAO0ppUWeU4HU
JPmX2uV37c4RFzGkYqpWJ64d+oVb6kmTMUL8f5FpfuHhO9zdTm2P9jl100oarTZX
Su9hBzdFlKULXY33yo0A4/7IPtTUb6QYnhMonN4ozGQyF+MDs2Dnzm/o7iz+ctwF
6YEgbHWtB+5CVMTLJjl2hoQXnfn5rxXf7Ct9WCxig0uiqf0U5yWMbSlT/Ny+x/+F
SMk8Z4tMZLUWS6TDfTrc5qG9b14+FH+FVY4BJc9NqWfQ24qLEoyUYEAz3SDqSG4T
QXJj8zJdclTtWRyA9guqdnolBA/pJkfOnp1ZsQ7cVUwioaGwQwiEXjx5tO7vfHZx
evUKttvjPcH2NfNlYTpXiYL6QSfWyY/Msf5UA03GVUny4dXvAb/ak90kJwMmb9/h
+8lpKmlbrB0+ZqZMnnAseWRm3GMvjSx/igmDZY6+vMjvFbDUKuAZhcjhaOoiIO9o
x6BeyK1WKiC3rlgQxgHPGbQs3YbEsf/FtDuF+G62SQfri+lRFCfhBoUh2C7BetOf
QYPzAmKgZqy0Ava0CeqOu8vQGAciLVGlQknNP+Sw5I7JBX2WkgMi4fsj0fgcZkrk
2aA+5KWj9sJhBb+OeTTMOh0l2JH+9Wziy/2YS0K3CvGTf7DSh4jAfkFOBAYH0Tg7
4kOVg9prfWy3isU9kDmJWEDEoM5vRKvcP8d69CexXFj2a+clKixE1ghM7IGilPVz
vitqZt7hbkFAw9yxZQZSWjBYPpH/ypw/zRp56OpuAHzm0xVG7DX08CpzO7RIcD4N
fu6SoU13XlMY6dbqMBxquUYwRojLc96nPyPKL0tN7W5LGD40XS6gHQ9CkltKCgpS
HPESwx1F/rSIU7HkY8DGNZ2J5to8Nca3gCuc6GdkFnhBJkEGoG3KpC0ABMARMPOH
hxMAs3xpR3uXqjASwpyO+TLewkYXadArCLSN3wbmi36NWAxpaQdvbFbIjwmhUsPD
o/W0iC0GOeQGP4j4C41e7e+EWgthM+x1NVW5m/iV9KAFJGYhhR3OzaKO2245Kbkv
E5gpQICyjDPMXt8z9r0RtF2tCb604OWSIwwo09ydpm5FsgEiNiisoE+sxXwrFHRt
wugTO9aN+vspGLMKxI1xb45scXEa7LIKupfO90z0+ynE+/qbNKEsNsP47GH9oPxp
ET4gqjHlMxs6i9Qwe1k2UByGpNocDwo00OR/rxLzrtf8frLAI3O4UoeqXt2VNgX9
YJ7k0isorA5vxPciRkRuH64BJhTeRjo+txrLNP7xCPE5MqQFKNVDlqH4CUm5flNA
LVocRsH5Dt+XdsWsYP9ZgUdnZkiDVLC/OIZU2ZVLXrZavM99pRroXJSxABuhRKly
l9bTESLPm64pWQlN/fuBdRDkjiC/wTsJfl72XOV9dUbDkmS4c0qCt1/48cDAGuRw
FR/FRueXwPTvlSKdO4byhhKH6gumt5/D8pAnwLEdfO1trlG5hEp9xY0Kukqg7AoL
95Rq7mKFpHdUF04O2AABuZFzphuFUdudNlcdkyd6a55V6vg2ZGDoDhynSzZ7ygNz
IX2T6izzKOGAna2x9aokQ2my9nJIVuP9f9eYHpX+6cisIVCARwV9TVeoXn5x2WvL
qAVbC4Xqh8d83f6ZEl1R8TKed/bsxzSuio8ImLJutG3HXEldJZcq6X42kCtaKXJi
ogy7+85J7KV2NZ19Gm2jrB8/elaN4hFdAaaWgu1obohSJkTvaA7eItjqQ2ck4WJ7
M8v0BsEZ+SHLgpDIQulJMwUSrZl85kJJAs2qe0wcyYhiyitmCq9LuM/lo1+oOcV0
RkTqKoWi6a4snB4nj6MLXIXUCbSU/zJOXe0BGLQbocsyi6qnUXZwuVrkxEAhCh1C
U9u1pJrBVR3B+lHMSFGACWKM1Fhg9Qhw6SpcbHCGG9WAxENmITqWLMw5mjsM7btR
pI1/2U3lWz1I+yVf+Q3MNO/A1OYXx9RRJOackGVhoi+tTH/rMFsV8NYFVJR4Y6ZS
U2q1y1NP4RAgXLnEJk+zdT/IhWNWbA3mStDsb8ERAAg5T7LRBjwNYbkpJoLPt1Pd
CqUhyyoB+CAHqvyMM/OONVKtyT/MoSpCN76fmaPY4EjLYnHL6qZ0bgKA87PXNKzA
L7oaKn5AICBthqmVQ46v0KPMvneb5SUjzO6GVbFFkFHifqTmjmR3rtCPbuPyG6Xw
QhPUVROzYNwycUURqW/cijkfig8S0e08ureY4aU03rXfOk0QpVQoFuAdi0Z5MILy
PQgK5uhEC4jXTFEZSPvre6CfYrvhGa0Z7E2gYP3MJ9E9TgJbJ2pnuy6egjYrJFr6
lZYQfsfmC0l5JsD1zONmRzaRgyWev4+DFXW5BD6EZdQI6HLyoVWORIHABkIb+7Ng
0brYDqhDvrzJFtiZqp9fDKNLvAcvViTWy+UhDC+moIeERkp4ADtOuqYxose8MR6f
hbXts7koqi0Xvw8c7bLX4TMJZ8I/pD1MbuOgV99XSllggpqIqUKT/UGfTmtoT8as
+JjtPEPha6Pi2thJp9zQgfENXhsBeLzqX5lRMg0H70HI2Kc8z9XhKx4A0v6s5u+Q
RbLv4lq+fnRmcD04vAAVLPE4hELjEUibVQEOz7OetcMzG7VQbCyG/UVCVN9zhYCH
O9kWlph+jGTkCcFYCIx2uzJjkk3lvAWEjqxncu5G79Hoqruc68P7jY1GVTkwzEe9
0wmO9bWmyOqQ/DcSKCXA7yS4KvyGj8di5bcv46ViFBHzzbAG7M79MNE9fR4yttiE
/n4PLNphdPvb6qEn5c+mnffpLtDnawL5A91gqgYb7SogGr4Pryv6KkFOcsyFGnz5
odi78GJp3S8U0U+wKOV60cpLOFqn+bK4yxlXJz3b0NUZK3Zr7TuU/LPCMLXPcQ6O
XHVoFiM8DLu/FrB6kd9fMdbTm59vI/JGc+JxwZ7RAo++vSvzb5HyczU0AWGCuwBf
nRA9W/AAoUvgveZUvw3uRpph3AbsDtG75OeSOQcK+tF2uPebxZYCgygmCROgPiUU
V2Jk2QPvpKIK/nGGqD4xKdEnEzufHWbaFqpiRKCpILsjSDnsfspEJ1G4cTtCPWa2
+7cgdfQ1PD6ZVmm7YN2BZUwey7BPR4THE2iiT0asBrbhbU58GWNTMhxwFtCmeAJF
bVni6EBsRGzthvuIxkz/3+MNXIrtKQThQQcFnM8MeTWaGcok+dAHI6A8UyX52RtQ
DLzW/Ehk3yIQvUDUQbAz0x4vE6kNdr6C8nDRYNmXMTCzMs594FMwQmKz3RlltEMl
AFhG6aNwqE0SH+bUaCW0owJJhfpsemInmlrqb+MjwkF4bu3LcCbTEZhnB12rYoKk
6dnugcYXtI4mQyTVUmt9JJcc+rTBPgw48rgXp0ggcARikKV5+dQdjkFM9eesaDHj
/ukOickrCORnz/1wxPwxCkGh2eXulzEBf5cbFJ+V/IQsWvMmzRbUIgKOp92ZKLFa
aAst2ZmsSM/OsIVQuFzdIATyT/CD5HuGO381Nwf5KcZgQwszl2Cr7hH5XOQDMVYc
BRnXTgMD1SXm3RedlVsJkEu2bg43mUBOfh0ghleeTTv2Gg/2yiu3D3b7TZRj23Wf
DnlT12+GVvtkafk/ZY4uV1x2p3DCykT7Zx+qAAzRW5VoH0oGIkJxyugRKu0JkIkp
IcHE0eQx8PtygHO8vdPhsPkFaSESRTBj3u+AMIifXk3+iUbZ/deke2p2l2Dn8YTK
m52VJaR401QGJ+rZfiD/6PUE99lNwGK3NgDIqm2MwduwGpVQc3JwPbJ2bUOClAI+
2ejmXy795pvZ3tgvQHMkalfbcfvuHKEyy3bBy+mbN1Yrc+LC9LXKuODJgJDNDCBA
arGxEO5YkfQzZvuXGWy+sEdIaWDLtBXWGwurkwtW9sJM1i5evDXVYdJBDEv0950f
jlDGWLW/EK+vjjA1hhSUGxLjnV1f3EP+MhD0I+tVQsDw8Gr2uoNx+IGpRS6ueF7H
doSzWOdZOldisqeg2Ow8KjljJXuKCrD9gUXXhqx+gCwOA70qeZgWrYIENKBfa3Z4
PtCLGQDj0Dxs2+a0IGlTDgqfMKZut0AbxQq0/LbQ5zYmjtDmf+9iBekYJ4IUn5ri
fMW8CdNjw6G+4fCW4uv1eQ6Hd/Q/HgEBYOgSzGEZHn75gOJ+qGfKPhNTM/Ucs5ss
5A2zpasXUlYsTLdbPHkEIf29qp3CwNuRPH5uZcfAoLy8LOPWwNz5lQgHDCgSwVgb
ODFJm8WbJ2JMsOn79budyHxF/kYjYIBoe+sjJCmJrkJ1KwMLeoqOOnKw//aRQrLz
D0fuyhv5O7/w9evIjxDJT5/vRSVNaqQPTv+GIOiVs3RzSROl8vhPeKYL7Nej1A3a
6O/ZfKaNa/rNAAWg+sjTwSNf0Ti/+XdaDf/3p301pnPamLl7js2jOH0XSt3oVivx
rIbCAQrtASK2Gq7147SHyzhiDmkdrdTpXE4T+i4vzKJrEhUyYAqeYuLmNaZ88o1F
lIRHQ3wLVjBwtUk+2FeOj9ZSiA3/tc0WPb5ZQuNSGv2kvKytY4PgOhYVRvgJZZGb
icsIbSQYwP6udY3XiQNAg3Wz8ZpRvIjYp1iUwpZeVmGmqsoju7yfPy4U51Donx4s
v1PPhhmqCNwJlwt3O1HXLkey4Bgmr1bvrIDrSNugewkZ7bRMlt9BYt3Yx4B1idCx
MAIbOgmZWKqRlNLyHprXwkLWNBWBNfyzG5uF+Wbs6O4+WGrJsbjogmfvG/eT9iun
VUa/wiL+nOhelSMszMQIzKraFM5JckqErqPA9H0HMqtVdmXZuAarYC2fRCNurtoG
UWm7qGvCv0Mr7P7GkzWL2SHwpmIJbJSAOCVwHosJsrSyFvoiWeJSpYr11YSRumWw
7sYT7NblG2TyCo3AUex2exQSHb+ELPI7kSRyJ/si8HD8Zjr/4/VVMKNL8PXAK8eo
ve7QL2BOfJHRfRC2bUoDsmLdMrZ1zTkSsb1jls3WKT1Ssh30ixffgNi5obRwU3PR
lMK4Tbzd7xpqx2RjFinmPErPplN423qsIi7+ieqgkTKI57VBIr9VDmkI3BxitnYi
dM2MoHQ79RtVXhaPz1+4SfvcAUY77OKqUfat2Fwx00+b/R3gFo5xsJHrGq/dThEc
TdT8T5Q0Po4ZumG344PtuGvCDV3vfZJ6e/hQJbPGbUY5bV63tc7tURurKaRDOfgD
cQzOu51RFxhNwEK1TIIGDeK4eCSkhnrk7aW4l9ibGzZGyJ/oylk06oojE485YBjo
6hf53CZXaY1/TWJ2IkDd4SjFa0qdi1e80iPq+IWCyQxEoHspXyfc0HpUmJRzzEiY
auraVULgrdcO6OxVEbak4isbUO7t7iIz33GHFqdCAg4O9YCeo91Xrku3Ri7ZmTB2
MOJIxLvhsOsnRwcqhGd7SWmdiOHbdupRlw4jyJOfWIYjZfA8Oiu9kbwLpDdahsLD
8vGGJoWqtR4/yE4f+IQi1VW9NtNaXCrArXzJJwUoa0LTD4yBV3NBF0z4Z61pAA+/
brLz+BNsyMr19CXr/pvITbVP1rO9lL5kCTCTDOd/x+OmP/1mk5/VpT8mczaSC4PG
a9DJq5sKNiPmfS/3l0teoeSSrXQQ9DNRQr39eRDfRmVAmOlHhLSo7j8iQJcdtKK3
uycBdzQse0bAkLYw1wOOgL+rtwsW2qGEYx7sdPJH7C+33YEZ1eObJhEd4yUfF7cS
tVFcVo4a1Uc3QNeryf8imbB9zxDfb+Ss2rTYbZpEy/VhZS7rfbBvCJ21d405Z6Lv
X0+/0NFDeZoWtLZNBP2FR9iXTUr4eOu6l53IXsqHaJO6zF8n+vgP4qkamZUDMJPT
QxTeCa8eaoXMVDqoVkQKDpiq+wRAf6AWR786VbXJbHwE1GYBWk7XdQQ1h+O/XX3L
UAVJ/4wbSKk0fcPi1gUYb7AeNVnssFaL4hnW/DdgQ7cjSz0rMHsOlG+c5k71+qas
oeoAC+wPoAvOjt3rp7OPZO5CIYwd9ofMMGYJJLAxOnNv0lfyrbjtwouENGNATClY
KeQO9D9TkvzB4Yw/vqKbMDE07SpfoOU4LBqqg97TDVxP25lQ27f/ayDTApJJz1KT
mkKOVuBcK4jL8y3KvcCqVQSt1LYtSrEm7BHrSyhRvDf5DJaLnIkHverdnd+Cy7SR
M1BfnU+Mi2bmIbzhuxEQm1JvTmdrbzqnreoGLIUkJrNbLWm4lEYY1FIGLLUGVP+N
Sr9H1f5eNYCqrvMXGIY1OKIX2X9edbyXFfqku5pILCIXrbyanVdvGBS6R6zKcmED
y+CGIOpvBoIO+josNQo3EUQvDmlvWzqKyydZO7bmB9VPfn8ZZSeoZYi2U04kCKzb
1ETb5RfioZwbOalReNkkApSCsB/SjR032BQU9zm9dbkbPP8GIBdxpqweJs7Vh3YP
xPVKPH7o7uVtYwRlA8YLGZRYV+8Fr9Ame2CAas3hj7KTV38sgN8AW6q1ZJlimHVQ
LnCBIpxRUdFmmoGLYU03T3/BdFMK66IGgvyX84fx0CWkcGjGiXHdcbL7s743M2X6
QtAb78r85NW1oAns7DZfmfnxKROa5YrMe90kXBma5gl96vhrYzRj/qmAEa11vb4f
hY6A9WsFaSgvyAXpx9/YTUEbeSlJ5NWqBXR4ynmMk2s7sEnxgpXps//bFrKAL2HQ
rI1kEW1cCfxesABd2Z+JQIa4V9vg4DYoFEeegLiXat5ynq3FQiYHbytl4XZtWY9Y
v4yyMaSE2yVaCLPaRwgmTda/6pKeuBebzvd92tDIb8YrniftOQ61260KRuxfpxq9
b+o6OWpZyvbbYC1TBjEj0VSBeccWUY1t+hYXDUHYj5PXB9y572rKpjb/ARbqE8Di
PgxApAoi8ViGSG3igMY2fk2VJdMDk35LmpNrrKCXT/sAVHDxNvgwdVvYQ/yIEXR2
nDbsachte1OEFDkyar0xW8erVMjHRKpLVZB3ySZxubnuzAaR2LcKg6uTkpzg6OVn
EowoiRNYV+EYdswIhkjVALvx0KTYWcp1jTqEdKkC2/WQIYw6qf4BOVhzISksAXwH
ca4PQEavGHiXkKU5gsr4wN0cDV1+Gy01Hjxm031nhQaGV7aueRYoopG0fFEy1z19
j8rBSglfnkliUG/ULvsPRAv14tHN4Mkt4ACs93RDknYIsUpb0jnSWYjU+8VX0rFs
F7Mr0sqrw/qw6ghWjBLczD6Ocmnrqq927CryUwt6c3uu6q+dETuqMiCjrCJeZTui
7wYOaaFi9FYPl8EfEXPo0DmWP+vyl2jTl4rbF7Fe9qLL3kLoyXhkkKdFtXhuQXhD
uT23xbJ0nCjCp8GdxKuMBzFJChzNF1leKLibqTCM8AyO+wCxjC2xXJlmxJgMoYjh
0spOdvkiTucZpP71w/itHQMPeNUnQOvwNmEkfsRl2NPiuDjF7vidvwJA9fgQCXEL
QLHxzhVD5wf75u5Jy3DQz8NmmQWQmj/NCN5mMrMtZb4W/dOq0LbFjbIs/zYAuYKN
FKR80qusr3oE9TNzbucBUCLYjh9kEWXU9P8cNb+OCLW1oQA6zstN59QqjicLTuIH
tOPtqTlhRAh922tQ6L8u/1wyUD4NafJvOykBQ00fsQpwyRS6/kap4gHoBsy/vA5a
ua+z3/SaHiJAlyjv8llAYE4a6c7BEMhcpu48qwfAfm+QrSakn+Z95eJ5ONlrmEBg
3W3lnXEIWAq1SpZh7aVG4eylt1Zvjw1KvBUzBlTSCjR+rPe5D6JFGpHSHbU2OQH2
+VfKS2YSrnh6Zqt/ryDl3EI9PMBiA5b0Y134qmGGSl4go0gv2d81qNwS2JngHBB7
FwpWWnt3HEF4YB3jH2DT0OK5RsKrVBkiAsPyvUuRR65N7C57/wIsUy4X1xDtJfiv
x1vbrE0c9tKI/E9Y0ksohuk89jB9nPngazk98lHaO6cpgJjkr8K1/I+CyZu7Hgoj
YhiERZ7CN/Kl6TidWQ9gr6ukLWxeKzKYw0g8dB7ayUGQncpvko/G/LvP5kZstg+g
BY956vwsZwK7v3hSrKr4s2aOPHVLcpLChTlliSAkQ4xMjLQ/5M+NQM4+0FNamhyA
CDlhQ2FtEls6IFy95fSUKsT91fWBszsP5sIFQfOyCCaEdorLP1psFHhGgq6ooZud
Cw8iemKKk/Zw8IzgNz/kdIGH3ExUj4Qhe9KTG08d7T+9rUVoas4Vg57z+gc0Z1EO
P/dFMpoAvjF6b95QhaT6/l/zPG7APQSTMqz8TRNMWKfXQ4xADgu6Xmx8EVrCFhYK
iL9SArGpU77D0KgEOjtwOs1iSrZi9IGyKhNmdUdzooSnWAM1v3NT8pk46TjGd369
DaADRZfVaMwEj4UtIemJAljLwwzmy0M3wc6guwGvX0ToZyp473AecgcuFWSUdLIw
7Js49tJtvZy2eEDa6TJhiHdn/+PPM5HmXDptcR2qqG8UMgpALMosCYfCYUyj0029
k+i52FAdc9qEw182xXwNbr6sxczoioRAun8muK8inLq/3RvokcGLVK9zwfmM186B
jVVcPBPJhp0W+6sp7nzxBOYRjW7vyE7PhAH7g8u3cttmn5N2etbSpfkmwnWuON/i
RjgU4Ue5wYdXTy5N8xD3xpzc7W8Qk8biJ3xBG3iJDzOps2xnR/24lFiy4z4BRik6
NBfQjzsJk8vE0MoBkX3ajfxJJxjRtHNb9bz6AaDqGOIXp+/21kAoDVAeU1/aQdRr
VsUr2RA5gU1/XzfcrNjXr8SeWLfN2gVqD/OAIkhY3nQtq/cVXFeQd9nfGB/3k16S
+KsOFzX28PqMf7bawOhE34oAf11wwT5gn1dUu8qsePcJyC+amrOB8y6YxoSGmzDt
Cy0tqJBaGdG14/qh/1WtR0B5u1xbe3J7j3o5y3ElhyvrsFAeMuBS2KwaSRP0q/zh
/Oc5XeqTo9bJDNehoTpOXM70ALUHXtyhpU0bIFFDoMfuAk7Q9d8cPCQUDkvWtPKa
dCPOqADuoFUVhYf6Z9CpOs4uubwuYlp86SO9KlZ5wKtqLcI420eV7bJzOTfI0At5
aPn6q06mjyywq5xTf4Q4xttoAjATO6/wF2oWNrDatL7Ahs9Q+9uVb0wwE8s9IwY3
wkLVVUsto194uCS02FQxmrm3RLbCjlZY+oTSsjw6W+1QaIMObU/gTFNmlqDlanU3
aP6rfYtIaVntIKTz5YE7gs0Eo//DjZgTefFiaMzERwK8QNhu9l2UtGKTuSkot8ec
xU7Vca2U3TE0RNe4ivsaXruejsHIHrTXN1XH2zjU86IxDk+wcNBqT88jVwmGAduQ
qPGx+g8vtQB/4me15LK2bI1iSlvFJq0vR6u+jTSvCUw/R8Kvm3vyshyPJ0jmPtb+
C74Oq2OcJvIKgmBzR2GLzEcTw4Nc5Uko2F80Epf55ou4F5nBw9K+uuenK4c2LNuX
gmiAN2xtDaYvriw9MeyBU8q3DdXoUVDGSZClWauRx+yv3uHqBRsw5IrN4TvxWqsj
0TZk+J2LZdz7PDflBpUJQ49Ov1OWPVcYpVOedfKLgC4j+CUodn+9vcyZmbVXvxf5
dPlH642Jxz83wXY2vouG0LvGfJwZXjnrGmgIyt3t2IpKHASl5sf1/IGFZWS9vpLd
yN0HEWqLuQFZCVu/SQvcNA0eUQU0YOEhS5VY81Ed1UNpxjAupQLeKt5Oamct4eR7
87jdEWzzAqki8dnF61rsjl87yOJC583cWI73kWCPOJkKrpTL4KTG+LkHb+2S2cz6
8kPm3zAldus4/zGk06m0MRzGcp0sAbPXUtECgNX8Dv68YZyz4e7eay8XkAnPUA30
6WbISz7mzFRdYhVbUFwW0fpmfoCshvLx2Yq3SJ1vmKyruoXq0V241A+2NT4WvQ7b
MzLvsK/Uau6CuoTUY9/Ke0DV+z/Z9RUAuzB1PU/nt5WkPyBqwpoAUeoc2gGM0kFi
s0RoxrNmicgI6e+lfdhOlh6xDBLQbWrJikrqDyOOlboLK9eUOJ+krrfx7EFOOXUC
b4OdbBbJyw+Fzxw9H2gnH1OaZdEyvyZvQp4Zn2QGZqfY4d0gS4FlUBxdeFGToYPS
1Qwf70hcC2frZidtNgq/T9vXyZPgSi/BlfJ6uiR29+FCwSj7Iv+QKjEeqCrbL16k
a1Pjfoqu52D3yPSR9xvMRZGnN7V/eXvNVhLlW53lQyriZN+Won/wnnblIKlZdH8c
LVMxz3gnkT5o64ndUGwK+P+3Yjj1H+iyHL9sUIhUKCaRNVzVuwZfF0NaG6oZduHS
7xQqoRbn/BleLcXqKt/Jhp1oUQnlZyr3f8jmKnBaDP6oOmvHCuWXKNQbmWQUg3Om
wLf+HI8HynH8LmOFw+Rr/so07tGhFAy4osaiwPBoYMf4YXC9dmWPm4OuJaXUYI7Y
p8lC18dB1qROONIAS4F17TtehPqn+Q/k4Q6oGmL4z2dCnmrLdUpyUUihxiotGP7W
jWyC2xiJdHvlRUtiPWhcjkkI4i1sDzaskvPHJ9EJVB7XwUXBaoEKJf9pEgXVJn/Y
LQ2pjAx0heAMXtAB78ZewUCo3WEtP0uWJ7eJfD4uFKQPOISjw8GBwc7Q9SK5LIBi
r7oMT9MLlCZWU6ASWuzmZOgIuzaA4uTvEHy4icW0Gd885YEsyUjjNucmBgwGc696
LJVW9cXqMng1Y9k2ezTvLr9f3RUb3HyxxObo6BstfoYXvY977y9fKdF8By2HhOqi
a7pks9BK1rl0XKUIUzLCijv427w1j1zDNKAVxqOxHRFxD6gWrsfpExcouArWGyTd
no/AFd3jSwK18JpTZnIwID7Bp2mPI1Ubozukntc/KNzIEP5uKeEE1LPL2N4qtNmp
A9wK4o39c5/M6KuuIPRvIOMsD9sD++TdFfIjGnAEh+OG/sbNhi6Hg12lirML6LBH
WWBYbk3sSAuof6ivQzTCrYk4Dj5OoC6Rctqni3uUGdeQb42Q3FiIvWQeTtRCxN+H
jbWXE+B3xYwBhirxusqiJUjXQurAivnIYdEKGyLhM3FYR7YH7D767v7XJpt9vlCn
nF1kyDmNaZ+BTjNKN+AM3lJhINXkY3dOlz9SAHNy1D+x7lq/kH0mErrHyw6QvmKN
mzpbK6R6A5X/3Z55g9ENR7DxsF7ssEPqgNs3+ZnVdkv+OsKYwS8LxZ4UfllC4edu
vvwNsAXQ/Kv6F8faUx0yeqwDeToTbIQCWAfU0ZzZqoLv2EilYmVIfTC5t7Ml2IpI
sqFp7+JWlkHvSDNlzzLqBqdUWZ7dAmn+MKkPq0ODpxEeVpR74VdnCWsY/iyXRRhe
XVrzL+RWIEnkdqtdNQb7dg6Xno19d/JH9K/jPPDZd61O+bPqvRhuIsVB/hv5wcWl
4HxelcjPr6CgAL3+XYf8k/gaj+M0geZ1vHC8Ju/GLdwRlayMyZUuBbI6SDkIw1eK
1m6juk0SYS4/cDI6CcqjcF0VDxOAkhpFcuC+zSDGXjL7HcRK/ZgE2ax34WpnlMAm
+CwnbmLAh7g5I1/8ze6DctorG6x1fDEEImc+KddSON3a4RK+KpHjWsoIOL6gcZnb
T+pI5dx0rZH2ZHnFO9nQhIgnZ9PeZ7ZsoOciby/+OlClb1rURefnUUsUgZYlgYvR
QrXVYo5JMDEaKxa1SakCivmyg3cdC6jgeJTwuUHa/1C1hBEjIXgaTkncOBLv3UfK
9HcXGbcR8jGhiTG/aGA01epJ/0z+oWO0t2aFVainXDDjXjL+wVSVZEoz7OGOFhE+
AKzZx57F87i42C5aNl2OeZBLKtYWXlI9kkGE180CplIevuQqcEt4nSCL1CvwWyjS
N3OPthqKNQR/Z6kmThkkOr82hEayM9WAUab3a/WdNHI5X2b0L6hqF7Njj9xNoELU
a/cd4wiogPbBbUOeQXdQTnl5hhesPOn83qUJG2P/Mc16vjRZ8n6sriNxchheyWgn
kREU4SdoFALN8Gdd4rAbv9AKS7wnMwHnl55oUk/Ipwy34tpHc40x1tI0ALkdYT7G
TxPxUBCQNk/eU1o0uHx5pXVP5RBwS4jAZv92DsZEaOLL6L5SViDDeKbx3DdkxLBb
C/T7Zm9wu3o9Q+NQhC+oyXebS6WjIRyLZbal1l/hkxkIJN4/GG4q8ky9P3gJmQdL
hlQlf92Uv7hdlvERFHwXhIcViJ9V/Kp2mq411s9kWhIdatNzfg3BMIraz1S3bdHC
zUU6IIcDmU7zlGFGKOENB1C+Ial2ZwecYIPXAHGQLpIqAxD1+uFDaFyqfSk98Qhm
jqXGzCLMvYedmaNxF2u0Yn86i9OvOdws7lCuiYfh88+T3AbnaIZeUNmfpPTOObPU
iaT+Pb0JS+t+AzreIQaTLu4b9Oft3pNZRfcG8LmXrvaaAlS3c4JWDmIDshoEr7Jf
J2ypUNTultiB5DmrdadvQ9mkvZR0STVqP3AKSNX2odCpA9SNDHfRnA8EpPhExP3e
6DVib0+nN1p9/jiLjbQgavE6Wkie645Ua9HnogPrN1hIydN7qSG7vG9VysEdGetW
zfHjzAyWeQWe8ZazJwpnpLF6qO2/TlEg7L9hNOrFAi79bzlJ2AEnEYwEaf+4C3Be
KFoRbIldZuDTwx7Jcr9NF2uTqMsG4I7HS6HwpT2rWq9ywlnJuQEyW3u+zsvwffoN
WCOSeFEfdBfbe278S+MEP8ekDSVKpHpy2bl7b8lKkAMjZebeFYn8E97+4euiuxGT
8Zwz91U3ZE6/pNR1riTgiF/WxCTJ1Py52IpT4l5kMfAncWXeASPpwyRSOVCtqKSn
1DA/OI5rrAYkXlTGtKLKzb77RcenKTiZUuJZbdrFcos0K3xjJ05qfqcmUEyK01JT
+92kk4PMrfh5+tXBCFCiLeNfPjqjYmF+sUuznwmGja83zh/o8cIs+uDwfC7K6tLr
0vZKMEEeWunmxkqJvjjSgN1km26P6xuqlYqqdDAGoKYVZCaA1V0/5zFPdy/3YqY9
/ZEegHoqZB/ZHVAorqXxwocoYcXCetMyCUA+XjJT2Yf4OvMxX4Ht91UjIGkMFZeA
+EOOn6zkzDe7TzHS0zIznwQnrB32CqseKfd4eIia2WImioQ5rY2AkhcMKT0RCNrU
eYzRpWdSMAjlmgjWvuQHESgZXhBW0URlr32t5+kSkAB1S3ZduaT+OZHfjAsm44vm
+MA6M3v7WlAJCz+kqPv13GsaS5PSbkr+ArNmiLxp2EcjQC6ndfKdqc7JsLMDZLt0
0ldQNlQLgLEkvsnZmQlifF7bBiw5LFwjqUO63Qf+z40QFfXdUTYzpXXb7gtgJClp
XVq57WTO1W/IQOtg6cz7k+zJp/tP7FPDZVIgUGjnDAycRngUu48ttmO4wqz/W4vq
UckMPW+KODi5i/JOtnulogP8KUNxdmvwwmwY/UtXTZsXXcTFLjlqw75EwNkz2eMN
G9/mahgmfck0Or2X+w2NNETJnaWlu6sxP/zVz1Z/AGQLiceXUhxMHA9HCb6aDtne
wzoTzVfkIXdJwHx/ymNTHxrqkb73jyiKbHsJelgWEHX/lllNbGxclEXJKpVn1XBo
448n/x8yN/gOhEpIdfcA2oQHzeuem/p+fQCucpat6pYx7ypGqXxcEFEUH/CDA9di
l8phNp4N9ey4f7U1IAtpJrg9hSEyJ+9SiNqwcxL6nYTSoKGayuH7yd3jqsSXJSkQ
DglDV5KmwVUjvp/arr0ts78/xPZnpeU6UVF/ooA4hQFFYwrL0ObgPDgcQP7+4DSJ
5cjyGm4n7LAMd4D1NebWxR2fh02b++U/FRegrY7GLVTDBAu+nERSwig9qY4kQN1q
ta3KlgtRvWmVmXg2nCVYw/Xm/6ap6AuUU53O0H3CZB8cHnUFLSPPwAHe3t+8Ieh0
N1OF7nzKqyXt9lXcckJQ6D3CQYymm4GVuystxaSZYn5K4f+WqOPzxZy9rEpp11/P
lKT/vXHlfCXvaSastv8T7kz6+aUlEuUZe0xqML/jW9k+n+dxKaULVmfeFVzCzzQj
rUyn6XTdmsVV4UhFSybk4n8/1rzVN91EmkrRhXPM92lQGNXxfWyuxU36ARsExJoB
5dRxY2ZliNTQNpr3GlP0Q4Dul90/37vgYv/wNFzLRWVzLCjtkQC26JYJoG0eNGZM
xdID5CvmCjGiQpR0E1c1kgVZczFLrLhe8+PTlDpJpMmj5X70zu4lDafo5mEJyK2z
VobGlHmVi6QH8fUlbgZvM/jW799E7eRFfaRnrUfPfB1AMlvSGXH6eCMuXDjwQL95
msqfnsWnitjObhNTIrPX7b8SMcJ+0up9HHxnUiXpSw9VtmKJqB6vfcrtCiKSZmyO
2QcSkTrsFiau9DCKC7k+VrgWhMNxJNb04eyKhjtn4EJodCUiJIO5vGbqkY5l8Muj
LONiVG55GNlP8wuCgBI/pfG3wtc/8QItuX32LCsTo+8e9D1AEFVtIAadQX6rFD7B
7mdR28GMCLr9LR/om0Q4TfTkbmRtf52opXZF5winXQus5CuajqE+4OUoVgBzz/Lo
lfZKslAf6Zxjz8REZ+HJTO6bAz/qlb0EqD8FK7GNWMvocgZQxBRfAsNJkyYrB/dc
D2uFs7Vw84ng7Fe0xGuXiR/X+0B6lqY5OgaC+WFxc7txT5i1IhnvEVeT7eKokjuq
7b+bYlg8UD5So7fA8vW3wk1zxl7+kqc38xqMcIE93iH/BfsFA6iloFOJRV8dgwGT
z3tch3mWo69Qh+GtgfYhhCqTXJX7mye4N1L7IbuFop+ef4XmlJX4W/RW0HB3YXsO
6N2P6lS/FFsZP/syHvq59l4pzKH33RSUPGVUpP0qOiY94Mlk1tzlO282lZXrsd8U
Nb/L5/meMERwJ7UgDWfQU+NXoOToyzVWk6/KncHWIcFqBHKkLNaEZzRA69mdvEed
k+LEZ1JBJJ5wSsRq+ExADo4vgZI49Aky5eKutoH6bQcpjhjQ/D4p9zybhHwu9lX3
pII76QuEqID7V2gbGDFps69um6uRtA+EVQuEfVJj44cryWNd6scAd4yFOzeBENO6
I2J2Ut89T8mqCDybOq+W047kWN8SJ7yARk9s707LLhf/lLLMupgRJMQOE7mB7pTX
/fbYlMeEGzAHxRa7pJUKWmxTOKULIuFKVY4rME8FjsYdWGE1D5oYmAcxs7k2aztN
djxnBv7IeQkg2ykbBnbs12/q5y0ia0L/fRRYOCOozEY0H9K4P6e+AAW+6b3wVpUp
EP0X6Zac1ZruFXyuZfEQWzfjQa5CVXZu+h1pcLL1GHDJj72UadRH9uJFtCq0Oe7o
RiyTXG2jzgLtBEwUO1inTpC6kvbEADxYL+EeAI6wT8ba2Zzt4dKU20LobOwSmdsT
AxXUIq9yz3DfgdE0/pWfMGfW+fgkS9ArEz95v8+lavSGRvBlx59hjfOOkkC/w0C3
K3DCd+wjrdY3mIJ4+ifRDk1MUmirR5f35AWg0ZH1UsrxyU+TtQfw7JQBV8jCX4A7
wCBbE54ZSonwFIFyhsfsLw2PG4mgV23ihA9o/pwf0C7HrtN3UFdgnvVoAS+W6Tef
Rir/c0H+uP45DS3W3xrjklG7fxfSL2vinjLdB3V4dCb+NLx2rDKl61aRmxFjuaO2
7Asg/8DIbWL5WHdUoDCNvqK/Ig3rCTiFuKqv/DiJAKPF+nYqyrpjl4cjWAxtQCIh
Bpwr+XKYl+VsaCx8E0CX6G2ueOHPixdqulfAexiTGtHulaQ6Nr4YbcTCD/imld1C
4qn1JwUJQc8YYrB7s0yQKak+82x2Fxwqy31ilODvjlJ6SbjHdLYR1mbUM21gHziG
UoH50HrpmuPHVthjVpMnOifkJneY9F/EBG2Je0ulkI332abxnlYn9Az+MPh/Ys8m
2BKj9dbq4m8plj8Ml2FdZS7XM7gsx1Egv9QpOd0mPrBLjGPtlZNzVyxaf29u4240
tDTTmuW01UbZXUZqHRIDS9UHMwbQE878HN3ZQChtYV2wwNzv2BqXaY86zd8dzvOZ
FfRPy4X1Fcs9uIJWMbpMjixRFzjjaDfEHpSintX2d3lFSvwO/tDBVUfmO2WBlKD/
ol88UZ6v/Le0T7ZV0MeWzpmlvbYxe/9xH2XAlOC/XGiOmApkaDZGStyBM7srZW9q
VnvLuiQAiTYVIFZxyqdNOcAtjQBlKBOFrjeYNyn5BmZBoYybpOo8zCVLf+92wnTu
MA1SBe92M0E254ZtFnwYzM0YJs94lVhyrd34D8SHtzxNSKLn2zaThKP1kUgiN2eT
jkWqP+kFJhqjjFZk+Hebo1xeixTejXHnQGgS0yVhW3frDn6seP10yNwvsPrZskEi
mbzuBfC782SNNcH8NVjOlg6Yi/EcMsP/Z11+1WUgVrcGi0SOLnFbi0yp8fCB3qUJ
IoNgp6aVHeqHciHpI8ymDpiCDKCZBbdnBA+k5GRG+oAS57HF9HId/sMOgrT7uhR/
/w7TMW7kjbEzsPykBWtcXIzXUID5QvWud5pr+KRDT8FVocplXDtczNWpm+kD7hui
LM1te3I0mAR1F+PDdhV87Zw5mRndm3NOWn/ASFzoczhAeg03HNEHdL3zBArnCa/Z
PN9PTI1QPbX/NvX82O5g/St8Ej+GgciyNH0wtbUQgKh3soBKY9xaLFuWbg9Knlkz
69WeCfIwlvc4WwbVmBzqDT32imkIxqdKL76eXLsQa9vokml4QOu/8IZS816lZKZ/
6FPNDGTAc1Slm25oZwr7iTBTMfpuSawmP38IpYMpg5m968Gzy3FWjpt9HYvlQeS+
ObJk9mR8GRPaA7n1M5vjmxb3h2ce2e4cBZfxJXfnB24FYsXxUieiNsqyaEAsOVmv
ILWZVxQyD4xPBP63/FM7oqkFw6IujBEwC3/Xq/nmvDHrT3woitEExXUSQXWGxT71
ooJo/x+NHOIDypsjLvUvMbVmw7tFTDWEwgYt97ovCNm785D9W39xKeV96axbrxGN
krSgsiTMGxC86qMyQJS6YxsAsXqHRbekEpY3KitZsURgeeqFUilNg+tlnUVVAfsQ
bWfyrRZAIIq9NzRsxJYYSMspFwvypZ42g7SCGwreliCPqULycvxnoaAzvBELXKK2
JiuqjEdbnb7OjfdHYVT3dLdCMEUKCVVWT303jg54hwWEyYSClyagBbFb2PuSwgHF
JKLgpIASx1T4M3JuUPNiUgSx/laiuuR1zHhpKxf1xIBDwO9nIGDBCcDT9sdANSQM
of3L8K5JRFv2Gn8MkBSoQzTT6IW1y3+KqPFfzXve1cvdkM3tUUDPADXunrJ7XU0E
FLTonjV0OkzgLwZUEdKY4rlRbxrhWab4Kcff8Jd9KIWHJtywK9WfhdDT/H9QBMev
I4zhtVSRe6Sz3i8JCpqoU59ekD7S2MpzkqxYYYLpmmOLZ6x4F8UsTH8FkxhCk+Sa
TCrZQ9SbEVKuFd9E+aHQafbNLsi1Gvgos0eMxuUJ7gJCpJP2mh+bS6m7fO2/Tn1H
U3USYAaAS2FwYdBmMcQCFDdRhaoojnvU/4Hr+cszoAYaBzSTpX8IHPypEFEkxj2Y
oueLY7uVDDLymLkmRYmgtObLIvOLvwykJn9oZn2/o83gj+wSJQIGrAfjSyqPE5BS
pmg29i8Rm7chbp+Jf9Q034rrpS/UVGd6lSZm0hwJBpd5Y+iiZlD59lA2tRfbjJvs
x8kz9aWg2wKvsSv6wH0AWcvuIae4TJMU7uOq7ooYLfAI/ap1VUWjfsWok//mwhR2
ziVpteWJ7E91s/XJcR8h0YUNiHFHYrsqe3NZkE2BiHtR9W+S3RtEmwFbaljd05Jd
N/EY0qIdydqbNJKNbsq31id5t+xt0D3hjNQR4aRkJIv6cOvsl3AnxLL20DFAef7W
pdN36lMY1iGbIrVqGxnNMQYGXiqtjaEBSDJ1haAujAlh0/Jm85OQwcC0vW2bqfug
nyemOGIZ1XW3qRHyMTa673uCFH7GQ3ePfeT/4mtn8LPSLjN2ysxKB84anWKUD2Y0
VGWDKkMftQVZOe8TkAukMbZa7Msy1/LeptD9LpTE5wjtWG58n7BpbnaCkC6HByTL
CehBA6g+dTIXiFkUB889kjDMrOmlfo6n9RdNgo3D4HB1hetfUqbPNvCPI7m/qLDO
Ort5dfq+X3YlyQYIvYLxCKJpuo+K6Z/IqP3auAuy620iOoSHyJ13gzTT34CIlDMz
uHBEygHgDsQPmeTnp8Y2mRDHf+8m7//QBh8B4nkD/nFTXwQYOKH4/OULeuwdjlAa
6QPwLuKx4Wi1YPnjn/FHj0LCklQK0h1Zeo2Y9Q1oRySVhTBJaSzYvKbZCXCsuCGY
/zPcJWCREXlW24IzYTmnPpftCvGzKrprZea0sRF8RYXrr7kAMP1ZbXl9BC9t3z8m
NrXzcGKew1X1UKp+JwqI4btDIFzXDygWgTc9ZevVsz8QQ3+Bj4317/GJcvMj/ng9
kx/kiYCnrkRC1hZpotN6fKD5ACJ3N0+L/zclu2oP4gBCQ0u5PGIgZFoBL2zSo9vO
49c4UhLih1Q3TCYNOmWqoQXTqOGkyfMFUWgnNmapjNfZ0I3rFC/J0nIZZXkiHCb1
zozoWcWxGVwr28CbqcepJQgw+TmH4qnTdEae19nG1nVjXdBh1IohG3QWj/BXxXSD
cQG+Y4LjJjd5+XHudCorGSgArSZEaownxPAhioX8z1GQiYTI3YZ9MU6c2krk0Lya
uixSm3QxgmQN74vuKHooOa39Kbp0z/cPJ82p17fUD/Fp8E/yXA7+EcGzVLzjjlG5
EPbgjcoNbSxMbX513CcTKjDMys34kvlnEHurv5xAkYyYdkb/F6964QMg8EH4gkVc
cMB5QeFs1nptfoAB9dFlstGEQhAQI2Uw0y4ImfbQm9V9kuW5ctoPeKuynJGX9TEu
histmGUzSwWbokLuGRv2isyGnuFtGP2Il8G7UtiBN11x6FB5mtavXClWCIqSv0Iq
XclGGULurzdVGmolDraxU8PtAsJGb6V/dmbYWcpwx1+pVoCUxAqX3HqEuntF4tjr
EKsTuw6Tk6EJ1soz8KTABimqKmlLdZvB/YDJV7L+38uLBWugmcnTI3vTwKPv7oLz
ydV4OYtSkpF0R/LOaiyT8vb0bBCgRriIMWJLWZ/P/gtdd96Yw2kaY/ACibgq89w8
6R+ClnqyrnJay7BOkGCQrcvsYxhUBFvISBbojoQ+p6PYo/WPlyi6+NRmgzK2C52x
IC05GP7NBBLDKjdjt2WQZJcZzfhbPRN/DjDYHT3btXaa+OWOnFcYDNMrJHyjJxCI
26yy4XVYbmcE3zJD6IJAnowtsFxu1G79Jxygp7yfKmLRH7cDtG31SIVVL/fMNip2
D2UfzymZhqeTBkTxVStZGgXYPCWjJENFyihUwqjaGWx+CdbkZQ9Fwp8DW1ybKaS6
5I16sHHBp0KQHnVoECHnowJCNIt0DOZbZlUEanz7GJHstzMbaEFyGfIjnLkOWmIl
ZzKsOejR/zfqJo2XD2q1jpAupKbl26u8caXC/EQ1wEiqPJut2vzEqfTiDZSdwyeR
zE4m7q22nY8iAUf591YjTVO8fI86/VQzSV0MfwfecLWLEIJWymmBHYoSkx5smh5D
j6Ocxu21ejg4orhWP8oxqn4EOCK2moJSLpM3jExpGAB36ederKLDDffOEk/BlmTA
9v/DVxyHWfbpMggkX4+nySDDENLSHon2ev8iXhXvS98Ttu9kf53DqX4Xlbi50nSK
tY351SgrR+d4EdfauhTxcm55ujBeIX/xNfKrYuMjhXeBMGYM9A69LEJQ5fKkOK1/
atWKXpoIi2hPRiM4cr3w/crE2fDhyvK2loUqf9ZKR99sOZOlQE1HDNKxBgY3kvGR
kahgfXGJm6fMC2sXp+XGfO/E9c5lc+mRa+9ny1k2S7MHpEwggzTNW56lIemxZmaT
1jQ5lYRbJaCrS31X9SWGCvQDZuLrkMKArrdDWLvTbXBTLlwXFNknU1VKuLtnUZrj
edVA4B9hfc7kRMjxBk9whIDke9oI8EKRAVsn5O4+QL3Vo0ImJENdKYaOORs/KRNe
1dTtCsPpapuCNlak0fdLgZ9rrGS+875L7AKM2lWm3MSOtdYTIWDsN8BPH4BeDwHj
iaOo88L8I/B6uq/cBoItPFX46acyxxQWM8e36S40X7/DJyOwtrGg5gDrWe3tsNkj
/2amzFGS8uaETE5qVWpKw107SW32qgmnag8qwk72KlpQOYwGYzXP5eUJ507ZrVrk
4c5mG91fxzthcZDVTQF8McSyAHutE0RlhUlt3vwxJqw3Dr1lJdcGfm82Hljm7yB7
2JsWBhnZvOAhL/cVfRcnIXeXYeO69QbPY/3H8j9QaGYF7+lMiTmtHHJklV+zKi6S
wt521NAbrYuGwMLrj8zEcXw7Ltqs/mspF42ipc91YdV2g+77Bd2LMbfLD6Pfeccj
M5yq9l8Ld8BanKqSa1pLNvCLL+FEBzpdyhI/kbr7uC/9CSSCKo0k9XgzoNEb54YP
ikbWLqUG/vJbDad3es0R5WZgjszolhy6Y0Ghy1Y5PlPyG3Xqqdmzw4r7zLGLLq7G
z6MJdfVCXm4EC2R3ecSSnydNrhxL1IuUZWSEjW2l8SogsjK+lt1969/Bl539iX3i
6Rk3Z+Cyd+e9Phn9PjlKxqUD7sab5Tlup+Dg1SA193Pv5Y4OA8EelWIl7Wwl7nan
MmCCXSZtBx557OL0xDWHme7Iy7lU4WLK0R19XyP6cEWdSIZwp/mEV2zEA7uIdaPQ
Gw85NQbxKb0NkxZQ5+oBLGFnufdjTw/IgCYJ/i7698qFhwVIcerl3x80w7UiBk6N
8ERlkCzcwxpAywU5Qb+I6/RpPyLgF3lEGE/tGQw0q8RzDCnqqxW0DeCwNSiyXQz/
AX/dK8kO5+J0JSBNbV13Wzq2CcXTBvQOL2rV4MDr9egH9HuDN+fQ5ghhANoThSsU
YBAtCM5IErM7IXcaXZ3fkSwbHiHoF/CMqYsqLcIk+t+UaomCFUqLMkFwoR5cxqfI
/ozoJ+NmKqCB37Fj1B5H7MVOSa/aZRFyiN0STO+KAm9mkofHTty6DAbnxD38TjFo
s0kMcuPWnJNQhwSz8p2/zSUuv8Gx5PfpX07O2dWCXJNyn2moFYdkSuOt8Wtv1Aol
uOHzbYUFT8dsnOerk5prAoX++vv/TZQVUgj13Nbvk+Rfv55Tk6jJyHnBn9AEZVWr
cGJS5uCUNao87hLL67uNOjthg0xL0ypuaBoXmYF2p8GvjJlfYTD8R4GzGbzGqdV4
sC/OErJQT2D4/nhPmUzaH/3jhUMFVNrQuy5RTOptyn95W213bT54NkFuH7hiYiGW
zIjARpgcm1KbWNUQlbp5rolWXgNReSekjbjcrIrKtfyM6ZxZmMXZYYn+CeT9yp/O
QMiGDM2bul5yWOUKfV0BhFAcA41jNt9w8Gjrrmxq5xUwFq+xfsdqeCmYOpOVH54c
SjBwmEYhQAufiUZzloXpARwALPFOHJ+1+6SF5aSd5s4cWl/08x6QYIok27QL6egK
fUmNmk5jP1l1zUk3tZHJhVSkID8Q38iybBhVBV07N9Rcko6xXi/d2SMhQ3mNuCrP
NXIvUZrHRt8N16RBruzKY8ZeniODGJywQbAPg0QYVX4KGM/ZPC13kZmtlhZR27HQ
EqDR3TJaJ+fYMDRZ4Imv+oFsQWtTxNVhVomnFfgPW0inZvl0TvKy9NCmBR4kGnkS
Df3U/6dwaxwEDp3jxE5S7BKTazTdclwAy1tBPx9q9gCqL77VTkzCb3hbULpk9Jmo
iOyTV2IHgTIc/yAfLgKKg2SCECW7QUQtb2G3miedRA/px0Z1+jVJctr+ynq/sROd
fpltmfVSH62bwcmKDIWzaWEy3AxpFyd5xzIylcNBgtAEjKnQ0WuqaHMni8HXoIoC
ZGta5MbggiWrZ1PwW99Z4EkTA8CgbvTRBE/KFmXyPK1rk/YTqv7fxdYNhD9TLf/Y
2WSEDZeZvl8zGFdQZvC4PZ1AAuadSYsz5IkAziMnYqah1kO6DqHUprACA5BAyWMX
eTlPPc/xqYXwgE3EwMF2Y7QjXw6Mo12J33WM6qg9fxG5vhFBHIwWTn4QJeX4nPTq
2GOyJ64BVOaSMYeUNcrw7NRnnISLZHiskybCzzvFXwSw0sEpSBa6Ux0cZBql8nUN
xrhW5xjPhlRnw8pu8cMpdu/DDCxHupeCRSgrvfpMn4aT+2GOzHIjoz86G7HYqGGS
auDaEmsm30SgOD3Uzg4i9991Ta038LeORN/ue8TJntP8JcoGX8TxZiHGquRbL5D9
pA9Z37QR8/IvAyFmCzX3SoxRK/XCKbGhcTm9tX2JZ4ZzrGlUeTD+BpTB9E04aIOS
TyxqNePG0rD3pKHYdA8VldVkQUG8/lqQVyp3grxOTTFkFaWyidm4RDUNt2xNNOi5
5wQ6YJ1atmr8Qkz0Doni1m+G1C1QwlgawxZ+XbPNNffM7N4u/a9yXspLvAYZOdm3
SUTjKtIZgz0SdbhLUf7nx6jT6YB3yhYVhZjv4PbkMzAxfEm4iVfXTXi1A3OlILU1
hhe16FfJczxY7jCe9WJcjcYpwUeNN1xEHrED2hpUl00w3URy1tCOYalnaN6U25Ol
3HbyO8ASiqu2p+CPQaoUVNUF2T1nJzwA0Q+C+2/50yKgSUJsmxuPZREGnxiswAWv
Yk3xpuoBNaafmm7EUdaBuCPk/R+aXjlpBX0ZMukkDcgQD6oUTp1Pr17VEuI2MTAm
sBNpXN+dzDwjws/Hmi8TU0Ew1DbU9JfGJ7XdWoduMpEn6LH+eBIaZwYlWHLc9S6c
qTDY6X30QY4S/XJqbGmwBZB25cUxtx/9klncnXUcDBOzuxarM9DZXt8h8JW4HDDV
Riy6gnFjxCIQ3nOITSey+0udQ0REaHzZCHOYHCZqh4UWFhwlWZlrEUsN2D1YBeaV
DETR0fhLZTWOVZdzzOJ36eMqwXSp62kzd/gz4SM6Hczfed4nO0e7c14NlreCUVPN
d4BFP75nTeJd/BymxGdlzs3fReyZTzjyCBUMaoKhiHePiw+8KxZ3OtdQ9h0Nkn8D
uV6IKviF+R09lWkKUsyw233HkTCpzJ8wfDjtnI3P7vWnmhDGHsR4iWRxP4hP9ps0
ejyLmzqFJ2k6E07LrJFB0PCKNl3L6p/RRiE9rsc52XjmFelFEvURJIHb2tCc+xtd
UpbgoH1OvgxvpZ/86+gk8ZAjPgdcSUGY/jdbkyXweVx7DXU/4E2fQySi8mvj9iI9
nQ+trhQZepVY2gE1atH0NWMmSefOAGkvvos0DrHps1siqrwpGYWVpNlhzn55TRpz
AIyoTe8huj2ZpZsQzEl59Q9k2UoBFc3BkaObGsFRtkPxxyMHZr0hwDEznuWa8VYG
ugrJdk1nB/odvuPfbpVPSNjyM7cJe3HTSuU54or4U+Wv8c7gdHAlYnz0EAAKhGsQ
oZGLlJ+vHg+47wkxbUeyfV2Ta05KB1/3jMBzHRoB6y9t99j4T5brYbczbjOtfF4t
+POn1srnaY8rt9fCS2WcTCA7K2aq2nttpCPpXZymYxXVzpRi7vlEHJQtMDKQd0i1
/rbyMMAgVbWOnmVo6YnzdcbgRvgWrQgginRZ5D/7VMi8CpvC+U7G+xdDz0XP9Pww
XS+b7169EDKbRXLMo4t2qBnOyCsB0nEahkkblILeW1F5ZMKEnW8QwaOR23Ow0+vV
BfkYF8LqlkzORhQ/3Vmo+eBG8ifaUGBUUPCfUFeT8uNLsrp98tr1n+3HMoBKDn08
rrcwdzXJOeIlwctrA8dP6o8K3utrmDslALmNpidpjXT1csYinWms14PXJmq9nnSQ
fVQVfX9/yWFRzsRLfPaqrCXULf6dBDtH7RmBA4oSl9TergRfLPoP8F80lnEymFZo
wHbNTqFP9kR15pMaf6//Ln6fZklrWRXOMDEwW4W8xPcv/CICDjxP0vtZjIXa15nb
lMGi5LkJSJPYwoYi+61mZc9H1qF72ztEOuhZApwmRg7du9bd6NoiQgTjHMDnJuGA
u8mXP6lyui840AXSKHN1KnF9blHX75aoKym8ZL483yWeVSSjtIuMQZlGEJNVizb3
HK4fi+I4aKTr7+hlBTgbJ0BNadjWsFcmTniTfRf0RTaNPQcAY8JgXstjBskhMQ77
qVPWLTQ7BNH8xcNlQuWbu2XkS93rLJPhYs34q3Vk6LW1YNljfDJE05GfkPrVW1SB
vK1+m6KCRjQ/PEUWXpblhVSRhPS1R9xOXfhc8OfNdpLNDjELnFcVfSp2TRu6UXAm
KIXkMJlmEkK3DPoTc5C1IbmLBqJqm4NXwhqFC/g5wSyfemeJhdcR1iBVSMc2UrOO
QL+sppHd9L9HOp83KLomNihZwkMe5Ug9zQnYcrkKQezN0g9XTGWPfLrN92ZxQWz1
Wlw6lMfuxZ6AmcWqdEOrLHbi91K/3+0/FGMxsrws79UUovA/QfMH1ZpMqwAvcanp
9KQa8tbqr88Sa2sFP2nfAaPK+rViyiLs0F/tq1YkJnS+J8snSwao2v253BqyUehe
p1FGCAW5Dtbp31jTG0vockd64t7gp5OLr3qEtBqSKgw+TnRg4YRGRV+akUtfqbHH
fs2qHVmCd3EiU8TSWSwgZW+UWCVUbSt5KW+Zu9mfkwZEyXkT5zzCJI0GKtPwMtRE
/URZb72fxAjVuGxNubzXljQPXDlWORz7Hr4/c2sVCrDXlNLzOTahLu4BkZlJJPse
Qq5jyhNX4ifenEaOLT/qKl0Wmi1zoku5s4v3AGHVBqNhZ0y81jICQfgau05z/7Gh
lN9K1Th2DD6BgeiOFvzpeQMKRp3qAskfxUnIy0h9sym6gIuV2SAkiEY07TOGiq67
QqbjxzzHT5QbpNezuhxlHn5MtFTIRKmBzfiL8I4qhzZet+sCw0jEYWLk/u+MHMwi
bdKaQ1w0X1eBIkqBXau+NQOWHhMkm0ZZcI97AyJRYNQMYfqMLv1nsipm65g1gZDj
EvJe6KXS+Im4vzbVMPo/x5xFEEfRyr0pEDLZ3fA4A3uKXcPwEVfVurLUUYQ7e1tz
h2/oLLLsCigE9nvxHoqVjfmRhI3/sxCCiWdrx0hVJ1YBuy7Nm5JOOh+0dUsdj57I
dfmOiLVnsOu+ej+0zNbwc6nQJgBu1ySzEKDYxq6Ujff+csCmvs9oKMMiaN9x0Opc
bzDzZHo+datDPVMoi+cDK0th/xs6N1ezfMq4jhtTvLuRjJUu6IF0ASMl7y9+CwkF
Z3KS5xmrdOfmLYN0Zf9Mo+Wzvmyv7K2Zq5iAlC8O77Pa4VKA5CYzYgKc/SMht6f0
4Du9PAIxseoqRo5ctuH4NF3rkN0qH31KVY0PCFVpDJmL41mpHrHTuGcxdYweXrPJ
r7trOgHMfAaRo7/5s9X4GHS0IwLfXwuG3LDW7JAUuGsuF3aHfq0pZraD9Xr93xEw
RQpFJ2Yi1Re6iqgg57eHVZuA7kdX4BhISblXmmRD1giv6rRXiP3dvi4RQux8P7I8
rkx3+oSLAvfDASkMVu/1u/RAoqTh7WzuDdN4/q+Wa79dKCyQJtYJLP+U8XtPPMKa
Xudpv4aM4UI1RkkEpgHS7kGfttzmFoKIKmbalo0/pg0EmTNW8IAy2tl9QzxUFI9e
BQ//aHZpexOwS0AbpQkDxBKLOGANaLRdnqHL49biQpyXbxSEITWx2ILNF19ro+ta
61VEeSRcE+kYIpAwKeS+zbQ2KsMhoeVHkJ7niX2JyWtyfqZGqO1FCGOH/sT5W0ON
6FXoh7xS0sXPWM5xYJquyUqTAdHQdXap/5MjMfzYt7fL0G9sHT+bT1kLnMO9ufiS
EnLToyhWjD5j/NmcWWcwQlfnKqIiqG0/pZB1vS7ICAoBk08IVSIIs1B02tA1DWSq
2jnXHvrBCrB+H+Us0CVRER4XStPf5ncVX0++7OTY0oNmm8ka7c/SVEeNBDHss59V
N9IHQyCMqlXdu6KnBpAWc1Io/hedUWYCRsI6l5F97mL+l+3luGJtNykdZ9ZCwUa0
jKXw3JdbCOxhwkcFMxBc3ZHIgAPqNejny0EQBz6nYduop6Ws9DJnKPikymoxieaQ
7yRjP6+vBRmhZ9ow/x5KuHQWYFLOFbmUlZvCHLbNdnh3Jljl3L8m6WZE4rWj2ypq
KpRZTwGQYVambAoUUHGCapNBN9OCM36UqJeq88cLAATzIdZ3LorQgTbPxJ206lxo
1bt7tOXeGUmyTiHM+exBRhML/MyrFXJdXoXgtBmCjAGrRu0ZLYO6XDZxYYeOrjzM
vl3XvTJR15ezs7En/O1/DPIgwolpkbepLONAQxAoIde+KtwSwc5hD+3lE5HxNr0+
dmm+QAXwSzmFcDhU4gnruuVlW8ZbEHf0Gc6Q3kO/XEhP9R/B8zZ09z3gZSGIq2Ud
qw1cWXIu51HeDz5YIBraO4rJt30jaS5emKLtiLA+CwhzrQ6fpSGWFyy1yxsv3Cml
t6zv61xSY6+RyZQ21p5Yk85DG8UngKegcShE16Zv/wNf3I1Yz3Nbhs4z9DmvsrH+
1pP26YUvXY6qiI4QC20mS9rqMaVFMUg5waKJZvr1wkXWv1CZMZqvyd78IW7doYeB
B6W3e+Dzp07ljeT5ejy8ou5b+wtVc7zlQq8WqBeOHYl0/jzJV5jAogLJbJlLiFXn
og8WtVntXCggT0N45VH+0LtcvgV6Wb+abK6yQaEaj7NR4iK3CSoegnCfZwrPZDC7
uqWLwxtcEakVmHVE0zjMzQ0V33MltNC8lMngT/r9sOBlWLjmvHJtl6EiOwzwb6rO
x9Qm57WnUwDS/lDJXX7ntDrEdTvBD6veJM+8Py0osja4Wb/gXIWQLLCO9L315hLu
G49OsXcNakcquGHmj5Z4qcu9F+Ocs8AYTVDCrzYegLLwyaXI5fwxtGLqlBx5lZ+3
+/XZrL1ZTwmGJeVmUkWHEnVa0ro/J9rkdoXwMa4dpjZaRrKcxRe4liH0vKvFtB8V
hrpDQ8uM1lr8CJjnwDgbhH1EAoTznbr+MAkxoFRAOqQZdTvf2mQzrUyEjWLPhRJB
GqbIg7S115kWb8geVTqyXaZALhh0MwkP0DNtk2OQLZ8lv/6lGdSE5JKGoOJg4Liq
DOkMsVJx8hYvHDKFTPgupB6+HsXcvsrIbds2RvDTH2/nNKEjZ3Ion/FfLjUNa6Eo
VnAGWC46/bNYqHMQrjpSeZZiWa+xjx+gCTqnSOvSnMRoV8/xY22m0yx9yJXF15Do
sPDdCvtJIlxVuGChZJU9icCHifxTvYPr8ifWGLWPTGSuCQc7swpiswlXmqdhlXj+
pZUc5mz1kJldk4RkyQC5FttICbTzAKfPK0op6re6DP/I3GAz4bWoapi6FTm8CLC4
902WnQrmzVJz1s+WYPMSaYflzCXV/7Pwby/y86n0YuKa6OfZERlEm+Od/jfw+Ebk
3MWMXNw4xqIPbWM1f89SqJCfgSkRj54GueAYG0TdJtzS0+K5o/tcQeEvbmCiMTYI
H+yrIweFCe/lPYN7xmBgbEbX7hP0Gryt7rBm2JyRwMiQ+t01F689TgKfg5u/gBds
VNbXLAfZnQyGZMo1pYOz/A+yrig4yDnz+IXjAerQUS8NVipjj8Dl/1lVB5iLzVnG
yfmIgQB2cQVAOFDQ5+Bk576FsIXOLeG7HARRZvQaZ6G17hlkDK/g6vbi1XO202CD
p1C7a2EiJIWkNsRnhc8aKylPn2vBZznjj2eAJ1b3jFchF6nXol5Dg5AdxuFPQxfI
xzj2TZilVK75OcN1QOI/bDND2STVrcEaVv8mZUi/FjlLa5uRQJmvpScp8dZfdFG4
EG69zeZlWHSAdANbYMFMzLJta7L7ubld3oBNpuDsLSNtkTe43jZYGFSVzzUyN8ca
nJt3kZ3jslttFvmfrKya1hgfGjbTdPFGZYhbKTEVtBuEgSAU+Lcb1q53J+RH2ECZ
u2lfw6l5VkJs/KrXs8lVhql9mNp8udAhPxnr0S3bLCxI13wRSZBiaXviLyBHo9ud
rW5N0JPbfU3l6IN7R6XC9MzvfX321iOI985dm3pVhNVYTgKKASxt+1sHaIVKlKiH
WeAU3M3XEHJXUskaJ+zhQrz5W3duVB4rzrBn7mtxnQOxHuGrrT2Hkg5MZWKMiPtG
XYL0xW54YUIPQ2tKD3mT+OzC+tGfVt2Pwbs9b+dphPqr0cQdcW5xVpxWwjBuzM5q
QUDkgrpIykG8vaz97e7L2x1EqnrcBP4BRjmz54ACpbhB5n4+OICOuCxDB/koLaW/
pizLubTRbqmm6xDyHjSaS7RDbqPVugbM4qL4A3obbr2jtYoNQiwYWyB6hgatChLN
yIFd6zER+4gMzBSqxiZQXysKt9UxLgBg/D7NHmwmsT/9uQHmyUnTy8fD7DKi8po7
BlK//XXX2Id2Z6DYxILIzs+Ey1BxbKRS9U7yhopeA05vAJ71YTwYvZ4m0FKGDpJy
PjI50J988kHZP4KEZQRGiBjkTRmQ8OqXfpdR2aigzdmTAtMuyp63l3Q8gTroMJTS
jKeyWvtpxszar30ayrgoC1RTjbGgDEhe2q7+3yeaR7Gg9BX81TE4qk0CzqHR4xxM
SpcxI9x88fFUFC5QPaewCykz4+FZoaxWOhBHgGb8oILB6EqI12ZVdCZMxl4QnLTM
tyfVU7nOOFLERF9RFtdpPBy2zOY5/obbGmn1GizOQ56qnvr4MXf04h2NcxZe/bMY
u0KJU25xd3YZgfem2OURbOqbSLvgGuugmahmzcPNIJe+deY6wRu2CTf6KDha+UlM
TianeTDPOlw61/nSvuzribgG39kwpgw6thghNcOSlMN+yATAM6rSQc/6+G+CgoGC
+GV5NkimOTJJbaR4RID2o4xiPDOxvCWfrIxMBpZbeVyfI85w3PqgVJlYfXhxTyo7
42gQ8mYZwr4djIzHrD3W9WiuT34uRBQaN53ywfASvj5ewANNUbfEWTnuznkZnRCk
ImngQL5YrZF7NvJWJSGp3n2cqB1Uf471V5F6EPs9F2aYbHd1FL+Lm96OmkGZ2/cV
o+k+Rq1bBa3Gcll7Dmf8fxXADUNYaXTKmf2wXnGqBtkm0JUnX+ylY+sTr12AFETb
mkcoTK8a1hbBJxscr7tblDAKQ8pVC+PoZ/QgSu8jT0IIl5+2loTLBoMZam1DSLDz
OH+lqbmPhOH7v1L9QH+VyHQ4PWeuDZ3dPTO5l8KMaX17fKHS2dqVxlvKtkhVnbiq
23Xgzsgsr1+DS8QIz6QojTTi5MACrrG3yT+NRysxBZDi3tXupL0cP+VKr15zqRI0
Ehu+7g4QuS3x9SOSkEIi5+7ue4zUSCb1Y2hg1dWAnOAywNB5yL5boEeBWIV8Dfmi
GWsRPITfiImDWqFtekl7fcTq34DajU3FqunaL3i31UfUKgOVekgv+OSxooBpHXyo
gNjwg1Hm+V83IH1n1JHLP+2cQp+wW4pPDXA+Zjf1sfE/0mBUKQ/4+tnXRBdaUaPt
kmtqMR6UeblzVmc0VHq9gUPE1+IcfjNRd9usnsMGhKbQ3ONfXaKXagsXiNwaNyYb
lY5n0gi/fsbQFYS6PNBAhxELUS2QOyl33SpMUzdya4EOs1jsZ+1KZm0S+J6iOCOa
mhS4cudZYmBf0eDI+ENnmbv36oxq8+1z71lCHU9vg2btJFfC1lPTc/2+HUua4/t/
5utEx4apxR/uZKM9UqUTdzoYkWm97mOEmE+ZhLtKSrfIt3VmIGAVmLWBXhdqqutD
5p2tUc7QkcpxMua9kCIoeNNjdWiR3ZyeL0QXDqh709zv9TezlV++X3eg0ZGOj8j1
nvAgqS8lxyGdMA4B2LIQLOFwVFNYrZeaReTmnaFI38zMX9E4mpVUlnQZSEABtgcg
DHEi3Yvl4u4qMfaBUe24/vTxvnLXQmkdHNmMVNaBXGD8NRM2GWixaYIGyQNcr+/m
3GLFGTqamG1Py4gqPXLRy2NVMxjfnvVsd1HTqZIYhPbap8OZVqfbt5SmsIWBCPb3
OLDWddzFEKblmcoDHBnbFazGowJowR3Xfg0cJMGc+xyODV5lcUFwm90KEG1PSgLm
rwJwOUgArpna96yvmDDjDR1ItLlPYp/HeSdoN95Uyxzj/joBALMsHkWgFl7xvNcL
SMpV404R459DjsIPJHExRI02Su/45iA41mxguEbtrN4JVhvs6hCPqIYjzjoQSAvt
Qj5Z/a4TNgn5g2ByQyTC6qJ75AWGu2EWc5Xcz8+XuOhOzBoZ9UQ7EsRpObnLpBsi
GD7LGggglfcvkGutMhlK7W8GhQL9MkFvV6NIzPU41Cb14rPpGtntssgVXkURKanU
uR8z13x4Zi9g5efIcKKGDMNU+OvkLAQhrxmdzMN1ZAmtxvRrASX0xBsipjVZr4/O
2lCbJzhejabuhrveiPW++h1kTLHxYr5VvhyIHC7o9CVMrllkom8tr2dy86U6uaEp
4rV2Ic44gRk5Qw8NHD6tmXLONdAAptW36bYNvYwdjRQG7fSOU4Ar8+5ASJNjYw1a
9MnY0PddBsJJsQT5mRgbcp2atifF96kLH7IyZZRO7xZKw1Z1H/0rDtTnBBRXKHAB
arWzhK9jzWyJYny1PGic+Xpp8CI5hTEU9GOmWKqoEtdxfMfcSEJybfaNeUB1GqtZ
bfohu8GHgOLUTWXA+ansZUqn6lYrMgMWyJLsbszWTIorm+oO005qXqCckyUupETN
5DH5zTfQCARLpKqMGsxV/2WQHpyegJo5BwHXWDOEeGep4u35q7DW6fABsNaSTEJi
gq5j1SQNpBCb4qSmnNU2lCHnia/+sQbkB+cFjXQ0Yr9YNURKAuTfkroPgvO9UNnG
2dRNrR4ZmCEBfSab3LOjqP6Q1O24cO+YZcDKb8O4YippLY61LKZHl+cuLWEsoShk
JZxoFkK0X9Y2VxHSIjNeS5eeVr5w8k38UzlRMaXs0pIZXzhF2B7BxAF38mG2U628
6ENjk+4PzzUeeiu/BaxqDaw/eHwEp1HAI8TbAusa7CoXT0iFcdVf+gvXMPlp7L4w
/jWiTf74esf68RHCipj06IKg0kQrdtVl4WkLCIhRQuYGRhi19tdlIZdiSo2VTykW
NXnDxCy2Fo9divRh3MQzCzv9lQHbGsiUtdv12g25s9PaCQulfyNyoo4aqKFKqWkR
omL671+1dm6LJ33/GWh5kga5wO3qr67AAoXSXjYk4BO/g+DlhnUWbMMP5el2LeRb
Fr5feWJfCF3ChA6ZzG50PCWvjNS4QKFJB+Cws/hlkqOb7bRHL/AkO6NDAat5x+bY
nK4e+q+8jXvj6RrxSxQuJnl1nuMHLOinfPgTfSVXSSaa2AQZv9PHW8e3zSZ/zlAX
H1WxCxTLT1WTbFBbQHg9X4oRpy0Dg7EdPWY7Lra3DthmHwbeilhIJevw5IPbN6WM
0qNsW7izsALcj8ohNWj9o/aUVigZ572rN0Tb0RYoeCj088t1iSLTYdEF9dm1ACmg
/98AH+Y6bEFx1zDCNu00sRpfGG5hGC+kza5qzOSd2x8auroicFguBrYzIwaqd2WK
NYiWf3918enkgpJGDyNSHlpzBiFb1Whb0VhNaThb7284SKc2IRt9FYmSkCNLMC8F
oIyVJInrYgmDDlAgA48CENrTAMFBtpawA0euE41rKelh6tKxs6nVgZ0vCAnuXGbp
rSPBMEJEnNFvm7IfZxJzxEyBVhiFINTsc0kEjZW3iGI7XJZWc8ZYi2EpLilKZTEb
+u8H7LtVmpYOC8j97haqKkdvHwaY4XZZgoR7WZH7ZmLuuqDwiuzrSF3d4f3qh9An
p1RIDR+yGICnb8d4A8lBzDepHe9MYfF/Rn6JQM7zHOeq/Tv19FKFPYdNs9IQmkD6
Sj8OytxH3W/XpQhdXboI8RWT7UFqNaGsXzjBIY7DX0iuZuKcn65lz3QHWYWdmj+8
znwDFR4hyC0cjBp7HFTNC5i11SCSGu11RbGYjxUHfBPMboimWc7kuBtSbxVsHk4P
0mfRf5S7ywZb3gZLsncIAKoYpxraYKoYIz82Qm3B24psi7w7grP8mVry0nI9JY9Q
ySlSc2vq1AE1ow2Qr2qg+m06gBuWdJ61t0YtZjRanKgbo+zRverkfGbYPoLHI57Y
KAikxT1kFmnXU4M8MN3LahqlENELzxC0HGJZ4ZtWVLy1xroPSJ/VFg4Ex4Kfhlpf
1frKxN+D/Ms9TGKrUBmR5k6maq0Y0UYaKwTG5hV+f76pxMLuApOn+ryyhXR4vFRx
Zpor7zZbzwGODgZvue6L0cq5Ox61LlPfkxT/DJZDoWi5vLGIsrTmIR67B7vitKRY
bghj7oy+qK/wWxgFzHdgppxfY+O0rKIqyvKKbRN1/YRroHZrBKsBHhr5/AKqPnkb
a8jooTdfsc0h1SFWY7XA/rN7GNBGps9e0LP3wbCdM8/D2jMIDV7lOVUcu3LvhW7i
Ucmz71U/rdej7sEacuyOkU9LEOyM5TArPZ2XY9fdN2eynrBQBawJRM9pjqLivlTe
rjtT66ICxT8zN8R8Hu0Ip40rUUU92AAPPXmxenVjLAuBcrN8FDQyJ5LF4GYDClMy
X0bl0JoHbCLQ1sOCG6WDircyLPXSoRwvsYPTM9nzO/cQCFLOXAibZFduOaQAHUKT
T68w8R8AQuUJn0QqY10otsy6Bp7j8FFoqLKtsTP1RqxSfyOqtpHNDgtw8RfT1beV
pxug/9ELByUbsfPp0XimL01KZnKMbHewmBEWU0okbzmmSQVI221e7vl74DK25CTM
RUY4XDlQKtbgWXYqgWrtMqqSdgUGEVmMbPOqGFoO7MPa5END3dLwC3hp2l/n93sE
gr9u5h3HzdQjyGhBCEHOV4CvFBiqvkKeh5A6ufRSUy+htwGcWc72pH3HIwOAshpc
4qTY13UAHsFI0HkVcbyjozetNBRC1VkGUO+cr9ibH8Z11MffNB0h6IqNVHp5dg4G
R57zCTWWjLO3vo6xVuCrBrgqi8lPJ7v2XWcaM0F3FJ0GHx79YssPhmj7mtj/CIOq
VstsTJn1hwFaRXZDlcd+M4JGzHqgS2P1xowJ+Id244nkYOf9MDf47lXnqK+kdnl9
ChYHzskkR5SfSl3c2mI3HJUY/tj7uqcHzrR8pHXKe6FhObkeodwJgBcJGELWFBqL
T7E0GSUXTKhrzAU08DuNACL6LCAM0oXzeLfy6j4kP45Z98PePLKLFCI7Jr+8oI8k
v/lRhmgaQHo7th1pt5SPMP1pCOol/58ew2qKFTPmjLCY73ZSXtxTpgLA9kQNDBbd
+rpgXcnwi5pk6TKZ7f3xGd35oC1bYl6WuaghlG3hgEj0Jb7nfbEaMtM/zLDKoFmW
HD20HKIka631gOgWLYkRM2z/A8lJQTwMUnUEvku0X6ebxEinWwD7ZQXyeRY5v+Ac
9ZFbSLfnr11g4vx3Z+AeeZp1v/V5U9G2Uf+MyKn6tA27qtOofeS1UUd78VLsVlBG
tR38Tk/mjrc1v1z3xhw/Fa8eN3A5wfQlAxrGjvH4LIHTWId7rSyRM5LOZNI835v3
oxrt1lW1Em54nh8OCkgJZzIqZ/f67Cwgd4q/Ti6/ZlHoINSXiFCWrDIbIjmXhjn9
wywg3Udyntunka3mv565wFGZfTL3ZfD8CEcHJwGzcqdVs6jgUIdVkD5wwZl10Ii6
uOdCUOuaEI9G62sV5HE2uWBuIythiKFrsOFJkDbqKncZpLQgCAXyplXkor8EyUsQ
RZOweRqJPRSD7p+EZRk3hFMup8hUPl+bP6RJ8/FGtcOtj52LLP82HcJMJK5BALT5
+4qfWBuEnZnUeA+lqZXTx0JkbLnuBE3Un4VSp0XFf8Mor9rPhX+uqxMXU9UpL5Nv
1NCAY50Dj+0Al0N09zkGb5EaWjcjlOOC+Rd5S46/RPNfz1p+rOJY9QnGlpdmJgKP
sICXoIodT/YxlELkcJ9H9tXQWnEe7glnLgE/TEUuV/7pFkOJ6r0Gys9jgTMdImi9
DFJcsACCPdY0ZwWVkuv0indxTefpUl8FuPUrrEvjybBVP148GUWhr1fwzIHRM+uN
7c7fbuSlBvBZREE6kNbMJquoVXIiZsBzQp2ysdA4Cc10rQ67rxfNW7p4AdvAiV4R
UjOXNT6xQIldHfPR6W+ZXHlHiiqzMGyM+tEo+etuXaGHKkT2p1LpYQ/DP5tU8YHq
aMbeWyRs7QmcKdmeHGciqlF9rIFREGEBfpjQJx2kaT44PbyC+8+vZIJZCiMxYH57
6ybDKSBPFXvhi0qIDuDJPxXUK/Oz29b8T4Q3FEkggn+edAHqyEvzTbQrek3OPcj1
7iwpeC9PnZL2cyQTiHOSNXrcv7aw2ZuKpS82dCKWEifjakjxVpRxAwTgUlhBcjFp
KRpe3KgZN7B+EN383TDZtyOwmcgu/YGCdTocEvtmhE7nHnAWfPeCvImaxMmK3cCA
Jxud+IYSpVTGLJuPxAplTz288jcqM9kgHHvq6DP6YSeNnazBrixtb32vlnNgyDDA
NawC0ZD5XOecpUZ4ryMkvAdscWCPgstrCSDxmgRlfB2PLv9yLx+EpTQuV/6UlQJS
UF6SpakNwNSBTqqWOPaoj5j5OGYFHChleHguzwZUMwXxgABvSupNwcDLpw5Hw5jK
/eIy/SGRo8AaWjezNBxMrwG6c3MYs3QU/0ZL4BTmnHV5j0EZmgTHFYaGrngzTOPb
BwUOGDNDSMRkBd/8K7/Y6Qoh/Sozugd+UWQX3BJUDfIIUtc84gKse/u7WWcqYzyY
KWtzplpnvn2dLrP1kxVJDv3LJvYs2h/H3sbN91Y8CnQb/1cjKfCKL7MDvd7HQ0zD
oThkKr3IOIMgOMni84BkzN54XW5PZnC4rgebFTKHwoCk0Vi4e2Lpz+5nY7f6p1aU
qnTydoL2/EeOhVPVpUi+K4tkvaNwg4Tr2dpeUYbMRdD9ocDkI9NmIKr7n9WmeR3n
hOrtHSKhkkenIfnssJPn5eg40Ds1aj1IPpdrwwAl6mjfApnPYFX6Ar6Rr/jmO884
dALh1gdWR74e+9kqERmbM4hHjAyDtZGQXGFMBelfHWgRcuJOc6/Qjm5yXyAbQAiG
u989y/4Ka20F8aQD10dfDNenc9yxsL2n7sDt+mInZ/sp8PNn10QlEdGRhNXETvGR
xLanH9nKbLo0d2yc0UJxcDUlpBxLs8TZqhoFcn9G6MsZTmLOfgUwHpuUEFYunHiW
gwVZgNsyeFQOHM2wR5FkcRY5Jyb+/uS6Vh0aeY2BzOXKCjKE29iobnJlOUUDXiIV
/RG7MP0vRuyfRnqYM6lSuiNO4KMUig4G/knEnw6H2aRTcDlwLP48uinf26KY9EB4
TSFwsieYsh4VfKCN0bODXSyjb96xTZ9jOVh5CSACQmXy4KPOUTdzc1OMbChQxBhO
rXLYr6rfHrdX2TO9/0svH2oExigDSb5cjh7rVh7rMuRDQrJbHk7DlkF4QBkMiZaT
OAycg5miH90wWovjgOJbjo8pb5NubdavZOSwtTslsgLswft9BZg3GPcfdgnhgb2s
5TdbDNy0meZEe1pnpd2B92r8c4UvEhdbnEt+5H0hz1DrJxoTBT7R2kdTgIxaeD3M
0D6gK3poAEFm1f0xUrBQeqEiLiviMaKhX0XGOlL6xBX/H+wL9abTne/f2JgoQ+hD
QJ/XX4cewYaeGs8+4wDomynZTjIzklDrLaU2WZRXNcyoo7iaio9LVCAFo9AteycW
nMdo6mr1sRMPbLh0JC3LjwuaFF42gl5zaC2vGh9Os+bvv5nLcqi0MAkrjfYcjuuo
6/ZPMqrm+Nl8WuCorHyUXuLWCk6HFKN8Z2/1d3iHRM2FTaT8qcAYFy3O4zg8gAH1
hHdolNGDzTZKGuchcDkG4sVt6j06gayb5NYurrFgvR5bfsWGMLxV+TMNcUFfQ1UB
WSaGJkL+l8wa6Y4mRA2XGDnT+wcOkH0Ayzckrp9tcA6+aQ+TQ7kZ92uez0wDcZz/
PwoyhX4+4bs0qjsCiVSJ93IZZeIqZJBzMZZ0iAeKDVuISsw4wCVFc0C8Oj2UIegh
eL8u5SpO69H7Snx0RtZVLeaZPANKPBqpkON4xztoYs3vnsgfVJLbs/++oN5ca4fF
DLM013KkkZ/At0fokOQGISev7HoGJOKYJwqn8ZG8BbARDVZC/LRfbbEsTHb3Ltfu
iMPgbmc3DPqZpwq8HBTDbfP3t3qv3eEQlkKUgtiVhBfu0o2ozS22CBnPzXddUdfj
482HYIVSk2g7qqJaV7INrzzk0z0PHJv/dMH1UISYnyDFRUfgwvN3FudFaB5xoBlS
52Vwj0mbE0j5BgwHptRGDSw7le76SOHJA6DyLEoxAvqZiEOnxDkzK3Aqlzpb7FCK
SJFRQJoVR94xl35XqEEo/KpzXEwadLvDrEpHX++6p25vPDjRfN4+O1AnJ9bj8kkz
vnPjJ+CnvRdWESeoe4ckSoX9HEVXD1x2m0Dhfbi1f4XWl1dM4AwbGezbp39xl3u7
o5TWak0P6l/DFyUZ4u8WLOHoISyrauqGVP9ut6mBL58Jq5vU+dpiCitfLrDYf570
iqYJ7HcQD+fo9FGRU5qq0DXFPQ/dB1g9bxfanuLfZr8tWCx45Mf9eeJK6gBW8wP6
hebgDi0CvNunS2eZ4c4ullhuwOFf73U8l9gNrREC09FJv2xB5n2ltkdLmN7/WGre
Ghc2zHbqpR4KMZX3vTHAxMaTovLH/2ViOCqwqkHReL4HygE3liFirIF93L2b56fU
aKGjM7jKoMH/iZ8tZQU8BOLlUO0Tt4hJPXzOG/rgHBQ1pneAWmFRLWBz1mj3/Te2
vewOuIMw2JPbeeCBD6p4UKNumG7YaTzF8T6/lb+kg2dfRkDMO8zzy60hLxk6VvO6
i6b34Haa9+N1oYoxCffm3fKlMOfAhmvRmmw/kB5Q3/GCXugf1Eo72cPZB+/rHN+A
0Azd+dQej6BbbHCyF4VRdHHAvRxezleWjflbzysjw5Tvedlyh1hxoo7oA0PooCb6
BHzY7t1WJivJcJNAxnl6RXjT0n0LkaTxZlR1IMhkC6iXuywDbNoVNuF+Sx51wAiu
Ynz+x+k2u4yFoyTSR8kUorJUlMPcZ0zsVBxLqV54WpRPql+Y6xq+TsTJe7MSBtUW
WwKcxPYfHTrRXCpxo8m7vB/Vp2SgX0bbdHH9XQbocmci0mHnlVxoZByLJIL5+zm2
asClNM75IUhMgAhe0e2rY7DDZ+lhrWT/tLv65IeioDL/1UiTI7ld/UqvkTy5RXIh
S/fKDrQ5CRMDrfnQoPSqN3ojNItQXfZH2hXP6uSyHi5e1sgd/DKF3iN9fFmbHUc9
TeVCtSHCXk8E5EqY++jdAjX71dNVnpPMhUSblF0Pa5e2EdkMM+tUBi0gTnwTwWHc
U/ahaR41GbUtUKh1N+iV8Ra6cdEt5geU3DZp93aE/BOzO03/xiSSCX8+dYqrsIcm
noXCC/5BOHHJOA3McZfdXl55ductD6/mIuAWoS8r270Lkw6l0bpPXkEWHTqBJIWo
45xZuMQE8L4rGgDJdOYTighUGT1ZKkQbFz1gkjpeY803RbXDDUkVa0Jh/VVi1HO6
E4PQWUpoRM7m7gZp2KFOLpJ8m2mnD788Um1KUWuQmnnfeJ4iriEFezBwKiui8c8X
tG2l7EgZTw7wUvoKdhz9Sa/ahlUFbsY76n7KemiwgPV+N/YMPAyV0v4ft2J62UNC
abUwSn3bxMqEIdHdQ34RlWEy6n2Yhqzvtxyc96AQNPKqcIE1mer/KDA4K3zy2vkb
7mJMtHViBPO8J9ZnoM7i21Y4SN9TCPNVQetevGC0neyokEj8jUWZ+/2PzsVmEf4N
TAJ8URPu2H3VtYxkY53EDvFzuUk2X/kDbb0f9ighMpFDJteBrfMGilqpMlFc5861
+W+UnuWCLboMi9iCXov1ye/a+GC6dqLF48eh9J7pyZ38JyuRPHLmd9g13RuALMCl
rT2peSZ9uEPXopLXsItTTLNoSKo/Uk4ccSnc/X0NNaW2SLo11bSBOF+n5pL26ubo
PgzRHnu1/WGVV+Vi2k4K9/M31KSJjSajeFPxvOiqJfGXZPG039epDbz7/Tq7Eoth
Q9yHW4p/qGOwJAntTJ5c920BSVz6JxRqKcEKB0RtMAtjHKQjYpmGddNf58DVbcxO
1q4iHdhFrViLyktwAymayt6eo5bF4J90QCCXaPgFxQahosRZVexALXppTFiCYV0t
xoCH3NnnCtFwdC+4+Cq67oPgQNywyCWb4jH0JO/Pe3qQbFoLv44+d25mx3czp8se
62ocwnheVk0rKPpzQ4R7doiZcu+WziKrL1hezaZ8AiVz+WI8N5pxK3PBOqMEWYtU
R/3FTcB01xLrZ94I6daM1jOGQ6iyqNrk96PIYusyMXk+Q8SUOMf0Zkefo3bbZUZR
ynYfEi8/UIp2EWEPoAMXUD1BewH7y2bc1ufUyd16jnH10m751GOohoJNCJpuO7dh
j1jxeQ1U7IpFhqNA7b+XT9LNkTgTZU4YlV88TvVIp3vQy3Rt2vRbu2xB7N1tLQ1n
EXm8yzVzVGGmmz3B7jcm75SaXvuFQgkCyj7k4NJGK5PlG/431KunuVkMKH1FJyOA
ZZK8XVjhw+gaFNnruZ/wCFFhuXeRBKQjAcgk3qD0E/JpTe1rsCUCeWM3PxvSxwTs
hi1zxCx6L8HoKDj5mPC4xNGrDggKaUyQ430b+VSLLlH6lcTAmTlF7EAuGJ3h9gch
IracB7Yfo1DUzr7ObGOU4sAJumuLLO2skcM7BtWw5kCMlm//WDCa2maTXxKhtUYy
iCHeoElLahGPr7CEEf2JSofNBNFizRNQFS9659gqnh0yVveZ8BTvzai+/W+yF7ow
kttvMnDgP+PdKaFWMOit+PWzMxzCo1uaT7CCfKN6x+WQE9cpKMvXW17vXu2mqwVU
/FwZJBY11ZDmwNUuQS4UgYW9qacxV5i//Ewdo0uqVYPaW2kXbzSakHtOYm914Sz/
KpxBebhf+rRk94C730yqnfW0rNVB7EsPcV2+Nc4RvGqRTpSTk41blpnsANGXiih5
O3+zARGuDtEsOw9PgMKt0+7P4a8nelmOyLsU2nbLeM6J65PihjV6BqasJmfCEvl0
ShgwCsIJFVY+DsIvHPzasxCLBDkf06c5xbun7yy/+LViLoVz7tHteSWLgAlFruy6
ZqogoQqZwovY8vQUYfsONwKOqgKbuywt20D0I5/uWi/HHnqkNcnwcoHxOBfzYmqP
QbIoqcJf+EsrCR0aGyA4XaZN0UweGy3J0SrFPoOOmH8Vz/NgFp3sPIigxfWtJ+MO
lO1FoIZGGz9tHKKrFRBt/zBIfgFCqY+xqeLkZc2SojsvHjMRzdPQEZJFrd0ANrwP
snU/woVh0jaYdUTdtM/FdI09/qjr7mrwxT3wugjrg2Cz98XnJ2IooMTqEPXypLfy
pGHtYofAqiEHnmDKSoGoFKCAXvXaBuuzRVdcntW664yUhhj6UZupB8H9hqYyei2Z
z79xEFT3+FJgWu/GOqA1JZ2W98jA0LXMbrMp6lZF7zsJQSOBYNYFf6ZJasWu3ixe
K559HKYvziW54o0URJlLN6RGhkB4LfFXMI68hlJI4128TGLcnzT8MNEKk/zUS51b
wZ4yxr2N5h8k4v0xYKnIQyfof2EmR/6yW29aDYWF1RlmJ0m+9p59iHPBs5pf/1eZ
VexyKSUllYTC/hsqVGtI5JVRZ8Q2UKrCV3wWhcWDjn+iutWQ4JQEVdGboaS80+Rt
SsZzIUfJqJIplSWBBdYQ/xmQT+uihEobUuWLna8bIFIxFprI52QLPFuak7jnlnQr
M5TIv4q31c4EGyQaM6dxDcQRTXn3BD1CpfLuGKHUH4AsJS2jTd1uYaulh0+xi2IQ
56zgfgK9F/Yc2zudiNH1bfjL5/p2krq4KnZHlFpoyciVM9g8tdt9n+w0WzR044D0
UeFU8Q0a2wh4g1pl9TWzT/Np39dWFyZ5YEZ8E2O/8cy2sOkNHvtGDDZXME2YiXPF
bbB5WkUvkSaMIkck0Zsjju0EqLvaaE6AeodHWZ27xEehfgY/FJ5Xr/42IeH1GqiU
U+JHV5D2lYp8VEShkabavCcL8kLHzfWhgwfgl514h47RklpAC3VpxfkTRIVXd6X/
D/JEVHNKSFfgDUwwCSvfYD9zx8NeWvR7uzuCSPJz4FuEe0wgULwV+PPwNhcT80NP
UfRLukLO3p2LiDcdwhrU67iW0gwMIOPFKjmH0nBsBpcUr5s/8oLMqKXQlsW9qFpY
qy9CpCiWS5C0l5vGaalZtpIxkvzb2oaNQ3pDgTB2wJI8sorqEPRBKURd4FoyXsvX
2fP9QqKSgIc96j1nvC4C8GySbRMH/gJL8Ef0fAqHef141w04MNNz0HnEhaL/kHtP
+jiGaFnR7fvc6pYzjuFFHGZKNxO11uBm3F+YIXo2TQSTahdyEunQs5iAHjScal4G
oSCWIzUgBeD6zzQ2spzkEnmhRqqo1rYZtobK5UE6gOAvY06FiD0powqW5f5rfq6E
X63XRnci8y6QvTYno3dLdushEs4UHhVOVooduHZ2bWMAC1Yg/1W2eyILIMD1NbpK
EBf8CVmpF5z3fx/75uDoWhpemB234cQc72eI7wPMTt3QTo/y16kYmUXsTeAi6Phs
w624MgQbKMdA5JdIbz1RzNz3Y6y6NXBx5KtKKUBuntjttWE4D3+mng629yrlbhvu
b634WRsPS7Wp8ViqyM8VB3amAB6wMLY2ilPOiAStm+Xw4PM/zJF3+oVA/AiqLSdg
l6A4Glto20hJCHwkv5nuDiITR0123sKAMqoy7mvJVmERg/YHVJw0NtVMYaVosmmq
Y9OapFJVbsOhw7wnVpYHQqc8CdDa2qat3/Cz27kC0GOB+9W23/+sj3bK9G6ZsMDj
QNoNYJZHGqa6+rTIKVJcnA44Wok8wxqkmdtOD4og6HO2dlrSV2L+57sN/7736j/K
dm60xSt+Aoe+m45/TmQv31oOpN/g98OgDbY2OV7PRnPTB7iCKC85c/yHzXjA6KMz
1RG/Rtt+0dxqOU8y8x/idBbg4fsTqn+zaitvYSJCy3HFdU3Xpup+itG87Mi8rzVE
9IKktYJreXJaLbZ0qPpvVGWiaa74qgkDcEgnFNVMgShzoOfh02mLPJnjRgIAl1kp
QSg4EDUX2eCaGI5BbUubVcTsDpcvx5Rd3KIJxQUOfa7w/2EQ7TFmMYF3DCcwdBmN
9ofqrTYETEvK4+8/d2MlYyO1ey3BYE/JZvhXyTiHnC3sGOQdZebcVl7iGTj5vpzt
QUPsnlJ2qV+MKxpNnlQYHdEojmmfg86GSOOII8clueFiNw2UQBfld8Q/HELSyeCr
MVfd7Lhp8tI9Vw32BXQ49xNCWqyclfqd8b0cKFtXXh/M1965tJZld/ZAJRBDFLLn
cGgS8IMPLNyxGkFADuMpqH4E7vMZsKZkFOAlfoDjPKD/kWcz7hJJtIfVdIWi8LkD
V2CJoQvFxHL7PaQQqZ0htryASUXb78H6WFNXgeCASGrBt4Rq15gdLrOB+U3VrGpB
Q0vW2rsYcaLBlN4N0FPas70uEGPpA8l8xyrAL2naLzpf4IJ1lwRewf6iBTH1Gw9C
2437UTzOoZUHb++PtRcednq0hSoU9TMaKKS/klVPYP47Ock6JzI9svLzsD3kBhQa
O6Lrk7wdoP1Niee8Do6MA/qbseA9lyWSrjhT02okhvb+Z0pE5EVpNiJXCP0JbeoU
whMAzordrMYFZ58Y4jfrBT+FWQ5p8n8jgMc2yz9WyYGTxT9g1etNVmH+VboNvvZd
XFxBVCDWVuRgQ/xcJP3MvV6gwgYA8hvll0gP+mppob3FLUhF0q0ILlmDBm/yzgZL
zVleqKre4J+xTKo7fH8MgTCEUQDKRQJA7HUZcUIp00CCsay01X71shfnVtDqwBBq
Tc2v9eC4BmcV76wt6zy7+E0A7Z4D2l3w4swdB8ClJ9GM5RnuYDZpLoPWpWnaWu/8
/aggKOVSHOtRHoPaRInYAsstn+wJen9nU9FeshN6OhXfJn8yEB/WGYc1PdRs7U0w
y6isJSb+w0oK5g9yZ2HblqpyBDmTHmIPUYVITFg/gFYWmV8oWRc6UFa1RWjI7o9U
40L2jCq5LA/e1J+u6RP+Xu+uzKSIfxn8hGb7Zni7D7+Wie69s8PUFGiq2/kTrxub
RX/LhbqECTFL7qYORqrq12FH6IE43PXTcFgBa/c5IOGOFYTfe/uDWe8m0yx9xJWH
5YtJUJ6FNzr11uhRtYV85zWkXoHGwCO4Y3oFgAGKtNm8tY8iG4J25MTGFqcvNxpC
FoOBQarUICzpFJvWl0hoaFy6wRnLikGZr+HISEF/jkQ31vgxa9NeZz+5vtw0e2sK
ssZjBUIwxfBuBkN9A5J6sYs26AL7hVMbeXIVntuh3RyVDdJyDerHyWJF+HAaVZbk
TQ4Nvo6opb9QhpV4oMWG0ueQCkS59l5CEIaYCDZCncxpuDR7qvS3yN+hy2HGrOGr
J2KobNuQYZfkUUoKRt51leTLXNG8fNHzYMowSvf9rcl8e+nI3d4JZKgbRhHjKJnP
zPaQj4ulLz2/0YRCp/DessPTGRe7dhusfu2YtIFCG9waLlkP7cl3t8vs/YFWg3Ad
tlfprcWljEvKJyal9FgdL7Op5x9MpyEHrnyJH6ldpDT2Aym6Ulj3StRzmvRboazR
LacgyB8msqhx7Jsbd3ILbRXP2mmTG+ETDilBfE8NS4u7zC3BDN1hM8RZ3lm8ljkV
o1HO6TEqC9spDud32Fe9FZMKlCCGd8CU1Rn6ZWRC0RX3zwIDjb5+mM95GbAogBLD
JptdOlUcpbYpTsDqWzvtmajnoveflgXx5B7OdS8PxpceTySw2OOCNxOVKwEUDHyY
Cae2JuSd65u1cvTqxLvLtir+Sq+K5AOxKE6Yy+5g0WedNbGSo35Pq5YBTdrBXsaN
uQKFCM4jwy5Kli0lJqOLepSUfwX/5cv0gS/j35QoAcZK00gHaToeAX4L6TTIxflY
3gdb48VB7WS7uNGqYtmhIyNuWrmV31a8ZSLYtg1wURKHI/kD6xrCl3s4xiLWoszw
BH7uHU/w4vEnJHidtVJrapmwM+M/kuP280PY/0w9dPbiOSytw1LIM3UGmNc14gzA
YtnIyYSDtAxyCBYVcmHT7g0Ff9vNAh1nDK7aK1aSp3Q/A+xGNHP+HVcupu/YHPtM
RMrjIt8z8J0ybKSGo3bjGUv/1BnM86ncwxvL/6ZcqsU5G+p38gXcoCyVHhRjS6OO
RG+LFgQYufwYGJ0VKIPSpLDaxVFTKDod4U2TmMKwrWDUqWH3AkgrayZ82r7tx8uJ
mOlz4LBZfUOIfvyq0NgCLRCbVHWC7tNrzetxzZOnmrS83hDn0qEYY0YzuZJpOogM
C2dZrC4+OgG6auyU+Pd5JhuCWyv3dl54PJAzEwJ5AVV9uqnMePKHCDxyRxBgRY5w
jnY5YhiXRILe4DMSI7mY+Mjm+uYkXQ6iCAY3y+bwd2dAfwiSkvKNZ6rrJep5lecU
8YgAOBzJ8Y0prsO82ySSUysfzIqrkdoK0IE3Zw4nM5EAJkIqWd7QmdeIl60MIQeb
Ml44tpSGXmxWm+oOzLZSKi6tyW3j0sDznGuLc0ajswqL/Rt+QA3QV2q8LMRI4JgV
Gzh0VF5OT5GcsMIZxhoa+lSOTE3zQnGriOcrhqs9xGJqamZvEO7syOsNIJgTAzh8
Wm/MTLF2RpkRsZv7Ihbh6L8bwXNkKALCWuhiNupBI1SuausTFaFjgHays12t7VCK
SymvqQ3fe9Us8wnKeiSfeTKXUCjbKS5D5ppVu5HrzNXaiCT3+50vC9GSBRHOpzSa
nAe4GvGYGgIguVH3q0tFK7mB3PLdIrLXwctjePhnxZwjJu22RKDPN8fAiA/bO4m0
lfWb7LpDKdvbyWH1H081Hziz4VttU2nJqeFfUrdcdGgLnb8AmBXvNaOnotXL0DVg
QAYoCfmuw7OJHU0Iq3hDPmqODtJGCdHjGiE4JY/Mlf3xU+0E1t2N1VPvtqcfPDOw
z5vZTLk8e+GbfecK/IWw8J0aeIaPicPol24sAOP069M6MsOgxSjVcM6/D5noVSvn
OwW46ofhtycsobm1X930W4n/Lpgo+NmS1SJX+SuzckiYBUKjuyq7heEWXgw5bVUQ
dIwAVsTXNGzr5GH3tJ6YCLswQy0XMz6qIIUE64o6SkWoviJpkUevkz/sSPK2i2b6
EHMyrODfTFf6N7tTdCverfygDzCo8vdDqT1CggIfqwaLt8D2Uq8ZakKwm+AgWie7
pJ6tKjdubXkaN69G4Qa6GYe98tgeUZJAg8KU+HGA+dKGg3voXvO/ROYCeZpW5tjz
FA7MBrrTG+dqHHs8SAX/6RFEEKeNlipsBeMFNcDMmqtdYwabHYWSPWIiDDTKbi0v
xZm9aNo+xb+NO6V2FTbUF/1Tv12HeusKVaMtQfvhGN9rpauM2boPLDuq1ujy9KRm
zMLwWF7dZkpNtJX5iFj/kHD4vfPgb4ms/0HrXz5Ht0qbZwYapCRI0GPZtBNOkblB
MPyDyEmqHwuWSxnWsTIpgmr7IdURnCluG+wSuHvhl+TPLa3vhG6obNmSwVjJkZk1
owUJLBs4szX5F840gZnqlwTNXmxx/sqc+puqcuhCrANxYGRf2HWDHgUOpXwYqpTn
ipE1E0qhQP9N/HinpfrZPi7Ta9/vzxfTjlwUAXgVg+DPw4v0Vjlnad4iJW7YAsBz
bWmYDTE12GV6i+9o9uXJ1H9v9wgXpAHRqeG5E2zVomXTjwSPLP96uIFd07Dszcr4
CcrXrnWMLkLIb4UVJi57X+HKTgCxYqzGY3Elem88KFg8CkG6RIV8a29ckYtmf+0Y
aKM5Qf+Pl8I3Il66AIPVHqtLgR7osGUWPvF1dZ3myo8thCBIoTQ3Mt+MMVhroGby
boR+tzM7PRkpWHiVOtnTpBv7cZ/6Lif38ulZpval+FtSEpd8QK7Y33pUq9MqAFqS
bLtLpp3hQaHLX90286D4q09wrN4WD/ynQ2cysAH4EcBmwU/a2DTDUsBUNVEx/909
4IeljvFzsPG3RfyLjVgNfCUKbSLLezYAdtTXEdq54Hk9VL0iBJoD4cNs1xiEX0SP
zXXxwHoKGbz53/yXnP0Ur01W8/nVKPwV79EqiSq/vKvYiU7xHTUH/mhvFojrvQ5f
exSE+JoSEXizWNwvEZAAJrRL0rK4timNw8AtKmcuw+trWgDw5sjODriCk/i5K/Y7
CAu2diEfr2L1OZhZgYfb0+rLGo859te7TGILL9R3gSiQG1sluFm8/xj4NWyqDyHi
hhLWWVi6If/A7LesC+3EYx3ARrFizlFB1ksRXXLAVjxX6SOY/BftzOlvKWrt03iE
ng+cbVcKFIaRMK8lTVGkGBB1AD09m2VDp14WIur2lU7aK7uRJL26jB85Q35IjJ6x
jFtmfeEHwRjung2GqrFKb15mnhpoZt39TrOCQ8GN2RvNeh2MIHDyb3PZFGFjH/uW
Py9a2Qte8G4YiqRpipXnEmih/uV6BC4F3rsa9HhOxA8QYzveCW+ZZhreNhfzHeOw
Va8RVzVNc08J1pntOJTe2EfDUXseP9mdhnKG8LiXZLXBa0EdI5CZEPbyLhFwS12I
4/wK/k2n4j7HEgReEAZoMi75TbcZiSZ6nIz3Pvt+yNnjCnBPN882v2Pol31+5NUE
tuQ3LdEJtaxgLoPIgY9rjNgwGc4y9sxYplOvAYdWXWpiGzE7SZr8QUEEy+y4VFKa
HGXPBECumVnwZNWpGs9dInxcX91t1b3l4MnMEmK7ccuF8GciEEjBcDHjDS1kgxce
zVEbildeHUcrURfjnGmWC/hRrUNB7mQfzAQn2LT9OA9l+MWPg9pVnqg4zgpx5mAY
7DrbH97zJRJTLjPVz5AkXg5+f1HiaoCbAD3jU+LrkhKVlP+raKYqYKNplBVHgNcD
yLau3wwF1wr6ACNW3s6XdbfPftzdFDGi0Bo4Lg7L5ybckvLRNjzaYG5n1VBdKhbi
I6G2QTVjGr+MbDgjokqa7DvF70cy/AoiPsPVcRB3ROaIBskszseOMUkTB6VlVAr+
hZqGyE2gXHr7anmoCPDwf5oxQvUGzQ1QadC0EoCBoRao2kPgKA8m6kKpUBKhsagT
6uV6vz3H9OfIcEXijkJOd5Z6HpWE5sAQCwXltghIPvTMNbUsFWXykSifXjLCAkOq
+PyOOUuHBFJTXyh47Jdw2pI8voWtT+2GmMVMfZqoPfBhZLlOwYLYXOIqUGu49xuE
37Ybz/DaoMh202Dwvgv6sTjTevfDLAZjm6Ztiiv1YKS3s3LLfs9BXgHA/WqxL4Ws
gQ9jQO+iDtNgkmRizQEJ57gycEEr+p67hn7Y+tx8VHaSjuMWmlcEdSJb+FaFlC41
FhPm4aEQFSebevvy2MgTvma+ezu+NzQUHb1weyGmSMVdUWF+Ky3cTkNWim964czr
T2PFG3lINsnxVTePFOUTqvyloijZDUAiwZI1uK2GlAfXbdYpVTyk5rn6ITxxsa6f
V4/6+6sbvp4yBH7l4yXSg12uzeRdf5oH7iUh6v7UIrwCPGjgLb7oLBRFtgNWoN8Y
AmX6ntMF6z80j22Srr1PT4Jba+8g9M1uJsX+Zasmioo9UDL8+0G4r9nRvjF8pg/x
sezodnWS5N/5VYIgcjTlZzAGsq3n1hY+FJvZTLzCS6Gpm8fcq7OEgGg+1Isr/NIS
u/tBvVldV/N4HtJzCzHqVz8AxgkClKFKmcyo1SU94ZYN3lwHtw9omXBBmBwyRzSX
QqNtgDM3tRuJYBZPjUXTVfoAFOK07G4rgD7Ii1NyGXvUitEXO56H4mxCZQIKO+FB
zysAOKDIDpOyvp9IyvdaAcEtrHdMcdS52XWf1bbUjvheJ4tC6mhRuGsHXzUQg7R9
Xc997ExoKDaG004+IaBRrzpLRp2m1dxWuXOStmTg8l/6tT1PiCdQEw+QvrTj5nQD
uGf7JXlL7kSPYOvxadabxN6tKZ14Xa9CjqCnbMMABmCWcglhROujBVLmxCli+1iX
DgPgm6d7D2SrxL10dYLMiTDGgKFp3PVNxTTKSYsT0hKuzNrB/QRnCberl9bRhGDf
e4mJcp2fHBOeOU0jm8V6stSAhY4oGUj20lV7/0Q9JJkB+j+XtEZH3YNOcCXU4eOe
Qt9R96yswVpSL5CPSNhrhCmTOX6o+oI9hiagRACLSXIkLeFlNe3W1IOES2VFpnf4
/yLVvNAYG+Zo8GPxD+aMCOCcOi8bHtrhi6xNgsMuaGT6lZx0Vn3JFqPH+tiQp1+5
J2lHXG4oar1aF97ROei6ngFo4RPfDMN/ud1273gvDhE2MyotXC0Veq4GbS0WpLQ5
NQOVhNfNvcwTwzNU7cItGKLI4//YYmVO4POfujomNK6GfWpQWTGMzPKnArtTxFge
KOYs2ktqj5zHMdeuNI0/IZovcAJsyBXZppGQqT9MAqdISknE1cXeRbG8t//UOyo5
9Zc4m8m1BqOJ/fo3J3qL4LivCfSfIxIU0KYgUMfHBZ+mYrFNZS3tQH2NT1ZzFMS4
UHWxSN6Ph92onDV+BYB0U4H1l4jJGjgUDuYTlnXifMJZrkz/crRhkZAwigHthIl1
wYQYFv4fSoyF5Uvbu7oDU5fW3685ja37ElbsZME6Q+CTcy1XDK06lEr7TbcYK+jy
mgskSBj1m3kB/CXVgzgt83MduPObUlnzF66/Unf2tx88R5TvhdMlFSiLSC7L/Lbv
nqHee4nhOi6ishPGczYBAP8v8zHH5IxkYogp73gBRuAXmdfVjgjGqB0DL8N+34aP
akxXDp+RJnpSPVu/lBYOf7kPYz+7ZiXT8HFbJQMmtTrSH6bYZfV3/dBDTJSjKVHS
DCMbZT1BxpBEDH2krmmfDr+bHgKlLVYBuWr/62aN8BGGFSgFwSbZxjEHIJ9TpSQ5
DtIbZrCs5SLltkGEjjlE2OnkKgQjx0z4Bt9Gx+h3MX0kxOJ01/Z9qg+1c1eeH2w1
DT/1IIgW79xVWPZMhmzFOUAOAYIousd5qd1wkTWMeN7JdBps2XWyWad5m72+dJwj
QAAbtcsynSWtPWzG/1TpXjpL4ZfJG52Ty85PIADPYALP2SqrYQnRnU3uFb8J+gqv
PLlvvVf+LB212e4NgYRyC6QtaCRpFwkGX4YKzpGd0gnPGw+Cjqb371W4UfaVhSG2
tnRbMb8k9RlSo2Av907FWCiVpvxWbixqimytlnzooswwVnW6UrTDo1bJ8nh4mKBz
ZMoP50Di8XyuTFd5phHb/IeAYAw+fKj3obRw3uvUrrBG3QcH+/csymTAfabar1bb
JqLvaQZwf3oqTRklb718N5TIoviRO3rKeJ8HEnz4+sJNpyN0+kNU1YAVZE9wLPoC
j/8QonPfhU/dEd9+GDQwm812yd+x/T1YxGLN41/HZyk+i9MLwuL9USTZbtuJeWnm
RF29eQyLBdDicqLWOKTdq5IAvGafnA5PLnLKkFPGHDgcoLQib73yk5pRvxDw1c1m
8bBpAb11dtNje4va1nT/gIq548EURRP+spwGVS06mLVNmPjv8hB0+dEgLjEw/OOy
kXaJCH5K7AW5MkeL6JD6lhYIdhTh3ofCcWL0t3+UEWlqHtkHIVxywtwWF1T3bplJ
buP2t73X7C7KBsEfxyLimiPdK8fJoBPc2qI10VTNrWairR1Zv+60mUETNJc6PDMj
NRjwJsD7g7FMU19vQgPnDGUE1rwc4M8v4MuixaMiFbWFb2XZm51SO7ONDkC1Pc50
QPRwbC1rpqgYmI1kjTfRSz33c9Zv1wkTo/04do0xLmEBPrGU0Xa4UOxNPh3uOtex
M+/5BQTMgQ/smEicrTHvKjDLRDXgFaINlFqq5SJfPYSTk+l+aAmD+5ey4awxodz9
OmRoAmvF+ieHheH88lS5ypdwkAyNfEVdWSv08kvfUmeHthKIhNWRMH/WNJ/qFSdE
zAi27bT8wi1XXygweDBtroG8JhUnRGK31fW3H5AmsCrRaVfAjFXCJG1SRyWQO0NE
XnDqV0J/1vMIP5blKX8Jyi5QJbofm1/JTtDhvZgagqHLhBnH4twfJasqNA4FqHE9
d/I7VKOOlcYxDL6dLhW+adcfjM8vW+TnTDbC04ZL5imxxXZxiSIXXoznipffMnLV
Q2eKf7lUJ+5xjnu8/mTMLVhfY5t8I2tvxN/Eku8V6sKHGYHzJq2+CVXvfaObM+6r
BOpolFLoP4rPycNq4qYh2qsY9wdosh3aZIhjKOjzSXIc7Jx/LH+YAG1mvzPERNYE
BGwY80tSNCzz0/206nBwnuK8c2skL/TdbACwWmfRVMlh6W7nF+ghQzntOlZ1vFUU
9mliHnpU2m1aiBB5R1d/zYwvSgQHLQPeMba73PynRC309HJJ4b1GrXAhmHatVXgi
E0eyhXaSlx8NNOeZUYFgsp1ziqWCwZM/Ko3azt5yyiC0zXBz/u536QrTp3r1ruYe
WWLW6MQwEPi9njz9td8pu0+aD/YUFdgwep8sLeiVa073vw8FEuzPG9bcMheUM1AS
xRoxXmMVDrgSiLrNid8cVNJIO0s28QY7ADLoaj6Bq0XnGPyv1EFxLQQuTi5lTzCT
4QwvGqvS2kc59zrMhGIXtYnuwOL+nTlWAGxP2Z3LFVXaeNyq1MUE48+lsf4GcFmy
w+RWNpkaag7n6eO+dN9VidOHpDedvts9BEZlQsFlXurpfcANlbdHqb4qMaCE+SxB
fhlVSN2RauGeF7O5UbqijmR/LE0XwQiLfc3bsv1O1qAkurZyJ7e1q70K0BGK5xMy
TbDeLrUspT4nWtBTZXAbcB/g2UNa8MxGex9LiBWwHGhI2p/QL5vnnYOWFoy4xaFb
n62HUsBR0vvKw2R7wDEpDiIwL6nEzQXKiOg+2/GPp4ogBfnBHf1MAfZKcOey5XdZ
gBbvo88UvxSw2CA8mbdG2vdydaNlfH7fufmGPSemMP4yYAReXgIHCkKrmn/pD5Ej
vsnT6h+MpeeyYv55bs22QkD9ti1u4+wgFH72RZnLBOIKlPMskfjHe25goNlE4mky
8S5GzUjFFLdzKN8rI3N+mcy9IS1oN5WhlHUNvfNS9SQpsOmLl8Ep66KKU5UO8LBa
FdljeS9i3LpIJrLBpWdBi1DgZZp8sDFiSN4yY6dZ6j6zKjiozLQJi55qap3ey2fD
63l2C+RbGJ7SfjHOvxanDLr3mqSRpW7VNX/Bl6M4+KAdEUVYXR8T60V1nWhMILgq
ZuoT8op+hnEgOOXhlDY7UIhnqy18FGeydiLahtl5Nc/QrZZsFHBlPWEI2SRqWYcO
IKJXd1a4+r3/SeX94hnd7xmQLBEhoXy5/oYivN4cVq+aMQXc5gW5qmwJhq7sT89o
t0XABdhERZrjqZBbJ2sFmg8YRh/dWpzBCystpqRhyc+vPsvJcuHxeYRztjPaAWNJ
MHACwQb/rXY2FXAQL145H+6mA1hP5/Crm1Jd4o5j0rlfbMWyiTrUgfOE53gtFn5M
/yzRcAB4qphLByJLKnRovmLpTF/hw1apIgcXIGjB2uko/R7hgklea9BwS/VVL/6J
i2MOEJSKlJk2/6HM3SbjY+5VFmD/3gDHtiYCUraep9FkXQOPepXOfxpM8TqJbj/m
M7oH39pCIgi3R+cniH2hk8t9OLkUsIeJe/LCmdMCqyMSE7pT8WolP4FK6C2EtPOn
Nhdp8dzx6IET8HoPLjtXHqQkOiAoPdVSMkuINx98nrj6TiQ+8HX4XaifUjE9X/tf
pF8Xur5rnl3zgVhAe7YX4dXYfFk+WR8b/R8X37oarOaz4hOpfEcJUYLo3vH8qSjC
Te15xoefq0+rK/3ldTvAENg1XGeHLX7p6W5R1BKM7OhudeNJ2Ce5iXbxjPhAw75G
sf5NEulD7Zq02woC6lI1MjUNHAw7W3rO38h4MW/FrD3ID8cXfUGSTtoxY1fYjFqQ
uZ5BHI9Vvu9aQNiniKZ0zgmF6ZXKwvbxsV4iF7+/5jp1BV6XOO+ogLWibV8VZrVJ
AGu2ZS8CPqxvc8DaQohmurH629kbk1GSP1oozsRtWfWLVA11nGIdAi6Y4uIrKrK9
MlyG1qYA7pt+wVy0DFtSRlePzDkofFBT/B1zOsUdCmmvFHFFbdD00PlnCAgJKZVL
OtGGcoPiMoxWt9YQgzMov0cQQM5izpeD/1pJ7y0bP+ddUReb+miNJhIaFm3R8iiH
rq1lQJS1d6qP5F6MObac5BGA6jM9Vk534eXiVdJSNfcrqBBMEU5hIxMQWA7moM7n
UUCIvVzFHqUcrE8FR4PDy2QOB8O34ZRFMK8F89AQKO6Sixfivl8G3y0dolsaExs2
dEwS/EpwKSD1LW3Sh1DuXtKLyykZQg82yMiwhWFliupNobiK5xWDxj2363KZb5TK
Y9wtFPpFbRFD0Jqi8KeTqRGFdkWjQojdH1YA4Zxk2+pjaIvIWOxFz6T2LJEyvvcX
Kdl9HLq/otMzy1o+NxFpgiiWFdj0ZihN/cgAHehCUU4hAR2KP48iTqcJ4M+QmHLU
fwxrQtI1qQMawrRHeqOTNxK+IuhWc6U0vLs0Uu9rJj+vSB4AUXQQLamHglbnrFvD
hGccFeNlWfPjuv91zElXEGkBalLCTsAbBGQKHsxhIRn4c34nr5qrOTbLzwPAqhG9
Ku167wGsE0UfqdyMNzXXbwa+LohbllIXL95VV2L4+SW+PxHkwmgeXgeoo3IHKGGs
F89cpxasIjguKRuvDg6fbOLilyfVdiMR4nrKRXthYqX6/F85cHAYiFZ3JS6PNzX0
eB95UE4oBe3Rg7wh7Ec5xyHOsWNcpkqY1E6gxa6iKfxWnoCowYsD+OYat/YSugwL
kq6WRr3tDVTMOBKbIp/KsU+EV3WU4k8jYPwU7acovel+XrWZlQMwkbI1izaonANy
oxJvNwTXIPzq8EciQ0VIS16U+0PHIC18Ckhfo8XMItKmnFMWSl6T46+03t7xRnyk
UciX8p6PVY0xLfMl+7xqQ8WnVzc2Cjq9Navu+ttnuAal+CJ+MxbTdYkObE8u1DLU
JDcCcJq7c7dDrWeZ1u7j5lF8A5kyN4W6QY4APpyqbIs1KeKzszCqC8m9PxLdCJQb
QLjUbx+EzlIZrfVdz42w2NHhGvJ/W+bbqaFPK8D8XTQtITwPXY9OMcMFNPNON6Nv
awiO7jowh8V6N1LaDCpWc7oDMfX314zXu8Jm9YLRDHJ0LGzB0A8Wf0VmpLjiz+g4
AL7UebRDHwgFZIIeppy7GCnPUbA2Dw+IDC9a4HZsqZma+O6yHJiDLrCInW//cjQn
DSs5aXa6O8dJWSznLaF6xAV3s5pCgAMRN4k29dROVcwDuqzj4OG5IAKLth43QfEd
OezdKmr8XHQY3M+8oEMhUckMYn9EPpmdPlbGRVB5NPRzRq6gFu5k8UAqWAvnR0zS
VBBtq9lWednGDfNHbUoegH72emMQ++HUKinax5MowlK7bZrnJhH4jhMiLpDEdS3Z
4NyEHVtonEpCvpDrf6w1P3+vcHo5BRrDwQvkzOMBS742jE0uRJg+pKyFbZWw7IJ3
VxD88+2yiSQ2m5jWVGpD9aNtcard1SnMfnafcFmLE4QbUCUmHcnG/hBa2KWA0/Et
RIn9xP2LVkKne96ozgBcA8hf84ZoOF3banRdB/uesRLr0Qrinmr1AmPyo5+osP2H
SiYdhbClcBU5GhE5KE/cNpsoBs3w1QEW3u3I1FeE1UYV8XQcIeo13A0g9whYLgOr
Nt5dSb9SPFcUjty27Tk9F7LvR59BtVRDawT+Roc6gpDtpxzCPi3NUlWRdp5I2vcb
BzypY32ZemDxDjqA8543gHpZApN4dIBkJfHKlyYJmVdBB3Xu3eSDOyubyrhcqGtK
EYN0+3tVSyGHT/EXFzJZ1mzaVYO0z0Mo7sIF+SgUNx+GgqgDfII8rvHt/mN4+btP
g6X8befabBc1dzN4QnBH3evEVKLhl1agzcKBsb70YoWVtN8RIMQ+stBLaxAoFHJ6
XxaFCJhTXAt0ggS6sfQMB480Kfs2h6lMHvVvryyTAp2yzVLyS61NsBhtpBQXH/ao
xkDgGft3HohKsh6KftlvtFmSX6Tqksa2hpE03CxguVttLm+3Cc8NLWr95HIGfqub
5aD4HtHAyKF2cusp7i7yKLRxbZdTEmw+9j0uT8O0neNBMrYKxneAHpj5l491OFX1
i+TsxWXUReahBerY0P85wDyzGEp0XRZAiz3VDuPy8Ys0nMI70YSfJW6s3n0YU7x2
8b2H7wiQD0FmzaVHUf2r26K+NUChyWpUTjNa39UjEoofQPp01DnSiUNd5cMZrRjJ
wfpohYTiP3pW0NI1VO17F8UY1HL9CfM+A4b6x+4WpvhKiqT6KgliWA9PXVWoJqv5
7aEa96cV/2PxWZC2V+IonbUdvy2VZMEDyHIYQuBLCPUKjYz89oiyKKy8bK1Hi7JT
90iJ1AcLn1Rq4g2KRudaDzdXjWOzxr73ls58PueKIc1eH7lWJdV3P9fc1TNzNq56
4oqTfIBotK7ooFp0Rgkv/+V4kL4rLCdbgSIhh2Jnc8nSWeMkEb+680hH9rXhxMNJ
bRmRligulg4MHVm6UJuZ5iPttgMeasxodCQ2Esg5E5O08a9WuRTZJuDjzCQLyj5t
t3rrXcFGv4WcPe7vSBXp6ObYjpmm6sf7mFJDRDj62Gs7ZwHSm5XPL1qbZs7sU3rU
/4FyWET06L3z3eTjShaUHmbZlAqH+nK8lKUPX1odTHoHFR/ghIuos7pLkQMqCrgS
zrzRaxN1z+FuP0B8XatcLWzfKgMgNJVyVgLvxZJ38zA8X8AywhrivpDwpv8t93nE
MNvw93S0oVccafrVpFh10Wqoq7DBcoFk0Vw4uMYXfEk7idfU+QanwokjxqEUcVfk
yNJAJc9ZQ3zN2+GsbULTYqyVkCh+fXyNr8Jx066l3o6xlAQP32/Rbn1J49yEU2jI
iivD4ZFYYgUfRYdYDaJLyTnLmuavPhouc5hL7M+tZUxC33ulCu5c/oaW8cfHs9p3
4jYbLWMyzefjdGO3CVL4GCXBkXnatpHx4U8aAYLR59ZvTVkWfCHnEHg1HVre+mN0
nDtCwTWsdP7XFT6989/HzXWROON8lzxRzjY6Exn/Kv99615cECjQcWsQyEJGSkjs
xJujjYI9RWuGtGobYsVlYOcei4MMzNh/oO/w4dvrnl1qcgK/8+ElSXkQbETINN4E
NmMXMguJhB2J93dMaJcGK4imQl1mcqkbfMQtCOSv14LwTqeKMsOKw0DL1co0N8Vj
KXUudZ+LARXmBNh62b5Oc4TQMU5SuY10C1lbtWmx85+Lt5Etqlha1+Sx+Z20o7KG
x7p6V+S9MbyzH0XrKkYy8gG912yE+3izoHGER3dpWd13Wjpgxe6cp1Vq0monc1ve
7Yvmo6NeDWGNRxNFuB1X6TGPDAfXVhyy/ToibiPBZYrWNhlWibYLPCj4ElPtzi84
/68TRMOBcQiuEKhFs5SXL36zWsgRpHKfLUCOvR58nokBly41Hqvz8PjeqzUXzF27
RrY/UQ3OmPy0fipCK4iKRZFwaQMwH5fe7rYP1XqrfjnpIK7jefHTZAAd6J5lqCAl
umwO4Q5rhZ3o3Wlyw9zyjRI5IdY5oHfyGgFp3drTuGvZLVfqQbjO+27kDnYs1Cma
zCHh9bCo44KykHJEXLpDtkHPLFK1JxUPmOLy5UwC1n99UuahBxqudtaPLK8H5Quz
3/ekCBUvmP0gKe2eRXYWOMFI6UYHWnu8LAS8nl7w6oobMcfKfAOFh5gIjOpXsAjb
uGNH7ztoO57el097poHD278awCVjhPF3suWetC0gOhAaaJ4xRAVViJaPqdugqEXO
fdxjwCiA/KYpEoW35hVwu8iSQnoZwCSrgzWluUfPlbD9YvVQzSvUazTKxOXhb1IS
xvtAlyQP/Iqgnhx571oIoMHX7KZ05eVRFQ3owQqQ7iPPdqpnfucDudTtxE+y25ZV
AHykhnbCZyIuZ9zaHP5DvBX786qTQCxr2IpQbYLBzFamRlCPg+LMt/cm1FIb7AMe
w5ieyd88gErrmUQyx+rf4+yDr2Iajdr7xW/f1VoY8tKYKEABSuqCgnTQ9t869gNb
Q8UHlb+CD3YWGKpW2WM3SmVJraagxEoj0V6g+bHZICTuQaEQB+QflBWfUWiNTMAd
2bHTdZYMYIEqfU1+Ruo+KmYsA16ihDqDSUurhmRd2W0c+gUYK15WdwoUdjskbXgc
40hIrPWrIENZE6g0hfno0JepCPuQK0kV58xjbaE0+eq+vZb6kA59aGT3McK9B4e6
zzu6GKElXKIq20A9e6tEQLYLcws20dVz4mz9A9MDddZNtOPYtXhLOr1OsppFlUTf
Qy8Nk+6KKqB5HPRzURd413hmosDGpuxpR5FeXzsWTRULkvh7mix2G7XRnBK4zdFX
C7r9nchbPQHReUJrwmQpii/N99oJd4JI98ce761pOsBwzVICrkkbuJvNbv3tmA/v
wutWVMwxxGfcEeDEb8lMST1VCr6Y/Yzngo1zrQBssyztuSKC0h17RD4kGth+THyO
5h+kmXv1l8xVuQ1qXxs2s0bixPcz67A6GMTUKiYxcMWFLW1irfve+WQJpVNYCY04
pGon7pllEXrE3b4fWqEZhUFjss0dQhCJ1TgrtaO5o2nvtWkzDLj12h/+uR2huqAi
E++0ELkiQoob9/RFrQordjDT/zJQkZyMi/SX77Ly+tqSDT2Yir2pBYa6ZaB5hNyw
tdIjIniJPkT2OyEdGPQhbc7ufctxRAtmUPag1rag4T928iDFmX9ZW7pO0P9lkjO3
Zu8mwzbxbDV+BbYY0vgOnc6DqEoeKKLysT1p+ysK8WJzqJfHKDOuoxCIrToYILqX
fPl5KmrArZoDVPxnnBbeAlZbq83FwPUOa8CqPrdUwWSscU25czoriZthaTrXEz2f
0J7WP1LktTvLYYvEx+YmkJbD2TJaOfrm8qqF96kzeWCpSJC0TBMkPVSTTYxwbI4B
XGgVCkxnLs/m2syJsmIsPTTehFZDDXrAj4Gwy8anCFHJGBt/ZDe1OQKFSNwdGRCz
lU/2UgAzi/NNOFpPibk7a/++3RkTyXqw8roupz7eN/X/0QeYkuhh0uul5ie2ku8e
29j+c0gtLFapjGPMrgtbpcgr1dB4NM2UsPfpAjvNRPs0Bwzj9b9+xSf2GqXoCBO9
gzJBQXUXn5hpuM5rwc1IWPlXJY1MFuGLkcJ40glclK4Zp+IHZww7QL09S4OPomPF
fEZqjSLzbj9gOQ3bIJ/PC3wN4YN0oxGH5odwk1S9IT9X7tfpn/sLpaW4zIbk+51u
JvMUn4cwrYsQ+K3hg9+lBkYWlV+VyutgQeLaQy4rlOCGKYL3lj2FN60v7a7Mf/Rn
RFkpMHnOrNIgHtRVwmHyelgu7eFYkOB00auX03k5SyH/z3vMEKAZiAEGGKWQEKpL
MXk01EZGBDKsMsU5TbJncRFUqCMyPGToBS12RByKrC0XMTf0Ys821dJOsHo/AroN
TjF4m5xu1n9ZFhVTu8Uldd9kI7OBGY7d2P73TeHb39wQU+DuJ11iYng9ehYk1bIr
GR2lDWhe3wle+zzC9r38nzG8VGsG9gnwku22ZqBDIw7kJiCkdyLj/WeaA/MEPoyM
mLGPm6Kb3U8X8usyWxNXVHYv+JuGq0SxKyF6XVovIsU1Pa0cydZ1kM6f7lgrqRzB
6wV339CElXrCENaQgqseeF0iydYx0d36NYjZ3rzutds9iUJ8409cSuGt7e8p8pXT
wuzM0SF4rDupTaRmgfpS+g2iyTJKC2OFGc4WxLTwQ/S6SvivqTmHX2wkupfqx9Xf
QCve49/daZ4K5LGPQa1BABzAp9//dCMqAeuIt8Uzgl/UOg6BJ5ALVXGnWXHEOeIP
VSwpoST+ZXur3R20KtmJxcF1xsthiyOzlVHHmz2HAu54VXcmxrIKXvE2IAEH40gA
EJ+xTU8SbP+VnF1SfeH++HeECnyZkxUds0MUU5UrLm+axUSb4Z26L4LpoiCPieTd
nCaVJaNnrpZuaMGAmyF+IZEZadIsdleY+TG4BkTqwsw1KC9M3bHYDs1CxkIzg42z
nB6pvYqlgjkPxM9U3l2Zr3rKq5/iUPWUGM8jRv4EKwl/zucA5jL6P1fvwU2jz8SH
UhUagcwvLnMxf1Hctoe/Sql5wmP9oEft33tyazUqv9G+6t5HR4sSFFXRnSfnseXt
GPp4bhwbDjRbHwpZxGgS7+AtmyL6btcZVua008xxSRE3XPVxmJAYbkia68ywLGfH
GbZqiG7WvRfZ9Cycp6dLiM4ZEzjz+YMpiDEv3CoM2JZk1PnWgAIKzSpSCFjsM7B5
FHBdynWAEJshOgWJoN6tXRXfL7JWe1dZ2IgiNou3Cm9uahmgK4cqd3cjKNcNRT6k
WHMeVsmHAiEZjCYpn8pIjl3ifP88ftuIOFxsWoRosjuXnznkFIk4fVFAC0V+WdRN
NCbldpY9gwR35emoUMwkU1BkFUb7TfskLVL5zjztfcFQDSmwO1lmaDXbbe99Qsea
vZ/9pANOm9u0hZjiTmxFqorcPxbjY9EtF86VSerZlimHsSZQ/TCJC6tztkB7IZN4
k7Z30vV54Mj7+s4Y/CJcXCMt+yjKXO/tdywx9X8QLpcjTPJejCjT7yxDfZLKLa3t
BBIzGCzN4/anpW9QhvA1GXzsq/0Fi4kY2EJPQjZsUIf06XLUFU+8e92QtP0dpT4t
rGd5dZKhC7hk7M/f1CjfKsedv2BxdgEqVFvsMF2UIFi/8C7SHL4oohUYnReck5eV
0x87o5AGiPHlbxOIoT4LA9bfqc+obHsSSDCrsRnoplVE+TEJGoo6iR0COI/pMdah
W3Lz4x1K0opFnQi1vT8erDs+Wpd3Ds0pBZvtGg+n/QOP3utTTK0T6+vYOEsQY8WN
nTS305Ov9ClOUsw4tCOiq8oYFktHbIRTOuNT/ooHzZSBs99XNvmFec8TgP6sSiTC
VA9GVWlY+kdNSR7cJgwPJMHILIPJWIi6RDiR8NiJ0mSW352VLgpp5Z6ZV3Xy1CuF
6MZYP5+legX2g5Q5CdjS7orioaUeJ3RqWTrKEuAYFyw9EtRRJ8dtUMEHnpIVF/pm
ejfQIQjJfHnp6S5hicucFEsU/q+r5gJowYFEtCjxT65SCDA0YyCOHcR3SIoacxUa
TWJbc/2s3IVZaX88Au/SXGkVBAcYrYHdiPuLXC2Z5NXBqgvADh7I67ypxVW8LpMK
Hf0rbHO3bjT5i61P7wXoUDLcAHId3BnMcJeigL9ToID0X9lEqU3bXF1qb+YYnmac
hFfnQ7lRbQ1RRsVoNX6YH8DIbnASyvdo4jNk6sj2tKtMnk31+Pt4LX5WzBS+S2wP
x9ujRw2bLKNbOx3JyJXItSavSs6qg/NP5G+Yqq3mbF5a526H+3I2C829S5orsTF1
r4U/Qd37CQLz5uZjrdZmuy0CvbgB9Jj+y6X1L3IHypznr3kYPu/5eoJ5J7rN9ZvP
T1txkcW4ylt4ptLjCguwpMnjDeVKFi6CE1TVzy+U2fejhf7bNP1GDt+SLu7HSgRn
98yHe+sHe7upnyZM2F2HcYfCF0AoDs+C6OjyKrPDtvgRZ/mbefLnid+GFdOSEsoI
4e3qdiai3dLwgUgoX0BICedc1x5UHpfNVqLw5QahsMtPY+nAcPrxt4PIdKrCZICi
28Banteju42oWxLUWrrbudbca86Ob/qCt1Mum2v3/F7g4k8C66WlJO5KVDbgkoZ3
hYXEDFGYnzMx6iziYwsfGKSrJwt9W+pAhgddXboAzvVUWUkr4KI96umhUiwRco2S
fCXNdqxTU0q3EK42a9kUni4ahEAHx5kr22RsvVnGt418tew+jXmc5iiyqd7LfeNV
NXfLTqdknFmgVky6Pfn0tTUtepR40kIsibYmyPCJ2nrq7S7T9BlLmQwESTOfsLlV
hfFnMGxbH3usu1336YWQ2UVViwgebSh5r7zMYtLpSDDFMHbTtmQiY1RAqz0uAJ3h
kI/95kRmqWsZiZM5rdNkcti1NTGN0R/JMpM7FFF9H31muwiRLgqHhX+TaPWx1Tea
od7wXte00CUNHA70mqAlhW5tztIqaGRlTLwVp/u17v7hJ2yc//jjdVV4beCRIpAz
bO5kfXqSXBTpjlo2dwY5/DTdI0Ncm5AcRJg5QvSNpo/YAQ0Ji9ltpXuDoDVzW6/q
Tc+kwQG+3I6D7q/IVE1R0tlDkoobaFdifHsVblR4JiHmndhKbu0yuhMNfRuZsKaB
ndXge/TTfpzWYkkCLbuFjSdCj32SDGxI4hSRmuUFtJXQQDQVnKKiZ38TkHGMBjxH
+BJ7hnJ1SZM4+WcMWV2KLrSpgXDTuD7g9zPCE9ZaBpzyaMZmiRtszr4lV7PR6top
i/Y6cCaKm0Kcpum5qARO0/VzgL9+q+Asz/a5LrrSUkkU6LowBtCGeVV/dueOc9/7
tZ/sF/QuXnMqUf9FMwtD4HbHZN/Su40sKXJGH0dGIYdGO1rOdKf2oKy/QICpLnR0
opFrcMw+ydDv3vJ5DTV7GgxUoRgbwWlRQPKxjEgPIO+E1P5UiHGArlPC4Y+lRUil
tNM+7KWhi2Kx/KlEjKnfd39T1dbZ8ZOJx36p8DTIZb2UINcZhU0WP5rLLn8t7vzz
aPlclFyG/yFaTAe4DBtY+5KkyYu0Y/+OkrqqcyORkMD+G/2e6nsyu9dL6r/NKGEc
rBpbdEUKZkYMFCKOF0lLUjQ6fuBeIKzSS64z3g/hrMTmzLoQstgpaBoUYNSAOGqu
7XbRcrQ3zzfT9fqD6qeSUdVyVRoKhvqG6JyvoFdvL+lgsQDwC+cuuFfuaNiUzehd
phnYnkMNaBFztHPIsixtdbgbWWdSiYeWd3vBdOu4C785Gj4H0cuBcdHgqVW3v8J5
6y4tw/DjmndUk73SlUVn40d9A0/EvLxHhd4wJAlXIQphsTYuMJ86Oq/QG1kfRwXG
Js/in+969FtJQYqg6Mku3DAAeTCy03xdfIZZ4/ho8423jQl7RG+kb36yslh1DVdg
ye9cxLCIOr9cpoAqsT9Xen9wIm1IfKWqbVcOtEKD+MH4i8NJuZp6Mr4bA5Jb3EmD
pqUdlMSlX0vOV88fV5LUYTr+67FB6Qjgab5X8HuiYViEfGlzG9xSNnBEfoY/TMl4
XL1r+Y18m4jMAJHpNQIeVOK4CgIY/VO/rs9P0c/7xZ2TMTPPgUjUdEbvs2xN/FN8
lVurboC/TY5P6nCTXX63a8kMmxsevlHvDX1BEQheNkWxrWcA2T6F/r2QdbLZZ5lc
GMsbk7IWMPGdEpt0UYrTixAZRJ9VEhJ2yolDIWQK0J9bs3O61r7QQvGlt6/8uYNA
ZBHYg0YZDVOFvslaHk12NIZ7LQkXeBltdEST16Tq9Dv517Z36UCE+MTb9I/rBLdJ
mSSMDWfsagrwRJIjgJ7zVaAEJo05Ud0Qk8bXKB+PqDVqb5FRMf1rmIeOkA9WDDof
G/Js2bsgADwso5+IFGH0IQ9jHRFIW3lbv9w6EZDkfrqz4OjL09qKccBSBh6YLBHG
dCwUDHrg0ryUjtY5yw0xe1b2wUHEQVk/n1bJxhdmSJAj7fdTd8y25FZ6upVF2u8F
TQaj5BqXm+kSlUoRaBpCbZqqD3F2QO3UoU9dpCyukMn1E98K9Sj0qguQCq+XMVYQ
IetAYbudttECa8whdPpDRH8Of/7/rC4Atoq/21RWcsBCY98faFujg7bwo1e49pDi
sm5JLnRzeTsUova6SebuIb2t0IFo/nXYcjZyiYM/YsDmXKXW2YrgxKuMEJIwaU4M
UJ3jWwwxjRMuJShcAXleNFnNdjSzysGln5HwKlrdsMZ5FCVpkfxqmpZNdXAOK8vw
JOm/79mp01eNwDjvE0kLFoxLeOcVMvObR9Y3SC6BOrcSw1OOD/Jq2mB/zmIqujv6
rq36kQik9NRmZmsL4ZNA7SJP/diu0XDRJNMbvWH8pDlQBXruhdq+PI6z8dFRL1gx
hKcQkoRS1Pa5d9E0gy2YGL88mQEvTNZ7FSEu2idrbht/9XppdD1oqXIkKQvuHLk8
F+I0DF/T+cdVCFBkXbc1e70TMcPZMguEca6G5ko3Y0YaYKGcP/2bshuRBx92jJ1V
KP21WkLlLEc400Nr+5PLFTLHn9hvohqIXzV6Csuu03WTHbnDO5xqSTGehoqbBcLc
ybN1GVoVWo9KGVscgAUr+eSEZ9r2Pp/+jFW7/XCDFYvKh/V3yw8TZCbR/wCAzT8/
8cYhbgQBCK2hv4Pr1h6u7uo4D4OSeMgbZiCzw6HTDc1JXzYCheNa5sRRzRSo6x6X
nsOQgUBXVTc5wgSJEW/w+Fu8ksxIpoxF7ewcthDDPW4x4DxTJrd44TJaA8M8Ijf+
ZN/6Y0b3StN5AZI0nmcToilqSn8htj4X0dOxdeTtr2nLQso55MhW9RT/Jc6eVoXK
rjjZ8juSOOYRltfhsprENdOQBpVCclWhFweWIKvhmOB7JYGddyogYH+zzG82oKJA
C+WmFOXh5LnAzc+bl9aU3YJ9jNi6twnvWzazZwDQZYP+V8bkto+EBCB+dg8aw5y8
uFqT2eIYkYCx0Huqzcl2heNmiyZB2xTXzFRSk4mUkgOBMS1K/rNgKEF198rq/stq
6Ub5276Z3BgW67buln9LpA9D3olrmdn9PO2KDoS3i5BjoP/l9LAOzLl+49dchEFd
t2rHAHviSaeHZ0vk1ranjKhtbCQ8k8Z8ZxrU/ZVgLFYojR463wZOrBRxmQPlA8XG
Zd0FPE1ZGnUw65Yu5ejyKyfSJPfIlvhwpKmY5XMbU+kgUAtmwN4Xjt7ojfavm9DR
St5sr6h7T1PujoSYLSsrAOjKbyNn6L3VqZeOxlyp4tYnF8rE4jjzRg7hDSW4HXVH
N+ys8RUYliaVShbkAJ+hXhyFjC6MH33BbEc0cT3GojmdRIInFdf64GCSzPENtntl
4vb01TWJQayHaE9QamdO5E1E6N1rbjGpOIDOrh1qwihzB7sab4+8W0nRDl7E0H8G
UMUw5oDhM+xZ9vJ6WAVWl6qrOs/y55CEvMdzd5pMa8N338A8wRFfsCCsyedAox1n
NIBKgq7lQuw+4NZzjVGs0qh7vC/BmBeDe+mdgmM2kBBI82vkldShwtVKe0jq7qEK
e3bu8+9s6ksG4tBM4deW8ahgks5fO9Y7gzZU2F+VPjAq+WuW3fst/atl/9gD2Ztn
nBqGV9Rkl7PzDMPDFd3jJ5xBQlvD56OvE1SBtJqZR/YH+K+XUj1IhXt5sttAnIRT
bfeVKFfPgndbVoNwrQvSC4dla2pq47g8VFgmaRgD6L7GCYsxPeqef6VAt1J6lrvm
SvnDj3AWvu5OCnUlX+UbQbx8MkYO6J9Oik4btE1iKRTd8SpLO5hNB+YkF+zQwsBa
LIYOdVMj1mGuZR4TEZAnnnPcVXtSMyx7QOVNhsdDcJSzJY0hmUC9heoIap4drzH8
aWpeYVVPQGr6nGbqji0e4VlvGZxKRTkr7nLqPG0znWREOTmZ1sJaBxbXVjCdXXUo
DOTeqFM1oCvfFzojjiYAzwPrOpaSdNlhXFfOLFnwJm7iTMpymGDwgdOVsg6VoTXL
Fbs6ikGXhdnWKQQ1fMl8pysXJSepBSZya6kTP4kXiopp73I1J0k1mta6Hbt9iSYa
zrXYim28VUlDXpDkdHLz6CYGrCfNSJqRk0hu2KIi4sTlB4K/ux9evPFh3EIjUoRB
SJN3DS0sJcDVcFBqpn01cUPKWT3Uv+PCBzM/gW1IxmEIDqglzecdyA/HMA5eeckV
cA4PgLus0maNUhjkVZm7R0Pjx5KUfeKx1ILfqv1eqiST4Vjd7GE7cjkWl8eueUSJ
WlSkzMbYeYN2+P9lY1E6FR30VrO3Q6IplD7VIGU8blyCcg9SCX9QcAlkBCaRu8v8
+wlseQmkGvpCuAKaNasSFodZNRAHaCwt7oxKJCKeRWwKDXX0KW/egEbdIc+LcI6w
4+TihN+Of7pYkAxeggQ0LL+TDOUh7RSEp0RmaDxtUwRwfhhSOaqfZN4XKE4IeE/5
HujLR26/IIunrhtzEK+oBWO2jFscN2VBwlMlbGvNrLJzYGv82Kmw3F64aT4fSh3w
/ShbtwOWIcXIQLmBVE+09BYjWIy2xmv/PiK71CokgWwWHLh7QCyoSu/OPUEU99hw
5awx/Oq/gHfCI3c07+r/rj1sSPSVaUMoSIZRNJ7PyQw0iu8jB7rRz/q72J7xVkCX
0eMJhT+xxS9PuJQNM/JrwHpkPbEvBTVRESoQtABzHqiVHmjCd/qle5uJRdnTbxkB
y/UEjL6MB69OSjy7ST/ys3XpATe+9XG6fiAkdvnRsRyC3lmHDVgC76Z4sjAWWV87
vN4tV3mmGZupuX5FfqElNq1aqZ+OaB6GPqZY3qMFdSZyCw32+2fLy36Y6VcEhlci
h8sIcY45+rgAcYYnPmFJRo5kbTxYBerBcuf6yTMAJRYmZgpBxKmYVemfFHNwRyTE
WNEFgPOBb+1UhnPzo9eFRtYZWHEmtMtsq/c/YtUsAfSMvKeKgItHs9cSanYAyY2h
T2/4qX5dDZRUZtPDFsjQxDiEFJ4OMq6Hf83hnOM5Wgc3PHj0N3pykMIKit2AbLL7
frQborvzlipaq1QZZP7fX0brXvYOnsYKbM/+W0Uzm5+dbQ8dG1mqmDMBv75Xg+n3
4lTrcCZc+GSWxzyzGpAh+NhbA8nTsceW98iASN7/9DGaDuXqOQoF3BWQv24LuMLf
TDFBwZE/xyzIStvybLd9UUGez6L9QVXQ0dfx/IVgG50lpwVI0OVOYbY3A7VAIg2R
SRKrrNyqAH7YS+miYhuP2ru+5BzWSFse92DTzPKEkmc+WwZqWjyNkkL427ZaW1Go
SChZHBEO3/RNyd37dHypjmneIe0ii8Cdy5/CgDCu9bLKch+m0XFZ+Rb3iQqqQ/z3
kNQda9m5zyymlKANjUtC/QBj0EYln+fs4nX8T6B7yT6mjMEMSsfBdwFd9pWDpLQk
b5MLmQJWyLtY+FaomZHTYdfAQStjpaSqPF+YWNAukM/Drs+280QVjuiQbDQ9HQ7G
krnuBM74RqeUWP5CGoZ7HM9ajJUW3RoZn9JSHWIv9PnBbNaciZutuTo+g/1iJV50
sKvvUJcq9B0YCQOiwn4Vawj4NX2qDm2R4Db8n2NVdYlxsoBZVM55KjbGczPP4SE3
AW2q+Aagvgdf4BDuu3dK67FAQHKm444AZ/6CVzIZUWubg2yQx08Yddq9FD3CZ9mC
9M/2MjzAvqJ+fqSn/8MFXBCdj3wI+9MrMmXUbXkjAb4WdIHzIDa4Dkq12+LWPmuC
NzJfTe/FiNliynrLh2PSoVdwjGvXCKpRugFyws9tvCK32KyO1lPk4fsUbo0Si8Wo
6GWO6nRKaJYrU9vKU/tdAadk028mFDROZBrIr3kn5wrDL3lOjFi/dZ/vTf23LPCB
8zifFRkC9r/qj290I54T22SAkFuaTJVbdTpVYVXbXgHzDYsZV7kV24SCIPLMoeO/
qYXAVVhe31eZ5FScT2sGUbi2vBq7MGEziz8xf4OlQsSYIhQ+okr25mpigxlSmbvc
eX3H1NDyHkYnt6CJpbviLknkoRDzADh4j/V5Rubju6ho5mnRrN7q2p/N+4k+F6zF
fPUdp/lc4ueoqH/ZPKIsOrQxZRPyXvW0pvcM275qekAMmta/ZT54ycGVfY6n5VG9
zetyt6vhHPUNsCKzj8pFu/s9g4eyLMdWeVi2Gem2gexOwnjJn8jSEUf8c/gtfncN
rRLJca37e8Zo0M1BNg1iw/xCZRUMj42aG8eJUFun5t2GAPHZVkGi/vl4YKXRIMIq
BUe4PxC1N4vRt/VSwKN1IoCv0/cnk0Nn1zrKPO5ZJoxp/lgtcOeX1Zq6DgRce0WZ
YIJbfJLTaNaciTclOrzcP9Jp7QWOaj3MVkTMfOgEOIHRheGIDgdjFViC+hJt0AZX
RXH2Kj9Bc6b8MPUF8TXC40KrX9cL1BPhUKDfGXmF3gZ1HnuqE0gmDKKEJ2XMv+H0
HYQj2+marO1lvFY7rOky+1N8s9yRdVRly7I410JW41MlSpHiey+eluWPqb6LKvl/
oyecbTXdfIPngnVBUOUJGPt8FcwOXadcuAVRAcY3TQ2hMieEqxYCQhXXgCGFYze0
QrECkMLD2kKDTa5QfcOIU8aVHK+Dz7z5Hvidhvv5MWtkkJyeEn3mgVoMx5F/uSk9
pIHJ2W1eNC+/RoiEXyjqS7gTFq0t/A9ZCpUrhEU+RBTtZkEgh0UF26ggIM+ybq+y
60oyy80wWVPwZR2/P+jd0KVKK3SB82mWYR+wOf6qJ7Hiu1Nql5qxs+6wvfmbIvlr
POwO1ORK7Oe8u8mijnr/+4+olWNkzoUDzIHcCM9uiQGNZQKqvfx3rYGtLHDkdCPn
yYRc5g7UapZR+1S2pU8cbVf7HsAlU3iWqwq0cVENgq4hr6CrP/vsx8y9CHhxTObq
aYYdPfw2nPvanYJGxQfnut3eLYwkx1hek5mtW7gb16rNpCD66P6Cs2l14CEm9SC/
qxMaLpakAWIInVVLwIrshUhtVNnvfAnjNr1WRAFt1GsVCSh7quRyrh39rbC8cwPW
lUmc922Q6NU9ff89jQHMne5pVgq6Nl8PYzvc4i9WkLIWdD/wCmshD122u76D3zaT
V8dxCpm3PvJukUjvITLwulF+UYRxLKp9u2bOrckLpzxeZ0Gqy28U2Qi3mck8CZft
+0T9JubX7TnCYcsI9gQjsF/jWh5syGVD5m5RgKBfpHVqThAkxu6ES91S6smdcfNg
C0oTiubOhfWkL7rHDtR8lnOpruBzjCTX3z/QjJj3+0MMQ+iKhTBrtAvznj5/g/rl
sP9VspIOZHOIK9/u0vKs9Wp5eBLOQbligxUAcnD7rjnKBuu/DC8XA+sBCaxM3rkd
Vb6jplg4PJrjy2t0ZgPMeShc6/h6k02zrF059d/mROpRvVAyu0SLvFK28bDuyg3P
fpV8tm5mtjVtHTTvBfEzv+Z+S++UjiNGixq8y7+DH1eP6hTwnjal9xjuOpOeDMwk
wdsC4Wd7Z+HEmmlnqdX/HOX3zO7RH5M2Xg3p8/X0Pw8eectmMscrtOjfM7IcUKdI
lHat9agcD/lC9q07nIewQ5BV5KS1dUXptMHGdVYuE1XTw9giEAHxL1p4X6UD2PXX
gZ2jQdzILXUf69n0yysT6t1fRpRD4V7auRiYDETFvNotZG0jrjoV4Vofq8wuoMyn
iCpcEEH57Dlh19J7C5lYYD75DYqo/kFC8V2Xm5nLkuKUNsixEY1WHKg0G356Bxep
+Uagzo0re3ZS8ldKi7guLkIAjJtunBlaIiob2mkc44YpeyTAnV8so12itwErdALh
0fz3+W1Z2hpBcFB3ujJ+ZNcTy9Sv9gi0MPLzB9TSYx3C+Rcte4vT1R0y3hXLF2sO
ZnLW4UKzdvKAx50UQqMCXngDA4KiR/RdhrV2jr/WrGuOhbH0vOcTFckoTHzx6igG
0qRj6vQHHhuNMdi5zgMmI1bCqzKtifeqPRe0yIrLgPs8gIKlfrJLuT8skpBMx+Fy
m07L/X/DClpmhoLAYjnnK7BuKxSyzpFS8Jnv5n6+XgLDF5DJWnvsUlfvqVX3Zg5J
ugRYeyx0EzkhwPLGLhU1QAU9ALt5D0UvZgUhSWwKY7q/uOAsVP/bUrpK/bR0Jtyx
lO6oC4csdvOC6/P94JffsEsb/Ap6Zr+mSHNNFRjAM5ULCGRQnpvjk4k5Vni9Emat
pRdinfDUPzQOtW7EGdXlA9ObfSmcMm2d6F46PYPThe5vkadQA4hYKNMDK550OiA+
+5s/0utTME5iQSr+ykVSiUipC4WVIjF/QxejSYgxZfj1AQ/jlZd1xsoUKtRTf565
eRtUCimADDvQAVPBez//V92xuUMSB3hT9DLkR1d2q2yleSqOiz1EPB8RGfrkw/vw
Zz80gApdfTO3WY+idYTyJrd8b24coeYZiOu1YgGbkISZnnWRRcj3thozljBezBAu
5ropmVSAOxNZHt+zwuyDHoCHiixV5aP9uA7w/47JQ0Mg0I3fxrOC840kkmARW22H
d6X2Sjv3jQ+kddeMJVW7+CiTqBR/7sjNV+Ny6R3zz56fgmDcZALtj+pnzkwXZd/7
B5PSfQQFoIuTqzreLV/a4ktr4/+J2GLH7MyZk4SYVnGCu78HE5amvrYvuKpoiBH1
3JK4Vjei0Zce4y2Wl9zzFPxATaKCYzu040Ztsgcn7BDFQy2mRt2x7VC+SLtbefvv
unAVKxhYA475fEq4tnvKl55JHEKkNzNnk65f+TvPETLVU/4rzs2aWxhYD3zLMQah
AD7VCj2ATXMTGwHwOrNtsmEkrJi8a7gz2suUhmLuKzVbDK6//dNjUezJTuhfb+5Z
jbSoIevhO28+6zxTdeEwkT6vGt2+waec6Tg9ybJIsOGoFDXyhmuqT5Y1BS1n+QXp
o4AeoVladA9oyo6hesQvXvvMAEllqjD+GpIe98yMF13g7Jg//FcjkPsWOMNq/Vve
Yegiw0/fJYKaQ9IzxepYsfgW45/LmfbsOELNCjvmsqfDW09QHDPUyEH5UiUTfXi0
kg2IsvFRYBvRHW3VHj/n46+nr/Ocsqd5oEvaBLwahA572V0XBuV1tTJHFpyTPM0D
06+6+QYo6Ajoal39XrLfRMdZxzgAwJGAHjpZgWNFBy+GKI5VaQsh2A/1Jod8pPCQ
02h81BLFJ+sTvB+jiainpNkNm7pKAQptJJ8sQRYpudPL/TCpI0nXbcZmOzKA7Kkn
HV/eRgHSBcjMUlT7esCSa0UaPR8Z19arJ6TsqBMaNpt0uY9h31iv5WZ4540Z6mrU
XhmsOMUFDSK/NbfRuYYLZi+RuvlWJ5zlpua9q8vRI80NSjhE2bUZ9e4OMomd2rdt
Qt5QhQBmPjWlN3+ujYMS8DdCE5mRvtp649JJQo0U493Z5Ny/hxuR25r8GaE+skiC
NfteHOeU+8t8eawrimU5DOfRSu8vMQr8bd3907GuiMcVlvMz/52nV6bUvSjItPXQ
7XE1fpdvwGR+R+P2G2H10qZCJM1OE3u0jhTmb+t2fSBRIwFOOQT+z+2ofBnZpFt2
9ptcLm+uFTdrB9gV2ZolfxPfxlVTxP9HhXr/SQip36nY4hgqwUV9uC7U19PCZ5XZ
SkF/23JXcJt9Zwu8ckJK9H6fjsp5Fzioqj4C8+o4/qneo7J29w9Lhfrfa2ULEcSM
rrQ3me8Xy9zHs4lmjFvlnWYejyHIf64vAy1VbHLqrYQlEetj5TZfZ0ymhqgfIX9h
2VeI6GAU70MjAd7Zjc3dCU24J+ZPD3t8ZUy/nO5GSJ8aGqSAHL6iQzh4as18YHYN
WnOnIqSIxOLE9oEXKoWh2RyIOKA2La3roCzPK3Gsmnfv8RgCwiwdwHGj25zvZvnx
jOVWVkBuMcr4ZhrhKS8UmwVpFdhdpcqPXIm36EJuBVTucMt9RRFYnerJb9k2K/XR
zIIIDxKdotwnIOJDJwlyfHdrjEjX436jv6rtFZQImNtoASOXly/yTUdlK4XytjF6
Ec5LtRvWXBZwbdfPqkHFjDAfsruU8f/o7P0YBredZ5SRcSluISEw7E+Z/oWrC9dH
RMT06UC8NQi2zI8Dyk1rOiQLYmHakUy/gbyzlxhLv23VPDKXh4RRomb/R9vEZ5Uo
6MKs2kKW+fMdNznCAtrzy6vosMZ7E7ppt/HHGzCg9ko9z4EAha7p7nU9Z860QU0R
/uHbfLIqLCnqNyob+uGpHLwlbh691DayE08N1oWfMNNlpHUXtnJK4Dzpn6b/lRoD
gacSN+tzzICuraQYw1jMWzq+xp2Grryl0sPdaKPn8QjdRxn2aEfPJMfazvLxtcVE
jonN8l9RNBRDVlCsfxNGueKDnPp6uvOB6kehBT5jn4yjZ4dCdhC8QvnZQvbA1sQr
2srOgHIhzviIzUlnyrhwaTWt+cPkQjRcvRlWVzzJqwmWDer0n43AOfISbYJODHc5
JV+COJOYH/cf8mcbMVYsju5SLlyBJ2rywpctKYDWK88ZGElqyUkm7I7/HRveY9t9
ZjBCg2go/LTV6g6gAHEsvi2+HdMKzU7tl5zAgMwIXpFYkzP+IURHK8bhfTRd7zSW
Ett+AJrDx0lFm+JW7iPqYR5Q5wnsFvV/UliFihvCYmbVCtiuV44xJaE104giHh8H
1UZSnPVs5dGIZ+y/APS0nALQWqSv7U/ME9tX2EMbGA7phLE31BdwkWZXS/mbCOpl
sOcKwkZU5q/OfKjRVE3kurezsTtnK91fMHUarQf9Uav6mh4q4ZocHLwI3DZyTgI9
ut42dNeNZvwiD70aXIVapXdI/K/wF5t/jKCWYYslFWVSfraE7xb13JH7Vc0+lF/a
EZ84Lt5qhzpmFEps/5H2lfbbzgY9/8jKBhPwy9vhNXzKTqLLfrqspj0I9XaVw06C
qeRBmfHxE/I0LdVFSIoMX4F7Z73LH+qjC0Hg76hff8TOu8vjVdQ+qDiJjYRjsy5u
2rVI+WRwwMgjlnEGGoySA5ImYmbLd5f/ZQM+LVIaysbxWKfc3snx4H6ffOw6FXug
OI/wyBvt/DnCsU6Ne1eXvx3uvNeQDlR45Xt7ZQ6Fo/hXXZgRNKJsW6VQO11MqgR/
g4xomV4BsWO988AJNdYoJ+qw0FXqGPTgnUyBj7oNFB0MEJ+TvGuTqxmx6hBMvPlm
cH76wVM8XEt5eLewFbb61Y754pnq1WXJ4JkiNapK/Y79x99SW2vqjDEM0L0Fyvoj
dEos3NiC9GXtj3uqL0bAaKEBKB1i23RP4kmEk6qpjR+CiJVBiSRZFn5xWsq94du7
eShDT1SmJovigiVBXrfutzBvXcUzPXqUQA/a2pBPDaC6B+PMvzWGuiZPO3/pd+3Y
FtF+0hfgLQsIBg1m0jLjqDQh3kTilrElH/KNnylETyBfhkzCGxAQgcAS1J/DXeL7
e/3Qak1DfMbmd2bQiTubBeAA6WbzdaHjWUF+1uTWhpg3/Upnix3ZAQUTMkrNJIkT
CdsmTclkRl4oMpW65kTfpMb1PpH8RpA+dhC2cSzrbI9KkTvzercrWovWzQjo4vNi
YsUK45AFtwgQNnTODeMZ7HoDAvGh8l9Q7fQTFQIowBYeBM1Vm+s+3HjLlSvAVoPx
amIWIzYvLxY05c0OcwgzjO8L/+WpX4rxRNBWu7yA964j3iq6kAyNiDffN6twmRDn
yCJDu4ZoO2xXkDFCNm5yUWcdVIYTDFT5WhEYUByZsM5ue4MzrrWU81+9wH42h/bB
NKX3MnB0zSATCSyzGnYrk0BhPQ+3/it1wZVrp4VC6j9dvXWueaJCqxFdQwBjG58/
iLohdq/hgEKlxguwtkG0H37gWKtVutOyHR5VX4aMWFsOMTxtiGCMe0XiyqKfehAy
nycxZRksA4caYfrGH+D4xxpKzjgRsuQsex/lS7Rzj63OwA4oCsiFuRkv6OM3gI3g
5UJ3CEVsvaulVZtPfDf9yhaxfNROBN464y19kxWeCAkTPPSZjwTco8edCG0fQKVJ
6SCstMIyaVvXgCYpzxana2GyJrbTLi66YXD3mlMo3skKfsARaNDMn2et+x+2a5lT
sUOGA4ioqKHWl6riUeKJgapnqxNUI1Wc7My4B7R7wfKbnJSj9KjoaO9qQmwKfwcF
hoCRKWKOIo16TADBRK0oHG83Vy/FfNNf6TZ8Aj5RitIw4ArXCKTt2t+W69IS6gtH
8vyAG8PW4sxTepADlclifzh52dRjc2MvragfUQhMvrqOzpC5wp6dPfpDTH8AeijY
0iKzyE4U8xYX4zTdeDUGciJk9o6CI3Uz5Uh2U2jhCxxtPZvL3gFAiIvo20LdcCYD
hdmQdelVaj3ia9m6RSVCYi63v8GRr4MvsGBiZsjCldxTV0t+D6Kzx7rTXpGge5TB
tQuxRxsbVkFvsguBGbL1pP4bWZ0GRWDoqq2rl/cgJTy1pWyojSbPH2tMPrrAxm3/
UGBj1vYWja8N8TLDn7SL/mHMcNlJ75ORyhfK5FRYFQL+tVuK4zDcPgS3PZ9GukKM
X6Pe3vuCx2XcwOrtu0xOkGt8nZZ/Y16yiFFcvdiJA539otL5EWM+6VE++DjPN4RM
nY68FIac4c6F8b21kMuet8uQ8o7bC7B6Gx3kNAmc/eGbo/Zw5wPMTIYbg3MTOmWk
yt3a+RqilAHGYuwNhEwzpUANS2MpbAvbOPPZdYvKm0KDm6/CjCxebjO32yW5uNiD
NX8GXagBzJSUUtoKk/6twASjkz+wICParxg+yVio5lxWjmLLIYPpY0gzl095CJ4V
H/dc+joN7PYtz4PJ+E/8prCl8in9636c4DQET5wU5f6wAoauL0XXNT0I/rmQKgn7
MLwuKfX+ZFY0bgwQpVGJFJd4jmrjpfaJFpTha4mdR0Pa1xvh0NNpE7huZgM9rhxx
Us9EEj/MWPfgmrOi170Jb8lL/2XMQLYX0QYRIA82owtqmxmYvzhqxWXQHDMFzFli
bb3k3NSLLUgxEB2QmToosuWsfTHaQ/ieczzrCifFzja/0QO6nFCHiJQkagSKTajK
eElKHc8cfapm3h61fIOmY1Q8qDNFlPK9bpsoVkgdGg3pO5fCrssz5usoGIrU+t1q
iSmVIId6dsXBVVOwlvjk9JHk/4jexJliQMvmuSbl+rtXrkh6V2RpNUdHA0QuJR+g
wAMGtwPkIWAG0RMN0iOjsDpFgo42Ng7jLOnDf0g6ZYHvhCnCHyfqikBFWmFh30pA
UOPRNBoZ/WrWQzuvLeBSj5f1N337Brzu5RYAI0fNQq14b/iIgWcjfvub1haPkAWD
+WgqhCfuE6Q+LOCkmdrH2bzzCGKT6BTu+soy4BXIdA/t8Ll/3K+U8PwMXse44VKE
1onDdSRc0w18MMMxvMfwib0ynKftggtuqOBJwDpj6AE0dLJZFbQ5kbs0kBcI3/Aa
/kqWMJ1ll9DazH4uGX+YuOHAWl3J5nOkC//O6Tq2xGzjHzFGOAC/X/nShwYSpG7E
RsRS69CowNk6an3P3Ifp06qLdsl1mWOcoHAdu8g+iu1yIlEy8bkEdhhGRxhMoWK8
kJCZEfW3AKzs8zSbwUalu9SrXo6Ea8FOO62/YXymLhDMBmMNZ+gAfzJ3iQFNPovH
xY/s1zwi4acoZlUZeB/TofzhqlqEOV1E6tkmTzWPyOZz/yKa9ITXH/z3SpcM3Kst
oqQy6Smqq2O5jmKOwp2/aefHMG1Hndh8YzblwVGYT+WQOqv5uKgosP1ZN55ox970
2MaYYGETrHspOFf1dDVVqY2w3o0FciABgHFF3Q9xGjRx0v12iR+IxIjGuNJ+qr48
fxXFpez8at3Gq2EI/EVhZLRx3lkiBW+iFkJUlLOuhVhvj97QR9Ot/GsIn3jIsd8+
c9G2Tow2QZjGEsx09BVDHYLXzpnGXv+ctNyUyXQhXPVfzVaCRcMscGlVTPvNbd4s
IdxXVA+fVrgJPtnzdcrDBEC4EUm33oQFgV4SVZ3F+6Ai0i6ZzzLVSikOapd3Xe9r
P+bUTy+mZexJGPr7n0nRI9ttA5F0eWUjr3UCAADZr07rTC3cU7JKLagdiWuSCyJ5
nR455ulbIxkYQZvmIS6fJLvF2NLBnYjTKN2eAWhX8WELMP7y5+LrmYVXtnBJWo/R
76Pdrpuh+wvHIzshM5OXsOcR1Hy+CKRYwfrZ+kcffWa7+wn5HUNSxdjW2qtB4s0I
mU422FdR0jOy9UfcO6i1wPInRexSeip7LWWlYWG3UcTlbCkyqZiKTs1MDr1BGJlQ
4+dLDyR/uXPwhNTf3sDiJrOuZVFlpwErHmM2QkmCi/6h8nmDVriJNNnnP4ehHp9B
9B+5RwIk0dObOfrIFSdVbdNiQ6sPD1Urm+aKFhaTY9KozM6ZT/MLuTJU9+/3AFlz
tulhh4Q+NDztA6Ccw0n4M7l+vf4tnDBo+oRKYYfDg6yhswPNtGojI6579Th+Oq2L
3GAMC7fOi0iCzBzIgYJSXcpPGLE6pfnb4I8YC4O7RrZBixMhT86s+TyZb5jSNhCM
VNl03sBwNs4rtc0/FUun8t6MRqqYEbchsvjmtax2S0Md/GEbM80CV1UfwpHQb6IU
+Sx1+jkeKVMzB2sGD7xE4sq3mj8Gtv9ETvNGW0XdxSJq1cxyeQ9WVuOUqm/MUvDt
Y5qF4LEC2jwpzzpTT2KUsiPmm1b6TwWYyLpX+k04gGTMOdZ6IVZOgOGr/N3QGQk6
qLWZv2k5DmH0uy0zfF4A189wOYBGbvGD1SxFsBv4F4NrdBIy6JYZXWk8xe5oDjHd
dePYJQ689h1O2uzY+Dwdkwwo8V2RvZZyyHNL4kI/ehBAuZbD0vgn3GBMB+VkoQK4
p+dkgq/CR7I4aNHQgbqwTTpvb7T02NoJqLydnk0GL9eTVtDHcmSUTaZl5i/MevF8
8w33rwXPt2gDir81v/qd8HR+bUPPHtuWmdxuooXLOLmQJf7ZOKdRsVnKLlZOVNTC
RiYZx6G8JsHo8vxuBqVm/C4dk9+jusN9INNYl91/o+mqnoWBG79HgyDlr2ELIqzB
17Ld/VuDbp2QelSj0wOO6nyjadFmmpr8YuPX3pVWdgDKYRgtAaQyAxnmdlhidnbC
3J4e+T/LXi1kLo2En3RG3Pi3eRObvAYh4xqF4TofFIqpLkwDbv2tROSooryJmNiG
bTBUF2MgfEhvOA2Yn0E2cFUqChmIB+nFlgFk2e69azlxFyiq1u0rfRMPsTOZ9q8A
1TTLtDzMoElRU+iyuLG1gdOzf6nT587F4jmQaNyoSXUqzUFTl3HoXGXJgTYM/yUV
ubacazb+/7OwMPS0UTXyiPTioaLM1Lq812zPA9NRB9WWXvVaM/hF/BVLX5SJD6oU
+AYm2CXKArVwYzI7cWaDBzajvrcPyuc9smOM5A8BJ806ktv3bqur6hIycsXleNNG
l6FpKbusMNALJZ7YffC7hW1punxW/Js4zBCd/TAi9pgm7+gN/B2jcvP1H01dMIPN
k09ycQcs5LNBRLg138bGwqs5Fzug4JK6daEv8T4GwNZTd7vOFa1fcwKy9s9oey/k
6BH1JJLqrQPdFCsN0olHJ60WHapnyOz08XeOu3gPyRJafvqOZ7/nnxOxrkqzPNuh
ecdugeJUuH7hdnfpo6kT1PtMwuE84I/vScSb4dCwklEqqixGgjB6hSdCx07YTJ1n
a22Fd57lnmx/LCyFVngerdP3Nj4a0CWr8s9i+5/IV1hxMf+/rhTQsjt5fxuHrBf0
8pJ7r0P8dZPAko3Jm/IbzlMaLoSIUtiTq9maG1eoaQSDUJXQQ6aSl3Pnm4/gEWni
4jfckAL2sl2l2S+ImGjB5pzxEz7OiVGcUkjoZfMcWndgfnd654QUs8BDzQZ8FZA+
HrCLcVMSZdPIxHv/MNnwukxUm9vSXOf4V5KFX20fBu1Z+bQF6xrAV7n0e4o324cZ
Vr/chjnCxXRmorBRXHvPcoD9jD2YAg+IXwEGPe0rG6MnwGLW3404DMapC+dzFX2M
Y7v0jmmipxsuT27DOwHtpXzUFXBd2jE/iQF+ZrQOND0AVYXgqTYKIoqS3ouHZ3q7
X+6PFTwCDHNGY9aA5B70MYJltV2h5YskwsI0WU7R1fDOyUIlIil8yv6+0bJE+u32
+DjkEsSQAI7HZn95t7v8BGPiyR5G2MpmrmYBPAifL3qFlUHEWKLERNhZOUYXY5Zz
ZEXr0809I3lbgFPGia9Mjo76EQDFC3Y1/2yv3wXWFZDySOWLgFQU+evXnZlI3SsY
1UYDF7WYEnFUCpybVfvO3zALPwwTMgLXpBeXUmw+/4yowYJNTynv5B3jljR2rycu
MCPvRHKlMw29t0GOHRDlllHU5zol76o4fVdejDdrGGn3urL02kraYlm12jcpEnrW
3BS/2Xg1nla5E7W2k9VSMuD3pzUlgn7yy6n0CxsZxTqY+ErQlQlw/zakhLwfPShz
J+irhQSONgB0IJ6y5n/BoW0Xt/xRswlghl4YAh/9CTOJ+6GMxOT6/vhcokkzSACB
/WD9l7iYPat1c9xv3gLVS7ZRgGIYmNtLCIhslz94kSnm6m4b98/z3hsjRHY6/bx3
DuUy2GnuaqH88dH6NH56fYtn/J/haq1SDcnG9PiISYslrub/dQIZL8eIS3yZZCLq
cM1I9vBv35lUKetc/G77w2dSEYMp9PqPkrU/mjy5FHrMB8NsElurs+1w06dZeUzj
43zhnVIM7+6Ooj8XZWnbiuQGO3UNvwwjxc2UeMLrPELnAXhJQJodhHR1LSKobEUh
fAHTatKtAJOovnSNcHLyEaxolexaGbCwUTtr7H2B+3xjI9I/VgVty+DXosf7ycqW
e2X32M2cHeCAAVnfL9AzmGjfUmU4WkFHoWEoYM60x7I6kpee/WnB5XU2KZn6IMpx
ijYrFjy9iL1MgOxmhs1Ox9/czrxoMnQUDoNYRiXhEuc78GkCTdle9J0nhihHShvt
BLCP3aivsaGamAgI25lQb9+HlpDrxFn5AKKTDXNxE2q3SFBzCuDJnVlUPqH4NvCF
ZqkYAr6xMqjlzx5C6jqMq0uTFdQcgYHNdF4+cZvvg3DcZ8v/sqIMRkKO+Inb1HFw
ixhOjJu+7Pdf/zT3CLRSY3nqvtifgKgmj3DBKxfwsQXp6//0xym0TO2LC5pyfPjp
KJRnW+GCQ16t7Cde5iUTOYZeS9QxepWdTJrX270mwcXR8uy1zyZmdBvb00gv9pLi
ggQ/KSBYt4Lfs5sQlT+h9KCzmg6so2/acLF/0NHhlMCcNZL1sIRxo3YcERbvfy4p
qQTVtMttaiyeCGuZg5fnfumz+aQcTXU6de5KB1KMbnYQA4zWB5hTucsjcNESZz/b
OTrVEp1HUjgN8TRHSInq5m2nm9uED3tk6ebebAWOCDmol4MlO3c8UlEM6oZ17blo
Uc3BXt0UfPkNyz5yuyASI497ruNzA1cdfdDH+957xfTxFt+rfKco6BZZG8ebeMIk
cVdSNQmv3lbmGGl7n/PZJzN5qao6PeXn4qEnpZ0Pp2kX9/lcRGKUzFZUJb9FKLtm
eO8KCr2G2oMyVwkRQSd/5I3i01xEmtmbQSMTXHneLS2WPWiqVr5DCDrZiep1hqed
cnWJqnwu5guBXUzKixmv8Miqvxu8RF+Gkv9vPM1+cKZf8oovNGbrShAvEsRXc3Vf
93s2+54bMWqWfW1P13UoY1U2fhLUYel5mqOVe5CjY9fuK8vSCTGwWmJQzERR42sD
Er9ZkYvkAldWpJgswlgHbPS0MoYx+Siyhh0FAb1YvYLTyDoS176PbmWLGGjWuhPr
PaxNgvcOziGfe2x/36KEWosIIyJzdrFrthVJiZ4BBWIfHGlVDefWW74kud/QGNwq
PiI6MyDmDMWbqa95MAlyh0Z6CyYX295W/8OkrYE9uGKjFnwc+jcu2Qe6/tJDgaq1
4W5vuXAoQm5h3gzuoBNPGCmAxcUrovWnRVrm9240kdiJe1oZU3f2TVhZG9G0GUbI
xs+yUFTmWTkcpIsVJNFi35ubU5eA9Ye/7Qx4R8aRyZNRvDCObJ0HEOFMHvCYm0uE
7N8pChpbFm2bvx4YHz+JcGewOypRyA8A1l4fVOp44furDHc7Rqnaz5zuC/d0UhNv
+M+mejMDvyfUvP7g6wjcfVW3/UAo4UZj/dw9C9R6yXaE66AWHpYDCIkpUlH/oDuL
dLQL3IkRt3s3/EZAUgAsv5P1zRuuxwf579xhKBltY42Jmi/jSZmqv9gFHD/U+c8C
Td3JDRKbAmaf3919wkwY/S2oOtw21Jsx31LyvbmyKs1JfMVk8pDkf6HndmKepIVt
LVRifw86jVg+BCoihGSI7YN8t7OuZsonoUNIoF4riQki1SdKK3rUUhvGAmd7GpLe
JF/efAJwtfgfh8qw99jGeGGqZl99IIKRFlZ3mfWr6sfh1waIC3O8bSYmdyqhobM0
U3fz5usZS+FcTuzwRLLXZqMrzff56stDDjtZGTiTLC9//d/x850XjQ97+GvMEcEC
pibV6GusWU02TKfuQ9LZMX2BIA0qDIeBEcDVOUdhR0q6wzWk3hCI0A8NP7y+Vsus
XL6XrHEIrm5kbP9Tla7Cuj1m3zzAlRmJmNSLhp89QZJkEwVPnmLDkQR9NxKYE3Yn
C7vjdokDEbqq2nJ2Pedo31H9NK9K8n8rM5tVJgbG7Z4K/TXLUZArJSdqSwkC+mHf
aHbw4Mx5fb8fM2ht7oeNppkz9tHIt21PqB39ArffxHcnwTjYfoIivd8afxNsYXNy
DZ9PoUNLdWEg82xIKdOg7RPmcq7HWSbXdK5Fyd71VYXiTcRmRnyrqzmMYuLJBiHS
T/mocVCkqcmGnFI5ldRT5ZS9qGUpYdURsAzFCPnH4k10bjFtMSHO46dDCpBDRsZl
ZZTMjpnJA9aBH2WJjFIa9YIy+XrGEtzVimlaUpIBTFDlQLTAP5y9Iotvuudu2fgQ
nemVF+W6g8nf6gkqsVBJJ6N6FJIkQ3MgiThlR7/OLE3WO5fynSbiWJ4dFOtql79/
l4Qk+1w2IOZvZgif1P+uFVyzCYBz/eW9QkR6gepvLB4wp8yuExMrWKyhrIrQpATy
rEK/Y/CSoUhS5CXvFh27fkwkHbth/i5DsILCq4LYjNnfj31h9KpTAjeiyUh8y07X
lgbODaawp0tG4w24eNZ1Mkva43sJLWgd5/K7medIqjgKZO3DHS4igNlelKC6I/0+
DiuFRVj0j13Gggg8MrRUA7bTckrJItBEkO8lhaDjenXDJU4R9elKUb16XllOsynO
ECky7Rb/+qnhy54w747Vw+fUJoyyxHzm6FyFGs5p8D58h4ORkyzSgXgxA35+5+/F
NUHpb6hu84ik5cBoh7ygHViDmmf2lYkOsigM0sylpvXgrFOZpnGHjbGK/Ky0M8l8
D/Sis9ieMq9KU0kdA21lhmGnaGqx1uGMs9BH0JHHYSeHb17xcnWiXnEF4JnbqH9N
0Nm+gZrPi5u0ZoNi2wwbUDTlUOzlkhwLQZi6AEpacA5eSriBThvoNrydFX+4k/2r
tBn1Zo5MU+Q2OyqqUwpDJmX2ua0CV9YbpOYdbfezYbkmE9qUpYbwB++VdccKpOC5
uK9ucXeNIckVR2UrYsNWVEMHkLVtiGeqvBjyPsxqELdUqp2UJFdaRbsYm2DdO7oc
NEnYa9yFsxi+VG0pdiFyPn4y1UEm4dc1g+MsINvHswWWaAxYShOMSZvYE0UURk+O
rCGnW+WHMxNUEeEL7srl9uJLrqYLsYHMp7VDejgYppRYK47GrTPtbh0kxVEFMftE
moZRSpmqIk+23eMM1vFgp+eoKxDzzfETjVRmweKsZGVkP7kd/fk7K0wzM/VOVz5r
iwuLEnmDOOyQq5FB3P9sQxCgJNMJRNzU4deOcnmxUR0WIqmhdoy1Jffr4O4qd/VR
xwwAFFbpLq0nmiCr1KkM+bXj123T2k396xlpClV4bQHjcC2AbpZIH7leyZ49Yx2i
gWPptDupeh9EoaH/hSKW/ourvuFqiHhvE2s2XhSZPvLj9Cq7Kx0TqBhyMrwNz60q
WWSuXyaXCYzYLSeSrM9AImm21p3o7Ens4kMXFUDhRqowneM8vTVQ1XAHxqsa1ilY
FLP+sCxwG9bk29svpCQaKBTsyQNYAWhH2MVp3S2bkZ93FMf87MC8Z6zTOcs9txai
90HXQSdUyED04dXRCQEOJsB+wR7sO3fYwypyjBnPsIsPoLhHkDH9eqwXdugDQeeE
7DR13FkokG2iU1UrF6oM4ws9iSd9V73+XfNJxdn42GoXdSVpMcCTdBmo5tA8++IA
ytGzL4CPSVAg6xsXHLj4kPDMtMAUaef2h1H52eMnSlT6jUdAOEQVpPkTZ/9dPE0a
NLcoOPOujjnNd+A9hoXc4lCi9la+ePANqC00WoYpgeCWPfI1VaxgtVHQrsL29aL2
57ZKsRA3y7glFXhX02YWrYk395mkN/ZMoYDXGduJu1K1BVhTNdN5GS65UziwwQC6
Q2Eu86+e7dhEmpdbtfF1sRTdqz3GBrfcLD3OGYJN+9X/VCO5jftFajKWkqqTPBrX
Lqghr1D4vwF5i2vJHyHpXn9Vj3Da7bVzO3eLsZ5iO2UXwRANU4BaEqj6jHyWV6R8
qhhY0Q5CxVHeJHEGf9rAXoIapA0FoUdRUYE9Yvr8KdNXxDQR9hp/qOMhcvwq0jbw
8mPeZuA1wIfha5/QLRQleSRrfEaTGAOJPsm0/Iv2POcv+zDhJo8U2RpQywBX/s2w
EX7lzXQujflTuXTLmHqaYRUt/L5KIHLtz8Z0L/usI3fTtAonynesL017aRB+nbbv
KLsyjiS396BjzbQ5RX1rS1yBIeFlnBqCEfqZ9iSCS+kzCVEdM+qZ/kJOpiyM4Cu0
9hosu5/UpFwTAwPzz/6W23bta5Xm+prb8+Q7wEaMPGyp/iOTOEsH70V/P7R9z4xL
UbN0kzj3E1x7/q+Cc3Uz8LEcUje1xJUtl+Nf6KV/W+kUcJ9HhbC/0EqG+eNzTm0K
PauFDUChKJZ8EB3DGw+TFou+LyFMmQ6wUd5jSq8A6hEXdSn53CE78rvFip04BxHg
wT9zKZmNHMqc74cQ2gjXYSAKj04hhC7ux8UeVeqYtwIlmwrIZtxDY+p1q85GFsvD
BeFODp5cgNGw+fTN35ZiD7NiJ+difSmn13uxebiLE0W49N7TQiCHMzbWZmnFbx/6
aeWug6hWQPax11xaXkuLspzFj3IWHqcJfwTR7JQ66lO8Ph7PdhDz2m9wJaIx+5da
TVzYingVpuhUaEzW4mYEUjJs/qLMYCIjZGOqVH3V5yK1bjJVxL3iB58fdJySdmSH
hZdekp4gSrhRx8cNEwch1+bTV5oeMFxcQshT9defpJ7pCFvBNEdbllt3oYl/yth/
ZfA0/PPM6Kr4qhru7hHiyciICpOdh4EFoX4R9vuzRFwPsaQ70eiv2sKA+nhR/9Sl
QzTWB91m2kJn4NFymXZWXj6j7aHnbs4HFKW08o8ZBbCzvegN0zCTCcSBDQ3M4sLW
qBkunPJ2g1bIQC7U+506jTtv/+Lnp94v9zGlUrS51ePWwK/Gm3652A/e+V/vCxFx
EPLNv2jD9lsWSkFHv74knZ/WlD/6EHIr9rK8RKjq9zAmMt+K9YOv7lgEPvlH/X2Q
I35SPr82OirijRwk8QVXGOMGqiu0sgBN6Iz4yknHXvsCVnMgLtXZELqxcsicqiwf
ppY+NkJvTuMKFCiKmlnnW4F2akT/Ku10GXEzhy9v0go8y4GbaBeb9Pfneb7dSdTP
kGZGFbd0c5KfdA1HP7m5NNPpHsNXLXXMRFSzi/sQCLYkPLX9MvY9Pw89iH3JDeEl
NWzHBPbIbXeds8VGwYrTiiLAmzif3ZawQeEcHE6vd16RrojZfL4Iu1J7HbpERB3O
zn9/cDYyFQlBb9eeolsAO5aQCVTuhYTjpaaXy4/CLjICgkcLIN6lqTRRepaHaTyk
yp8Ik79zYCQelc9/el6MwXd9NayLfMGJsyLQ96pursS6y4Epp/v7RJQZUc+ZALmi
iGsULDDVWDjMn+5BiyABC1/SQkAfNSWj390BB/ySvfhP3d9t5YQoRCGrXmWNQOmq
sifaavgvoI7Db5lLI/64GiGJNy2574106EL+4VFvC2/EGd31rVh/jNYhPRteuMtQ
aunIA1J3QnJeJ7MII+7V1Kllc7zyaoDORujBIowDdrOF2ZXY1VHe7gMd7iBPONC5
DvhorFTK9s+MSkdcbXrol1+dnNSUQQP75QIOPFbhWig1bCzyh1HcqISUkOMrVcYY
+g5rI6xxkGje6L5pkLQDYqqrgtjs150KPeSKU3d3EmL2t9G77FMtwGNaunbHJGzG
tvlBGcAOwvz35fVm4eH7qHE0BEHPFPrtKm3HJ/3PSX1ag85SY2ed2v4Gy2jl1Wsy
djHVTxHzed8nune2m73DiUGAhH4w9bICBRWyOZ1OmuROnzqbEYu/OFIg68K/wO9g
Dk838D2x/pd7CPRx9Ac5DT+LntNMCs66jOuX6j2KcHBFQOC51JvC7AhV2V7Rc58G
nJYJcNQxnb6Im3HwU1M6rAAM9iAGD3PBAaDuk4fwFdbSdV3NR9c8miiibBR+jzlY
KariP5C4Fl9TEeEFhenH0pmFApDtJq779q+GHIkzZ2y96ATt9ac0kT8ac0/NF3E3
Gg/M+Nr73LhkZb253vnkkAS0FaAov9kNIpn3+Cr9UlRYAo6tfFszkyoDuW0JlaEi
eCGvSbPl221dSx4T+KjEXDNtaKQ/SrguELzQfJv8vMPUXBzpadIoNKLxFyH85P/w
tTjh63C0fAsEBWMABfH4ZcBGmfWkxEquSGAwJKzuLlzpNOiQcDlba4jkc7tkw3zk
cOZzbwGQVuey8SDZueANP1u6ZNHjU/Wgv24/WKBoEnSdEaxJ2RCRxs7OHBSZ6Dvd
SeyyrXHeARhxb74pLm5ePvmeq5Ly9Ch22ES+QEUDzudPg7ZZ9lnoiIMBJ3Qe1YJf
FqYYzlkBEe8Fb+SalhzxbfdDV8mIW0NqPPVuYJx/5wzZ2ZjcLw2Yzy4mk9ux9NRy
zG27mzYYK3pECYxiJ7YVlSH+oqwz7WSRsmhfd9Ll81LJjqBbSXmsS00gZYWlDKEP
pt6GXbBUxnsNXGIDRVsnMALQ9HLAzBD8R0rmbdlwvy5S14WCroQKkhnC6byLeQk/
iBU50MJs2Tq7Tfvoz8An99mlsTDBbw8aHVIeRouZWZeBqfjkH0ezJB+InqbTmBzy
lyA3ai5ss8rC0sC5BRL/WYD90bXY7TeABB4FaLS2gvFHLwUwt9XosLjuHtVmJTZ/
R25r2lDey8SdmGzT7UixeXarBrQFu9o7zXVr7ZfYkv/XgUrOojspRRQPcxunF4HN
5syuSZs1ItOqaMd3pjAiWbZfYjh1aLpI45a/glONbgqMZM0YtC2/Ca9nsKKIAC77
qw5Qm/4iDP3b2HrHa6L7kprGSRRbY0Pp0wwqkSZ8NN5O57TbXUMuMC+Nxw+RxfL6
DaTJ0vusXzV7bxA/fe4V9+od6bW79i3JPPLxZJTnIs2V929oZipHxi3322HUn+3E
LzaGYwk0/Ek9vcDFj2G2xpFgNPwzj4n0YVbkGfrCCMFwKFAOs00XjSxz3WNmm3dE
RqdYkWfCyXbjypS1T1npXFHHg38SJP86vAtm3S8rT8IVMb6YgW5yBRQpLcA02Fi0
kN3Kt/kwEaiusOMvpLUzzKiKlmn5VJF8eJ/NdW/qelyvlF2kyYe8zvyKRfZplzkM
sgmy0XAouoRdBOQUHIOChgH+hwtMSthoBTZGeAd6pmlx96y39qmGKI7VZRAHcBTO
4Spef0PBH5jiHTYt47BqMjM3Nm7ZUYhjlRjbfORm7n4Hcyrt015VbAe+/zP+kt8l
IUIlqPYnWm7z14ksErtZ43mF1XRm7Q09GcJ7Uf3SMEYQcgyP1Q6SEn4e/Jsb198y
2QK1ABZN3if+kXEh5hr6OmEH7Gw04IHXJmqca7cy4ys6Fz/vCN1uPjK8x2UUKSQK
eTiXJckRnTwjwLkkRLIKu+xfgcSbpodBLFqh8LbY1DY65rvQQTZFbnWV5r4bmISX
SPkxy1+fNvmznxv+uFJFVbLS1dTVh4UUIRcQ5ZqWzPePQrxhRNXG1s1TVvg2yENe
roLRy8EOqTyWM0hJtbFg0xbn1GS05AXIz49icTyJrKlC92AOt9s7TIZTXfRa2J8Y
YzHe9XjZ/0ut+w5J3K4nlJ6ExdHpZOcP7FSjNjqprq27l0LzGJeNYmveI12qzImE
OWCb0Dtl6goysguprkzisu9HrT2Byt7xHg9aP+usi0i6mty8vr/s8XX5y5kD0PPT
AscJF3N2gyIIsPq9XDUNlKmVVXyqqHpoCQMVWdoT/UfA67dBjh372AasQsc6C2jL
cPyxw4Jnc93Jc8hcV7Jch0fZvdS49m/ESaYF9FtJ6c3MEaGXOk2lE5NhjbU+i8xB
IUahMB9gj39bIJq3+DIBBJOz4iUlpGLwRUbkVVe7BiwkMOnhCTsS/WUR1hidfg78
Fvjaq75gPwAVz1eUXBq+uqU65H32eWFKxdipYd2lYHuduCNuD4KD5s+vAzIny9ne
UjGWWnx8myylSFVQVtJlYgVFpTkcxO5sYxybVl4I23tUUhImkQGuRDXNcAg31PLp
F2yLWfNMky3PdD7WJKJHpSHz4e5ScLP622y/q3jufXGccNLLqyktSLDiu1JgOKzD
+ffpCt/YfcAFJAm1yx4s/R6w2oWMp0BkjBJHUAbIIrfQ91ufg/dM2ago53dOiROo
dIZMLtPKJM7xOf3tK2+l4et3fZjeFm9E0EXR2obBJLcF+mcEjF3HVn0m/C5rqQdc
MDBXCYn5d+pJIj/og8K+3ZNSmX/kJ4VeohoBsTVoHpGH2NWBOXA0CiwKORT86VzI
k5QIt5lrQTtkZW/IzvfgWZPapr+JBPkzPcus3Qr3xo/TshsK3cs5ltaT2DJz5VgK
IBv6P2ZRzFk5t98Q6zkInMx7F+i0q/D5X6pxpmGfWSVCoeq3Et7/QhMO4PT3vYYw
grUwGG2VkjUP7NPQIFQmqSR3zwCDhwzJ+lUe4pY3HTiL+zmEzxdNWRB/xadJNAaT
LxG10z8ZVvkQCLt8TdhyPUwgzckgAp15lG6VFkppN7U0LPiHczkmI1FWlxb4YDzf
HxE42iYTj9eQXqPUBJRl+vmaOLUkVURhza/cD5Cir81PfVcL9eTIVWJZciSF3so2
deVYYmhU32ohdgooI4aZM1tzinvM0u6gc645CTvtn12iic3Fm1qvW2XnCLEon7wP
w9tu76d53mxRLn6vcK00J5IV3fnLZypp7tgmyiuLG7arh0LN87vLdPh9dyREMzHc
0FL5rPNct3YmRL95V6ENKdoCzA2d7E93HrWpy7JGVIDpyUg2bDzVHuWbCoMLyInB
rZvLlExkM5/hf0bwZeD6u/N0SHqYu1SvpP8zBio9RZnfIxJJFJobntzdwn/xNvgY
d8WrUXcWHmcI58gSsKOucSfIj322/x2d3m89AuD/hIn4jfvK1EjEFN9Ql1AdMauu
nvDJZw4Z0NZ2SrFM+h1p8ZiguT6It/KucOlyeyf/2ghyQ7Ez3B5zZKBn8D0dx/x1
eYUjS0/nw4L/+Uhe39uTho/d0ramN6go5ZL36C6oOSMqTyYxmN5ErlKtjXbQ2PkE
T43O5/1PhUbtgAzAIzgevBovArWG2fmLIG/MFuL6WWQJmjpYZvQrO1aW13XGkj5u
YEs5feo/GCGn7byO04Y04H27pxJoiWLpwmpErT685tqo6ir0wK6he0ciy3MyPfwk
gqd8GRu1h586Kewpn++mFUdVE34iHHjxWFUze7r7i8rsc7NQK0/Z1n4M2/3/Mjeq
nDDce5x0L1lyo0s3BaaoOGMJlRq88dpqVJeRhPE22/4OSydgBoKErV6iynyZD+l5
D5qVaOno0b6mod0o3kL4f+v2XvVKC1TeqorJJOhxCEJ+DVJM09M2kPyc3zF9zz46
hqeCDZkaLAaf4T+GMhNn2Z+yC701xxS7sQk7s7FGUPp2Iyg71oioyxIe6Wi7Dipg
ZEAXz7V4bHNYJ++2cRFbt0tG9v5Zyx9T8zNClWqui/TZ9jDFQ46AyTCiETjyV9ZR
tWzfrZ0wrDeEWyFG+7nlD6WSTI5fX8t8B9/30Py5yCzw+Ti3gtr87bHfyVyJJmYr
1JawsPg1tGbmnXAx21+0kDalpYR2DpAcxlxSXctKvX2j6axQma5NndNq/aJEc70o
6g6GzJiv9Oyo/oBUkc2Y/xZ8NS3oj3AMfVJrvnlyyX7D85/3MJ8HmhZxXfl88ufI
bx6MFjkbGerI0seZe8SlA34JhEOuNyq/gKLIbDLUN7vyqg5ywqksyNqH4pfbiQLl
DEerUZLyWt90A1HJDR17cbzQJsRPTOGSjowNZkJR11li+zDQR9iiryENiy6juu/X
FXoU2bLV9VvWfcZdzNU/ukF2KmiEuztSYO7m5mHujJc1xccE/vp2/GTcTM2CbL4j
g7ATYRIl/DJz+l2ZsqhBb+jjgQKoEGo3uSYQMX3LHPCPPnJ+ziTwtYKsepeQbDqv
DZWtXP+Yj+HwE7nA2VrRUBX0KKE6MkaPI49Y+hM1SKkV9CikUChZI9+R8jX2FwNp
7hNvvNN1tjdsNqGBjTQ0uqHSdJYGorAFYXsd+e53DSbcW8wQnQKWT4a76Cq4DfRV
XnWyYNt4MfS9E9ApVR+e9XcSA33nGxvY2rvbeQrxa82f8vsp4eAAoVUHAcYOrBkb
840YpsEW5gXVTeslLe5BEAFseKlhHd61DpXX1DtEwha6wwH99tnlcdg9gvj8WDc1
SWN4YoYH8Pp7ZfJCZxgmLE6B3wQaGIOHDojcuLilc1jxYtaPCvMZSCkL5hre80Iu
Gj5h4aV8xKsnRgUBpO3fofntHJhAT47lx0sOflESIE6fg7OmMeqbwnD+aW3zxJOT
jdpGBdu2XwGJE5Uu4Lm8TNS2De/eakssjfHwNCY/ORQU8/brI21HsAHzXd9OZ11d
hE+1M9MD87O4H/n1bz/dB27dp78KB6ej3UxSDOk/Cvq/xTicNIA19OhZWHFevOy3
mSAUI8pueilcTYrGev2+6cM+OIG/pnMroh02wBQfW+EitGnI4UZPuXDuHqQbn/3U
uGEf999WGTc7hG0UWQwQjoVQ7mJ/O2ac2bzwUJ5M59KI6TBA6eKg0U/qNkoXsDlp
IcqTStuFeOMDTJRLT462ydBk9uiDvrONbSpPmlJXa/FSxhjwN/SWSspVAmn0BoKa
Eo3z3WRU4XJk1w7LlP4J+VvA6+TuetjaVGT1UihGneBL7Bi5ExiI6rhw7CXgdF+5
kS2z95hQUfXJbGl8N4fKPrBOUQEXbajfkFZTCXeSAOVEEnAV/hkNHoMFPPDux763
5xWfz4AFYQy/U45zsXsQHNHx0E3lm79a7xSXq4P92WzQNWwvGSXCYpTZne7h1ik4
Ipw3o1pc64fF393KvjVqL3V3a1vacDZwWklSIz2VqGL7/wgw03Qbays3xfB6ARs9
lRMAUSCcNOobQdyYFhxXqU62xiYDjwRbQLpt+50HUn/hK82oHM5A6w36mAE/p5jM
xIGk4CdVwNkFg8h8OBDCarHOy7YcP77815PAJ8ZU2zVXVxpRPDXz3KHccAuCHisN
Sb+ZxTDHwUORJ0vGGatuRvmhr+ZBMBBu3v0lpNJPEnsGCJ08SPgsAblSH78vXF/B
nTMCbkBUeB5Fb+F/82VZjFF9LHu2qaGbSbsFosHmjXBrTYU0+hQwcqdznOJ4NOx9
CzXhLuiN0a0rglSHfrljeFggL9aouhTJQvUQaCdu+fqt4hxtW20Gr+7A17AmjtNp
d5d+QFwsdMHG6n1BPhFeKLm3fr/7Xhwva03+8Vm23t1hruVSY+2I86mpIUner+id
OJof+Am6O+W+cjYLi2TbeU+Oov42IqzPKMNkAp7nQDhl6FL024e9nAXsQl4ccn8D
QD9G1GoNrgUppT0c1YvRQzqokY9w4BO/2SyLjlCmfMCTwD0gPwX/cvZ6w+O1Z1mx
8VFhBMq7ccMK2jCs1FeqBuuepIZuOz8aQTkjgBzZkh7gqrUy/eUosiRYV4+vypvn
nLFseFq6xIAIBouXy1+Wba8Y/05On1BGqpgbmnH6uRJY1Aq78imWdF+xWshr4OfL
AZA2QTleL8zLYDE3A/uGRVaSQteCRZrUnThhBLu7+/WzFqn8RI0DEnmRqXC1Xmh3
dKPDGy1wh/igLJzCUPxTjr/krgVcidpOSmXnO5T6G+XT+XfHMLAviNuw5V3NP7V5
zrMNMuIYY6iV6jhKzuck2aHG5hf4VEKhPgrmIIXooYlW54exKqo9cH50j5r6oAge
qk8hfB6AyGngIYXmm0+DeQNLKQZQguq8azRCAk1+gYB+mNdXeS2M8qJshDINh0BX
XRP+klpkc7sp28HuByjZIGaAf+kFimivjdv7zyGNMfR+stxCTxC5XbRGlzjbWEt6
q8DPH88qexdm+0wqiDbsb7LwZ3XJpzx5Zw4fpivu6oQytg6qEoRHlsAdt5qxFdAD
3udRe+t6NL4dWek1M+/FU1iCqjmVNtMAvonR/idfJ56QcQ9YSorTxVfn52cv/rfP
2fcQX2/mNcp8V2gkCi8MWfjLlLgWiBTCNTi+qrwijC9nx4jq2vFwA+Z5q1lcqGej
potXja+eAfjWnIAx4f+tv9b0a2FIC8HLvmHRZcZNKgKx2ZsbLMPX/yGR5JS8AZ+r
ka9ORXrBIiJNlYr/nQOoS4kWHztvy2YZuYhRPQIP09bRgd5TA5lV2aYvVinHvvX/
GQh16NNVtAH35oS+LicYn01/BjgDDrLChgWjQ3Rs6XTK7HvphIjC6yGa5yfsHjkC
9CRnkLP9ewiUtN9gzmDuSxzr7yq4mzG73Dw2xWYt0ne5Ofak46DbMhchElrCbrKH
27pBnQH6xw1r0qkYf3Toh9XzZvMlMFTJkz1HzFiAMiIFSpLRBZAoT4nTiDC97iMg
FzA+01+ezfuFoFeWfn7Ji3MuZv1VU8NcrsYfxa+MNpH2SjIgh5XlFTzMx/Rot1k6
Nvrbp3eMchozcmxuw8PVmoemQ2kube7veSaXFGYH1gDepZGj0LModlj+knXhakim
DmtkmKUFWcoJxFjC1s2uGO+xyxfXPSfau5aEYe1r0MWHhLJCbZiVOYhL2XrdG0m4
VN6OvVsLZ9D/3eit7u+TrBQXlk8cJWN9xOS/PezrZU1dkZt1yGflUK8DpFWrTmUk
I38d4FJ6GFEvGnmxXb18ltp1SzuswAVRsfzGt2HOQLT39NzmV2S7kOpMea4Ztqpr
7RkN+bGvm1HByNphP5snLPHhWja7ITS4dc8agHEpT15s+nOxJEkRHRRVgwC57NSq
tkowgRi0uVkZDNOuu5N1bukbs+cSU1ObKAEQpq4Kvc1dEm8PJjSTIEo1PeGcP88i
y1fM22VWRvzJaLnl+ewoXDLFq2Saye3TQeR7aFJqKE1Jjd7Hlg/M4tawqDif1TRk
qPiT/m5c+YlUDhGtTNXXEv2gAgWXTIAnDzHL77Qc4iyJkrOh7Cle14d0scSq19qN
S/Wic4mUkSqHLCVIyhsSQam9ebcRvBVe8Ob+M0p5mTfAfshHNzO9N0YdDUEZLJrg
Xj/VGAnwzpyqKztNnOzWAdzvKCNVVI8jEi/w1Llw3gDLPn1Wsaww7TinddOGrPBC
72OwlirtXEfoGU0Hojx7RTtakDCJMdOpDYirj+ZKAYC4bpO/uDWLe4uSlt6bO1X6
CFxRsXQH1BoPZrk/GLpASmFLCrJbj5/If3oDkqRXkJ37NbyKGPJ/z55zA98VcCkU
NqaaD9OTrMNFJwRWLHHsYJ9dvC8n1LzhC6uZDPaNuwnmLKBoj/Eq0QEuOPKJeBOW
sig8ddCbR6P6G9ZxF9u/EbtjMjxfG56GBVMfmSh2vDSn2HbeXcT/Sjb+YdFurUeS
T7ejTyFecj9N8FfgrL5PQwQQaIGxgU3KWyoy+TOR1vyNfZfvz+OrGvCb2YS8WRxF
JcN7Qf2JzKNUZAvzwL+x0ukyUByOnOB1PaeXuzBNnwZ6gDCKPqMcNcsCT8H2nhRq
NlCRo4gZJyzhK0IvSr5CggSZ4JU1k/5MkiIv9tPwJZrXWm7/9T4ewi8mFp1di4Sd
4XqvAcxCcQUNcQIcaxA93BaAurzZ6ljumzCk78GJ3QJ6tYc3EmAps9xeQCA45Xrc
uuQG2QD1CG+uLgLfteU4Ipc5w8rsfVembc5EYzDX3x0XJcdPJlAq9+CiyGT+T7yd
DwwI6iyXyEzz410XrIiC2VYj5iwIrLkmIuta9MZAdO4BWUCxSNfmkJ+2ZNeTSs1Z
QgStVF2oKWf/zqoRpWenNyKLd+Er+umgPbGxCv/duxG1gS+rBk6+su8qNNI5C6d7
NpdFQbelIWIbnGCPmYLgM+viHXv2S1sTvmmZnhwijRY0/cJLeL+sFmZViOvwiml7
Sosl/Oq+t8QBlRjPGKQRDl/HGl9qZmuIJSikKOzKFXNrN0fI1CEPOYxorJQ51fq7
LVb9uQyKDOlN+VCp9MTSAaxu3AV846J/S6O3O2THmbYFdDojp+G0YxZMr6h6QZIr
r1y56k1LlPSCaV0KNvPlZ2ahWc48TbOXJptJwTkpRsN6j6wJEUrpNbZjr+BRcTwn
+SEtY+cm7lk9P4UGhrMjrGBPObFJQ2SAa8aT1pwMcX5vKz3gZc1WBSLQl129es7J
kgRwEN7CXq9zKYUjV1b/lgtBbriH7FlSqNyZqy2Mq4UWHm+XWRi4B0hvHneMMxYb
oYeV4ysBQxxCDGnTdi+FP2uk5S1Q5Y7p+CV2YnvpWWn8qn8vbYH05rRiYJq+QsZ0
iua+xjuP/XeDsJDjmXrgUihzDdQniLXhuG4KA6KvEOq7dZsMb/iY9sXws+IXgSil
3z9NMsa9PUdr8BfOBe+mkk93iKEYAbElvMs/qi5c4Olj7QwmLfTApsXnBmwAvps5
UaOlgPgzHyBkWSqVNMmw9QQvEve/BGvGkkubKg5I6zOeFT8irMwgyzwV6867UZqa
73k2DIwrN9CcaQtQKk3h2eQqSNS65gSOek++x0Ljqvq2tlnLZa0J0Eqv1jFxzW19
eW+ny6+SKhaflKLVSlcn7a0LaqvuYS2hd+Fx4Kr8qvYUI3y1ZsxLgditIAo2JMVo
jlnlWq6d8Qgwp76+RxRB01HrKfqiFQAbp0Hq39tpGP6Lv13egQRWZt8YzS9tQE/z
VwQIAujRgomIuQd/rS9pwfs21qsBG7cXaxP80JfbjlZ2cMK50em/D2XYK1jF2cCT
BrcyGIgjqp3r8zTtxYHLO9L+xvUprlzZkpx7Z8rnS3vlnwG5P42x3iT5xWZVBpu4
NuMZHS49cT8ce3rR94Gw4K9WJ9k9Ank1c6ZKSX+xpi3IM18k7Fz/wkv/Oqg6+Y4+
VOTeLA9seiyDCnFAJ28hBR18oaPz45uUZitOxq6br7eSrlSstFrPfiAfSyBQ7cn0
w9uX88k4eO4saaYrX0JCexW5dUoMipaaJhxVQ7yw9sRA5gEgkEFv/3qhg3BZIrov
TofuPMtu/hlCIJoSc+UXPRX8R/6VmC3nEeHs5VGCU7VEcncAZCdaY1TpD/IHP/aT
3hXl+Puz1Rz4wxw8INB32dCdrpfRKTMyajKrLWs6xOGhYIabmay8S/wdwB6qWiqg
tfCtctlYzRf1O8ustuB3bVKNtwBq2cpjDOsasC3P2ktEvaCmJ6egllPSfUNOrs24
BR0WlbPS3SUOiNGtbCv2JqUVqW4+9ftrzI9cnn/PX3qQZZPbBFVcQ4NhCcPJg02F
uQ69fdvYGf8XqSfPpH4c+5A+GkK7n2I9hYVQ26othf4NlFqY4WAyMBcdIq7j3qAv
VLDTS17oVlJG/cP5riq0xZtTyAUUvJwDCP6az1guSIxd+k8CUIYOp3TWooTunWNI
zJI8W34zuvQcB3SOZXxCzppLvY7OhZqYVBk4lZ+iKc92RXh9K4t3XAcJHsPYOObs
XKspZmDJMiyOL7tw/jihdZM63aVMFD7M1rF66Gkrw7d+QpQRMYUngVK5UkptSwy6
fN4d+v176LBuuUJk6f+feyDBKsfyTotc1ilR4givuxPUPzcRDRmO3nYZHsnX98PG
OnCtS3VQYkI/reFi/xIS29JV8ZfGGBZkkceJHFyPqI3HXo7lN4J5XNkdePSRIeBj
p34RjwcPAtafiQ2GaC3a7ql3evEMGzv0IqqE7Wij1hJbHj6notwDl4WM03is/NXR
YJ3XHe7CCzDQnaoUXKZt/VMn7CtszrsV7u+3pVM3rPUmjXnY1c1cCT5mZK0ZiwB8
xQDQd0IR58aaYCaXUXgg3Oy+sMKrN7tC34TvgKpN5gjoSdkCQHUWpFat6+NF5i32
AHeu444zvU7B/gfX0zGM2wcaHvjpIJ6ltBimlVL/VNGLKz0gcxCPLGkvP8/y1hUW
2D2T7BvZ8XSvJNuFlwYgYbWCr7Xgn7oLSb7YDQalsk94hQXYgXPOG2SRJbJw2PuG
LUur2KvMKx+FgGdyppAoTwroYlmbsa0uOLH/oJ5oJhy8llQqgEBtsCHXqD2aZbQm
9fOuxNrUwu5UDbZBlcrsuVZqZmxhWdUyxzKOumpFvksB7SQEn2lkpTqWq84byZOh
WSXk0pcZlabIXuvpKJMtlfRzoq2GNzHX4xy9EcgRh0UItsB3EMnpJScZC1nGW6Lv
VGYdhHvF26GhQQRWzMDeyOja6zDMZWOW9BytpJAunxHWyTL760GhZmy586wMSkNY
n9ODPvICZhYrwxqv7wlSHGPyrwc/0IidP8RVBSb5Y0ak5oOP09eseZnIGj16d7hD
DfRSc4QYRhbs3Pscj2wuHSWvCLrxV63pXxqtAhznvElr8t03Cs1M3jwVFwSaKm4s
Kn9MYUMtgnUu/AEtaBjFTohFaX8R7nngKIHj1kILgP+BhV+lFTsc1tMlGckUlR0e
C1koXD7saaOguCsBVXr2GIdYzRmZFkk0vyr6Ayodg0v2v2SEBxBwGY8CwWbXBHig
YJnrYHgXEXFlv+R9lSNlC+MxmyWd6fo4U/ZfQAUmLtnS84RGuhxH7BZdjc8OD+yN
cPWJhVqHeHDjnh/8O0Zi0auWM62lFba2+PMluFx/zUwZL2GdCNmkf9GWMd0OMeZE
1ZG+oEoXtSB1t636PawXJ/br6qV/dZdisnuwidhZJ7YCxe4eKzZvvmce33qmPmQx
Jz4rKk7/S7XKuPbu4P2jnNMhcw7/BzhPOWxZJYNtqR80ZdejtHnkvH6Ke7Xkhiu6
r/Ctg3Lzimzgu6VvrmMtjAvS+L5bqW4/YfsNNNnlxa6wDsp3wVNloWzdemypUmIA
8Fd+6C/knJTj3Ij0yrA5wbogQWDI+3B8iTQ0WDt5zMwg/ywhvHhguoc4SjzoFh7A
/CxcXJ33JIkvxbFzkTGvgun1VaAGtPLmMMZvQL2A4sKet1naCvywTy4ZVFoYobko
v+mtlgHvKHKrjUElSZGyHFiIuX6gpGXPeaGAAOQd9Oi1C/LEe1NUrj9Ae2ABnWD2
OSB9GINNWx7N+N/b4mkawn19AY2km7EIrDkhxXLgFHwDR39DzYtxe07/e4OJA7NZ
gdgelBvgc/kF402WHs+nX0SxIZXYzp5gMPu7QRS5jPyuCrrhX/Lh6n81c9lDCOAn
IAIDODbMUBAJOWFhFZwcZchQXdqTsAn4jQeTwY49SuhID6iw/I14s/ParzJtUPO+
WBOED5sTnb2rl5tO6iiKRKU79ZUhNBWvwhLeC1WWo9uruPQuc5TYpTQ/CjUljHNf
879jEkcJOXtlNUMc+I87/Phs73cve8IARWm3yrviGwXS1evUnfcaoOCZiDDY05QQ
QtwVhnClGQZAI7YZIL+mCF0+Kww05rHwl1c2Cf0FMt6QDogEgto7/QkIS9Z5m7Pa
/vbW0AZtPfaPu8dS/3NFFKH5lIRqPp/TJSrwfrfJbFR1BI1o+EwhRjtybZrG87N7
7GIJGVILIbcbxvsrioob5cHkr3MNH98gRrnvkDAuAvrW/2KloZtahjPUJb0LFos6
VMlVTa6WnItHzJAZMpXxh7FtYa3x5g3G5Qtw8Ur7DfcqWl0oy9mOr/1k3fhzEw1l
myIca+k4smxofpvpGPaDzjm4l7ubLZxKBH0T5MMAGH0IkL3yGL7lt7NLWxXOcCQf
GxF1UDHaLHXW4irLrryMvKA1JO+2XBZNx+U8Wj95sNIsw+Yw4kCmc4vtZgqZ9Y3b
vagmW/xpFmD+NTz9Hmxr5pediOh0pOzTbmZ8hJnjYVjt2VWCmIp7LrmDta0RMb1q
qzsOb5dTRK5z66xgGVG6xG9WoRi37M3Xm5P1RpPxmQ5GVvGkPgAhFG/F3BtfJqjp
svBiqFILtREAUaM7qDfKX4ZYjqC5jABj7b/8WphZArDQKC7FouLIEzMHIxm4Kh8n
TV8JCc/Jf9hHJUNPhbBMrL+oECV51t5PlbdwOD31GHty6DXNvgT+rXytrZ1qnd41
VUImDQ8hbx2n8roxKL4ZpR90NWRTlxleuzfIqd1ecHnLn1Vf6uHA6UK8nBqwXw96
lv2uIwQktdjdMzVB/o3FsdMxNl8ptEIUqAQnUtP1x9So8AE9uA6C1tY1UKpqpljE
/6xJqObsbrwMAY8wxyqt/D0GuTQu71qKOWzvP7l2n905hA+jKptv+3VKz6MnmwCO
EFBzv3G0jc1ik6l60WLRmSZ5ewTqYq6zHo8nefFLAG4JN8+1foIXuGBXb5xR9dMQ
tSWzGnt7n2eo1M4clBlJdFExSzM8fVF8YHShgls6iFtNoZwkRyGaqIIZg3Be2dSL
nnDuuu6dD6IRV19WEEKMl50MwEl4qM9P/EeLRtqIFKF2iVIulIF9HtzJnPie7ViJ
lfQlhk3yqMjAJbT0mQWXurFnAzhVvOPHQpJsbXkdJPROfyf8NXgW2lGojpizLFDT
uDvSGHkYBZG+z9XdzLKBJXP8nEeHEQ4ArUV5z21fJK3oFIpk/3DYefQhlWf6DP6I
kWAQJq7Z8Dsj5IAgRNXq/vkUhnlKU/nnBzBZaslOH9xXpsPz3n+j1USRbpJF+Y1/
cRcgn+danwjn1OYh/fdhxW0jnx9oTtJ6yoxiT0E7afC8SfcQQo5KX5hxCZh7ll8Y
pGB9RkeBb3tFzzqhtjfGyDkquAhxChENy7I7H6XydqzETyGmCHndlQClBGEhlqKc
6RzlyJgymW4yCcXUj3fsuXOPejQYoNmaEsOnguCslY6cIq2X9SQK1AWOko1zuKYb
4AwQ76zxbQnks4PW237bmgCVLu9MYPuhdhqLfR/NRDFMaU3BM7QG3p/oc+Ofzwny
/x71UgXsDiqeUgSC449XGxKMFK01/8G2PrGM+seZYP3hqrMq+unWSGtlP0uBEFML
DEHMowC/lWrd03wjSFNPI3vPIPnVs6L566L9kDmlcN+Vp6nCj0qQW0XPgTHaqc0O
8ME3/1X+jCM4EFLLCoOyg48D1qldTdgQzoA/WCmrwpENr4XE0p1pfLvsjvUY8lds
PN9pKODJf3A2AlQQDL5uYJiQGKNJQHpaqHosoCwSAA1rqkEdS2UKs/wa8iN7hPU5
Tx/9A/fC4YEu6dy4pY/PN9PPaHLE/E3/j+54dqcDc0jSAkLJmQD0QbVlg9aaJl3I
CPgwQOZFbE3WboviLNBo1xxToHx769jaMs1VkFOtBsYdIkD4dzPYpmDc7LScJR4S
oRf2CXA1lsntdMxg06v6BOh5+JysqQ75i8Vmgke3W4aM8KFBngnz+DsjS4FvNzqp
dx3TjQ9MQ1bIlJpNB/tWAXZt/XUNlAgpo2anuXCy0DIg8T6WONTqweSdxJ2ePUTy
0szUNktr9Cd3bDpa75HxSWFHcM7bHVDVlmiOf/sUXtZGpAAw4IFkwfA9od30+Gy9
EoL7rLT/UhyD/U2m9GADtvis4GdkBcS4RliCRsOokU7F44fDv299hrcqxgDOb2O2
AEqGuL/iUaFur+3ceXmtETEKUskZmwAZHqVqxTi1rIkByEMAN7B0xQ+LQTKDx0vM
ABriV8g1IY0/fyPU6DA7sllZKPqgI7y87pfOZZmPbBl8572VO4pHhbq8HZb+aA7N
t0QCbnEtRmmaUB+xXEpn9grng1ffypmH6KGSpdk8OGsRgavo8yo0LJ38Be27fvWn
L4KMCUcM0ordK4Ypc9wW3fkhVSDufyfMrUVAQCjy+1kMTtUIFqWgDBoF7ocHdyDB
Zjj9HlT3sVRkKVgpN09R7VH1v8KnXhk9lXCKBO54rrA2Z8cJn3Ad5H6u0PLCAUC1
AVCdTg2mh8EuaN9O3X35516dpNSKKxgCizvrbv4iuJq57QwWIa7SoKxWeK2nVB0x
CEGjm4ECYWRQBs1eA1GPmPPfg9V5A1hgU70YSovA6oNF+LhRV6IULxuoAoJu3l09
BqfiH3InsnPZnmfVC+UNfKxiF/kNFzgtQLtCTQf9Dj6MKmytNuaVc8t68BAJiSj5
on+CG1vCcm8SijWlYukWSttUmbi9tra8hc8Afa0fqMDvlnLHqq8RSaJf0rlmE/bG
QEPk6+qMUpNwdhYZ8G1qB+Z1Q5EHu5nx2hJQI6l/scU2Cids42Zm5lHqtB81V69/
FKbHpA1/b1VkRy7F7sgRPGDmDbluXZzwnoV5Ikl/doKb88J+EGULj+naas/P6wWM
I7lr4AT/jZkteikHADPltGIVywJSLCKqITsA6/3DwH/ytjP5s2hgfJuvcJEfOmgH
cmBg/k278hr2xUszyNq+SszGwCkmdm3huIkY3PYjWPodJURAywoNhwEcwEnOU0xH
owGCMtwnQnNNXBVeQ+0Vn8iKU4wz43mQd5Q41Z3FAYyC8fNoHk9Y3fSbw6Bsl5u4
o4P8mKSPvwj3Ku2TugUbTV042hXmkLCmjPXAPpfoBXrxeWmeJcxVnbx/zhd8rnRf
zaGSNSZvQNHpFuusG7HxBX/EocXfTnoIk/l+2omd6yTr1EQ7kLkWNi5CJcXb1dtd
NsUPPS9qR+t0LkcuEhMHrbGLRj2bLHR3fLPLmVKoGgkZSdiafl52wzZB8BB8gvcP
o4Mk+7CmU+7SnzzP+0cTu3IAQ+jC+Qia8uhbrJ8jx/xFwxY7DJet/dC3js9utmi6
UWLqZQO6G2fjMszx3YpEgsUD44Oczc4SPP57n3FgrmUroGWOEVIl7+U0sCukCnoU
/8o63TmRTVMFMrX8hURKF6OFWyl7y2rNH4kJsnXWUz1nFV/IEt94QttHxXzDP8tt
lbtyYT8dTz003DMy83eX4TbGubCSxs1/Xvy9x5EJeS6JEFhRhpra3Urj2fauMzCs
4JBRhMAI9onwLnHDmnuQ59P7EE1Z0zbQFLKGD7KMb1Z9V8kYgmEIeCE/qQ10v9jQ
jdh7I1mPCl1xf9nyYHztqcilch6PosD3Co29/8akq3m/Eg0jwDMU2eEeT8snnqrk
K/ZdVufNJRcudhi1DdLzFlUdYaZ+AeS7B85BIGv0/poXxGVdoJeXK5EaWf3XAGle
3iFD6mcBwtCDdas54qXEkTL0F5L/YtfVTFIrR4fQ9yx+e9ZMV6bcvYruEtNtKOwz
1Y/P9WNKNRS8eGOGfz6ZPP4Wy/bdVrTmhDh/oVHxGGYCi+649B42+aVsQh+/vz58
ACxZ/vkIYF/7F0/6ICYJ/Lr/GSVEeHdQSH8vVPGtOdUThME2usqrcx/G5uGiP40Z
xtMN7rh85F3KKgoMwzBDMbTJ3smJi3ELe7gCEB5AhWapDvrXKUfntzj0PXxNsC9n
9cSaUMuaudty2rgvmXLFw+6wSsVbz0fr4C/REaRLaZmTzrH7bz1KgxzgyxkWJOx7
E9RIkK43EBDx58OQvYrWjSd4mfzN3OQG66ahivA+3xx6k50mgF5hFJ6e+Hy6BJ5+
X/Ny176m/xr05CL5KYt34dSw1gi4q19ZymlcZfnfJTsf/4nKfWE8xBMsGaiLehPR
2c5N1hMXe1LVoaTkD1l5vT861bvOHGXE7j/yfP5Hpd6hh55kMy+TUqG4sFi0f2/G
l1j1MkwZrckbk0ibOXag62QN6/bmiWKJPsTJgsxvjaCiW9RHhmdflUQjwMdBv8TY
AaSKlf5oz4oyKRDQbOeQFDtm8EreatqWAE4nYcvNFmIWOpIbhLGcimEhkUvYMYyq
GNYeIRdy5Mj/OHyVcxED39k5yxeshhJCIbdozvfc2i/cYoF1R7fMWMrYvvHiJbhB
Ad/XVQo1KCOPIrE1E6QymRA39L5/8q1freztSROuytFKr+CT9evrgnnYJ8hLiuJa
r4GDSlu62hFa/36FJN2+54bhE3zcpDEny54/J02mqFnEz1rf5baBv542m96Y/3A1
NjOyv1PVSBhjaSlMfUGBqjTyPxU6PfsdG+rezHMEAyCxAIFQmeeWAhZkBJLQDBvw
KU/NItMTrRKNOg4ukzrQYPPZ3EZyDAOt5aPbSwEJoQnP+vhn7I2QfBNEK0ZUtVrl
SK801d/QmqBEjlG4kdqT3TZbi4xlkjt11//FPWtSL11BcsG+HmS4IKY2QBqXjMCj
vmYqzfBt6eUm4vcIw6ht8Zz9pVp608Xrwpc/cURyxW2F+HX1BpBw11flx378vYiL
RuTwZYi2x8+SSsiYQBphEVtKhIO3VzzNE2w7uuYH7NqssEu3FzWqj3LEd+bAFhSO
RoKKCTjeDYwXlZUfKVzqeI0Jh3DN6LqD9aW01TOE0BNJcFEVnBb1f39mjqMGMSxv
U+Y2gbBAMJAxOa/6EFP7tDrQFTp/pN3FzayiE6QRQNx/4iVKXxGoamKYTDOgQQOQ
s9jjxgdGr9DQ6hI8f3BWYRIW5fxdQCu0kMs5HkGoRJEa2JRF4f7TmnALgJJ9pjt9
BbbXL/33PSzkIHXvarA++7YmmXNCjttGQ1SdHsuFdmTBl3iZZv4dhRvrSPPCQxgw
AZfefxrept0pshdeMSqh0cq/wPpMO/dSy+AI8Q9nvOpk3AjxLmCDD/fsSaP/UTdP
OiY9ONmJizZfULWXa0cxJM3eWLwUXG5SHGBaEpeYmrUstZfdmRk/hGjbAS3tc0++
omfMP88YKCg8xZzlPObD/hFXXHBhtwXHkVAMKw7cRFkYtq/QRHaymTqAEbboBweq
OTwZlKYunpU58ch+5ltKAs9mMZOwsFOesMTObVYKquLsgrHvUFnA6iHoOet5Piwa
wFqbuh5sMmFmbeaeRlFe9DWkuFIt9ArRVG7gwADOVQM74fN6bDUJi/G+wXVB5qST
b8jX0WmJ7yuzCA2lKlZshW1eedO5p/0QwLu76YE/lAYIwPcMEqvHh8N70DbV07bB
JTD5JylJQ4yqnTJE5scwmNTj38ueGb4NNGocZB5ci4NHQzu4mEBmnSuzCw8c4IYQ
w9va2hzZxyFDLLOMk+bfN4SsmAWwP34FD7i1Zn7aFPM2tIlYw3nD7ABiOXKwexLy
tmVKRdgnj+1r4nCUySqVZn90S3oOGj7/5JmJOXrvE/ueJ6FcAHDeLuXex+d3YnX+
O3rSrrcen/MPiOtHD/JRT99Ig71UU5PUvqTnn+KguMOgSQe6xJWf9FcESBcIbb8F
5WYioI43SBasNMwzLrPFxPljE1a3iEk7vG0VcUAvMAdiNBjXKl/GyNRnZzh8hFk0
UrZq/364z9IKsiCag9fgO0l+nrnlKSklB7d77izm2UL/uL4vtHKoScy4wCzl6LbT
0OMDU8E8mNKUtnah6KLMLA9qRtQXLDPn/ulCnYxtf7l4gxjKdgtPennQ1zpPywU9
uSVWXby2tt7rwAv9wVkAyDd6sNdI56RpjxcY2AztfB1DNEiO1yQM61Y0C0zlDv8N
lNdGhblG2isH+sdphWatYuQEzt7N3TydHw6ShIYCW+2CQvzZUJoGpQjs3neQ7MGe
SDdZAUHRe7wLp7tKEn6/vYWYUKKbsjvLFR/WH9xP+P0+Ce6XQbKsQiM4nIWIzz0c
NvnhPLi7iRXbeiZw1Q+rg2IMF1Q3QxQtoeQyRqbpz/P5P9bgjplskMEFvbs2JMSI
DBKL51pVIU02tzeqypJ0Yo1CE3JaN2j0ZrrXjqTk0c9AZc8Ep1rrtg5n/kUNnqeT
1vLkM/oFTdv4rVtQquYfKTbPMBnT+IAg/5/qzBPRCNAKHJxgCOwECIqub7nmvv+L
OwiksMB2DH0qaUGJzCsxmNWvKM6XznZaaz6oJdfXn1kcdOlDcPQMYgL72FlJsLnE
fudLvboEwBz/zrpmPCoIDXNgtOZGScfCvhLjNFCTGietx5BBA38LpHlmusq0qwZZ
cK8BSaLnOfvDDKLb8e1mQb8byaH30Ct8xFUOfiAL//KuJKvqH36EP2VHUVDIkAC/
2cJihmW7Yz3KGsRI8WxLHyuShaCcpdBE4mJWPXvmqunzkiLSkqGKDdfnK926FTch
4xnMYBexasmWwU9jWrxgHNYSeib8cUZsrzC8pcn2/eIgk36ee8InfmzXRSMOTpg4
2J0ahHjMXj/3choMi+IOeGD350PKjdIRTs14XWezHd6GIGWa/hoV+iVLMGWp1jBX
oocQMdvgU+9IEyYwMS0CzeJyQBxQjqjkB74ebfrvQAU3BDhHeraEnt0A+zKvwkoi
ma6PG1kw+AnVQ0udtrx+IsBdZEVN31GS6v4qohOLuazJM/C3G/V6K9Xo+XWBgc1F
GKXdrRKVx7QYC8MnJt/IyiYcYVEEZvJELPh+GEeA8+GbZMOIrnYfIowMthvoUM0I
DitC7gcBL1B5rX+HDbC3xqb1XGwitwAF0OFKXyjifFbG3wVbYxqH36MOJStSVMqq
pwH2t/2E/DX3gx006rBN3MiuXB3lKiJ0gkzzXzznohkQAool6xtPHwZvhrCiifX2
07jSnkrlyQe/Bod7AB+Wu5gVm0Qm6fC1/sDGnX4XmkwgGAdM3Y35IzuEa6aaHLgl
ISIB4MqrBfMGLp4h6SSeVuvz+2lc5yRPDN7jh7EIJ8QH0vflBgTduD4vCab4u0nB
B3wYOqwBw5tOp4O3KS1sbJEkLui9nnO8x9GFoSJPFz8rT+VP9jErQOLzmnSYRiqU
4nyrTUNhnatzhDoB3VUsNWLgydUHeT8ayE4xhkvtZ5mYbGjyA//2Vtsq2N81W6JF
eXyIK3zOoXGP9KO3kBd9nTIJylY/ZYSHCQAhmEx+DZi8wOLDGC/hdN8domtQfWI1
5NDcLsW9dzYdpQZaGXfIRn5BbBQJXF0UrONuhfage1NlnKxhACFiWiLi5d3Q35R9
k/oQvAx6TBi5RA53dE9bjo87ik9lGXTCIvFWmku2ol/ktaLHnaeQgrUXDlfiqt8d
RN7QZFJGXxoenjUJH8Bun6umj6I9HhU2ykXewHy2NCS3EOJkDfP7KXTNPQTSLTAC
PFM1k9+MlwFzK2qrChVi2bBHtTFil+muC88rKW/Gr4O9W0whpjGTQW0uEvyUSd89
k7Rxf3Qo3n3O4iGayMOVr3oY7q7XfLRBhnuzOwYQWa8Yv3D3o3wmn9vPOfBiTVk+
K3wieDGRAslMY0D1BKbKZ53sOnRJxGiQZvRygzr/iSaG381pPIC1T89RSCusnGXC
zS8aPXdho13W2hKov6Q/6CTloiGGgnLYMzNKHAqM9WuZnU2g2IdJmnFdEDomKS2Z
KKho/28N7D35iZxVq6VOAgw7vuPGi/zwA7AdvdOjW6He6MJQoug6f0Vy79O7xpoU
GRN5q3b6qfOYDmk8jud+Wb5DZC4NH9Vf7TPnauuH0GltoJob6eBfOKWQWgyIrhIp
iJM3zwt7/VOc1i9iNbgrjzQ6HKkMx8RfJk3qvQ7KBq13D8HGTEqBLgacyjoZFH0L
V7rZI2hdINDIgG0mu0/Y3zscq1EMzd/qy9thUE03kjnL3wE20TYm1fvuVrXaqHgJ
65XvDU70efAUOe59E/TWi73thrEZZCxKfnB7J+90spLSSG45yke/ASScBjAJfAzJ
vUGbKPEIyXveJc+NIURPzlU1vu4A3UWg/A0kcfpVsri1mElq/qPbZujyh0FSb27d
0wvUJXobqkFx9LAsG2js21S4bKFmgTXJIjVnntb1JfIjvvbcOhDg8+PcD7xz5bdx
I9q0nEsVxxU3WGPLUhh64ENnwuriktoGdNfetYaRB2tGTX7Vzuc6uduYlgnyB7ac
EQLIy1rJh/I0gz5kIf0nlfrvV9lfFvCYGuH7o1Upe/WbzLvnrXmOxEjQidbqkfxt
aM6ZqsBksiPozWoiOfiJlQ4/i7VZN79XPJ1z2p2RWIG/G0T613GR5SuNB5MqEZbj
2H6/rsD1WVsdtwnzbk4xyHGkziyqX6oFRRlzaIXeyfpyCEkwvCa722hS4nbYRs5l
w/l6iKRX3oZRYW5b4AQmNDdhk11X2BjJxY97ZjPfqk1nUn61HJmAylPjw7oH/6Kw
04TE5nGFc0XI1kIWgkTFFIbg11NZo02L18a3V5lsgQuclrw1bQTNtjGpgIFKjXcS
wPU9IwqL2toOD8OZqbCfKJ2FMF1QWC6ZC2DSJa/Gwv3F4WysnVB8iZYy8giWFmfX
S+Uq3oehNHtaklmadCoCHxe8Bxjvw3HLZPKdRqFWtKB2HoeSalmbgEdsvmRjuMFC
0pDJ9fMOfoY8EmurR8VqKCEqXPOrd7o+Yuk35KxzmKAYgqTOZ5Tr5gijyeuMDRUS
0uS7HtxyQJBEgXRMUApB9gLBKoHMg9tXhE6hMc06hvNOTEHBHScocbut6VkvmDHF
U+KfTLX41vqLHS5CNDJ6B6dsIwbRZQ2l+XFlj6122rJDT/CBnPbRS6NyENQG7zpt
dJQvPDc2EEZnSeI8PohlJ0UpGWCPT1vJYz8v9RRJmtlsi3BuO0/wdU9/RRxce3xs
Wgj1etAP34SY1SeaPlHxuIE3c3Ugpve/uXUa3nUbazZi8n9FJ3VkODm1+3r5q2/M
lKTvMQWgkfFVllx7Vz9EaAatONX8vE8r0ieTqBaIVdg8ffcSKiDse7ApRH4rQSex
Tiqy3d6O1mjCrkFy19SFBbvnoj1DAVaA5ArWor7yft9W7BmwKe0mz/xPEU9RFjmr
mxBbcyw7LDcyaa8zkUNftNq2cYzinsnLgkOHInqCqZ08PevfcR6zA0W6omSuohbT
C7plplQiKufKkyAm40S7CrEHl8VPvkWOmSnZYGsJOslfjmk1BkCICABxQJBr2f5e
XIZ5JQU+YvpqOzGqePMAR8egc2oTSq7WwNLrpTl4o4cYEPfUlBDYYooVAxslpOEk
PyOKGfl9eTdE2SYJhMBXUKEH1p28uSlTQvvGYt1+CUjhWZVPatAYKJ8AcrJaln+h
Kt1UVpvdtuQwRog3DyxO0dsVXvA84zwh4SHg1MmFFMsZQ/3i5dhnL0efV2dbkpec
YcGyxze3jMzeA8EOOIhNLPGukfppH4ONiwR87SY9yZzhrX51+yiemZhSqh8eXGS5
43OsqpqLtOhuBlJ638UdGJ+07/cQSiuZ3OnfpgjCtP+lg+xHwmYjz+yEy22WgtIa
fTLweLK5tl2Wl3ljwxDtRHzKdZ5COj61k7/yQogqwE3Pu4PN6kIp0i2izuaXlEcr
8j82aPdq0wnfw3h/INFZMj67G24QW35P7/vEFpHKOdaYVLkvbKuv5X2/S0M1fRn8
vRCoSrz1hIJ8x+7nqCJv4zjyg2iToBMs1sYidvVtWYsfOsddAp7GhDYnyq4x3P9A
EiW9lfP5h7eLVcT3NhxQ91Uxf1KmcZ8uXjgark8/hY5dwUkuBkusAfOP6WcsV8NP
o5+0rcczlWPO6nP5DS1Y5ixsKRIcFV7ZsnkGRa949j4MCktSVZpIOVz69seb1k1r
29nm2f8ybmMQLa1xmHnJ/d7RdAvwdvkAtzaQcB1W1GBysKKhdUHYJJ/+8XawcyeY
0psL1N542Ln5uSDbgQ3LYvnaclffeKLRK8MwL2Bfm8WGDSU+H32JI5kHEzZjdRo9
XKoulCnhyiENY6N9j4bmFSrV3myV3QH6ippO4d2OFIJ1qFUSzhqkngRFacMGycQS
P/0XzWMz5DdPoyUJuaKMosC/3YddBB0RlrPkRCUYqod8jOPmDWDMbK6v+0ZQSGTg
RhGnAQs0x6fQEfAY+va2jqjK5TzD7ifanz/kAkPfxGMcOj7rAOltybj9FhgXh+aq
ZmzxQGCWpw0ciWPdyHlpIWZIwuOSStNL6PpTsUwdnikTXB1uiTytDPyixkgmYJ5r
VJPMaChFYRSKOFDjr5DNNhAPShzjkhFCzM1wddIOE9LkUqJBmvRwSjOdMsnbV+Cn
WCzGG7/WAKOkZlrT6LCqhr7biKzvFrbikVUht567ARLFsVHVZ3pVieiICV97lCcZ
GBmZ78H2jLgSNiWSsQIo55UT4h9q6LUujZs/rouz7Ftt/d07RqnSH8BFHTaOOikL
yHcofHTUCdYSkvxTH4hZ+HgKOX5pX99r9bc3CmyKt/Jzk7ZtTJnI59a3YMomFG72
nCFDR+Uhco6AN5GYtZiYkvUPUCxmGjoLy7LtrNPBdGYmUQG9vXfEgmbue03sD+Jm
lEMSviU4foWX4vvmMcbDzUlqRl0zcRe44BS8ouJFysgcIe/3/KuKOiuH+c2KvG8m
jxjVHs7g/HzF6++FUJrVD0FAe0aVoeQsDApwMCfTH1MKfYPPsJ3VQ3qlHtONtYjl
DYg5Czlz80lc2MD1TU43BvAKAqi4ywe2rKy4fyTetYpCxLKUV5jkL9nSIHYH2OCk
oInkwAfeYl2BOavFVxQPLyIyOkt+MpW198LiPcWv8FBJ4OqGFNFIF81i+E7AaaF5
XiVnN1HaDCSgEoyyRa4fy+z4NZc4cuuLQjtl5FwGPgb81YQBfaA4TUR6PdRrYGCd
qQLHBgKlS3WgGQmyDsnyxbWaf5n6Wqr0fzrNYhUjnm5baxYuoZxsgUHndaR8lzV6
etEHk5GTMqAM8/kHRUPXgKbuHfN14heDDX5MqY7xErIZfw9HQ1o7UGuYTHmF+Gnq
6VP2EHWT99sx90e+uya0OgSH9uGjVf1/Y4FLyYoxR4fl/m6UwDn6PMXuUvbsfDWW
doynHB9rzJEcNJFU7/PbpsIKs+qLWLVnVpLQp7/GG5uek3d1zsmFujFJhSO1VNS4
nFL2vuaT6mRR7hu/ZAYXzvJ+hbqIOK/t2xLfv4mvSokDgiOC0RUuoyi8MHvRLqSL
rLY9cNaY9GU3Os7Uogk7pLjbvbps5PVmDfSBXwZrG4jvAl3p4xg3cSav8C0/N25B
5PNwqv/fnl/Y5J0uta4P3B7oE03lqXGz7tQhNOJjEh+7tFcgXdORbV1/CNAv8EgZ
j0lPutr3XIcuBeG81Hj4NEXqV8sCqr51qHEQj08iO9CnKtKMlQfR8ahvyw60moeK
8S8h6CzdUK1P1LSF3NtO0ZNJ+ukNj9kRxHcs0w9xNY5+x8tEluIsBgcdSGtGB8ex
/L/JKjz6zF2lUnTFPE4xd+Z+ssM6mbMxhwV7HuOjgzV7eHjYrEj/udbv1NOMV8ME
+P/vS8YideqWAHBO/X+zYeyLJ3fVw4K8F/7/oiGK4Wx3t+hWL/WZnRNdocCbpgpc
NM+d8ep+lCl8noE3eZSKusnWGH9OTvTBJIRn5D+TOUmNBybazs1R/0FJcAL9hq8J
dfHhSQqhBMmyVNZtR9ZxX3fJJJ4vUwITasQnIS14Fumb96UhQrT9mFsOe+N4YClf
6s8uHen2hTya5I+XEy1oGSRHQUL0C8OqTDZv01Az+Zf97Bw1xIZ+1lH/RcsEwtpc
NI2i8u/8BIHjfCBx8PS/YQagfTmR8h+uzEpCsTjCRj/abXkm0JuK7C+W+kAm4FcQ
NF0Xs2mrDgNJYmtyXMqoraw/ndb1iS2+fNGP54LklWirmJcGgU2piHBffQs6JYsp
H2S1F/86D5OHSIYjq2BWMaD32OKwQ6//2jGd8qf2gSJKq2+Sg1asbyQhso+jm0H6
sN/yW/LHi4ykdYlAPvNTk5U/V385g19+QEDDPZUHdzOyjzOt7iz0lkqbtiMYaaec
MTucsBlIljJw02miafq6AJWx26L/mdZeMTanBcpn+EyfcP2dcTgej+9ClhQSTefA
vQ/CrBFIM1tMkEdXG7fuovqFsFgaJ5IL3vO27SbmsiVtHZMnTwx3/GUZCeasGsHq
4iYFFQa1cPN9Ora7YtItAr544RfJ3p5t+DfoDGdUAbRhP8aAblGHyFCCYDC4FmMS
uoNw3L8njFAgLPyVdioGP/6mDXZPthmJsu7ANboP6m1vHZBqQmPyr9lVnM3nYntZ
rEnTDvM9sb3t3b3Sj+UjNFP76+0/y0uf/X+BlD5N7K7C9idsassTFAFnU1aIeDwV
drJr/tyFpoSho0gGbjkLzdc/SWW+shodRUcrEhm9WXmoVpG9KfeZGSgr1SazMoHW
/C/jCNDniQxQvXOMpa4p2gra3A1Yw2NJR8dHsoKO1RzyR7Z11HdCajKTlYuvQX+l
7gWPjbSEdqpClrtjBE4YkUm/4X5TUdurSxpDU9I3naFOqbbXZtyOZEAPbm9BNdrJ
3xWtp5QhI/2P7U1LowUiZA4A4MB7x/tRXote9z5DU33ZLw7gEYSpd2wV/2aKql0V
iilIQeszNyp/12B+b6nTTe3pVu/RTXDSUPy6TBBIV/HkVftChDTuZQUWAnCiAsvb
/SCvlTR5X0lo8SbQTL3zFDAFD1qRuKlHclm8xkWGBfrr6YKdey+9KZhY+uQkcHS1
2SzoJ/YtWwcox/rf6yxqqHHGpNG71VRZlo9RHwcogOOlUPCSbxXUn5WFL8NrumO7
x9jjmJ2SAzOgU+54iDM5fXVpVu+E7QOF5UOsWL7f4/9ekEUMwh9cM2pTlt536egZ
VyNUcV5RLUaGGHKg1IJ8HdPLsiKq0ivxr/qvWknSCGw0Bw4SZIrKK1x9nHMoc+t7
A/xfxfBFbpnfU53LhF+Ph45FqiqkLljYFVEglNhP5fTFzZ6rUf4wlr2JwPp7U/II
TRizYO0Ipjbkpr6Hwlr5f1ST3rZPvBvnjqkC644RwjoTiSndMEYXEa8UjBscYUpy
x7dzC1oKRkaDVxP9bcpj9QDfywBgt3cjPWIRr6BgMqlFMgyQN+3HkSI0U7tzI7Dr
TSDMqW5b0W2WKJkoGlaYPo81izRomyNojvGAbkspa3lBaHlInaXWHX6xex44ulN1
6nwMzoXT4SBsgHqNxV8wPQR+rAMZt4C78ELnOq5o4IjGl5tPtMOq82sGvV8d2Ij5
USQHeea8nNdg69a0rTvwutxbwL8/bEaEwM3A4hQ+ZadzGYnzWysk9rSo7LsnjYGz
6uYpiLIZXcIz7yfYFoMikuroWoKbh6x1MXSf7hVH8j9FIuBlOmd6lQT84vmaAsP0
PvWkXl1UqvLDF0nlKYDV1Fl6smEgmboJm9N9CMhKvPAIZ/GsDkY3d5xE+IosHuIM
dZfX5pS+2hcrwLgj5OsED2pG+ZLWiQ5gxFSktqJAEohw4rhywky0YjANHM+i2igT
h0fKia147n2LXAwD3Ub/JR7C4lwucI9VCdE8txfCTWivCcmSPq71fFSwEDtXMHyj
AnWkVNTFtpnwfokjdHD0NFr8xfqctKwJVlUCKJHbSRwbBKx6Gmd3ufhRMweYHa3B
MOohvTS4MSANNdQGiEROVcvolB890UDZXIML36eUCt+j1ZjN9ZUAAohaWwbjgXen
vsPPFsxsffSMupGMLHQ+bf6uJ1O01reqxUfe/7YFG4JqWih2FIXFOYNORoDyypaL
Thfzc+QP1vWG8tSlqJ2pv7q2wKy4hkmzx+eyOnRUXH9eYLRxbMhjjK4RpJfkHOcA
nMc7eEoWGwx4sZCIQu6k5kxEdMm7leMgSipvCcbHuFsuA7C9nAh2GjyO/O1sWYTy
e1rTQB3FBOxETdCjVXY89QD5BU/p8asXs4yp+9gbOXFkUWLao83i7S7lZEPCcnlN
3dtvbB50ZsxJOgIzpe83jrjZY+a4NqgHYA+nz/t92H5RmBeAUQCkGyWfuGtvIIqt
O6t4yNb7w2sSzeB3LXWE+amDrVccvrtKkmOmfdz7/dbzxlYx53ev55NXeYsFMVxd
Ps/mGzblqzZiVMod5mOONMPHLEkZuy3mPA3hUD/Ad92Sm55/ZZI4Ya4HhxdCaVbe
H0NvlWtwPo+KH0/XFHbvg8KlYtyIz+JixyIXJs3Vk19kHP/UuH8HvR6s3X3ZMOhV
72BguE7sK/5KO+phNDb97IsyUzkdt39HqeHWkzfs2Ms2jdS8SMtOd0Xv2eERMOMW
DXl0VyOekjY7p9akRvOWuhG34ONyKIiFSqD+WNzHL3Nx4IXaIaGbfMAzdDe80qrG
kZ7Uqu5hdrlDnc6Ttu9CIg1KoAOJY2uMUnzlWN+IcU4W5fbqQBt+RETDRI81Ba6M
4lu9GD19h2VESwiGz4EH264pbrXOFziYVUgv/iKykkOBKTQOfkVvwg1mrUxOnMte
ooxvcCyt7B2tUlFroUSUHhFQM81jgiu2Ps6fuzGbeIRh704vil+hKsTYm737uwYT
J0gAMdeu2x0xZcoyNRAraP9an8YtFb377lhvoJjg3fVauj17yRXzCkizVOrs60ml
rttxiWwZl6RQ4V7JYnNqCExK4l7SnA4ZwxTTNyOE0cV75l1OKw3ymWpINF0+GlKt
yCoouNsU2xNp7rxne5FisIk4TvWrvMr6otFLv/59B6S09hZykbx9G0itRnmfkSms
PX3S3SrztUIcz/DkAVEmOOrrmM6X2jHjVCkqwJgH/+mcmjr1DtBmlWrvtU7FOUyN
/cdRhM/9m5Zs6jQ5Gsqt0yn3i32DGTthhWPzitZWJkE7/7YpZmZumU2d4tkLwRrf
Uo77BXHBHvMjDLt15cynUdquk7IMciV85YQ3EeGHhAKZ4XYVbieH0KJD00+fmP03
46BmrccIdY8qQ+sXRLu+1HLlSzBcaMvM7fJ4pNC4cIarKJnAUd6wFE8dEu4CXDHB
8J5L38MiQPSdBe3wH5VfqpMia15L2VL0sOPh4n2zAo6q3glTAAHYz1a4VxPzUCO6
+e9gCx0l6ytnGPJvsgLP2RHJdwOpSNeyAQvrPWPDifqAMYx9NwhvrqJnq/3YeFjU
foeWcul5+DVvzE6jbbpfJNuvVDFAT60Lry1pP/r768iU+2RJNG0jsQ11Mh1tFLji
2HF1JqmSuxyFxErzXmBt7fOhTSSP0RFJVNl4gWxH93McIreEBd0UeuBJ24wQ2x0y
Cy+auVv0PI9wHD5DiwZaq8dlY7a64tS2McAJijr67FjeTfXfGelvRWsb9mFpn/1+
ZD2sLxVZHiq3QQsk3DHD5wdEGkVeggLOHB1KzTkeBcvmpXfIaq2r5Qoyo06z8q4N
b7ZThf8lAl9olW2CWxvwFHVrY1HshfK5zkGHXcOeTU9Mc+Jvd77Ios3YXs1UH3H0
OsoNnagz2a3zL9fgwA80QUABx2cZj9JDuQT/VzwK9ZEGDhywOPdPHkU0Lcr9+QFb
gF0e/0//kp90rbJJ6jGyvuS2RZKlon2uY1VQF40GU1AvN/KNP+uOgd7yCw9KQdhi
GrvgiUk1Vt64KHHnu6CTLa+SFiJ0uc3iXdbnw5U3/n1c6rXxmQF+QFcpNv+KMMxf
ziddxkOSFA3hfof8SZOzhXC8D6vJ1+QZPzQMs397UyaWmQUvvnqdDIEY0DYU7Etx
QwwLNCKST4qrC+zfc3NGQWahwwa4wgfg9zhakT/F3zAnGuUxvQAINwRVe4H6FRt5
J8/Jhv7bt9RafZ6zbbHJIQ4Z4/RfrS/8XK9WaQEERoKv+3TjhYU8O7U27GEs+SPQ
DmTZi5JXh5b+Fxl1KtuFLFEqk9GYllp3wGzC29MGoH1iuRznH7GvSei1+tkFhXOj
23suOmiINwlL0QBgCHkUqg0mJyGDQZs+xY1GO6n0qMFkewmK6+lbRS3ITMKXDx87
4W0xnhsAedl7k9/HtYkioIS9KR5NnYsj8/ZeSI0tKAddap+TiVH+v66S3zaSSONe
53hNDLBaSGMjed6fAgI4lKlsquo3nE6QijIAOb1hsEf0+w6uDk1rMBu56EAgj27A
Bq3QdwkPAjdM+qB931GzVJZLmwHzNaNdXleLbKtPc8eRdEh/FIxAw+I/EUGHUHLN
/vUh685j6sMlWY45uMV/8wvXspCwXLKiYDQ8TYy2xjaVYU2RyfH8gvbyMU0XJYLV
meRrYwqbWhZ0V2gkxfJFWiYJzxRsGrWc/mreeA9ZKMjDF70ftvW+LQut3UuIN56V
Z08MCyQAfhs3O/sJ7+2miG3GvzduYj7nQthEfRkw0t7elfSxBgRrTCMQ3LHvRFIY
Yu9cMm8DhDh0Y99Egpt3E1qZzkGEQMgIXnbH4Nd6+tU5VgBnixpnWXfzp7FXH8pL
1iqaC4DbVFy2m4xQwPrKhqxb0frWqJBjNswkbb6penZpuB7LTluDZ2+rUEG8i0e1
x1icxO1TNDd7tCmcpselhuXQGHBgpncG4cGRPghQiLukWYYSkNyBk0pLdvqWeVVb
U8Ran4qzHvaKv3eKSa5nV0dxb+tGeVPxUOeqVR6Aa4f6LV2xLag/4TtBEDiRtrVG
x/9jICt57k+jw0plXn1GJqVN1kbauy0X8v/UwT1sbpxX2T+3VCBlFaTY/Tec8Ph4
Ne6MKrfvi17HSsgynaJKq4EVtZcDSBCPzAJIvCDRjfs+na6JsMolPorynyM0JlSl
Pi4qbaMzUIbLrrwaWbhXF5zkMbBnjH6/J7PAc4fLg9Rr8cJx+fs/BbjZ9Miu7gHO
tP4LjutWIn3QjxeKa5sSUmTuTAeBHmgzvKhzxn7dB0r5BPP6T7qwC6ZIp1ZHQCVu
j2jItcXIef8Xa1nmKHuwPkGQE4dXLi8BB53QigCwbpM7XgGfBRHPbni/l2sgT4zW
20FdR/wPpnA7eKT0/NGNznFZgBwyToSkVUQ1CMABKzXhJ0IJ2OzE3wid4AmiqLEE
1rwkjjgDqUmw50aKge4kU7YU9RYKOMxWl8ip2xydAMtZIkHE17HVqSMROQvmv22q
/CyrxBMtQYgdntzg3Mb5zt0/jvAJCnVAObh7SC24rfg6oVDQgYPo+4N0kCrirfCw
9qpuHgP92FRxXOOPJORfuZ1v9l8DH74gxkfyHsX3PQBH4LixvPuyiNqQw/yUeOeq
ooP8BWHvtyk1rHiQIVBi9SJE2QAtKLyXbw4wQc6fG//Es3hK1cSSa0IqTX3fqae4
4iqUwmIHFfeqiQMiUYlhJqeLMG/p5V3JdcpNDcaqTjTv99aacWSGFxT6Dbmo/q8C
ASoYj73cjFIhs/BvYujrBQjrxddSeIRPOsZv0oMwRmLfb/uW4DE4o6YxVVbazDJC
yE2nb6RdXP3MYWxIFWBRMkeICj0ergpmEHLR29kydO/cBHqHxA+k78jFAS022vJp
zbvtlii9MNQU8LdcQ4n0VdWB/WDNnWLA05/9mWEy9rpXgz6RkOWRO0qMcjS6T5Ed
hLna/PbjCyxdfBgmyb3iBDcQ2gVZz2KtFHOeBN6EYU4pofv6dQJrCu2MgY1g7af6
9LMmMSigIzHEBTrnBl3XG3OUNmUPmwnwYuY4sl88BigenzASH2sjWHlQnMK57bxh
/mZCNwZJRvhqkUZ35w8xY3g+q/mZbdMN+n5F4Aw+dZGHPvyMqSnD6/83qdzFynow
AIl5pOxlkmkg+TtCSZOlm8zeMxjMRJ5BUnzmZiRdbqygBAiMa4Mu68SNR3k6YFQ6
mSrnoXvhS7Ueazrss3253IhPlb5GdVXMWVk6Z3vPL5pVYOOVzZ7BLQv32/QjH2B+
ovKSUQVZPZHjjTcbtE6FKg+0hEIqwP2Dj/ov/ErKRLqkyxLiY5unY9NB7Vdj5gxe
Yq7sMJhV5Ui0oZQdFf2rs18F5LQceYBeYn+1rpNxYrBU1OjZ4kP9c6g+VrdjjcLu
FEzt5QRbZmtsiu+Z2Yu8WVjrjmIq8P9J5cijUspYOJHp/EY2AQoCk64y/R91xkvn
cf089/+jkxxI58TWE+458rdeYXb84d3hsbYN9GRZPpYr99YNeDrilXUlkAIF7Zgq
V2ZQ8FBV2Zt26YwtGsqCRLeZWidVuRP9SGOzVhjhSlqZQvdki0Uy5iXT24Uz2Js/
MHPFO9RyGFb15Dg6iAbb9DypVmgqJzEIQD4O/s+8S8OIw9YYUtlMw1uxm2L1Yfw8
X7pvB3wfFPc6VduO7yiVoSKuonSTZFZ+1hPKmOxDwPzo+8qKIOl+rlU00E/WLWg2
mDCF8RoN5A+rSEyyrchxq/SjJWLIwbR6l+HjQnxrXdGPu2gIrQehvzFxfnxttXJv
p/X5bOBu2+nWt3U3RgGK/emKkUFJYLB8EX74xBZvCBhezXb0H4LyLNoAjTfR+N15
m5RqUJn5eBY5ROR8kfJFeLAjvcyRI/6w3T0nR3hwwaLTwJdL3sRb3IeuWVbzgBeR
miCSnNZfOu9tKCxuNgWq3M19ovzoi5nIbsDoJoFsFphOCYBDKxtUD5+slT+NaFyw
Jbu+L+A2M6QDUml3MDLerwcdOXASsLiegXMzEY+y/VZkZ7CGZRYmYSBh3L4mV/mL
TgIbzY/lEKHR31qIzXnrvjK0zgBfxWG8CDhOD4Vcb6zsOkE3BoyQVMGgor3c5rQO
NgxAp8UN9wcJ81Zic0p9j0UlLTx/cFn/lZxRshBIj0GnzPwEg396DglgQao/qZ8H
NDyXYWHiOS2W1jNiA//ukhcTbz4i9KyXpQuRQaxiSeKOtTaibBQY/4CTfoX3UmI7
PhQQmgZ8rkBZZ7rX/SQ/XoM2TcYKne2nYkOOmhKQ9Q8NpagHa0OuRnsnUhlQIZKK
O4PWXPj5buuUEgK+2PjTnl3wsBrxrKcQ+8EsZvjrbPi+6tnh3edkZSVpSRUexgwu
MLJaZqg7wQRogRKFR+tST7CiCwvt8qtiqQVwPYA6d4ToN/8n7AAR2eqxJV9HmVpx
HjSp191MaSsnE8WS8DuxrKcPwzuF7oDAhq7/31BPTFD/ZaptVJweRamaNrh045zU
qsqc8xg2r7ERgyvVMZuV4dDblfJmbdjRr2SbXWR2nLkRxtFrfTwkCgTFBleP204+
hLe/VD2Se6rE+m1z2jEtvNvLcdsGq/En3NKiNvcURw4AHVMtkRldraYbubk58BYD
GacTmOYa+U0vbwAKCkPJfFmNJgeuPyZRExrvxwob1G0gd92x5xZpYm85Coi7P6ei
nMHXA6z+snBHdsd9zaG7S6e62UVj0fdDJAPoZ8iA4M44jeHXDcylyx31kGcC/XzA
qSs0X6cWOe3lz2ZNXu7F24o/+YVt2mo+79fw/JX6jIMpOVASRwPok5w2EOh+mYwk
50fCmEM4ZdzlhT/GgKYYtYNeXzrH+26jnsk3nji86Io7HttYnl47ZQhaiwwSG8QF
BuKAv4JlABB+SEhajE1yLZLaga0MbT3AaddYRx4dt4QjbGBOUnZ8oBr+XI2EDInE
VRKTLhXFo2NuB/mqNWaJZYKSJSp36dLD95+ZcnUxLIGCmA2VUg98uv0f37whbhCZ
EYRe6Q1mJpY5T8cfdk5pg27/klcUmZdvapPVsSvoG1B4CXlepWW+VKsvwAkxRiXG
Zhsa08cZ94fTErgLCzOTm13AzilzEH+IMi96r6gHGJBmrhLqE86eqX/wcJzN7c7j
NypLGQSaKrhwx2nFbnJ6in0o4B/5AgZtwtPOEHVKsXBXELwlmbSYosN8skFiXl20
ql/u+5j9JzDdwZjDTd6a5Zno0q3VZi9en2UXymsLWcs5LLIbU8a/hPHhkqoiH02N
wD5A0Vv3Y9np+UKlXjZ4GDflJxvWgh36vn2DKa88cG/v25SVMwjTeXZzsge2pIeF
Mjnm7COT8embskm3a49YBU6uN0IJE1BO3u94kjJiuwPuRQ1qCkshKh/RpwdOJ0Y+
mhL6WzhGnCMW5g9/KdP6LylXDC327xcS8kKmeDMZAw+5Dh8tyfsPMTQ9Pa/jyYAJ
R0KyfUYf0Imz+2NXDObJ+w9pZAAU+95JId2ERhi2RtA3c6jl7feeYt5YZBLYCyZi
CfZ5dUZZY9GHFGUEVAVSGrbAcE97PJQy3rX1M7Ygfv53pW065LTTRfnCKpnUIwE3
gc7To2JDJ9S1DsAJv2U95FA1WuKTYetMiJiLi7CufQvZHUmfm2YKh/g/YfViF5Fj
E1OG6b+7Jb1v0ZErwC5Z8mWvfcPm7NpDseC9CWjsdT/4A9sV30apO4jc6/tWokLQ
SI/22iOOUIeUvWUlwPZOVvQqGuhjy/p0fzjdne3S6v7joKfwkRUvlh3Y+uYaWu6q
M+1siuyoNz7b6KKky3rZ3sZdb2Z34N/P53VxyEGpF/pV+nD+Zcvz+z1JkgGFxaPA
IHQsMes4h+VCKbsw/7GkS9tyJvROq/sm9LLVvCKM3762iYQU6zm5zYhE2lTndoFR
Z6RCriBVJqrRGMcm12rkC29dZsE0w0lXnNnCRgDhEwSjuqWBotRnXg2n7IYkEjU8
Ca7TJt7A8X35Z06RJNniJREPOJLKywXXnTeJxpqwYqz69nFUn5PpuraGE/iyPw5m
HC02GSO2SnWVmryVfpDgAPzNuK2Fv1kI5cq/JKMc4Y4VoK9t4uL5PGcV33el0vdH
Cwz4gkq2bOWEZyZyr88zJccoLQc6ceAQKRh3PQqEl+0EZQ4DpK9WV+vPvGRIT8ID
eB0gNa51XmPwerAClC6F/hMMYhJG2XgJjBLHsE+LZU3RcLyB5sotIU81YbNS9zlC
lk2j+BIppHVsqI+0HlsrdKQL0w7J7Dy1dIWUwdqJYP+gwkHBERcEz2UYjeW2rUjm
473MhGFyIgT2EvwpHLrW9EllkblJrhQ9JpnucyjHkaVTpv3trL3oZVrF91d+xOp8
wAE5S8CGszKMHyBR2/Eb93q3qHt9GfN57cn3Qu/rRb2pu4FWhK8g25ts05zbKD7v
y+mZoV/JRBo8fstz+8OrErfZ1ikFSNTloq6zX3xi9gb0AShnhmwrmd4NC5NUInO6
l46sArKYecootmwC14gFup7FJHkc/EUpXvAngyJdTdAwqavQ6sZ0X3x5LgILfsO0
HUflFZsiMrh3wsq1jjlYcU4spqPVw/eo5Z5C72DMp9DhWF1h3XCPpdNCc6/HpLeq
4U+vVUv98Chc8lBAuzxQ/SeG9tftcQ223HtPKxj2wsD5wguKSo2Z6pp8iRJT7/Vd
nwd9JoJCkvjEXaqyMV7rVv/PN86HVL8CcYk1Q/lG7w705Oom2C+prEBPyhJt5ktL
loMh6MQyrIxcLaKOMQHrWxlPoYz1aHkSTCGZbO9ANfKojt5X05f82NmSy6RuBes5
b3VRV7+QtwyzIDQnH1mj0xEiv+G13+UF0nKM+PTT1XdR1o6L5Pshx5e/hcbY1m9C
yXgPZqRfWAfGhza1P9YhFF7t1cg/HMQinidkLRFLZYIaI2thaABK7rjEwva75Smk
nEaChJVonONAn3C0sLU6sPf3PxYPD0M6VnWH9UCWzhitVpGwgfQOj8i71X8322j9
G/gFqz/5OA6i/T8dBIVsbvQxxIAoZ7EEhjsWLazDsvhaQBa49Lp8tCg+8f0Ky4Sq
GZRi6Ut1RvXU0URm1bwOpsAUR8vIFrq05/2Eq7YRMQd0QwrjoAKkN43OcSo9hCuI
olJRWWjfEhBG7weuuS4X/DnYjq2bhxKgEDDzqcCVftTOcHBpu3mR2zgckkMwE6/7
Gf3Mu8BssBWNDqVyOTd3KuKIScrUqs7mSLeBIXIZAatYH4HyvBXU1vg/ft8qwP7Y
xc3cGdIIvkW11wmAL2ygMZtroAGsnIqe7fMlpdu22Y5YbnLNlZ3Agde2kMaDaDEA
tvV05RNWyfiaEajjp1PBS8R0uNfnraQ/kJeot8q5E5dO/VNocmMMdROZD9q9R38P
ksPNmE2QIatpxiJD6VEsd3sy8zD4izA+bJ1vRJNCh8B/K4xryyJaJxjHGZ8+Tj0t
R9BtS9l6TQOWbi33xEzEgegoRJKqQzCaCuGxKx8obg0/0G6/NcDETerwzFKtu8pu
8EAtaxc9onZH/0Ki3Xl1YMASHxGhmQY/ec2HXXSB5JZnOmGmOm9uOS5NhnGokhvm
GlhyYR9X5cigwtZfY09HPO4+sdH8lWDJE9A6WXUH/rz429MgQ+YISFmR8AQh9p8g
pubD3ajzIVN0bTMvZbSPfth9DwRKSshsQd3hCZF5bUbOiXFimimVYzfxPt0e2N9X
XJzGYyktW6/w9bt8fcZ0m9HDqz7CUhUAjTXxPIDHLWfuzjk9mWkOR8gGnP5w4NPy
T1iECaEGUl8D5xpDk0Jiz5dwdLPzpOhXcVxh6U/xOjits1E9jXfGU9fXSeP+wfVM
Dtt5EtQIaErIxeiXE/wIQKb7tM7sLdTao0NjAgkeCzIPDuUDe6Sh9rZFwamY4Ljk
+pJnF3ubY/I1kHbGEpHIAMLmQECCrknMReFayW++FYSNnvvxfWD76DGMNAmmVDgE
XzUAiuIURYWlyinyqYn7FgL8/GxTQ6tyscH1vltRj+pFunDsXxK+Srpxb+CzJ5Zm
T6vjdSiHIK+5+D3CUcUliIyuakkVoHrl2Wrn/rpFAR6d6Do5rm7Ltz4377yeYuMm
7tlKKDQ8qxXp/+W79g5eq+824V2zo/kgQbnnCG9+Vp2H+seixIJ0zZurh0cHHLMI
2nhXKmc8JNzyhJBkeMG2pGqtg2gje+DtJpQduwWqVf1w218m10TuJg9O8VV5scIB
j+IsDrqOWs7MWkTT3TXTnxxGG5uUtYOENcqN9oMQlemv6G6Lyw01b1l/o+lD7Ckv
VD/zumFS+iA1hlU2eJGjHzYhJpPU7cf8+dvuSJmBtzAgFsxrr3AK+PNs2sUoz3M1
3dzHfVvQoqtbGyVawPEf7i4xklOKxbwt8ckPjc3q3HS2ipqbJ/C1KFLp9gz5vAe1
oENpw2l8/f9qo1PHT6nwFaTeIiPZb9bw8Be34DUHEoaU89MBHyULUrvvaPDRA3gb
P3oRz2qoxrbjUiTbcJuAVta/0ixAcTRboMCu6r/qEhd4SmX6yxYMhpRTTSP3A/TT
QaXSa/UCQPgd/p6gw1VLP0w2PthvBhJnV15D+qHFWuOkwwqns5m8KMKrsm1Exri6
ZMF56BqO/8h0jo90+6lVdue5noEWhXjTlJWSx67h4jZCdHe0ZRFgA7AjiN0IRSb+
ldOKEZGGxtPQvXs5/ZWw8jJjl29Rh4OQrWACj3Ugi0s+bJDTNPAR9N6EnD9EluHK
xG24DfJ5cWgcwKenDVBOg8sRkgAf9ZkohKG7aI9rcLa1BgKubpV2y0NIHSd9bTfO
XNl04nnbeKCZBgcsjR7bgSYeLmMIxTWwi9zL6LBErOW7zuP7v2cLI2QggIhhSLpr
8SuI2F7E6C4s7bOPKdKRCmKqcNR2F6iyJx7yUmEJ5aycmgSd7KFVZRCR4xQnjISj
SVorAaPtaioKiqh4KGxgVZGqwYAZcnaAhizoZcCfgUxHk3VhAin2Y0hLPa/D4IG6
8ukkgN67Y8GOEyVjiwCV2phP2dSNC2eHEBQK5P7g5GeoIvrLA2wquzf4xNKcZvFk
VlHBHS7vwEssFAUg83/sEsGh1XRcoxQawqu0RyprWOdNsDkg4e1vxyFTcNqWyYnU
xlhNtOTzOyVURbW5CNjo1eemgIzarskFwi/kI0JtmNWccdQrMRQs0ah19WO8+tn9
EPYGZD78Zq6CGjmSvC1XlbzmL4KsuzYDyVH/pmWDJuYCOHX9ywOTamKryM3vOrOd
bSRXse8fMVw7qoK61foAo8XxXsIhyHdR5N+s3k673Uj8anBXc5XtvYD/9sPHZ1yj
iVjf6+5DbVTlgsLon9zC5aAyyUVg57wIi6Rg8sPKHVEVboN1DgT9VRS3kQWNOGdG
aADwBemVkVHL9+6tivphKXcs6rWN8ppvNAhVdyc9bjdQ3o5hjTPrScR6gn/DcUNr
Q12JDGRtMhk/QgAXGA4tG/Lfw/f5cXXQv045XOqVGkNmawq213APKZC1yh5cKR9D
tRCw1Xb70yX5k9Az5aV5h/9CL3t7e+5GwXt9AzKgoCDQOW6FG+qaRyMyoywaJzov
o+6xfXGg7p9oPd1fQs1bKzM9V156+aVI8jxqg5HYZNZVGCMLnahg6RcNh+tkgJxz
UyDXQxRNvn3Sf7evZb85fJ0S/3SZsEnS/hR3q/VSe6282XLU/9UNJlzgmgsVEYlf
EWlXCrDp/XjKTWEDwoYA/bxFFHvl6CjN7N2QwDcGfV2fun+JWTSSyGsDEc4evpQn
eAbm5cu4PZ4a29Ffe3fQ1BjTmKNcQv2fKMfiu/Ga6l+47DeifyuajNwI0EtNBgN+
CBBGeob9a6RS4pitcqXG4PHUBxe3U9unR+3c2vuBn8I1EFG0L+uKcrk/ouOa2I/M
SE/ZdKZVU7JdQIDP5mmbaoyPlmT4QnnEDfGwHeNmCN9HyM3LXfRaVrdnimK+6cbJ
3aeoi5ehdR4740FFOqEEUUHVnQWdEjmmvpVqvx6bw3fcfU5tAjVDm+J8VBsKH0n9
LRwk9yRbYQgl/NO2+Cl3/TwlUdywBvptOKcAE9qeW+REiwDFe2+eKDPMLLzgKaMq
p3xda5jHXYNwlFnuuzMEFLe1ifygqomd6vtiz1uMxx6Wh3aMFepftjtKHnVtSKqJ
3b15ak7tuNFwB5hCkBRfK+RThP0aeiFXF2sQ/Say/GwpspY/l5/lA2ACDIU44hlt
cbMjqNokGhd1xHiQuDbvj953Xilouw4QlTG+NLUeTo98m1zZ23Uq3SYSisKPKy3d
VRgsLRLdttiqdAbA3E7fVTz7N8z1TyrZNFrB6aygWKA8vcvk7hAkW32hgChw3iA7
1m5Hgocs7KgsjihzVj/EcMmdeNPc8XEGoEilvSRTYxXipQPs15bTBVBfR4tL8lcy
GjsTNK8n48whjfE7G00zC2o0FDwj+hcYJxV9wnt2KrEOxYfCY0+Qm0fDm4y8Z2Ke
sTIbcllaCsrCvYKdU56SGCHNXlA2gVeMzwyf0QsgQtsXFK8WLO4pcSOnWB4R8pb2
sEDBlijQA1y4UTmb6VD6OvHMKy0hJ7ekWjFVgQy3NCq1yKMgbgglH3iclLj/fAH9
f7f6C6lePSmZPFB0A7DBrvYrZRI1Hhwb2kf6DmC/4Jkh69nXNylxdh5XTExRNnKW
8mXh5zP/LfUhdfyd2JH+ii7taCC+D6F97fS6ZTW6F2EW32p8VOFJXTDjkAtU48aF
k5NoKfd8qLlHwGg0Tpq3bQV1LIDaVbWljKThfSG6snclucpund8JX6ii9pi+DBTC
vwdXAxvK6/pSnzoKsAplBvbhUhdMnjouw1Lz+Mc4blLTbLv0vhy1DVri9dDB4mP3
zYhTKavbXRFhoC5tmZ/ipB6HhD+PTbf5Yx3gLKhOmAHEQdvxBZtHqoEkKqlg72zS
tLg76chG/C7GSTSIAGCRlZDMh94DaUTMSSNUKyZjk2WvzAxY71NXW4rFObTbOeQn
TMnxIu7xn4Z9Xm62JpqyqFjp+XyVWZubKALHN7v7rMe70aKb5XcO61gFQZbU+nyZ
Awpb5oIfALCGXzn1uK4IhyFhn+c5TsWEoikbZJslQknHnDgvataEwZ4UzHCBj3IZ
qXWbG8byiCAW0JksujqJ18u5yOZ5r6pdqtTw3lNq5JPFSgX8oR+CGseX5mq9uwMr
9wRSxxvNfSv0DmTuKSGgsf4hr07JcK3jGMd8IX2YXAkRt7HAxIEygq9mW5rUZwmr
qVSBTsco8H6QiyflML/YaqGiz9lUcVOZSxNxJ3oCuAwtPiWhMtRDwqSkY+H5Jgak
ecjFJwBE2e1z6o6bVwdI3gUKSZQn7p+M7FowqBFscGt75lMs9V+9yq7AI9WeblJ1
ph2yVcgX0riT0wJyMvfb/so7jDXOTpvaT1b5RP5zxd2AdqPj6nnCNobYb5WjJaLN
vqwaGw2iO4c+HpivRHtd/WQU/7Se8HEZ8/YDFhr7WSj98UrhuOae65udjrszosmG
ktQ5ZXMMC0cT4pZezZ7W98ZTWtv7xh7p1vl5tKcZBTvmKlVM2VrvWN9ZYYRaBMA4
O5B1NkagNob4hlTxnyreh/IJT4mZRSy5KzofqAevpJlUrOe4w6jTtIXFEp2SAw71
4cIor50CnuDBeUcvvO2fAFuJiat3qKqeXfz9Oa1/KsPj2/mw89Rv+ZeZiYxzRlaG
b1LjbB5NeS9wgjT//QGTRGyUXLQItHawurEuJgEtOM5/zNgX6bSqKyXcZToShwC+
N8GBeSCAABvEC4bngetRlWg6BP/JpUitwVWTMXuTqmuFWTcZPRnkqt+TipWVV2Rp
a5PRInRrB3Ov2D8d/p7XhEf5mVuGvAit/z0ryeaJz1aQGMI/OKmU6UTEK6L+JVQj
aH00Yv3KXnHPM3UufZPGHkWMoVx+lExI7vZ1zbhg6hsUeEZqkTZF8dbTgMz0Cor6
6G7KXPMTPZJfIXGVpozzvEokRgx2RUbX+1X7tyZH4wIJ3pwhOcucfadcZC9du/1E
+KzkO6CGvuSr4c1w6xxAJcyz4ycRumG0IdrelRHh3CDsq1sC1tRIxQ7fTTE98CQG
mlZbquDhjcYtUAFJsyAIhIX/ktjKh+XoIoypRWH/maRW9jQHZRgW9CudAn+au4Je
U0Dtv2RQ61XL+y094nJ+azq7oOC+Q0HRv9g6N1H8eHONW4iZjDiTIFkWDCmPLaQZ
yq4ZLjSl2MHLflkLaK47MtOQpyOmQFveDZ0FCyXVxMIdlDs28wKgGfm1Aqw6iWTj
b3Zud2PoWWeyG1W+dpL0WdeI3hpvL8SQcoAgT06DpYcMJPnh05tehjfhn5knPVjG
Qi9FPzlJf/L6zSSb1yRZjEGgMyA+zX3fofq4YW5YNUdVeZ/k08czU0D6B4+OKrAo
7kT3pZ5N+TFuq9zAXnQFDaYjd/0ZTtKZQS6do+a18CNilTct64U6YeK/hr1QctIZ
PhCmnFWGZ/WGXGWhNaX83ruvfU06qtb8/b1riyD1s4M4Iu8c0eoJLTFnYhlWEa1B
OMvQ2CcWyd8CkYiDPoqkiqqmSBthrk/yzRzlYLRLoV0T5TFa0oW1t99HFUZ0SD9L
mSjhqQyPI+qR3Uoil+V/dXhhB0+xRFrTwmZhq9WCnazFvoXs5s8Al0Yu/1RKsqWj
dj/VsTOZnaqrNeX36rWl49b+yjQtZ4AwTHSmVFdBp5lekfNWuWKVTHHFipYg+gd5
k2KvYcUyo/L1cfJ+oNg0dCxQMmRhjYjA0JTk19I/I3iCJxNuZvKRd37mCUfWcNuk
5S9GtZnozs24GjhwqiOlGe0yE4oaNrzlmfm49Ti+T+kk3GW/2q7+8Vk7Xi7iDNgZ
83xFfk2Irle3xr68zJlmpyXv1xlHLt08fS5G9EDNyeAHRhJpOpONzmbzf5LNQ+JQ
TUtBo5lvJPQf00RBs/YaXug3HwckszmE/WeSB+02DV/UmifOQx6ehUJN58e5A1WS
Rd8MYMkBQI0PGcEvi1eS0sWmTNmuBCIPgFZJHIwnsWwI6EnJWX2+mF09g6sV3srT
UAeI44ewQDCHddSIbQHdizpU3FzaGESASY6VZsHCBOUxMxy+7ChRPdtHSgNeWIlv
3Iv9onfRBp4ZQwbwGSflgfFnVMHcPDdkdPfvWnFQ72rKUbvhSprNuYZ54raheiQM
8kXgdGiQwsz5fZAp7/6uiTMzAIkYZWkLMFt16kDIgqmmr540Sy07Vokp48MC3E1A
H6fGV1pRQBiLjGNzxCCdX9422kUpBrq4CNEzK1O6fi7mwivAC8qrN0kQsoKMum7p
Ii3K+VwBBr7CEHf+xixhwF60ykHFaS6NjVN1dolPgXUG463es3XaB++Sl5ktqqBS
HhAeIbmRRjzjhl5nAwAYQaH/3/8VNAlndnd1xO4cfFbIT9dQjqy92PCJr+9wu0kA
0nS6d+uBGVAGYV1zPv6+d3cNIN7xJg6yqk02tuDAS5g7AeIaGL41H5Nep44TI/pS
SJbhgOOrL8cs7zmZWJTLqcjcT0xsl5R8bDkiMJWAqVkKF3pWEjsGrMmxq9aMFJ4I
4rmqrB+6IKY1utpEPT8q2kpbk9JvRIZftaCWTKgpvbnEhCUFX/JR9kZvjYvmCO5T
0Eq1AJWQXT5nIZ4jfEEQesn99qmNR+Oiaj/GVV549Z0Yhv/MFYT1IxjWY9QqtEWx
Xv77XER3rvdFm8qWslms6vd/M1M0NFL+X0ZDF3kT4Ke2Q6aI8JUFFPT0kV56MHI5
4d07/Hn/Ab6Oc3m3g+stcrKWlI5pv2mhp2Z7mtMTBwTlyCC+trmaEx9AiXI/4C9O
qgRW7aDmXC3+jAEV8EEJss2FifGv50cT/GShgoxb36jyntxQsldWnhG3+ygrdjla
mWDVaIjqgVj/gvctMBzvrR2OWeYmNm8tPwRXvLZoMdvzf7HRL5l39FwhYQS2UG4t
mBLYws6+KWeXb0oz3trSnkYKJotpdI6HsQBk8coDF+Pzw/7KwUPT3ENRvshFf96p
O88HnGVAVYV2lt75grhBnfZ9JnXeUEzCAJXh36s6rEjbfC3gSXaEfcZLUaNm47Nr
PqugqLlCcG+HYe5wsR03yRgBREFMWMVkVrUjcbW0QGczR1nZCuDt9Esc4nLf3otY
4mc3l9wPjmAhTrLIB4N1Scj8dIMWQwXOF2E//tCyt5FKynpv+sHNe7vaZ4RXsaxU
qn6CalVVpC0xfnYHBzsb0HUilBJ/UNwuraiiL6HLu9cuEFuNUzNjQKiQyG/jusFN
Tdlarilsa41dQIx5UnWF3iNy6TgMwYq6Tn+7uEsrUn/x1S0Y3tpgkn0Wk1R4W3Ho
UM7SMPKEjWj0IjFYKlf67cemUHaq3l5njM2Rw0ebN90YMM/o3uUiSMw//A9s4eRI
+qy6qSbgszHCdccFF+bxT8CuFuPQ0xOmj9ztzmCMpR1bsid84Y/juuHyVjWl2dhE
799T0XpH3A2g+xEzjI6rQKiyrZdIUrkB4KOdHOat3EpKo/fLccCtDt23UA/JOz60
2WMqy56K24DnM5/hHakr755IP0fTAkVBEhFYTsI27rLFkV+msKKICkysy04UkkLG
+5fzv+lPZ4fpTLJ2yHr5P0GMsjqezPfXQhvSLyZcayp2OZMWcbVIWk/t5auFTf4/
dQacqR8ma4N8CBdHfA8p+6XfRW98h7sCOdOaRb9qhY/BLYlFqG+kDetDR+hyDEfT
p+UchZGrlms9P3itGZh72NoK59blHMrHkFczYAMQukAAoRy1okNJeaTabeT2zv1C
hOMQHc2wg5TENF9v2el5u7jEci7hRIlakogUcatYEiflfF1k8zkchznwVRRjFs5W
k6epWOGcJ62wtSvLomMzpJgXfUDKnhsHiHNKddoP8NY2+wrKru0kltnmxV73bcrl
NMcAoDya8QwZ6wNvZwNYLcJ7Ahod243LutxoSRPjQGA482UF0o1xiCFL++uh/U/T
yAUYf7MzaRWzL6Vw755cPBtnzXjfuYW0jSbuMeCcTQu/3BJhhMYbli9JCcuF6Z7v
s6ZcxzlFPmgWOxKLKJL+MucMqP787R21DBOlMNkqugTq25tl24PWz6znI6/OinAh
wF6cPY+Id0EruT8yoEKBs9bKDIJCwRiCHEt+jakDcjbQNvNkSgqvuMij3RIefADX
gJrIiGkeU1cia9ohSxkDBDDmZiRka0pvhC+w2nbNLF1NR8u5J3u7oOM9XDxTalcg
LYwhtV/3g24kiA+Xbqt4Nc1dCNy8JffQcE+71qu/QZXYKwukl+9g3KzjPO5Vk+Z9
ywzkuO/I/0ZFye9YLqBmYwrW6BERKbpV7KdI6Q5bRoi8a53QKcqXmrLP+aiVe9Jg
2c2oNB4GXDm4cXvn2RKuLrQbNao4zEz0UAWjpvcq2BkKXMMR+L/MlKvkHBKn/lRN
Pg+vdIfwaiwdiX+xpVZSp2FUL60I7Ydr4UsljVf7ZugMkyuhGv/j54afvlA/sTUR
ccQfwhOPmWjP+GgS1v0RRUD3L9xGo5s5XHBXg+SV3uL4rChY5eIfThia8kuTfwW9
rRC7AnVRTwcSqM0TvGigFXO67NjrNitTMUysi1AVZFuEvRZzR28PCKOQ9LUFEWk5
0sey6DxAPfYhxPB2fLxO+mshXFbK119yD1Tw+tgATuRhjFc0XR65PDGRHyJS7tK9
oMJNfZuJRoQflsTQLWcQdXd+/MjDPClx+1ymrSz39iR5OZGCfAPndoLRBLoaR2Em
LI7qMhKXDqsm4YKW6tZxn+dip/PkEtaZw9GGTtyMpVCZ/8p3kgDot83KFBP2I44/
C89iYyzxC+e2dLphfXzAfixb/NEyGcY86Fp+i0tJoIAKwqgNqIboHFdX4oIeSU3A
UqBrLBhL3jFE1TiMPbiU33z76KJf9uMYL1ENVYxJFTYfeIYCOBHx2zENbww8IOau
yHzbcnDv+Mrmu+dRi81AYqEjpw1/b39YR0Gynu03UFvmhFJ8eRIoZlw3c3fO0iYt
fNWoxMkAJ9u5Dr1inblQB7QmhIFECMs5WUVL6WRBaCT9oSnoSAIsJRlJQ+Rc5rpT
DGreg4UUjixd7GBoRoyOFS3LDcKnR+Sa3Lhgvm0fGGwmbSXe8UhJFHqX1H761XYW
nmoNuBexH9Ram1QDnFBD2KaCoCs0u5IfV9EF4G8HKkN2+UZ7JVrCDVVc3evkP44y
G0t13jhSSWR7L5tyie3RCpe/cJqB4apKtlfHnTSbZFvdZ/Nlt2i3RNXIMZy+glFL
0aO+Qrvd8f+p4MyQidv9ZcCzdgrAKlZf4m84VHtNTn/kuvJd0is5s6QBuISX4Xna
oh9nvLxPahuDhouX4z5WmuztqsFrISg2mlOfQOBzvemZbUgYGzdDyR08KQ8GxilK
EnWGolbfOSCwxDBXl88xMBsInBb+TBNdxX6MMONtgxDt+bEfMjMSJum/hRnPTEl1
u6krs95ED6a5kt71RNnHcWmFuTWcnTSrLwyl8+1D7hDKj5TKwgWF6ZMoSjUVqJv4
l5tRDtcA+If5UWStTVyPXiCYWJlz0I7hAWk9jfXOBU7p4YYZ6ftkoi1aE0o1phKf
E8CiWVlFgKNk6i7wTvFqaaMKX2cQaJMWziBtNavi4O9z+c8KLIl7F/PyU2pM93wq
uY293X3tsR1QT3eKO9tB3YOFpkumBRjx/JhXj+mdO1CmIxcLwuOa4HRC9he/XrNk
p8p216tQ1M5XGi9z/3s3fJ9dw+yMGZd4989okiqA3DewI3DLY3BCdQx7st54erKj
+RPhDK3+lHPlOmFUjM3tEQ5UghzdRM83q62d19wqXNZfqHge57n/ZfXyJFTWAXDC
Emi+mOv/LMXd2X7UIMxpG4AuLRl9p+R898PHMQ0WSuYDb0k1tzirdfKBaBKb/yIx
3Oz7IUwE/FfFnRvLFc5DcCKU0ggZictlgJw/Lnz788dpYIFKxGlGFX9RNG75zJ62
wcJ/UGHEQ9dmuzqmkWKRYAXeSHGlN25ocnIYFKwSMaBoKU3mOYrySpEScBN8+Zra
fONN3yWx4V/fcHLwprPV3dy5MchqHWiXjy/QglFFbDHze6kfOcNGZH1hiJYNVT5D
nVyPpaiJ6YDTaQfMHprOb/U5Lgj+uk2Hisp6LCFnC0bxArEjhyVPPl20V74u8CXU
vuxPAPdrmpK/U3J+6mJhYGhY9U6XSHdvdWD54cFFBA2EAezo1UKeWkcSwcKwrrHr
fl8GhtrjDrf+LlAyM1yCDY66V77IbBAVAuOIowB3qoUZ6BIw03Y/7s1+JQVs4TSR
CC5FCMvuuz0SakqydaCmskzJwnh1EeRTYSCC1rOo2YuBYX541O6e37mNI2bQAhRw
Fp05ODJ9V/myvUcOuq0qtAKsCboW34ddQnCo9S51EGkoLYmTsQ++1iqHbpVfoG/O
oZEWR5mnxciShl/51aqWPbh+KEOHttxuRZOOiQf0/qpOwiNg8slDe1Yt8IzICP1O
DeKVtzgZB5PmqWreded9CohU/GEDL0Wgl5+fElgxAgoEg7ECz2d5gL+bE48TJhM8
kwcJZ5qeynGRCl7QDozDl60ioDgr8fgVhJFQkLQDuHSAyekFF21kB5ywrB5zjIoF
I4f8UK+/YOfXf5QQiFZLBOAWuPdK1q92y2lRkOaIxaUNh8IMqY99BbvifO5p1Tbj
FxwH8T4CVOHlQQiURapNna1QfsrlndUgxzfBp6yIU16fz5nvNCUi5lEUOs9ylDVU
uT1Dgdg8beBTko/2X2t2lmn3HxQODjCWaIai8OCQfdgDd0gapr9/Z4GD7fYWMbXL
aQ97VaD7wp1DEzNTJpSVnHT9UCUIpEKqoMCj0mbXUmnc9zFN9/7Ol7+MZA47677s
vWGWrfnDKbt2ZnLb5NAMCMf79QqKATC0byUJQrZJ7qDxwhxhM0yv/rOOiOpCA5LI
JELgdfmmk74t8CsVOhEIjuNyeZkHCmQaPd6uUPiaG1cKp9P9Rjqo35Z4VnlejFlF
/mA+xDhV4zAn9egoAIg5MwL94ES4T8KqvhGeCptgOartGNZjh1GC3mMgmDXqAqdB
UPxZLL1p8Wb2I2MjOfNW8n2+zAvxVVlm8rBu7cY6sgE1XDmxGWa6ZeEjZked4d2l
z5fc+CIynvDdgX8LYV/eKgsUWdCnklHSrlV42N+cs9Gl5cgGYftlcQzLAZoi5a4J
k/fMdEqNJOKlwAEqUC/e1oORT97zokpcS3IIRDG2gcoXL5qpfyzMSIoX4QiP0OQ6
t50HuyqjsDu8nulDpJhzh4EVBc2bsxwdtRsUOiBUXza3VmpiIIveG9EfnAkNslKU
zbFXKGF7jETXtOcvKhPTKRNcydjPzn40uFiCfGn3JNj4v02yPVWaISV4QfE4IdtF
EUyWaWgZKSygCHo4K5vbx5UFm15jpTo0rHmPf49mOLdyzM3349OT/6tTCsVM0NvV
f3p69Qstm/GVONFsClkCE5acHPqkUGjRfNYv68+aaJR0zCuL7fVLb5LotSZPeWEE
RhjOvnRVfFCNRhT9sSK78WFb/lVVTSIVUmM8wkGGpQPTH2fOHesokoikSYZmrTEX
YP+x5IfUa615nQE5WaWuSNikKnFJaVQwDxCOZZnLmwT4R2LnvkpERipnY1VdxQVE
9GXtYbbUVLx3apscEX/rmImdQ5JTk1v3R9HCe+oqxbEcd2ju5Lhxjz4vQiU47b7W
rmndXUerqNzVrMYF4UyJwZaF5Q/1zK7CAmwIfvgJDIP/AgipC+Y5+0AF+XPqRSCY
Np8bJtV0beJJ4zjb1+I9t6YaxIEyoEh0GwFsxKZPcYy57F6GujwBs1CkV07KUxAy
61gGId1EESWT7tBmf+hutfkp5zt+/Ows4SXdjtojGukrJptJ5Zav2ocBoVktVNHX
XDcgIqqCz5nhcTaW5gYlu6I+/6POBAtXophmEgoVs7IVORfIo2o1oQ5cUpIbIKd+
5peit8kKnAUJpjxWKuTLgnHyaV8ymZmOqPC7qCFj60QRG+mXx9IEJxT/qcl/ey+W
bAeMQzJSECAS2p4ghcvqCItsmt3XkMKR6HwTG5QYDDovdS6UJjFnvqY3UiFMJNYG
1/G8hFquYFBC462owgRIe2xMtweDlu7u9B6ZrI0RYu+SD6KzjHKRB4PkrM2SbjMc
R0+NVRDb19SGKbi02/5Or0faljjSCZrFArdV25x8JxnmPguqanafMCwA7b0ztw0S
MpVBqtUw7VfXfzG5aTIeMVLo7z1DZn1DVVGngQPoLxcYzSOwKClRyW46ybx85rHe
AMvSYtnQ94SpEPyVlcNYPs8koqNqcQ26fDyDGePUM7684BZBiHT/jFYdUuE1FWvJ
ynEdINp8/h0CsbDJZZXvWJ78/sAdOoFJ0viTz17hZ9NB9PIA0zIanHAcySnXlHO3
LsXhdP+ukaIlNYS3gLZ2txxNZhbjoIZVxbf7MeORK8e8ztCWPWrS1wRt4gARvQzO
VfEFNQg89eyXFRMEcPKZ/4YzmyJEq6V1aMO0j7LB9RoVJOQHDY2bDfmqaL68Z7BH
s4iuGCntx/p+Wq5Oa58lI9ujy5ebHUQD6AB6DnXHfJYLW2AZf7dUlFtWlrqZqvSa
bBXpRzF1LZouodrcRScw/sp/2m5do2bh4WTU4Rh1kGO+qg+TTbiKAxBYpW2H9L+3
b9yX6bo1OGkfqbDNUBlMjCde8hvkgCOnL/Fs7FyIEQD+msdz6xzpMqOpAo2SUmin
ucdivrxEf6OteZxkL2vjXnN8ojjMjLtY5fb/+5ZFh9eE7xp1N/GvyNucjgjlBrJN
OylgVQwEt5TVx2DpfwXP5ewJbtHbyX7OFjJE53MsJZgEA8jWNiNSg4F+uDBEgKPw
2QfrMuMAHaAcH0J3BEK6OslDjgKt4wip1yfBb5UrJl0RyXGJonJRNQgd2pkL7Fjs
BwZ8jL284VzCkcQ4fMfwjCKFrOya7lZYAFwfDnyFiG5RAc17CTxacZCAd73TzrdK
Jw9uu1BWTvNV0CMMF3TZp9l/ReETLZLkWo5FX/l8KCzo3+V94ZGa1h/eWc0VFVD+
ocQt+wtByVcIjGvNBaT8qyWPnQ7StE7+P5kBmtPWhkZvr6onBz/1fupOCNmr769T
GQFoEHvceAf6pOWpdQ1k1vCWweHymDR/9jzsxkYd2ALguP3Gf3krTiAt3teSph2H
5PO9G371DAVJ+Sjm/CfJNE5wbDcbcU59tdhr/geDj8dXEYfn9WgTIyWZTMmbo/9o
fnfqCATjoCkb0p2+McQqun47c1bXcU6kmLIbVlHL+T2dsiIo2OJfgfw7MUcjEESX
ZyeBW6UZIfPjK9B1i7b6Qme6acTC96Iyx94CwdSD8uWaXdUB7C32e2ojDrSNITyO
QIuG18Gb7WN1Y3Cw/L4jWcsgz1fYVaA6HRstLWsX3rCuSDkNWtKM37cdFC/J9Z16
9H/1UTO04K3y04njFkrxecOuOPPWCEaTiVvG4l+iwh/dTvP4NE+ks6mmQ78W7XF5
0er40ska+4A2Zi2bGik7Km0999bFp85HuA/4oqzbYDn+c6FxWUJ9JOSo7oPykmit
RfxL24F9doWQKQ0I4YBkTYIMILDz9TyDZUHNQIgp0SdGvYTryuJYDDhc8m++Z4cc
u8WLFIHFONvak+rY8efQNaqjXqKl9471X4oB/Syisrwz19V1OSdfKuhM4iacYvoQ
zqyf4aiuNALBc2o7J1ltBkv+92O57qjuiKop/berFFWl1JC/2soy5A+Bg3pvJJPr
6ObGsQQVS9Ut1GsXkKlQF1ModkyEANEO322SfJMWzOShz7Zbj/lgtsQBMolt3KI/
QiKzO2jPnjLZmMm1fhRLgFOs/7SzQvfceVn1a/kELpl7AQbyr1ZxCRkx7Xvpt+AH
Q3+QFytZNiLAChawxBwdOV+JqLOTQCUcvPLoSBNL7ff497cgso+y0Bge6t9OWwrb
D4NLu2xJ2oJR5Kr02nDRKyvuG/cbLQw36I1K6+ma0hZnm6NOv4xu+Fpg+mBOkz2Y
jNJ7j1SFEKPN9bkB1AKuoH5Jlt9ZY3hLCzj7MDfgsYU7Xvtqfd/ylNQ04AQO569g
3gzV3KF7Kcl2j9OOEKc0fEtM9XtpJAH5FY8r5WaRb7HnX6oqwb49VwwTMnqB6yaT
h+X4FtXQHVdG3Xlo9BbrwvWgN4knkHN4fplVlyyKuS3QhwA4+sGDGf13LeX4EKUG
XJORgmYaOTY48V2uhWyT7IkDA2eKu2FIMrQ+7qzzK2gIo967xJxo7UJWWmNkd4AU
eTSKWCP1PkhlvjI15Ub/IbwBNZhwnGKA7ypRLwAVWsQzLprCt8e5VasOwo45ExPC
FULvGCiXk1NX7CBWkYzMoCyXcB7rdlMtivzqZbB7u7JZ49JomqH+7+L/zlebHo/y
fa0GKOb+E3E2pNjzX4X0C/bzEEyKOhs1VbiqXOI4pbEx9Zk0xR1iC8/L1EFkShtP
LEZXALxbwEcvBCcyOTFmbYS+sJRuX6F+qeh4kQJDYD+/VtCN/xCTBdyKHv2/LXmV
HKWh50VGsxwi7sBsO/ISB8aF6MKxFXiXygVzQfgrjn9eD2f8A79vllzLXJE1ux3C
fPL+zOQR3y/5EEq8MFcGl+nmQHvxbbqsQk2cd0nBbaxufrjGE1B1Wart9oMl7Kra
B64lUbqGKH+5OQ0h97VDIMTc/qedXrPSVTeWpLvSFDyoiKnl8Xj9fV2+hsSBA/UJ
KrMe/wstv5j8ykhh2dzjIbVqY4Kg/vZ4v44c8FTXT+7iZ9XBG5+CIrX0EICr2jI6
K5hONkY/VhWSsru+ZuUNJr17TyOSL9kc/1kkkTWzhG3cJkBGLRdI/n6A2itIlnzC
gvN1MVXCw8VILwLdrOUWEeioq6UV7c7D6iBfak15B/5BwUMTZjYLyH0WJkHT+IL9
DrCDb9H2g+EPV06joYBMlJkvFg+ro9hz4nOlAQJCZUj1h3/pB2gMD+cURFphzbF5
DMracssMT+QoJzX25nUwsQ1uiBqhxfUYJ/l/N7Oe2jTVF7tJ1ltUVCrVpbEYU5YF
ua8fSxe30paBCVgLm7aY3fNwplBHfFIDs3bpbbZYY+4+KYlzQRW7YH0JJzC2gHKV
SM/7M8BE/2MdDnwI296CPsLnBeumZiwRSmCYK9XUhu+qMAaXOZSckFN89zW8N+jI
xvNd+PlXl8OnH9dX6Uh5vfGlfJ5BTux1lBdOHjCUsv0eNoB4dVqNSU9lW6tpu7lV
cm4tgcJtfho+WMZYclQH1JAIS1eYo/6g7UhonvJiEcc8/XJFOYtgEb6TYvm8Q3Tk
7BXhUEONQNcByzN8inbFgnfLEh38UmRWm7jsmCm4mfk36O9hqKPgSL6kTMALjbmA
GEd33LnsDJff0wN2F+oQOuZvT9eMLV1TKeUD7pO35sOw2ONBHgulQzymM0uW62Ea
1FN9FYKb7/Yid1+erNBt71SDv7+R8/PSQiG+eiKrYATZXfEEFOj2DQELQWDZrweu
LPLthKLXHTtPLcvthDwpqWNS3xk1oQee7jPrVz7rZR4ymR5pQwGyN0s89gaMqBxH
jjzBQv9+mdgsnSF24ltmUz0erPAzJ8SS0ctuBxOkWJPk2Xg7X0EeYIBKg9HVcjDI
B+n73JLzY3UHCci4juHQfX+pVSAJALGBHlSv7Rih0SGBO/EzC9I4U5kc9QzGDz4l
CA/b6RsmgLhISgywrUcTByhRDEaKhAIObdBc59eIfshYBNM8gRWmYZfevuJ4K7L7
uTDfepj9JxRw5pfoIZ5n0xxGywhQiSaarV6XJ2Vh0F39sqZL/sdY+A8YqJf3sj32
ORDIPiIYj3W02TN6PBD4xmK/LGSHbdXhM7A0FMqTLcmaCLsj1ZRp1J/0QNtZuLWr
FFpN24aSnmDNBy0lsaAOp47qckbhuzkV1Sjb7B1o4WyBRrgG0brJASWMke/CN9X9
fYqFNv4dgmWkefo9LwirL/ILvwikVEch4pSeg+lQyOmMR0BP7btQ6n4r5t1QRn10
LKl7Adw5fkY4BYRepJb4iutPKrhbbIp7r6P6sdJwC0KPBXf1nxP0k7kDT2fXsC88
pp4iXVShqBctQqgASeqdpa1iwgcE40f6n2MNDOeQ61BaIjB4lIKe0Ky1WpKdiOND
Kod7UP2+ggi8zdp/Q8xS+rLk6/B1DXYJJ7aNQGQDHGPa6ohDoGmvQO26Eac0VV60
03T1dFWWd7I7oZ8kwzUviPxBxIgVb4ulaWUvEgnrxx+OZE+8sxS4nT8FL6GSIpJX
W36awKmdBkMhwIwy0WV8DsURdlUybpjsXVOs8aYV/7KrQVROFyLgT4/DUpr+yUXH
4qB5m7o1JKLD6JAQ8dkHqrNmcKIMNImoQASNr3Mbs0kJr08JtGbfFXGWl/Gj20uS
EpeMvlA/H3I+X2gUiyZKt/7G+n+rX8VLk7PDPGat3Zh0abfWxRcaH2SNfGtjxCdE
6/XtGEWnbHM5mXQNasIwcZzE+Ji301FkNcu27/vrdRKNJx3vdg0+aWvRxOTVitIm
6LoNKIwA7bmqERY3qQNDFXq+nUWbj4bc3Bxube67YRK54BMYNL3QKeRGF5ffXR9Q
hYiO7GPZXiJMjOAvQQcP0z9JWEypLdM+DwymcfvmAvoIOKkAXaetzpDVG1rBu7rK
doVgDmBPz7M3ibaiorWmGk+UGSK02agR+zBdzAToqws8WOetR3cXujSOnlv1txvp
oydZk5w8s35BytqgAqC1DdUzgIzacQobfbi5oiTJfR2pSCkS20M0Kguk0UHoDWsO
u5Uk4RoDWl/Jy5P3y8mkWBolMu4J0P8qky6BIVLVsQeidA6aCxTBRSRoH7bhhW6W
TxpbLYo84Z2EQOn0otTPs3/XzayV78eftZuqwWW1b4Q0L2TK6bn4v+Q2yHVO9ccp
3xMtqaAVjlB84+o39GSXfmc3LIiXXQdNOU90G2vfs+VUp2FIS0D5nY5Sx7yYg47/
wwRqcucBYnJSpM1QsMrGuoswke6OPhIOtQ+OW6kubskvYsTlM2tP4ry596svGJHu
3IyyeGVyCTEfU/Kni1Lp0isotW800V7+kP/4QP3JA4vlyf+yIi7gj/gDyeLcT0RM
gOoJggQocQflwL1YIgslhdgsz+J8JpbUA80Ql69XoHTb2QxFUWrpwspcLZvJcjvJ
Ho4GxYRI1SL2TTqr5MgDTDR1A/BCTSi4MCBE+7N77epLhjmJt2n8I88VrGnRWD5y
WCp2eittNUjLuVeiSdpfVvQhSuu5l5KPV0cuB4duM4drusCa+VP+KQ4XImHKEkks
6K3azamo2qzGUwPQ54UHaujq8hQdxuJcscNLmJJiMpM2XpyQ3/VXe7uiCsWtsAcn
iHLu3ZeX9eJj+axP9Wq0Jdc0mYzF1jYXKxYcTRz/9O9DrnrMeFTbqLHtMHvUTNGa
sTTwpeXGqzbv71ba7Esa/q3GRnWt17TGnZ1l3pkouY7uIlwCC+3xkFzaBxhtR61o
2HcRe2GzyrYA3A+1T14FVPFdVCefr8s7DwIHhdYj5K8HIPXMOwg+bj7X1AVGwa9z
f/ofVV1LOX383Jd70hoq54drusgqsmf1MX3EJJlZjZRwS66tR8r5Ce+1tFTdwxtK
FNguRk42cB4rksZvQTVEO8Fj1u5W7cCxRzwdrDHHrWsBVL/fGIjnOoT4gSg0CEOy
U0uWAT+jhUzTN86MMhmV9Ys8CY485h0EZD3re5VZQEm3j8Xhv2a80Wsqi4ug7HFu
f/0kxTmp6b0WbwlZ9YDs5FT+VBYUMBe5Wzfs1qF3Ot9RoW5K1wvWh/6Tq6wj1RVD
chb5tiY3PIZWLPg8AVZcEnG4xspID9rQR/L2565WCDjWbYoeF5SDHsKVK+JG8JcH
BXu4/9obuIRSEfEY4scn51tqJbfd/0tzA81MZhzvUKiHmMPrFGCiuHYzJrCDzf6/
eOwIT5wzDNFZ6UeRlZFL/DYGqQT5gyHm5w9SfJggMHMtqYWGSQ5t398TEBFOuT/M
klX6pFsPhDEzmVqmgbBVfSzMIrBy4tcYgYbrbgGr5E3WB8FvybnFTuvgok8Q7RZf
nybWXH9ADUPbsqsEcJPGZcadmooU8ZojgQnd3JRo6Gc7y8jxqiqIEXCdteh7XpUd
W9hwzr79OEgNC7D4gAYQB016vH8OJHry3HY2brIoBbi+x82Qv6V+nPBD3kgPO+Jo
JQ9jTR4vvq1AKUEEBlCyNe8CAQBn+2bbDKwN7AtL5iUp1CX4OHao0DNVH3iUWpv/
syMdcGAsaTpGXLHxMFCOUbiUA+0xQBKVxUvCqkZqUb5PQ3cCRfnAnfD2m7rKnxjk
WB3czOqAEYHCEPM/85WG4OIo+fb1uqPMI/5nCsIJYw8nITQ1aK5nFLwjtZ7WTxPm
WBhf/Bqp+M3al7JmkwOAtAnMI9BQglpEjgbugtEhD2LwJW6+nxHvMt3Feie63pNy
2jHV4SZd0QfOgaIvgbtOZxPEuKMASPBSzAvwkgaUM/pvpEo517P76UsHq02ljrYW
wLnt4zTOvGJjOQiOG7gwMz5dZUIL2dliRJNtG9mB+2qAjBzbY7FD6XaVEwqS3Uar
xd+5oxa70kYvB+H7f/8YGEKvGZP55YSbFtPHeGUz51EMK+3ESWo2WS5iYhoJTCgD
GS++r1e98cDpm0OSTgLUSRhiAu5LfvOIisQLUTLNznoBSop+ZhX8LG4YwlodPl4N
hzErpltV7k9JJqXPCCeIylg0YNC6akuzgOGQljt4LGTuAU2ZrXvZsjXvtKoarHEC
u+7KcUVE1QbySjgS59Vr4x0wuKLRh800hm/A3kriBgwIQgSKM3j+KY2Xbo+JG6WT
GlqTErrffSrjty66mpSdng0j+CLAxMZBbmbIlv3DupXPDJb6ha+GTvLyKTvPWIN5
jOXjsdYSq7wkHo+iuHc4V7OeS7VDsA3XexIxUY11pT9c86VmSC6ernzvKEdMS2qS
ElrqhQihODAKvF/4tsstuBZpwqhGvQ/LZFSV+nLy22aASKZno5VGHfrJks45Ywfa
WqfSKbQ0dbuKha25uJ+tV3u8EyF4cBYsCjI1MgfwSqHdC+6NkderMLdcBDhi37cd
nf/rfUEu3lrWOUMef7iUqypc8SOFWTrCidOiLMvQZ2DgPqOpgPiJ2drAmK4ZWxRY
VobFMtw223XwFZdyWX4sXsLR9qmBehQK2yl4FYRS6nAbjlAKOwdNNPs09ExHSaIk
t65xL9kqSZMX7LRYveis4r7L8FEQomNkLLzZAITuIWwLWmhj+Lx8mjLCh0EWlJQ0
dUiumCon+YdP4LnIPA79e4XZNMMzvB27QGazhkFVn0jA9IXiabTSAxROa3Wv2drT
LvphBuO2lfX95GQ3T2Uph8tLxB+fk3ioA9slGFTGKCHhXWef3UeChuavTm4p5dte
UQFDYfZskZ+0KAfyoxwsCzTtQCGArcL647WjADOAu1IGq3bCRm50WbY0UZSKZgyn
pW2a1tgs8YMStt7MGTKzzkzb/Zr3W/ke6aeODhtZuwsUPuiKx2xci33bf/3QAL3K
Xth4/1TqNgHEEBo2mn7ZwTmPB8Q5myeRr79T38NH509s0fJWszfcEWf9L2eGP2C+
pIDuNpk6Lq+pgYfaBuYNQa/u5U0Wbf8yvS4TvFEYTh0M61c4epRuNgtyxDXfiqOi
Yo1ng8tdsNEyyUCB02+UyVVRo0qlj0g3+r+wYGCz7E53HMbPvD6Hmep0MIbKXs+1
rqH8srqtKbI3Du27CNp9ua7h6B2XEPQsE292kinvP46aOQyWkti5pjQ+V1TWfWZA
f1VN3N4P7o36HHr3wWcVkGshlA0FUMc6KktuYWGfAlVB1bQXrDGQFPhbdHw0Y8jf
Cz871lfkxdSKKKZXPMSprXt2WFCNd9HmnniXpy2Z+dBmwqgrSNXTmknMB/rNoC47
WzWx0TPIRtwdDcFjBFaWJ+8+nxI0+7ImaPeQykBNWhRDZs9sX6OLFBDQCcijORqo
O0JoeGxKHnlJtBIauJPClrO2s9llf9YyZhGF912jaDRbj+Mdl/mCiRZGUz36y3KH
yu4l/0GfQBbk8g6Mg44SJNJzb0nQ324p3890CmRmiEJhYUCUd4wIB3NJSxExk/gs
zzOlB7UNODqGvQkRZDnwbHhZNbeYtCdPBh6U6mYw+WVf94zdBFsbgqHkMTKKsmwN
NBK22KbYpttikVCnv36VqX5kBv9/t+sjZmRTRhmqKbLLLw7d8Fb9nBvc4Ej3js/M
jlFE4Cx75+dBdtAKa23dL14V8PO6kwj+qkSjggao5Sw1z64iIoaINeRfiGBi2BUm
Bt1N21lMM2+Anb48+8EqbUC4gCUdJNX4X/RvjoP6wFRaQWITDkFsWAHmYv1FeF7C
eYZN6X2cKCsRquajG0DociJDglCJ3E9dJ+MNcQCrevi94MfMGkRM5Mq0Nz2WNvfq
c7J2MDvx/Qw7TQBw5IecskEDN3h4tSKIHvkyYtNwrDgy803cZsFxwIWd6TH3EQKM
mUTy8jEGUHDv2b7bbNs3MfaFCZj1blGNa1cNc4A3gInxWhJ5tWZWO3xL/CvYlilu
lCxP8XGyP+RIL24rqwKKTDPzdJ+xdGRheo83b6397O8eIJqUqLnM9cFWkHo4GjHh
pEm7pd+EcXVncrwTG8DmMgJb6ZGhPEB/idrJJAWP+GbDgPfGlEyTZ/P/67Y2S6IY
FV8KFNbRE6lufJaOtIb7BhgYykHLmYI+K6gwKst8mcke7PFqR12bpxlw4lkR7BYF
MaM0qJQXMXEfcNSolOYguZBc/Zr0oKLCyFTbvoU26NCGuoQ1e8FrS28eQzmLn5sB
IOssJ/jfSRFsdCVdHtd4g1Gq3Rp5tgR8ahAwHrcMNGAer4VNf/dWTTsLNj+LFvSG
xZY/pfnbASRcSc+dBWkWdhKfn0IqOBgOVqA0b7zrY4NzvD+aAnhzziO76MJKQ9oh
F7p/EiOVmBmuoSp/6I9rIiVwnMoINYsyKW3Wf97O602yazJ/HAdeBv/YewIW4qZW
cYp6uk2VJ3SbejL6GBqDVG1kj59S3VT/N4VaV34ZpordMYnoOQkKpHJ+DAJ7k5sp
h0U6vN9ssN8w8r56ZYaurpFAl+4y0oQ4e0j/bdBdHtEhiNY2ajtwkcAVBCj8u72i
weuZlu15RbajMqttdM9FtYVX/481mclF6RFmsybjxwb/GTFCCF1Dbvtll06jBVgd
VVtENzG7kYk40GQObeae7iNDOj7gPMzpVHSvcfVSa1881foZfAzjLHdtOtXait+i
yXwEe+qCtviV1wLTKKJ8L2py5WI1AlJ3DYejLtM7EiNvne1VgC60NWDZov2unXsJ
G8sE0GFqnjUeG2r6tW/CbQp9Yrvr00MJB32itfhMHWUpKEHGEqw4b8J0WSRr59oM
Rrtv49C5pajqWYCq6NSWYEoWst1y83mY/f3WBysp3akqJJmYUFlkLaoW2ePeuM8n
1TEwHBKNuCRAv3OfCroTaTqM6ErPivbKMznmRC9g21qqi7msrH2d7IgmsrQeIAUT
vPYnwytJo/Rn4njvIT3FUctL2sPf/ih/ynu2mV0kW6XBJcpWOEuf2+sMjN7eckww
qg1z5R6bMb3g5ULXxo5SrpfCg4dY1x9riB3glFkrGpgdLHBQvfbu6kSc4pjl+IOR
JfVE9NZSScJddDAN0Ex867cXO29CtL2gPt3YgWEcLRzsuoNC+jfIQIFlQjRR1UC/
pJRGttHBmFqaPWaPIk48V/xqvkNAQzyzW26XtzXnq3QfnInySTbt3Pd3dy5pjZwZ
zonLTFyY6BwAeZxUbW2jiVtwRQ+ohPZLfsud30GnZKo4iMn2dxvxK40QiiZrcMXl
E5bGFJIJgncngOXh7FcpOs1SVL6m7yEsHu5H8lyDtXMEFy3rJL+Jb5NhqvC1YUqT
K/DxTvd3Rjk3Uf9FDbLGZGV+B7lJKPNrhFIrr7XKnTBfRwlj5Ul5q2NLitC8IQlO
38bVfu+7Kqi//3nCsyCtBaQKYpzwvIFmg7E7iTsKKD1yHPmuIJWfVp9EVxFasFd6
dZcJq5yFta801Ce4X+5IBYhw3w8xUJdMPdb7WCbGIHNtvzT+uTS3N9rY6LKeGgby
8+WSX7nJ50nfoxqtDZRrQr+3uYDTNWaz972+nvdMd+6/zSHPfyjuBysR1/uYvV+j
ZsuJ40zoT1ikU7BIliWqzTnD2qOcTfzc+Z9siRyEAfUnlx30CHjRk4qFHrrTLXRk
NW9z5c+PmNQaZnS/kIM2nQw77Nk+13jvcWpQZ8evnVfdJYEzyDwB6Y1oN0agOiOz
VProZ45QnhRRph0MFY+U/QuWpZ1fZJXng90tkGtPegyZRV1nEC3kULdpScLsTNxH
en6qs6qlp/buSJl0vZtG7s/2Xbptspe/24d1KHbBZjKBtAlDHPCyY4pP8tffTcj/
2EtuYyzGgaWZ2Mvw7HmAMtxIXFrSpWF4lr4c9SBOnkY94DgD9JlFLF4nngbjEw3L
suUmMWWQr7NPTppG3xX1/3RT0gMQoKkRwcSU75N2Idd6xq7IPfu+Mhbcwet5BTDh
F8Tyw6FOv/O3D5MKs8Ad7Pwi5OO+3NCxnH6RuUWSXY+ywpyA19ANuGHi6YWijrgp
/xooxw8d3vsaevHmtApzin2cjihmMcVZbwKpg3zYdRLtYkM6mNulugO8Huwn/UNu
gkQqv8Lh5eopu+nPTSG+L+gMEhGwdux7255qy7SvYgRNuUQ5CVelUFTgvrahwtIG
JdcjLj9YBdZUTcu+QlKZJFNXuTgcjrjEw788YxvMmRRQy9aB3kmGqPJASWhfvAhP
Zrz1O6bQlP7ctpobHUqFeqT12ivln+QM1O2v1+Q87H6C3N28CvALj/aSwVzpsTid
SSGFjdoUYStg7IcGnhl5PzgWHiPDg6PcHHDO0LkQrp6dGRhoDb45c0371NXNzSWB
75rfVTUWkhGgqyHDeGbPyKLV0Cku8J8BwPilKG+NIGi4uN7eGQQvsQ3/vKH7lXyB
yEfWf7YWgMIwRrrE5f0NASJb7VUaP9eF+5e/nKxi67m6s/idboDb1EyoqzKZt5E4
TrdvEGGOq/0BQrFS4p168bc7JWwlb5Kj+V0B89IGdR1D4Zly7SivZTVBfyH6lP8C
3+klsRj6Pr1rg1gddMrN9kZAjUIdzbN9SVJJ/GJs2KCSSV6SAk6mZvaM83RZIM8t
g/Hf88FsJXlNr175LtcAVVtw7KRa7Mp0LrUqQbjCAgm8LPOQc1rvtu8kQ+MnZWCz
ljNoiRLJoGBaQ10MSul64ph3iZuXQ7ALlDtpTNp70u+TTWgdcIsXFhC388GgFHed
aFzrTocn8EMf6Kn2dFrtkGFPx6mO7v8x2DFfWEwHdX3F0TKhaH1rY8sAmlPeX2OX
fQp2WLmWp3nlVV+4il17UIMWyUVe7mgFxm331VED1GKlk4puqi8PrJUSP5n4VJXv
0dYxER2sVr5zZRq1I+19/XCLFdtkoGkfCIyO/WMsns7Kvj+fi6WNmcZKxItKEwmq
V3XtGVudVhYf3z18glK1o7GVDPDz4ScoOx0x1N1bMz1ulGfzdwRAyFCjzaYoF7UN
osZV+3BQd7LeiaMm00tUERv+Xk0ogC2eqY3Eh4Cf3uF0tJjrRLZ7LHUZ9w49s1PE
R64Cjwjcy/fURDT88TINO+DOmXqjcrP8MRjunmVgW43t/wCO2OpXiI7Q60iTIhqq
L3MmMVrBtwlJvQjAU2rig7v0GjkN7qjxAZFNUGF2NQRH3o5P9lykz71fU89M2vwV
Lb/8Xm5trUvCgYRTGmOFok1IBRLdCthqiBzubWfnI+A0h698EgcxnqCaN7eI8VEB
ElX/YK0CNZQS0nX/mjvBomZZRBlndPOLcLh6xeK+7GcWhon5sHvSQkigV9OygIyO
l/NM6HloX/EtpymSTIx72fw8kzD1zHndzitnh9haT11QRuRkqv8Obvj9W6d4Va/y
LYSAK0tbLhGgQYYi88wp11SzuaoRB9Y8sPd9e1o0tts6Dp6HtLuG1sICFSK8CyjP
4NgxwKCqon9GwbomFvKBCi6Zg6SGKgFnakb6TMJ+jordBZFAsabbI+1PeHb2DkP+
C2yoisKvRHzaazpd1WMrzaaTARc4hx+JuwoWaaQhxWVaeb0xQRtj4wgYel93AWBj
JOndwhXCXBx4pw0puKCpJRAsQ3NFXcyfUr2IlvnZh4kHdjplVdW8w2z3zrjPu4z3
Ww5xlIuwXkA6y9pb7tSf9gmwkn2PI14EyeoQYlnET9Tlnn5DJT1jqmG0F2IhhYS8
F4V9BWSJdLzYo6YwSYwiLwjhrPLNQupk96xKSh5DKzGaa7ZHoK96BrZW2y2lWsQH
G4WDTzZDqDAn/e1ltVoBirhwHIEZis/MePRU/KLeqJiuOsP0jmdg67OmoZ1ZvM9A
swe0gtF5Uk3H6TA2Yia+32udm8Drv1r9sBcAt88qG9TA6+qaTR69B5BjozbYPIgm
i8IWz1BiF4YWgT6DhgeI3LApX/AgMzQKHb4l/S7xNL45DaZORGlWep/hSASM7X7m
0hlsalbrkpHX0gjvZNWFfbSZmezdKgbo4ZHFkBbS+X2GB22dhomFc1ntZmkbdhPM
fWSDWLW5zw9BaFv8I2/ywZEQYbOa1f8DnPorm+egOmym9ZA2A3tfYJRhEccZ+xlD
WqPeMWwlnfqSZ8r4+OmmxnkknTf8+qHJW0HY6CfdQIIkFiCgmSgBoSc5oAVIiamV
Jl12IWB+GOhSxh66eYjITaiVQcoqWLZjzxBJ68OxzVRB5kanEFgHgYEw9s4M0daZ
sJz6iDY3qEKXH2NN3jfiVKnWMfvwWwp3Y0bdbHsKxXabD0by/6Eq9i7fetATtdOn
hRKi9ctnQwUBIye7vS0nswKDWFKoMk3zQAwCNjI/eyDbuX5COjb+nQMH6yoMSa1S
k/slOPJamN96V2/vrbdILS/lc3EXlq+CP+iq9ryVw+JqMYNBi20fZeQyjh2NvART
NamEmJaRonuB5I6k7t4AIQk/sGmqczI9iHw21IDFWJhUdw4qpAW784NwAeON58sO
Ypr1r+UJ5EQZNNgzOAOgCUeE9WIfl7rYysUsjr7FgcpO33H3ao60CMMa7068YBPo
3BvVOWxeCtvp7ZkbdH53AN6O0zFNqkmZEVVRXVc6620iLq+U7aqYZ2lUYfDxvDNv
gtavtcll2Rze7AF8/qEwZZzSIScsqJ4VIRSJ25D/SIKlJp0bQ1Sbzxo/BrbS4uQ9
7dPd3fzZGliMZ5T/PMailUrn1/sBTvxsKOxEdL7yBqs5Rs4jH527djCCrYhioDDp
NWdE7BaEC5SsQfxrdywJUTdFoKCEjrtLhlWvVBKiXvpLMfOu084vK4QLWnndPdUR
ck19J7D1zy/zeTFjfivWooDDGoF1AmP0HHf1MXW8nZ3jio8cSD7pOkSH0/bTVY10
vVDh3P+WuDrDAJxlnBuNjzhQ4CKEShAy8WTpbQxLZfQebbq+CINfRj3c2afViAcg
ktuQQzNgpwV+vioCZL5oV7MwrGu66B+Kh+JueJaRngR4CPl6iTgTc8GpjVO4NGSn
tBVoB2ngXzrex3THIj+GlfE/F1tVpEORntglykX46tBwsEbwx73gSk2GGnwPWyWw
rgq+ODo4Ru8m+2Zx6KSQ3BjmmVgv+OeW641Ul0nqqcOSlnzoMifnh/9OcgpNq265
deIfzQYwkay51+VxayGkttfKBZyBDjZhkOLMDZ5fcHYo1QwGO2oc25BrSYqgc6eV
YjW1gpddvcgaLTmIPfZHbf4GQBh+a3prLpQ4XlUkIF3oy4cVHkl8eNxebyhyrTsJ
F2xSG8NfjKjryBg+ZaQbr0X8kPyRSPg1Boz22TWRRZFJG5h9Huz0U+h2/QhY2O6v
3dIvaVHDVonqtv1RmTOk3W0i6V6HBAfqaGpyUjy8DwPan8CR/KNggLrq7KLo9j8a
3502QEx1WG60OBP9NG+OvYCIU/9NtPdC9YBBUaWGkSB+7OYWHaxShK3YrQY7Tw/v
94dsepSaUW39+3wdx+dsxHAL8zsO7uFukL3LvyX5U0K3iWaB7PsQunvJNyuthDEO
F1PebcKA9C1g0gJYKWNFcuHT3jLKRhK2DDxXHgIGGJocKBp+niPtcgJxr4Eh2a4h
uW9QVr6QZBrzCw8OZggw4EXZ2+XhzMhxASkTpnXsAsLjbPHUA3sbCzLbZVW0k+pl
+F/nIrM6st60b2c5if70Jax4ulCusfoWnmob3dMmUBQtl00+xIMvioToOD3dEqWj
PcDr9CedOis1opxHWIulMkRexgeoCYSOj1OcP4j+bnCFm0jvYtRyNH6V9sTKDw2b
BPivKhQbTQJgOpd93q4RNQ2AhCTjyd0izPMCkMrfPBPFLs5YvALPrnkB2ePFYcd3
VmerZ1P0pwpHAa77DCvbUUCBbV+Kg5aVWZOB97tweVq3mbAoXYncZKPKRHMB64OB
FasE4qYSQ5oh0SPkGqZu4WgH2oC1ZR6deRH+RPKse3SuE/vkMqiwRghPVFdUGose
ZFc1Ez0KbDqiqUiiCWxBP1n5JrAqePDg3d65fTKM4wtis5Jyf2yHMk98ayFytg/C
0Pov6WZQa+eCvK7c1D+dIwALI6T4zIzqvyRnzuARTOv6vPSRysTrhWKY8TI0Zteq
iOASvlv4Y6tbwsWBVjLrtKfvrPSnqmqjH06QHGtkQHzY4uNWmEoCe81iahOdlKp7
5W78bs+rs4acFAivTLepmgi8sXgncL78/Sw0IQIqs6B6zMiIU6KmXDiPypXlv9i+
Go15Id4SNcZhxEn00lQnJV/stx7QqGVecZONIPmQxP3vfQ/xtBEWcc9fl0DQDwkh
/Hjsgl+7fBCAVNBlnuAY829Vdh6924GG4Pe0GXg5sxhGi4JxQMVw6ZalWEzNDFAi
UUAr6pfqq4YHIV1bJ3LHKLkBHMF48IYz6XP7k00guOr5sV7Hwu1c3vfjypMQWn33
2uKKB7whilb6D3GVdBMk19XnTSLPX+Blv2eMAlJOI9aiCuox4qwDGei/IRq/WQO8
/wTpODJ3uncjwOFnUOqkp21I+HbsX6PITe78zhME72oXbps8908ubPVqwwzyAhMO
4s8tbyWv1ipCVl4KA8J+X6uDmNbx+pxyZj+azlmMzL92U+fppw0rgeUCMZHaLqEk
BjyIFgFLVItQ/lL5aPjDh8qPl3LIz9HBBxCTmWANcRCXJdup1KU8a1NBlbT/yKRK
iVR1dXbWisUsXdeLzBrV7Jrh2LSns3aCYXlHPo6vSI9nCmt5gFRctVAY/D/b/ksM
P09XXPcJ+g3QozA6+yWzbLi1qeyMI6sYGeREqGb7cv90Nwg+gDJUaYbTOf8hKiTZ
tFXdNjiACMljUhz9hgMVLBnK8imx23JvMsqs3e29iDxF05h+hzBeiBtsQ1xfgDgK
euWy2gzO5ZGXTM0Kr5IWXThLWIpUTowP8GKDgT6DPqqFDZfXNEITQPGVWVzJq+s8
XfdOOzrRRSBvnE1BXT6ChuIr0jpLZBNLRI4wm1SsH+Bd6JJAXwnptuANYlHr+QDc
5nitUKs/sS/NJFUAMkJndkOABb/vfmpDlyKOodLrFs2ylwzJYVeU5URunwlmDcO3
McyKedKbe8i1MYkgFQCCN5QXuvFX3l2JRAiNTHIJ17Jk31E4PedoFh1k7gjHRo8/
yL8Cq+d6q0OlQwY0ksI4cZxhmmsZMi6chFwKSY3v2oGyG1ChSJZy/963eZD1n+wn
hVP9S5SwCmOQVIkeeTDPWMNkbTwD0XLIeilhZbmx5sWPWxrXYrgMB/hyBlUl6pJ+
zX/uie49i7ilKqG+V3P+mKSTu7V2+xN+b4C840ZOspRmSnHa7eB2PNEXpP8v0VDf
IbxDBXDPVNXjtQvZURNOAF4S78KT+Ap4FAAGk9y5KyXXjMCRnLe1lslhVQgpF3cN
w6VKTC59sffwrGbGoAmImZy0PSX2bo9pT0InNI8Qnam9uavm6WvunQdatxsJEYRE
Ct4hWjE4jgKBa+/EdRnSPJgk45p+0hQnOZVH1s9pkaGzRuITfoeWWc5IkRlO2Q1r
sXQL0RbCaYfi8SK9b81eQumD1iswcX+otEZ22YRNZvEryPbK6613W+EOQeAkOCUg
zehnvqlzaKArlDlz2+iymSpE36ggZY7rRyQ9joFx8nRiFvzz5A4T42+WZ2gM0hWQ
fW72LkS3/gt6zH9CY5wliUTBsplEsLxOnhFniR2Sq2rPSVeXO3/baPOYunhUai+b
0C/Fee+/zOwp3NF27l/tC0UJgARM7uFe4wVdBWBg5DYFBCKDZyW6lAETDW+MEKXo
HqlspNlefXuFZHDML14h51ZOGwFwQsvmnzShzywg7tK7fpEOjGZ6eSH2G36XVAzT
VKSGlrDeifl4d5pKGpg4F2uoNUanb3Ki4VuZ2AUIOp/epj0OYBlbIKRiPtNsz5+M
k1jXl+3rFph8Q1NcGXG9tElYE/1BowBxeHGCafa72A5iq1i6WrTDU0luISWhFgSu
i4LCqmE77GAvv6x2NedUCthq0C7+Mk9K87btHVDGEWsR4pECcjrb5SqZDFc/XeIj
ReCPLp54SNrRh7uTjH3WkAIiq430QlOzW8wh5psYzgdR1rXzJmoKoOUti/iCSuEg
LVuxshhmrq2rHe8C6QGyEC5OF3OkwBua6sDVvMOmiD1uBX2o6lNg4E1wiUhh/Zgp
FIh3V6lXTqUXDJvU2CgUDzvxm0WaOwMmTmlzO0ROqLBfaghzi3L30xEuv1rNwgKY
CdLEvu7dz7M0vg+oC8aVkG5D+9YYGdork+WLRL4bcznvDqFs53t6x/UallVuxelU
VF1kwkKz3y6lhKdQtMB6W5JkV1TQRPEjyXIHrGI/uwYNi7hu4WzPvxT3DGy0PMLP
SlU0lkEofdd2TgtIelURz+VSclW3euBqk3WD4KZaWuDnYKIgZB7Gqlg5hKdfBDPp
fUrYD4HSckU6vJEM8WRnZD5Db2QmPfcTvSeOzwo0J4Sho4zieL3HzJOxQIwzGpqc
JJa2cTqe4Xye8BbHyqrda4LsD5UrnGUMdc/7W2o/NbW302BQaUygvivVkYjJPTVQ
wQYCba2W63Ny1Bo3tXW0sYPc/6ofrnmvPAmZSqoYpRyNrxBe0/ONcOPQsY3RIOiu
2a8IraFAhJFgN043ESk28i53LbXC620I+Mbl/HObGlnTD3+V+PDPCr5slu2Q42sa
kxvY6keUk5iwHbVDT2MwlTaIm6f8YKWJ1uuHKAkarVzz3L56YCbqoIREKJ0ICXF4
6BriyrS7YpRJC5GMf82vK2lwEkp83Edswh+QWj+iXI865ZaRpKN33ShpF8F6//bJ
pfRsFTE59i4xuHh4kKlgmrhNSYCmwFh2jnAdZ96KfRcMYbRycM7lXOwyCZ9Xilaq
draIlvFNQ4zpOdJ6mx5mODZFo5+Vo/7AjqT7O7pUOYO1GdaVAWjLceSasaV7rxNs
pSU9Ht0frXkbn6z+kxbWnTkWem5MJGdr22aSHT22xIFvyYk43Ydt39doGYosxGMb
ouuTmTNrGG7sKOlmNLx7up1miA+fOPR/P37McjCP9xk5UMYIJm1C8+bjbr/A1L+I
JhFx240fSPmsHNSNx5iIDuYfiJd8XhtbmxLS61MmUGmEzilnfApCcGYwA3X/pUr8
GcWQjd9GOvMM1BL7BWB+lWK+AJk0VFmI+Ru3TWEE0aJKkdGYafmvTdcx19cWv28l
kz/pK0uqHLuiiw7BTd83VsgAMr1Gq8PUG2JNgQKxt6X8iK/kDbmBrHuI+zlWCeis
Se8Wbwxr7hUg2feb4tTjApqM/02fMn7S+nI/QeYJosBqS0N/4OD3WoHvtkngXzA/
EAWWP7T8NAr9jNHoU2jn2gfvloYWSjVnkKXzV8/HC2ahPLYFy5X7AoTpiwb4aB25
xpX1Q8emXp6n9PVLyV19kcUkGJI6Zu7cWRn5i4K1kvMWjc093+kECdiEgFpTS5Jv
LI1O7Dqds8d/NI2mVIsjxOn5okg4cqDNzMiJBQNdptK1csdi31tc76LmF7zwZR8p
rRuYtHu05KjJYFCWMiXX0bSNKqR4esMb2WTfQ8rHkKh96TzwXTeGV1fuTXF2gGkV
Mboba0/cGMXUpy5dV6wqN36eTmTAnquSLV1bLu3jUJkRG/fH5uBl2FOcdFg+YQDK
mo5cJ4Rj/PiOgA6ZTlh19X1bFMLnhw/InLe9lOw/CYZcrJ+VoDMUtQu+o4a7GBU9
jcdFdXwjIloOz4vn2qtw1+NfGkgR3WOFyhc5YnPstAwGszb/+/8RS1FMnRbio4AZ
IOGtrnGoQnmnPXDr4krDeYyJTkpFiW4KsnlM5pRz1cN1x15w5E8QBiIHu1xqtokc
3FleW3r0ohkqHl0bFYWiv3CHB+keDjIHs4HIZ2CrW6ovg9xBVCsAX5AazflH13q0
6O8gzIpkLwOwIuDsPbVhBh4hJu+sP3M/WxQ9vpyXgtJpX0cmBheu44rNI3gcZlnP
CNRdemhYzZe9YJ1hHZ0N8g7k58O4HdJ4L8Yb5TZvkPZBvy80UlrE4Qq4jRmkpu8c
gPTN4LYUo9HSev3y/8/elcxQ3cRBii/cPuc6lVBoJE32auOfOAj+phy6N+sgMm50
s88NK9WvopV8qCnTq0axbgtYBOniSmefRfvJHc/8H+7GZH4QdKe1yCDFS/plgdSL
5QKHQz6o3y3w3w2/nOI8+cMRv/zHCaxZLvFsTQ0JEN3oHa7QQENWsZl4DPWYPDfU
49snBPvntGxFBSKoX3lLcoldYCBfpStaQAzHxysSl8LvgjpC6b6uqDPNvxQd8NQ3
SZwKRD5E/6azMnvJX8JLkSp7sL607F21uAxnpmSCgg9X1VgS3JIoqjDAWSwnPBMM
mhxlokr9Pb+DzjaZvfKgRt8EjsWhFF5QIpvNcPGhXRcY2+kZ7FsBc+2dbl4ApS+7
OQQKGf7KEkn1nJVGg5VZ1FA6EjLLD3D1b5JizrAyIgPVaIF01d20f5Ds18tCRtrX
aL+le6N1JHjvNbQ4ElwvKgSuuazwXMxK4glJ7i9lCvdknUAqbKdbYa/KyDqLGSfo
jN6127wfh5NLUCZGdTWd7bBhucMkyyHc+n2ZyOBdrB6LzsxnUFG+jPVhg7CcRHe8
4jH4GgS2ETNB2Iu8vsoGbilfpt5a1KPC/DMn8EJIh3jRY1ecr8DbXA8DZmTqRXQa
3FZPpub+vD5JJ1S4dMLhHoTKZXDKtbS85JT+XrNslOtKF7Yek1322JqEu9nKutqa
SCdnNDVVEDtoZxeVseceiYmhPqL0wE9FfFYEJracOKXwoxXbgn2s5FfCpc+rugEt
GSj7Jq4p3pgvcU1STvSbfim2QhMo7upSIzRZrBr/Xb1MWJ5Impy4csbNWpmfrfqp
fmOs9v+L7bJgrummCC61zdIZddCcqBvmF2/SFFWYL3P89lfZDyzVg5+Y1Sxe9C67
WpJ7lVzNYSJAm2bfZoZBcu1R/pYmTxag6DIbboHBQ+8K97mdjUqdQBe3FE7KuVUx
soyprQTrlx7vfGUaNHAyCJq2MPa8y6dfESdmPSRWhnMs7kMIKiCYHhzntS451O9e
R67h3sFDColPE/8g1ymMZVHhobq5H9Ivk8fMbKVvVV7saaPwWV1mBHbMY3hWzYsX
np8R4dtsQBzUA6s1xAt5PuqFUkJHZmK0lVER1cSgFmJ0IEZ4ikuJh5VSLgkYc2UO
zHMZCTw2DGhBxek75pwL4XKNJwry/r8Qp0yLNlMee1KiJeuaPC1VIMPVzQ0NdgdI
kDneF+vV7LYwEfS4QsHwMjoSuinbq7i+bHY8dcyqPfqe60IFa9C6fB95Ig4Axopr
0Ykkn/WiuUGPGMsIXSdf2GJiIcMK2NG36jmmenD/yAEHUE7iZZj4J6iXyNgGEPqW
q830q6/lFouB5EdVAR2vqAgle+OChmSRtlDI9HwsUEPGh0iGEBPH60NF2/wD9HDL
YFk0EjD/zB2/Yhfm4lVCVl4WH3/V1SU707b7OgoIASbYXgFWkNLgrt2vp9scETVO
qg7FfKTXgdSlglNryl92+948ZixgxkKuqovXIIVjPBvWqSFA9jRgxpyb5aaIAVLi
1eGzF+qsG9VcfVMtHmAk/jw6/02l6CyZjVIClmP3Vw3b5FpCmFESLkZ1eBZ5cAK6
EiWLdqgLQJD2VkBZ52tu1XFmmlEV4V8oBr6Nz+bIixnvib0cDjCuKh+SbLov7KGk
12m7kSq7gCa6/E9MBzRJmmQ3HymEOcq+8eqzI/doIxtr2cwFP1+IwfLzQFJ/VEhu
iqGanLm9H6zX3j5UV/Ec8bFXN15q1LeCVKplH/dJhX/sMs+7uv/NunpXJFGSPJzR
D4D1cQZb+7Rv+6sqtFcrrNHAm9unK5nQzXjqN0zlTJZpnVtRgUsfcUNKn/qsk3Bx
NILIey+y9f5GdCADVA6qgteUN8Pgq+G6vX+R7MxzHYpQikmfOPLYUpox4bFGZPko
LdR70ZKm3z4N8lvEjx2igyHqYnY+o19UEEb3e5dycW3ZLgqVBbEn5T/10gK5OThK
wzPTnVfocjarTlrg2uyId2h/wP5QiBUVQzRd/h/cPHi3XgYcRHYbfcxQ9yfU5+uq
E9Dn8xCt2xcyUTGKlRibCJBJyRY4TcjiaGQtqABHmbtw4bUlSrI+nuvaoLEp9LJR
2T3ZQCZmDINlmmSfsEGHAwDYoEe7gC0lGvph5X6XmSRFE34YcXDzHyWvQYpBFYj1
XgaYjyDGXfqdPb5byutNMy4B2jWXoemlCp2gO8aKXtzK5PDBquEWPjaUhfYVECmC
LmSFTfMn6NOdmVLN9wivZ4N+N+jV+U5ceg9VwXDlHHCK73NBqxFU6WJBFROkCL6+
b42mIsquEXvdKXpYAua68YmmQB6eYB5+aumc8yihfgFgrplIhwox8NKF72I/vB/f
iP4DZAgw+T3JQhFdHPRmMOJ4hlqcpB9L6byvppVhb8I7oIrBV0Tlz2nLfI186FhT
lYnsPFQbKXNxBgPWHxUEOnBIN59hdFwzvFkSwjCYKGn23aezqRfXMAz2cZzSvUXf
Z4IiSG8tZkb4NTAUwhbnRGNttXI0MHemX/6A0J65TGjQp10Nqs+CMwkRxqzDcfqF
hmpK2DR1USZwlVxNKihw3K7RBsi8rU0CIwPMt/aZ5dV+m5N+wPYJwRh/WS2Wcl0s
bTUiHyivCZcIaNcEmqRxmgLu3jdGp/YmQO1op7b+eOIAE/W+pl9Ay0he5HZA7phr
XbKChaRBL6He05VsvMpt90nTJUaR8BwDykagO58pNvCEHCAPT5AGmeAnC5yEI/AN
k2hh3tDGPWWjugBXPEqyIXnUtTtWYNE40v3b1Ar39pHNoNPi1Fu2+8/jxispUCdi
Qos8jHqtLocJVIB/7Ue03NVeC5Yd6qa21Lnd5E3pSCdMj3uqhwl7LtOIbIgnLuPf
oc6iDrR2g6H9QHLj7CKS3h37vVfgPir0omYz86ZwsGprU1skZn4CWcbmUN8/y3pM
zNUdUvIxbT8magDa4s2Iq+uGHnoplyK9Yz7wHhcTrwcLqleUUsCyH6eLS/xleTLg
HFUn/WY9XJCdMcz7Laq5NVTCz693w/ajC17nMwGvq5Y0iSpoonOzHs3eo+x84HLF
i4pn2R/yfvipJZqa9RqM4R2SRLDckBj5cmp6EPyWLX+gVeV6LxLYiqBjSbN4RUHp
IzrsGjb2SZnjnDdWsKl2DA5dqJeSejwMsMYyLseZRKquwY2yHnPT+1x2T4KtAV89
EM5nuZaLOSkhpYA0QKXPEgtVZf3ESKhGNhnVnMj4p9FAY6e/zL7Mcb8bPiqfY/8j
sqB/jHWdc2PnLfwi9oXZtb5hwDGK7rmYz8R9gLha/lqNwWZhsmxTq1rDNmPqBEm7
rqKKqHO1ok12J0C9twX2znKUVNTABqqdCV6SAHtsdabP4Bc5/1VANQfUlKri/g0k
8y1FsdXLVZ70d9FMBhVr5zVkZ3zkmj01Nc9Psa3BaxlqP2lk7H9KuJVjOzEIn0sK
l9OVAuKMzrPwiDDHMHFTAdywIlQuNfX0g/0CkhzBLe/0dmhIdq+4pIPuon24sE7U
Isd4qvv/Sjds2e4tASjWq0kmwB61QfqZvHPMnyyhCC54fdGu1NPwVVCeq1YxGiVX
VvQXHKkn3eB9J+K8h/O9vOjKqv3pjJ77y1H5WQJGQWGw9kKrkMeYl+z93WmNNEGL
eGl8QT+9mGzPe38WjjlHT8sAME3fzEHw237fSHjBKY7MXcNuQoLEoxbY3rl6HdQU
VbAr9wbEQgFCrPOQWNC75sZygohqg7Vh52u08uDwwfptpP2stMgKq3G1hOtbXPpN
D3Mdr1TH+1s9fpFlQGeaayHtvz/mL3aN4hUB5X7P4Zk3EA1F4BdDWOUEkWgvJ27o
idf5F5fAMeNO51MWUKK0d2GS+k4BRat5x2Q1WT2vOsZ1C76cyrL/CUBeh8Vniyda
MM+ZLVTKrwTOa4OGUfDwAM2220P4zoWG6cSH2eVUHZDoYEO/7rcr2K69twyC3cgt
AK9iXl0iGAjmFCmZZypIkZVr8fOa4uvVv5vVQvuFmJPv4Une56MwLlhdeT5zy18P
mFdUoGsNhiiKDzEDCaIVgqR5B1mZvV9ucDkSvPjuKXC7jg1m2VMIM8T1Sag0XlwG
bY1CXxrHG0AaoOJ5JKAn0S+XIZeOczVa9Q1gy+YRUaAo6kp5q3N9R3kJR0IkWIy9
Zhqdcq0V5y4bjIu7d6OUJP9ajAWnysRvNqn2uSm4+FjBWNE3lPYj7SvRXlon94V2
EjWvMyPXw2jC80FbfYn8Ki88XoUMGzbaTNwuYfn7vNCI12xJpiXy8YJkNCF3BNv2
O4llXPi+o4DNRdG+lSB7P6ZjOhIl0/6/TI0O6yszOfAFx45YrEWji6dAdG5VqXX/
A6flAQ72EPJicLx3JNaXCygDzP89b0wlHO7Qsh7+yFtmc1Cc5QG3GVZGH3GO1BEc
QlCGpX0kxUaAzgtmhRIhb5laVeYOoSTNJ0E0GIB+lGt0GGfvSTAATA+S/rT7jMp8
asg0nfmqQTgXETaNYmpqECKpKeblv65MWn2Tir/lm5gSkvtPIrY8k6XV58g7YqOa
A+p4MDd1tqIfIG3vOHae92yDFwS6Gd8DRw3BgnHlzj3Za4SRgNc76JUn8H0+0AGB
EEDaAr5ioNoCh7WyXqqwE/ehun09bxlSDrhV42m1UqW3IMM72YT+jlnZTOTLLzfg
5h7wLb/aacQUwe0r+FpPVd1E1rlfncFF3ZWUfU4qQuXH1ajqkpMwzXmzM2xFk/v+
Xp9nq0RNqce730J97n62dWbIMI/d3sACjWR2rgXRmtSl92WRH1FRkTCiKGN5EIxE
zU3VHMwpzT0xvCJ20lkvEtvXq2yCHxhzJZYe8q8uL0tEUioERjI4VelqulvPsokS
+mY9M/Gw+3LhMnSRy9xS4tN1me+k8BrDpBoKh9/HC8DFKq4cjoOxWKXCT4h7eqrn
3Do7Yd1R3L+rkEAzjjXBIPz8Be2YEUeto/JkisQWMh6omBpSBoIstKoYPLpkwGLl
PeEBongkHh5sokuJaKALcgnch7gVuH96i2+uGnV/TsuYcyUB4QtnFKPlhmB5WfXN
iieoHAT6Hs+5b1ImmVhfsL/icMMyV4wztlhk0U7neuGcK3CqtwhQT17LrxYX4jLz
0dVMR9d3vHT7FJDJJsyRaCFgdQdvGgHZnXlcb8jHzJeE6sCf6GLjdCWOu36qspnk
SRJpFwjNz5vsQLo1wPgLCRZlnc5Pt3awVEUPsfvla+yn6IIazJqDkFYrO+sN5BLY
Dtr3ZzWNpTsCpss0EUmAddwW2v2dRrQ6r+w7R5PhFCUFqNPSdvWFFNPfrdo4HPUt
X71b6AUPwBlEB+yMMcBShB4wXI1V/w6pUuYc9XAHHl2btagYrXfrrfcJjFN9/mdx
0OY7QWChdaUnK0wu/dPGVX5yNR2QwYFOx5UBXMI1DSiBCmWI3X8FHCDC7i8JtWGf
7f/u1BxfpssOnYewacyGg2oG1IObUJmNe4O68Z0Ls6apCLnqjCXbd6/+x7r+LA21
3NM96RlesskRjNVrS2d6uRRPDuVvz4d/mXifneVTFJweD0jcTj1RWDTF2V87aKZa
p+oRbhZHS9heTVKeJ9SE77HIC6uPkkCjr3kQZBndh9AU03fUhT6NT9HJbPXKOqsV
lBA4utchfxIrrUbnR4/jPfHG2N0MjV9jiI7N+HVXRkl99O9hy21D85lCGDMWP4f5
8o/NT7Zxw3w/mapLzVvqlEwN9mtnvpoi8qVTMr6p5re2SLsoiS1NiAdZuEKTuR/X
L4gczF2jpOQs5wgxjnxgG0OgLTnDKcBYhVQXu1/9tgi6luzg5HCVqzp/hxw0nv1I
5eFoxfXLhrbee4qIBxkVG8I+oc3iyXCwVXFhqUhL7zWbzXZH5NgnZkllO2YPeFU+
dusmZMvqvGrPVwxM+3CekeNPzYBOHDkBlr5SB2xf37T0oaOc3z46Bt/DLglYyEHI
Qtl9aWLoZ81rZwXufYsanq5qdRYUaE3WtOaR/VFA96I9J7kIvKisL1ufcCmy1nKg
6ZGl+UHbwEE0tAuZtzFmidlk46dOXoFbw6vwEspFnTw5/Pkhalqe2OpLh7fJFZ5d
A+mdqJL3VZGX74sKCAmdj993TC4J4ci9yQ5Q4Wx2LoAzHdD0b67dYznvUDMS22d4
LnRHpDQTr9YGzsfUWs1qtIdccB0am5ZlUjFfJg63wXeF8aYZQ6369QP6RnW+0ciI
iA6mgLk2Pv9m9HDmQE5TDQ1yG2xNP7+1J9omB0K7a5HMLbVch0a/+V3Q7v9sAtK8
eQ05tGCo4mIOsiyaH2U9jdrrjvFdoKjYl32gOoQkodPKkLPZdyggbp849patZN5A
fTP5Zu3+MnZlM9VSdz9TDIzQIkGlqzje44elsKPpTJ0OKTeBe682aJRVbaakuJJl
CrbHkD3RJoXG+DhFn8HFT4g7YCNJxIx7a2hfQfZ2Ep6hOqluo09WJN/cMrZutz59
ZOnwFJ0JochR2+9ChTFr/s8nEpuih1tfOws7StgVuENRI01dNKXZZpxSCvIxE/jk
eU3kQea5vA4RAOZodaIsbx5kEsnstcSknMWap/3iw1J/LmWn9g/prF6JpwpcZur5
KGU7SmPba7Tnc6h33pPlP+7+AlGsrmN7aSmsHl/qFujYs+/4RW7xNulNb5w6VAYs
L6bv1D/t/1TxX5+jfBvVo0tLWXBraIemOamFxmY7VCMs5M5vHHjPtf23mi6sWc2Y
bGjGIWm449gtyGs0LUst1hHfGawoz182YQrQFC41+MfYloUhp9znIIJTl9ir6Ag3
2XTtiXVHMpCIJPf4z9KvXJrhGCpjk5CLOAlNhkjhdc/GD18WInFnRGuhw6lhnwg2
rDRH/ZXO3legZyclwlSIhaFr8fMWFBGnq5WZ7uaHdWc5rCI4q3w3qyE82fN8GR5d
Dk9D+4f72ZIFxoayjTDaw/dZHhRy8fRR72aJ2v0VBEmi27mmTEbOS449zs7I5f+B
G2soSYbZcpOW2C2Tnb8U1Po6yWhnp6Q8DVB3IxpF1O6IIseAZKbhIl97BpzmJRvc
hdveWpFEaKYu589x6a/KFiX74KmZyAbXXMCMlg8berM6hbwaU3FdwBDXFkkgFH5s
gXy2byvwpU3Nn4zTLsDAfch5vLM5GI7mn2zjYvheR8x5QlqsA5jgDNTGI4fTP/uU
lOR6TU2N4a5esDpe4+fiBBwMm4Qsb6rtbP+9fPEIBZbCBqJ/acyrrGKR50C/sg6V
lK3DymmluyHlIGaRY2Aj5KuNgqfQBQB77bJKRQMtTbIdJMd0TdOx1jxbdVC6FcGz
Okx0y+HWpwnKCXIZGrKaWuh+5iE7nOBMmNT9kfR5uHJfobhTD4jYYaP5vBCtpx+7
LICbkf7ZLcFi3NizqZZFfd/vyISs1W9rdlRO5/pvm5/vW/ijPjUXxgQ/pDV/zZxo
yjKdJz2UDIyReIjdm1QdWJFRWsHqW/hQ+ksUlFHQ9ki6R/p7wqUKrnYobGiCsXL5
SHiGWyUW3v4GRJU3McpYqyaDR4ad1+T5KtRFP11eIDm/Si+WywfIoi9n8v641rHj
hgf+exHd5R8ZJgIyzKzu7BgAA++h9d4IPGQost77bfTLptiNJl3atGTSKpnpFcgg
QE27vW80w4IHw+FeHaodxqUuY1b43l5FRHLOrgNe6sXpUtWBWbp4nj3YZUcnX6Vf
ONdtK9nspH1MpSvHtH9ETrXjcwuNAjJNkgX1Hh6EJsOM5LAT/PM0pM4oGoQ2H9Eq
tad2U9NEiFL4G6XF9AUVQsIlvL70ga56zPAVfy/djSjhpmE87TUR5Go4Fx/Wk0ih
GH4HTP8rWz/T4D0ueP6e7ZBdYaMPt3EZok0TGT/KGCno8AFCIEsjEbDU9AjP1eGX
hV7/Keqw3PFahmIylbWQ5Fy7zVMbbaYSN+S0nNe19VfPUp6070JPwIA87atE5e+D
n9TJckFapqvTYm5mMiRbi8RwrhDhBB38Hm1gLsRV7Se3sOlRTc1Z4D0ye/H4rZ6O
J8kYICs2uCmkxbNJS/7C0e8XO7q1CPaTkoDdJbcsc4r53iyCO8vRO/Z5AY3qNu02
SaIztIb5WPA+2/nhDkbe6zOl/jxjwz+FrkCI23SG7f+rwvfHpZ/LaVtI3aKAtEIb
dcEva+t7OGqOuLWSsvCdDn6OLtRhGSBh1wPQWBjW+MUvXsEY9nrSEgqyOxqRyB4e
dOI856M2T8ynv8qh+aE7S6XC6fYSufKn2OeRwGcdzVUtr67bhg7gbdRXHT82GcB6
V2tsKJSUxdUuxzrX92u4ZHlxsxv28e1M6nLACkq48XMn6+UPe+2hf899jDm73Hlj
rXd97po44H4X1Mz/IpkzhoEsHITuXR8qhaTGG/JmmXQr99gvoD6cOskTLuSXxyU5
FARSCKXSQiBc8C54KO2a4XYaRALqwoqNmDwlDPwj/fF1Q3I88knwBcqPSaT7zGAL
phFdDGJqXHFvXg5OdJJjFF4lb+gpx+F0mPaAI2pa49kbxKCgSfFp/kNpfZTDwJLr
wVLZ8yvvZSvdZ+Wwx6tiiT9DJzb0+H8M7mm36MH7vD0lYlkLA4MD1ybAVO4D+I86
HZ9+hhSvxctSATbpGTEW0FfhCs9eRyqkv0aQIEutnM4LIdUxRfzl+okqea8K9qIQ
P/6aZDfIlHF5y14kRcI3nKT7w0AhpHmnAZ0RS+/gKgyWYQnX/bUsasS1/5W+Y+h/
FY/h0+g3/DyY4lFR278KOJBZ400EY1pda5a+7BH+n/GTMTqeuzaEgGn40ctlJe7k
uaCvMPMY2EGUBSliq0tyo5NJ0XG/oN2ifYSeX3Gpe0tCtsxp2pH17UqvxPHi6s6H
N2+WHh5vfII/15i4YXWRcIRNZktanmF57Su0cfam5tgHQnhEhETOFNGSPrtJSxjk
oHgDggMPOIW4Qt08ymmUcWl8fUCG5eGpWGl8DX1E0eZF7srSUmwLk/O2qahzmJHo
AmYBKJDfm+LueuJXZ/WnQqlJxELvythD/d4YRuNBwp5haltydbj/ykLuv3AT8TMN
jZ4daY22Z5ytPWXmW6qZKuzahhYKZpHAdfmA1pMeudqLwhIk0n/TAAVzNgqd+YE8
mH8p4riM4ZNu+G2106JDyequmSSw9bSLxQ2t+45X0AgDjh6qNq35fdGttcPJl+jO
ibEnrosBY0tffE8E6Q6yyXQ6W1vsK+pILakrrSQdhptiKuQAFJHVsED4ky17Yz4U
yyyokHS7HyWZ3z3PFwfa7QF7UzUx6j0oXaZim9c8W6mkCbP0G23kT08Q1OcnvvVJ
mYeI+EDLJLHcIySTFXGLYu6NOj/QhO7FmJWgP/2TFLKuESuhJZZDcrucjrO7p6EU
mYYXIrCh6+juUEYqV/i81n+F7aauJY+X8ESXkO7pK03whLCI9Xp6k6jMCRJhnxLn
u55ZR03GnquXJNk9//N0kqgNgv17Gt9U9zd3PDp0vOXBDkZspSuslq62IVeMQE8N
B8nvOqFYPHmyRfoewh0WwG0ndTCBX9WNP8GYheCGNyyuRznFIYT+HIO5Fb/Y6B9g
zQJl7rf8uM45eca4wWiVHwncWzzNO3Sccsef620u9GP3UAaYFsmHtgySIRxqM44y
t6ooSvq9mYWPndNiRGF2LFnu0rKuTjU1DcuwBDmWs4F0GxP0UnPW/CD8+JxAMcnz
pbLqST/aNGkrGRl7yVdtzLAIyOTj/jQQ3tUQ+iHiqk+42YI+5xurTara4kGcv8aD
P/88G/Lsgg+qoMoPuc+1zvUMXLphsPUe4CMNZ3pa15NzIMXvE1qhGfnBaUkBcMtC
22KlQgnfKP4JicUegquyXTVmwe2SnHLBpfgNODPABv3jnt2xtBIebM4BdIPEDzqy
8zJ8M1PrjJ+Yo26klDPuit25p8G0CvrqfzKNLhtfdk3tY/gtBaPa3tcWkL4WN8k4
4/WWI2YupYxZRO8JCKnwnX7/hKMAbrIRzU5jh1Hy1UHzU21KJMXgslo3KPiTEU9U
fLIDCQmtXdbk8IVClRqQRQ7E4ExppjLKY4Z6cx4oOfH/46OEDtyzekT1JvTmY28K
H13F9pIU0SoxBWz6ZXeRvfhDMJWGZov3ekq6bcPz2aKfJKW4DWjlKGqH6vP/2S9u
AF0BJtSBTgT1ViysZH0mJ5f4rGzlJOFL4h9rwRpN7lwSJc7PG5O/U0eoGU64cDM+
CE8KGLK5kBE8Q4qMOHscpgydABW8mYvw0mCCSsapAxUb3Ma6y2pgtOyje2NDdDGc
IOLkCE+dw1H5EUcDBZfuujodQ2U/P9y4jyq7VEFfG9/0gQ/B37o31o9em3rA81o5
RIhReZtH0MLoRKCJm4rvvNDCFcJH2IQx55Z7gfazC4wpGBRvndnE3FRgRzYzcVrP
yWagkFS7fI8VWBmNdiOJnF8AnNaKJA6WEapbLwBpTGzWpQ6Lk79Yj544zHhRa74w
se7FujRiTDzUOW9ICwXG+Z8WNUazMWYSr2KOoFrIurw6izvcsK2re0C9HOp0hkHO
vNDfpmSPMV6D58r/+sdt6hfeW0iiBx+pK23DM3jNZ1NM1nPctX5jwNK5dOK4xaQV
Rkqv4n1wSoSnwI3yLoO74NwELWUX3jLd5KMRfnMeFA+jCAYRtZ63KpFhUfii2uwv
bSTCoWWdTthSTHcmu0YSHUOsuLIS4HVAo0xVL904oI/aYiOpMnlXFOlkSFlD7WPt
hv9j8FKfM0oVH0iXrvb7bj13UDSpQCYHAwJDj7fC9wmWuZCzO40nOkXDJHRqGAa3
VRaRGfSrUecCSVN4czRHVcNDna4qqWjcuoKvj4OKhazuSC1tjj78lHEFB4Vgnv1Q
dLgb5jTryaMy0zmR1suEm9NtN8gb0uTUMf1rmWZfuL7cLnLfE/BGfj7pnYJXS6NG
9R008tEoukVDSZWMocuoZCjrG/wwuC3o4GMwgQNN6JVlbCvztVLoTc2Xoc52NKXA
iBZbRsKCzjx3/UpM6ya5yOXhl8QRiVLpwXWL2vLxGA26/ppzFQ44nuAVBNTrc21R
OiN/NQGZle6lmaxCy8+QpwSAiZ0XUXIjYuAGPkAWylPOlJB3OU6Jd0NKHoHS4Qae
sIwo7Sh+MFH0Thwbh2uXFprJ0FuuaWRL6hRN7oD1mVwrnXzEdIv4PIQ9wNiv7Gyj
xJ9+//3c/ALxufSvPnL1LqM6GgnKXnbtBz3pEQPm+Ap4XXroowmFvgfdiW7RG54Y
KG49kcWNlYOPa77VxRl66BiHezJPl2Ib8//cSDzm7KP3bm4P0VVvxZ7RE8JrTNqp
rMye7LZV1BjKIGc83tSgvIDILzuJ4GAIumhcS+HqTyc1f0CHsasEQ3ws99rjrREC
8nNGHBVRHTlYay5cbbJ+gMiHbwkFC3xh3YItcCnxde/78aaCyX+kE4GqH1kSpBxF
DR43d770yxUMSX2Qp+h4u54Zt+yzVOaPQol5ur1oT6Vnnh72wMDjfgwWbgfFFTYc
eiNTXxvWKOc1GfSFaSKW7NrHBPFDFEQa+69SWnI6VPNH9j+vSJxGGTpb6Q7I5oGK
HiuOtBYPSNKObiMdi+J3xyKCG++8fkZyJ9IknLRutU0jTk6S1/j7lIHMF6KdGWLZ
LM2eNMQjiB5xtKhcEhUlz0rKE0i0kwYWC3HfdjloDb0zgcrY/5nLNyUVajS655qK
jiwH6RTt6kEuyKJv8a8WLr4tCTCC/WVtpQqmKySb5c79M6LPBhE9ar+JhN1QW2Fs
TcuIzWbVUEYtmYb5DODU+7ItrRbdGQT7et2ezb+5bZvu/UwBEpgveyrbsOvEvo5L
6qVYO9h6kWV3MRHwUcTFL/hkV2t5VckcvC7u4I7iqzk8rdeVJFRtsK83RS2SeQxd
HpY3Jc5PrDa3y039CO/qO5pvijaYXPJOUHMRjqw6H+/T2ROc/wNsSpvkgSPwPR4H
x8wZEKElVOaij91CKu8DDk8PzQdOPJTHjJuj0ZC5SUulNDjcbCjhn/cnsIos4VEp
kDJFxyfdESM8RV0xgwuAIMoERBU+7Ptgku53jHe+wNRaYWd/Ui3hGiLlx8qmZTlb
7aYZC9aZLYNuHXfRIshwiVKy017ADQLE2li6AXw2/n1luVoZh7KAp/RaCQykMPa8
bd95Y907uSIIPg7WxarcilyjcqJzbZjaKliH8lmEbSMl3YWinWiEsjPeoiyuAd2/
LZuwDO4NINCU1ULCf2UwWnRNbxJtrAr6XqqRqgnxeCf7gZ0Vznomo+NRzXsH82To
UtKzp4D4PZiyJytUpMQPWjvoI8Rbb93Lf6iEYChWH0xpX/OF/RoqpoQ7kWNnrzLP
CFpEtwK02j7ff/T7AZU2SYts/hy/ieICP6wYAkkAQUc2goeP0Z9TaAu2syQTqP5G
xu33U5xCB1vSDQBBpfFsdXDRiO6fj30BghyCqNayWxXdAPv1LjaLPMSzCSiQq9YS
H7GRdd5q4aO8NAWFoxGUuRD86mfC4tsHm6Q3SebK8GOmVt7HL9eILoZYuiTo0Apy
PCxSr2GodTorwcd4819gNbDwdCUv9FS4YhWJMj0CoIIbfoMMHt6HAOBtjPOyRkyX
gSn3nPA4liPHmh4Z6yGRWlYOepGvK/8fnYHNWmMdQwdp1I6QrJu9QRqeiPunWinn
UfxBWtY/VJQOpbtDtYJ6Y3K8g3MiVW2YOCOTOYQ1CEl/83m/U9gveePcWjTAiKus
lTv8zxjKxCm0jhJtHZ5ZbTyK4crH3BIrmr3ESqVBgQ+i+IjEy2Ubp3V3Uym4VpsI
hCwurHhbLRkHF1Ygq1i5/0W4HSPayZSRIDyGf1zO5E8jZQQqTWepPiNdNuxk3K9O
jMfw51x5GjZrUMWNcNIEaPUecVjZRrXFGrnC6rOMMv1Uy1Ws/rj+Redma3UfR6Tv
novFlQcyGNxZNxrtuqrjS7uuNgg/LM0FJs8ouV1tXTuc+8D9JC20K+WEASG+J8bE
lr9mpNpa4XLPTR7WK0DeGvubXdNYBwJwxnv5desZxQn2KKAdsXV86QSZ3XxJc5cL
yfARqRxXnu4KZmZIeTbPxFPmUHAeb2Yr5suK7dQYYwcRLjBDZ/frpaL5rcpAx0nJ
S1Mrfa6CI9Vena9p9gQ+mAAe2EWacn7ao1kIfN2Ge5tTp4ALta1rPgU2PqY6pJjM
3R+iegjrghheuYiBjFQK6YGXUBxNgvh8R/8i7VyWTmOT/f+YysIIq54fdEjGUKK8
mCBqYoj1g/sLiFE7EAuXnpQYldAmswR2hrutjfDiDVvWFNpt/ARh/FtFRmUaSbX3
FSIwvvi6PQ+efxuGtD3B7I4NTJkFLhYU1E/6FbsG2hiPHrGe8Zp1+/MITivBXlCl
lPeUyDQSdbQAQOX6SSajKc1HCknqSLQbeETJnaOETqYFBFogIKo998ZWMRSY7BDN
brqDREvnm6kwLk0LQyH8D4XjJd1PqP44HucL/oXX5o/XjJGuZS9L+gF5aSzE8FXi
DH3wmyJftJJUTucNhcIlVYYwlCfnhesIMESeqzCmTMWZdqUhhdg7cenrKthaTK9k
5K60I2JtoDzVHTutQCO2zLLckfUwi57pVeiOj49IpIG/9mLVK/fxliSpvqU5u/bC
7tzo8KNY0I+E1niNsH0aSwyjRsKsszVk103kG/TvaJfJvAOhARJSEdKR9/zHgv6A
dmCNoc1l5oa15Rk+GaGUh2ySgksFyJsjkLM/0ExAkTtCH0dUBUPC9Z9hLu3LRLmW
TvU+udBRuIaZAT+K0KGemNmMk+MPC19LrRVdHyha56RbP2Y5STeiiReBDvagG96P
KP/qMx07YKImqoih32QuvsE2GgRS+cjqus/56P2ReNIqxs1iAYMpYaMcnkkAxRmg
t5JxpFaW1MbWlTI0Hwxa6gg2wnFZUYCC99emotg8rpro78DTQhf/Ky4nuoIXqgyH
UbEHbqnG4JHPAndd2hHMTKjti4KNi51HFBdbWhb4ztXDq/pqFtmqMNAconA6LwTL
+KYXj9q1DzXGC9BtdwVXLXn8SvVb/CR/ztySR4pQ6OBqHK7DtAegpXP6/p36mmcu
WDrGXlB6CB+AUrnr4h9rZlmpp0/BMqzTnPkmkqJlmF1K1d9m2xxq759xeF7xgVre
4hPQDutC1p4S34EtMkWBdYpxbl8NE5Yirp+U63iG3QQMTq4M6clgFr1QYPRbYWdU
3vJnBl86BMJqCEMDb4RYa96iEEzWKjM2CEB8bluaM51/PRLFKxccyqkDGIjhn2la
STZk9nRvn4sk86gt/lorCeKaPdRJT9M8UQk+9XZs7i58pZgxFEU2atCnSC/RVY/Q
vFynkFshWT677+ZGrCYkdejMUk+qynbfzvBR7AdkOi3sB0waKWN/G+GpTSzMhh6s
s+eJh0Ne2fXrqDF7Mm7Ym0Jd8IVyg2JyD/WTH2UDBlDYP3cFy9Wc0n9ZjEv+Swu7
Mj5ySSTqCE2FTJIWVIHDPsAa/qtvbPuCJKmfzC/7tkiG5n52ZytZ0TYn4Qyuevlm
HQnuOJiKnTAozM0IxHQVd1FIBXlZWzd373FuIswIrPsKrkJGefwauj4e6zwK44hX
CVXx5geI9UXOO7HDCK6NAZ5maROv0YnvGM+PA3N6doNrmej/5+b+vNngkMSnzNFz
uvirzPHEOW+xEzlpx9uzKVVLJLrBdDJIFJgjdB/NmPBRHXIxC1VLJfxZQEBVHaR5
Fp8jK3DRHiLPn+rJvc1W+KAQFF9KJE9qfErP6J9B8hPLRJNskOIsuX53JCLwRmfB
fOwxL9CrVcX9ugG6bmpvqNSnF8r+OwHZXS16kF7BVdM4Da0gT8DEMiAdAj7HkPQj
eXVqUuuhn2TW25+037BMfhcR8Uk+b0iwr1Svr8Flw0injRuQyf54g7ykd+jmhzgF
YC3pEhTYcTuEZU2N+uMu1xcNOEemYbZdlJihHMUUvMeO43i0+oeHSewUSBQyhpOu
6We7VD6J27ssu1eAfSvPSyq5qvebrXFQhqHLoDlQ2y2vrbDiYabczKYe8n1muCr/
WmATY4ZysiQui1xxFGQtb+KvMLu8BR4EW4Eguh+me0dSLwmr1tHxFF1hgPWZhYRD
9KH8MdghSR/+X5GmduMs6EplPD+wJo59Z1GEu8F0nGZMiiKRd145s1/04cy779L8
XcIzi/ZUrlQeerVE+eKJhGenwGF8wDqxKkhOWiMFPTU72b5Jyn7+INMS/8sNUR03
GSs6QqQmqmtRvNHdB0oM8s5MPAkoBa5DuKImMMr1inrUQeAEfIKblt0kcgx+2Yjz
h53gINwzm4QAeCZaI4k413zKU5oJr0+JEfy2is/U5ZFzxyrBWzt4sfQs21DhbGen
RoWCkbVw2FDyJKIv6E6dJfmTuQdEUIN9YZCaI+IsehW47Wgyq/F6GF8CvUUTpdCl
CGFDoMYM/L1frdz5ilupNDT7+nrZhJ3LA+p74F1PPdPgfbEv3NF3VzjkAm+9HLVp
IIq/yI9xE0koWJOVW72xN+N2X+C8FJxQ9bNMmlisGFnayfRT+IEJ1hIXygjFerCk
mIjb6B6e1zJTni2t8WjNb9a97pko0PuEiagKRgSglSUPzMp9pVLv9lwabdGgcnDP
EIp8ppLoNLcFQFY0aD2vwckpX004dVqHpIS9rt3+6q7AJLNoZkLQZDIkmSlO1bq1
G4yT6eggnZIPDo6mV0nOjw+8DCDii3P341Eaa2tc7gQB96BO+lbz/LCKmSLyTCGf
3aTOuhi3iRbW/9lZQ9ATqEVJsd43MDx9efCl/K/gIybarx+mOzBCR2ltA5gdpOFM
aw78nNrLDJBKnUUMnWzfNapmfTVtNK+KrCmZxD9f1IFvo6isoMtuXH9vAwEtRCnB
uxT4I8g4Y2eGH1uQBw1rqcUk1RfgoazD0Cqu+Zge8ri0sOKTuVfVL9T9KHDvoUEe
IsGegFEgXJcP59qqg4T7WvkVoH47X9H8hX6MbnC68fF6O20NJMx28McQ91O9jzYf
4eRg8Iqje29JWd0Vl8nxq+lZBKzB2A0skzxdUEfoZoDDcjD2l8yHyoU4HvOVDwxQ
Aj2/eVdbI9nNdy7msALpcdyQISPv/Ditwndc6gJjRxrF4gucrY8hW3NWSwzlTYj4
2FrV67FpenjtXOI2FMlYUW2AxihPW+VxKzJcyxaMnADW5uDuOTi4fT7ED6QBib9G
lvIReSFq7iePWyPaWiXbsGObM2n1wbKonJmT4SOWhHMTLatr7bVqsKP4RugFDtXQ
SEZImr4amoY2lAggsegCky7RK2OqE6NSRV0icofVEz3N9R0tcqoom/H/otjmrl8M
AMFAWeHNa/1e3j0HzvatDG7l6GShidC/gzwXGtbeAUV0YjND1r5B3hudS7ATsLCH
gOgKDNwOxYM6CmZxhnSyIOu3/pez/u+CaEe1w+T8BGLNkd6mHp6GZsGf/meK2VB4
NQ4txPhLRkyVxASOP1aJl6i1+R/ZzG+m1H/XfmaicgiqxhNNgdH+OrWDpda2i/ES
8VoPKQb3Z48b39wfH1YxXpXewftZJneT13v5EOfZGRhmaUgxwe210UT0ctoxQ2Sj
JCkOZjEvhPNUMVe9ZVd0K4RKF5csfQaVcpzXGtrwMjQ+57aT0Hgk3QV9/Z4NRq0v
506OV9t075jcVH70g3911Mef7ehqG+ax1eLsfZC2Tia1qzM/gyHoI17fLA2ED2HO
qyVnui2WBO0Bqwmjh9nVO7106VlUbbqA9bDOhbURLaHeByosU3sUCSb+DkntDbAm
VRlb8rKFuwKMj0Q4BQzHGjIWo2qpjohS94XeOsr3Gmo/BJA4aaHEq1MUMuP2cd7c
uuaCgaOWYBTaSzIlHzlIXBW45pWfk2E5jM4/jsr4V/QfWKyeq49uCnaXnwYF+RfC
8HjLYLZde8qD6vILoP/VV9E20maR/9wYIpdW3yhXj3dwKNvAPkGnzO8Vb2P2zrO2
wVSyTa8yvburlfBispMJL1QmXikgVo3N/jiW/lXKf70YKIjWqbQ0KvnF/+T/sMoq
mXY06ZYrb5Nzrv1Vx+PyYjCgLifP5Ti5Ntc2MhQhu2cWybFcg45RHBYQDXbdh3p8
ex4XUmrT5cQw9EEz1sinV0h+NXRkTxg3RCGFZlQWCQ5gAo/iY+cvaU2MUWNMLHEb
cT5fzHkQWNwA5xGaEmaiffrhh/WUC2fTZOFt0zmVIcGifLIbx/b4zWlW9TJ1VDWC
dvO/DmngtSOTd0hQHe45ShneLKTs13aOp1QB4pVgo/q1g2b7A6/cKA2VGAEvq7sL
6so0P9AiasyiOVRPQSKtSVL4b2XadE0aBCR/7A1rLEoxVwCfYgL+7R43tHWdgbUc
fLRDPTxCxwAGWNN4BCMxL8NWeMSPRbD29L5YxhDc3Jg3H1aofnZRwK2mWjBHDpKS
bLPNpS1yCgafydtTEua6luz5C/1yMNd4vXbJs4ZUtrXvPNkql7ZTpmJiZE/8EQhg
LQmGV9oy4qYnf/QaNIFSfgIhvRgzN8r5jcDq5YRtf8PkGg1o/Os45/f0Bvq3tGWH
AqMiGzxqzBcjoXpW08ZTu+nzFYDGxyD37NZJS4f1GnSOpMa9lWn0w4osQ9YQ4XDM
1SyeFD21dOrbFOrukquN/FtRq/TMQ8rD+S/nNgOzHUgpZ5sxiQK06WXgMMpRiEqX
JAulpn/5YpaDgEw+lJy+uKNmPV94EP8HWyDrLxfHxqMtR5ryKUAzWRe4J7E/TidO
CFboyYiquP+jfVTH7OFO6sOcaZEYEPTDaK14KnB2gUztu6SFfSTu52E3P4GQZvpB
qsKw75TIQIi8U6A2QKy3QmxT8tTjWnHOUcLZcq0QdweugbEG1FWYqVY8RHHMEujS
hLjWMzaF1FLIibStN7SKdQW2XzKh9o7eSaZCC9pcv5FI0/WoIx5fOuV7NwIipA3m
xRxw/K9ZAhhjXoDieqTGmrTr1pQy9Lb5oEmA4OBKBr9JZSBu8+cAu/DkiyugJttM
KdLVD4B7euRt8m+GW5fItXb2dH4w9jDTjo6Q53F3O4r+30+bjucV4jvLc/nc3Q0Q
cqk/uycTZcwdGfKiGSVORuIaIZFjP9WhAYDU4DFmMdfVY0DV1hl0NmvF9qa8Se7b
g11alaWtzSm/cwGXYmpb54HGB0Ltgt4TBEwsURKMMYa3nQ8GFajOZ6spjT85Tkql
5CiOWwQCPrwReY/bg4S3aTrif+tYrDAUIJksbcR14nVmH6JH82C7ACiLtnOTy+tn
T15Cq3xI68+OZhCzQndpjOnAZ1Pe3uZ+jANk7mb03HRb97ygSiw6esXY+NzaTvbi
emT+W9nDgofjL35UPgSa/cKT9yvPb+P7gzhDOm3XDjUY9EzvRHQ2ZW5DK8ndCw0a
s51h40M+L/2czFml3UTgfhsL10GRqDnS+Ve0M4zcUhokQW7S8QGQJGHvFQweZ4ue
xmpfsDiRIb07QF1lfxnfQorbo7BIV3OkVsZn5NDSVF59ZxOOXfc1dANGR660FVOI
mNCAfALBWQRLxJRjsf6mhvkDU/6J8+CZCNpeGB6dxJdSxPfkaDqMG7BL0lAzD39u
ETQgooRq2yNz4MlrHimxChVRb1eNP0x+TpM3wmzCGoOEcSej/tmtIfXLChk2HXe7
BgPwSTcWc8gPfxJnZq5r5XHkJTZDbwhSQXE8I6qABbkiVKmpqFJRO0TcSHsBCjdy
8R1jzXGlM9jqDe1L55TEJRqTOHk8LJvO+lO02iZIIUoJXyi28RYv+p2fOt0GLm7T
Vtqu8zh3nzaxXRc1SplsMuyuuzNAkadLkMLUbvFq7uFJt42BbZ0/pdmEyPw6Fcvv
hA4eXLrb+nBqsyEcShqk7w6mjUNM8NComJhKo4kc83WpqK1S2EsuaK1gngZwPP/z
6PEFfRMUX9jdRQv81wQdd0na037Ck0enUL8xNjkv5vZlQLpQQ0Eud6I2uDIw/eb/
bMUq7tUOwpqaGY8dXXRk+1vj1yFCPpmrCCtm/iFl5RKr76epCvZSWLUgsDdM1vPv
NK1bMTrL7njy5BkXn3+Vwd+OotZnQDaC03PGpQFD4hyTwc9qrwM/UNCSWRNCivwq
vghjb2edDDLGBCJbJ9sRs+kvPnPck2UdToQNQwWgIfR47UH8097pxP0XCXFJxjYZ
dTdO/52ENNa0dqJhY+qqF0Zvuzy+Pcv1UfigGlEifWwHTZZZSR/gNYSo3ZbF1CPa
rC63aa/B4h1xETGIL//94CV1E2mLnImrzk5wGGHic/cpsT1vVCixhSGzp1N4njdX
o58wreA18t3WgVOkO4Y9duK4pEjL3faWuMH2zc6Jb1nBq+SShYP6ePU1aFoSDjj0
aRn5X77Ve4bK8lNv7/KoY6o09U0L/zM1ZVBfosbijXHehL8lg11T2yCnjeGcLpP9
nimdnBHiFsc3y/ksjVSvpRn1hoeXBOg3Ic3fTxJYe8rcV2me5eSIHyuZgxGzcBL7
1XGd0/hvVT0TuSzmY4zMO/ICTSUTZMMcT0aicEmZZAStYFLzFBisyQyJ227/zAqG
SjiraaAmVNyaed+zpd4tHY83A0kVR30whFBiPuFAvc0QTwFbdXymkxSJXFjsyspJ
IiwxuWeENFXofMzAHrWX2MBSstPfy5t1c1kofX9G4CnZz6n1Fy6bMyLDHErPaTOJ
rQX+dFgGOALSQF1rFKYS0ugVdXiU7mj/xwty6EA2Pyhx95lL68McBm020n/eb7hx
rNE9LgruvuWJp8ca702f5F2kzTIBOLKfJVpf9eZ/SUA6eSfoPQq6U4llJ4G26SC3
13N50bjwMEzy+2Ly9K5a5KUY67xKhEufXS2ewwFJX1P5FHjuti+ri6WJYePz+S0S
0Kz6Fm0TUQeWtsiRQE2xQqAPPeGRjCbkZ+tOnaOSaj45hReRjB8Vakq3hXr1x6LE
IO+SO8MobduBsslds8uftvRou2HEuU7+LTqVTqWfOTPXpCjR2ULH1oGqV91i0LId
fRngGFQJzT0qmeOqK2GLetDJsgT5++yQKv3eD7W1AzYe9v5ZkOQozpQg+t476Y3d
VnAPInXbLk2eP45/egVof8qO2C0fNHIb5e39dFifndnz+uywn3xtOKUlMTU1swXe
7BwGylt/0tPG1GzrIVFVbt/m4EcS1pWe7KM00QufcxeYR3gQZ3RBg2IJOeo8AES4
eVBII6d54WDNzVaG2YrJDnagaaVl+b0xmZDMowl9EESif9tqsJiGAT9eLSlYGgHs
ViJYWEx9ULmHjoCmYwsk4yUBHFjtpxQdDCxOch5wqtVwMiEEkMFEog650O4cx4LO
eJBPziBAS6g4BFKqfF8T6fv5EaEdTGGAaQfhGJh59/hIVOIRvzqwpqwkF1JnKLBJ
vhBytSyeouo7UteAvq4RKSJN/kcw78SKayMIl0SnVM8zLrkdW9LJiWHOosVyEM23
bTn+aZTLBPqDTzMJ1cfAYFBlcOKlDCcdvg5hnRbtZL6XM+S26n1Jh6slFl6SJ614
cd16Iz0NfDsTem2rAlDAvIM0YgKRrNlwK4msEyjc6a94q1XMJXnHFXKPL5mitNob
70f0n49VSqvNtVwd/E0oN2UgL018knLJOa8qdfWUhbY+zn736vGxyx16KJfXHigp
prNReXR4LEib5n30oAdtXDok+kRqxGZOmJGWYXJTdfNc4hn4VF0+yII+d7QZ61s+
/hETwtBG3ly2ilsVxe4xRMcFwN5mKb5hlgRwidJI/+aFSPHrcbE0G4LOkdyueLvR
9LSZU+Rj025dz2HRwoiaKmkssTlMK8YrNz/3TBms3DNCjFP/qUA++H4C33f1lq3n
qMAxhL/1LR8Y3aPKXmf9RzD8DQFI3rorS3/xHjjVc1NnQz5NRAvAlL4ASC0pICVD
Cp95EtaJHhIZGEXbmMB6rsyXEsOOOOj1jJ8zwXj9+IJ8xpkjT9KlARpLqcRaHtPu
wEh3FyEYTJSVdn5xjB+3+ssDSv+B1X3+h2Ib4dltmdcY9oX9I2pdcd1aPzGrAu8B
p0T9G7ML/GRvWcW2te4H8cMzFleD0vrboD36PXlYIa0csW5DmnTjzZajElEEVVCC
fdb9fvNaZv1QRJhV8Bc1LSOQXEXVM2bqSr8+YHlktmX4qblIYnzYhBalJMRmO5bs
P3OvTLifPUMEUiVZRxUWlge6yPrZdCkM22rUJrDCx9YEk8ylR2xplWHH2yNQC7Rv
WkqZgzq+q+ibJ6tK+N14xXiqFbL9ZV3juwjf9Ua++LCrnaImG2ybl6F/5KnVUQC1
5l2t+zX8a3onnNx0LP4ruGIlRmvxLo/67BBmvhuGnuft8H0A6cnzsK8558Y3E3wD
SygSYFh8f4qrVPOGgZb3x15L7ku0MNvI39XRqxpogbA6RdudiHSZlKuE5q7HSmnp
FD6BNTC6ZSIBAx+zt26SkceDN1t3HzSN+sdWoEEDG3jPWXhc7ApGfz8tbsF/h8qy
M7JHBN/2n4WAK+EL4KmUaVL5w46byEvwKF8RCW2WJEdVXpSw3pWt0pkkxDSTWKYi
7Q6Z5GLfkaNIa53OiMJE0Pa2INMgf9b9EwFKYx4JAk1zOlvdVpz421sTuNsBSYe9
XuGuL+BSTVBVqJOgvuRn2xCeeWJdTMf87Xwa0+XcA8IhLcmk9oa0/wfveqEGGNay
rhCjvKK6KLK00aeyX/Rz7IaY+ej/oH5g5a40rcVrMg/k1LEeCSjK3t0UQbFzpYbO
aAYi692kQ4ZCc1Rp/vF9X3KQ5Esy2mGnqe3GPw0n7HW4HFmumgoBhx60IKQXTOjz
JAJQmHPX3E0AvBlnCay5tPjHOeUyhS4c3+wRXqXJtEZGp1bc7yHAvFUPrTkmgSHt
qNavgkUjZ5WcPhs6DB4pfsWpMTkVqeovwse/1GajoGHdmhUakpQJwMDa+YAp9ORh
AwgwfSWcGGj8xfwzAxLHh+E5rxxSz0gSKceqmuFDZhIvoJ8QxNWx5QOcKaqZclPK
vYe4QVIYUJp9KYFrv4kTpBQKzuKw0M1JhV4ZQh2+1lM6rWHuCiA458F44Eb8LSML
niuaa4LzH+CAR4YtRUQRsuyl0HCb6cAORwQ7e7syGx9hu7XeobHfKo2Dk+WiKezw
5GocXt3nePZHWM1dJli5yNw5ETYXk8H2+QeqMtzpSoM55XpSlBhWEu2FZFXEVOof
6jjNaW2FeIAqXAdxwKfCDRa4iXYawslyeiFk55YBckkyOCE0Dhgu6n0/8XgAB1wR
zfDUCTbEFvj5fcB8rMXYbmZfCcErN0Obw4a4l3n8qQhoFu+VpXOY0/ezYXpHhkIr
nAa1ngHQPheRuiEjrU0CgtO2zzjawwW/f0UJKGjKYApodPWD+60WAvAFNWCq8bM2
/NN1pF617XyijjhmlJEO45J29uO6k3wGu39rdAAFcRRsJFhVnuzibk+ldh4JePjy
2gOtT9BM7/ACyImAmiLqeeXbTHI1D7nCWRW0/LsjMkjIqGkTbPNS7RWyDA3S435R
k9YnfovaD2dg6jaB+gfccKfTkrOb38lpfEuPGTdmixDSgb9HwdbeVnNIEE/9qWY+
inKIkt6nGozxR5c4fJAehFqESC9Hfto6XhUtby+alaPqLR2lEGbfap4qMvCqzkt9
f+pDVna9UZ4QFpvOpEH5qK6nzLoabyEOrjPs8rZE8fSrfW0G2eXGxSEjaCmPzEsk
e7cRBROB0EUwAuCln1IyO3T3Rv5lMks4G3piVRWFOx0tglLPW2yBTRKD48i6Bp2l
ycAU4UwZjqaU7VwMUQhPqTmmuxVCeLf2d6x+3++Ms8DXEEY7XsBwk7gGgTiXqrsE
QN4vGKilcYQR8hn10OkYwvA3LOpn+elcBb75u7mVnb8zqKvqUsSCEtkl6Gh953s9
OlsVN+YY4G+aY+jhEoa1y4++2eZL0JgosTMUCFGGuVd/RvOm2GoL0ISUI985gHZu
vKH6Yq5AkqHM59FeFtewHri9AI29sjCtfEYsKVqlNPNj5bcCj34nWmNfSMQnlhRI
WR4VYXdPYO2Btv5f82QpOcarV7wjA8iGw8TBsveWapJgqzrO/WEHAZ38HRfWNKQf
4Tzgus5DWQOOmyLdXRoCQGAtB09674LVUnd/P+qnNbRa/19hjrDyieWHR1AywlG1
zPmKn3ee8o8erjknukvTmrkXsJyWZtp54os3RX2CNmGXCENNXcmbdAHjRexupbRE
q3OL8QQmXJZfJtDi8QX4GpCrV6ngMUpvUwtVra5E3ETSLQerVZP4ufFf4NP+KtlV
fEypLDoT+dJq3c5LH8x5rGexK7AcMGBePjfVuwRLTA/QLbdxnFI5JCJqvQDIL/9F
+uqqur3XcN4rmIfcTh0/CigpEwJvZFBLKtgxIVZumBFo5tAMXyckxsU5hh0r4elD
O2k0FNNZt+uzacHKuMluzYDWeuL4EzJo5EGzc1usEa2Q9TXRQhCihi4qaEWgMhJe
TIXgRLUilGAOhBYVlIg+5DxkBwIamOhbpBrC6LvogPGqFPlxdyScBjR3tqwWelVa
vDOmHh1SWJMSmgXTs/XyIU7lJJU3VBM1a60a6RKKHDdUf3ieKzcuQpOp/60IcKEM
9dFvR5wHSTJTS6ZozsflKpUZ1RyxfuY5ZuCPQRMkSlNDiEFt3mhaaK9FncZgxFGe
fxKDUcsUGU8RZ+f6esifkRie+/Avkct6iQF0buNwcB/MPtM3BUB2BzuKll8DVRJ9
Ff+TA4kVZEFj1aUzn68UTSvIh90XxT7KPjE7/s51TlZfBSwM9gOG/S9L91h4q12n
IECdvITj7mXq4ajEwzFeiE6zVR7111jRzk1dNkJEVOt77wZxFhB0bPQkZYbU91LG
UP+PvmokpLB8g+anFZJ92epqTcHpkUDnMKlCIILRXwrmE1/QXWasZ1HGSKtv0Xxu
VgbekIZSqNiegjofT4zLvyy1kIx7RwSfRoHsoiqxl8q17hdzG6g/LnrvZDdavlQV
4INKeURzDoR6iudR5jQW8KFXeTcrISt7KVyU0efkKvvDJG/0z5chqn2IJNHRVvWk
Wn0fISdSxt/E1XRp70KT4Cf62hcRwuWGfarn2AEreaesgFGYDYWTQpXd7qh8gc1q
OjVWy45mBju/ULKaHEz6gBbb4ZUHHFNjbWUhKinWJpkCPQlTatzfYKh5P8JcOEvz
gSGS6KoQvAGmiOqlufsRNU0nSGHM+x9qR8rCvmbUVucTjlS3YgIOWTyKPVolxmSA
TPpIjNpFaFTgDPINo+hYPT1kd22FyevZEIx7q4LuF2ZClOGCool7SoTtcoUPvTWp
3HAw06oTycxkfs6d95aAeXZCiAzEnFR+/e89szTEXQBNHDMH7Pv1mkxSHCSTDPzk
m98UyA7m0NBrMtwb4S+IfMk6oHWaBZ0DZ/x/c+X3fvd7GD4+t7sh2lu8xcNtEXpx
1TOISHn721jCbyxwtyzIkh37HbN/xzICGTM9F6B0xU+L6Ohf69J6TvgH7LZR+BsH
eimrT8eR5wZsAKng6WwmjCVdHCX3csYG9dFrLeWnSTAOnr3woxrg+f5CJK8sHG27
MQwPFy9kyTqiVWsigHDGYk4AU9HG9+jLsQCQnXKmZXi2JP2Y0qDI019GDpMBW0Ng
ERF5vqtFw1RawoCNG57NpFJy4FM1IyS14xzWpuvxq9G//J7FFdimYuxfgrPX0Jw2
OKkOr5I2yHiWDl7cLZd78bNwMBw5BWgJL3SMrqGpg10ZVmsSQfM1n4iLsmQ+fihI
/2cjRch7y1D04Qnbodz8IMdvZXbozy5i1Y8jgszVSEL8HEYlcy07bCGGDS3NcePC
pAoipgaq/T9nwL1zhfvOG9cQzkPV75Qx+8EAvm1j8VKkdyv9YFgIbOt6V7hgZjJX
fgEgkLoSani7/JNGllaSYSD9DqQWRVvtcfwKku7ykwh0fJRuqEkJYl0Y6sdON3u1
om6LeI702ttkx8Yvw+esml3ghtFXt2sfbeTYvEUGH/YJx2q69aVovqQWlLF2LpWY
D4sBX3TWkloRJkCMSxB2dvcT+5FUMyvjfb4d6gt80L0TxI7YuNy+AZkw40c2cmpE
smILBTp1UPg6rznu1wZPx2qXzFHF+NRCYAAULAghvojMYO4XWaO8vDaZllbzJc9G
LrJNvt+SjpdhQk+hm6Pa0sg428MAOJJYzk59WTMJrOeOOFR1gjL0kwJXG/2aNg+x
AGzgyQrYeS8399NvjL0Wvp1zvmzT67zjy1GJP2ur8OGDgJrBDJusI341AjTcrRWX
xKsk+S6niMq9clkP9UZErhBIYXfS47S55QZPo4qIhLPWJB2KJIBtt+ZOvh+z148c
nydByXDt1x35WB1NcK7F1W9KJYhsWJps49tvJ2nzRfIH9RPs7WWLBkVsFMXXEwXl
47WejKtSatMKL1xYa5qwRGidB25UwMYgDeTo9052HMJMf2m/zSMOxGIMG2A8Y1eo
ypwLjThRzR3y19LsjhgMIgbb6dwPIJ8x0iflKH2BJFx6bgDq5F2OJvnrJLSBN/C1
/ueonG3CqWRuthMtDMIC1gfdxbC3vbsgYd1VYMiCxQujdS+E7v0Zxe2D4wk/gzCJ
PSa4DDjXxyJPnEODvdimNvW5mcJbg8e2y8F9hni6goMP9Lxk1vVH+LVwG+AToXNm
o9hXPeGQmXPlXc5xzi9VriuolNfGPgKR3zhi8q9Fo9MOPKnWrNmrIg8WqN/WoeBu
mDTUwhjjJXc8H4wzm2oevi7RtHy92dZWIZA8ICfKLcye95I10cjercRA4SSAApFZ
0Ac9978tfD42Fxd29jGvuuhHpOHrYuW3B1CyBk3H1RwVD0mh1cFkLCdCB2Dzsu3U
r0Y0pjuSeVu3MxswjMl8gp0stlV3DuJscwY8E1A+m9xFIgJeYLlnXzQMBTPBEnED
/hZGbtYvmG50Zc/FiMKnKY96scVaOycHjrhVjx42D4RZmoJCfPTxaATXj5P/v9rW
jkCwTUll3FpNbgoxPvH85x4+8jRo8t4RsAS7FyYAqv5eleN4RnMzDBR9y+Sjz7Pa
VFMtL1WFlPxo5uNiOCRCqbpXZfa0K8+GFJ0U4A+ZGkLg/cETL3bHmH3mtZf/QGLb
oIVwZjUGYYhpTHkzNLz28bV/XHGWf0lPN0m/nx9ddHdj3yEw048JcF04lPqsFnH2
Mgu/wf3t1j6rS+sGq2LfMdrlhe1SpOTNfsDhKkH8pIBIK3XguYB2uenOtJSjSeD5
0mycvPTZnud1S/yMJQHC3mdjespXtE0HhGY2+bLlbz28DdFubSNwH728ERd46rEm
ZMe72F369p3gay96LmHyPVShqP/C8iF0gRgkAUdjIqQ7Dv1ICfei5QHQ9lpH6Mvn
Fgn2zDr7wWnmsthdgFmv6iWA8DSeIneB6Mkf8QGP3UyYkaNBz+dLgp16JktQbpiA
SxmlD3Z8ojUXOfBuFJyP8Pu3Gb8BSiMqNPYDDI9Yzw9ih1OV/0efbhbhIgb79Uag
CID3TfhQFsnDEccK36eadw8Nc0iozdmlP3MsAeC0331CZ2OIy8zC0cONrNgynpda
8GHJPudht5hlLcDfoY+PUZ9omnBPOMRyfHe0o/N9/8d3vS+f5fAxLPWZm2DGBFBs
6/G8BW7hanDuIv67mTpffWcyBGxAps+VeeV26qi96TQQ5ZIe/S1AdzAqZlK0IcVv
hajdUa7PkuduJSu7jmmsQ89SnaFeaMrZohweDdxGeokWBqKQi4takE5xkU5rr4d4
xDP+gzD/016Tvc8kBHj7qYYRNuJ3tCrhIytON0aXAKnmK2LqC7CprLZKntQgSw8z
EbZ5JF7bk7k8DnXMtNA4qbNfNY/HKa14li8ycAbi387KyPUd2AOwxg2kXrcCqzHu
R+/jYgOheOnKemMmRMebiq0y7lI7h6rl5rDwjEHYVk6oFYiCabUeU0ri048xSi/G
eLx5y/xeoHzousvDXx808FgwoDtgnxCe7TCpJswLYZ3GaJ7zK1VqCKlKtI322qYl
H+/+qwg0cF6uomtqjgGiqxbhf0GClaBlemD/cjakPR9abQAHqaPWFm+opMvkescj
437QYI7t/dphOb9VRwEyDZBLbXkbFM6NSVhmHqTaDfBCXNkQelSGR/Dmwkkscnfr
44znRzMt7JwjOMPSRJ/SZlwaK9fclKPiYpOYGXm7gLGsouWujF7Q+f8Cr05KdZ1G
8v4+/gwW+RL83Mfr609honP/FnHRrj8BhGresafNjDhnzKK6gKJMajPDGyqp7phX
smjyDVcOzsXBYDw9+v2ZWa5VISqrL+oh00/29zU11xHfF93HOmN38pLZ/BmppG6I
pcBi+xuMAMBs73N48rc112e0v23wwmQ04g08sP7IRhI/4KA4PQjqPijI2nNRS79N
Cd/8i9ZSZDJYuzIC89675H/CSyUUr3hETCXdJnFUo4+uiTtmxba6HMm9ddprrHJM
qDRXBDFZMbZizGesQuCYXnT1vQE93ANJfBRtpFqDXR0+gj8kwspB3EDX/7eSwXn4
gS3NtY07vd1lcaMN5C7KjqMVF/Ytka6yg9wImHx7l6n1iDXhI727s3UDJ6oZQ4Fh
8Tnr+x6sp6qNYYrTqppF2AWBI9XQMMmfJzDpi7a/d15QCgUQ2oqbvyEc13cTg9sW
AAv/8fP5qMeTOuqXFmE43XLxvFTBm4FUfBNf+bhYMo/XeUGNbSy6sL1OXCS5GyLt
sYfoSPUWkn0LsQw8lIdDLCT6pfnryZssk2hw8OuGINRUL+p5DXbLVA8phFQPEd5I
rcOFaOZkRQ8l3/QEpaPgkKOgEPUObt5OO+t533gdKMCXm+xAxomzXO+Oy92H3Lmk
dtHpTb/iqNM3o42U7MSyazyHqb0rGmnhatRSimDWQjV/21hgIp5Ocv2PNjfVgxRe
YFlTXbKCj+cgqBs/ecrOiGHH2L409sKiN7V8tfnyUgWGmpo2zHiE8vLNi50KSNcK
KBml7U4y9T0yCx2VkZ85i4jyPgICwsCg7wZJq6ffiyIPSe9xefmfSb9A+sYEsH1F
nsTsnUqidlgisr4rXIL9LfYXWFouGAYxR0Rrfa4eIcBlo2p/gKeVKO9XhLJuj8kJ
pFbRq8F7xlqzuF++cSnV4g6OsE2ZiZ/Rbq3gnvss7mZJuVx2PyFZL59xkt4YIqPO
nZ/6zZ8EA+nYu027vpORrsXLasxG2w//PqqcYmx+EPsGqMHrnHgFIZ+5EUd0WuWG
iFHQ8zOhy2ZEO7t5hbkTvcjugM6PICrjPt+i+XgZff3ct/b8WVW7uzSdXVz/LT2F
iCbBjUjH/XHNHI2oaFzrtMRGh5Xe3V5mTULyGiyb22pgbrH2sbSROB58FohrULE2
sU0uOc21lHeNofRd7meVuB4dNIq8t6kb5Fb2LRpMiYtLKtttAS5h+IDhG9fOfJw6
/zQGTlVJxUb5/pUw5XQx5ku/8MVhxn4EmYOTOaR8z84Rqc/lavDoT4qokK4hhFA4
x6L7sGhwMBG9VvhTtGYbwzPFHjR2WMxG1KBu3esjwwgqStK/NU/rSdPJp4cbGeVi
FrDYOXlH71zyE66rr9FiZ8DWhLRQ0oymbfEYhqUnJbtgXB5+IaReKh/KJeLduU8n
A03LBEJatVbW+xcVmFsc6mAl0Utp+fTJtaN0zGSTfb6Zqs7MFOd3ONzNdKCoxKvU
Ka6GPgLBIjKvZX/EW+XUxOQB7yWDiHmmOM9r0zaurQ7gJ0BHENTNiJzRhzlRlGc/
h7sTGc69nMTdZVzKYWM39RVMGPR0LqBHgXT0VCTjnSDNaAuIs8jg1qUFMlFP98y3
APXs9TP83YfXIHxgj3YwuYnUQqJmRu5EP/Ct3iaLg9ztJvwC5XisDEZDPi3IY8v6
Zw6J3zzKoVVQ9Te2Ipb83Ye4MG30xzYHkMjJf98/Y9pCT6YzLxnf0x3DzprsfKg8
1BN7pZxQovE68Q0gBitsrgNeJhNt2b74hjzc08rYJPEDdwgav5YlT/jcTeyhA3fN
cNnkqCouUG23fSBOqAAjagM5nk3sGjoNTz1kc5VqDrB1BZeUK6LPpOTGuYcg2su1
nY2aj/w4movu3OpZvCfRKW59eRr+PSykWi8ns2cAfL6N35cZB+XRiGNlovXLBKUL
Cl38dpglYpugwGSyeC25+dakncqSQF474Qo4hWZ5e3eXIDpbldVw29IYWtHst6pv
MF48voew1cuNYnVv1x+cLRZjB3WNXWwf0oMtaEziZ+e3aCf5ctXFOyGqRXSRfuuB
wRmLeMhGxn32R6LmfvRaBH2tLkIwL1G5dvgnTMW/rL+/RLdtz0KoozfMTo0n4Msv
fjgQ+N/4UD1idpxPEhTzki37st/I0Kn8BPH9DdqW2cras1qXLQhUMtwVTPhLBc7n
tSGX4xleIuNhKT1HXBoGczRrl493VhkszHTl0lFBCGHsvj2G++kdjbCpOakdmwJM
ictpTM7v7UHDQo3fP8jgweAi9I3gPcp7MA3nBuB0+JtxtmiuvnmvPA1W3Pp5tFwT
nDjkuiQhv5N5yEt63EM3Ax+O4CZ66af5WUJ1Ec2wDRv7qQbcnazjrnSFsqY6GVh4
t/0/RfzZCu17wTElOkuOPKrSJLLWDGmPOW3dNGJ0Byz60o5GO+pIQ+mtpd5vm4Ss
7ppRmkhqR1Ai0CxOg0g37l9KJuwdcB5/cpUOItaggF34UVQSUlEaqQvZOLcnUX4O
o0S7WkKcZa1C6Wc8bKCG0NCAlkXAvdE1x3CrZffKj4mNPAIPCKp7kSZcTve0GidL
JLTQmxWPHfN/XWMrDXOLt+pZhXLLeYGNVeJtMTXdt+f3a1g8hPFcObw4strG7FFl
VZbXOPOFnifH6Vgjsdkm1IoaI6X5gZ/BLYtO0i7jxgUvMlZnMlRBOv+bZUXBeW26
7eX0S3jrRNky54CK3FmmRrtPmsHpKb5Pyp57QEjhxJIhlyGNTUbVWHxSj1W1Qb4C
2zHMdHmEa24GdIDU0okiEE3RUMJ/BVDUHMomkJnRpoQHAof5AgVAOEX+IDBBhkAy
TZfnq30OZKUIftvvZT9Wxqa62Lwo14mJdb6Yjsn4rzeiPWHaeSdDNzEhqgWNBxMD
RW6xhmhIJ3k2JeonX+pQoeFPavoq1iZMcjimW18JP+d9w1zGxjA+/1beH8M01PLe
9rUbTP6Lu0CsK5s8FeuMYnllF4FNa1Sj9d+Ax9Mz8kbDo1WOBRFpzcmBO2a5e5GN
gzO76btEf9kEcgh06RdEKlcqf78gjnfunWqrvxzktdmRg6rDPfR3D+HhjnnkL2aa
BOuw+g6ArcRKqjCegzva5VJb8qWoM0eZfaykyAjbcVCtuvZCshBV796CTHVskFe3
JOkMGQxmtlFvKXiwqfFE/zVME6sC07UrWTi7zeGSKkXoL4mF3P7m+aSD8rbhNSdv
4LqdVBukh8F8peee+WtM9ps972O1nmZqmmCaMfaTN9xxyHr+gbGB4mVXsql5Xb7A
BIaspNq8QVBBNSixdcI2XG0h8zMnfxWKZewIwd7Ojot4VFO+knnz0+U+H2pC6xrV
NnKcv6Ca9xLwKoccoIetUiRNwKKyPmBw7NZ4psixy6YOKE5NPybWf7RpWx1M32pO
3H+/Q1bbSMXDBGAeVPc1glFZQfsZSphth2uB3TNz16PCfDc5vlNDj4qIDypf9pKy
AcdQvQz68HjsaUBgN0SZlpgXvQScn1K2INE6HFX/DvPGR6ovespBpHKYfdzDKzrv
cU5fHCuX5MsaAOasWpIDf4t9MnZKAMQ5bnwUA4ZkZd8K2TwbMLL4sIDO7vBgJaFx
pzGeqFbcafUPOwr2JSovr8ZYhYwFtCsm552akuAurd7etFtyFKqThTK1hWYYRptL
AZlk/gYguV1BaoaL1Zna6DcBqn2VVlCOBIZEkC8YfGPMUgYz8HF6EIs5HxKqZ13A
8Dp6pQTUgUydD8KiOLhfAIWGoURVIDi7RKxBsX0c9X0MH+qVBRk+RRv6/C6uCOQQ
6Fx3xY+ZUYHfmyU3j/rC/nHMluVLnbb2/0K3gYao+xPzYLOgV9sZXJq/3rooFD4X
cb7ztwD1KCiysAq1xgOzB+dNya1tzi1dlMbvz+exmK2rYGNB3dpGqpgGubqSb6KZ
c8HMcF9H1HpLehOYN78Q3w/Qbly1qtMsFTWQS49gTKGfdNs/KgF96hKAMoRXnT6O
1yJYC0KjoPwvzuY8eU2HL6UZre8hHTK4VJqkzyWrj/9VUYgqy0zw9LMfKZmKa1i7
2zMqurBoFnQlAYfUGAYuibu0FegqV7sFE4jd8xV6n3HyK8/VqfK65eIC7EKfVUQN
CvJde4TVZITkKuVDEcH06ATUm4+5lq/6oWLl1rVzN32JEM4yHdnTrgTnHIUsPRws
eEHDLsIWYVSgm9p3Nf5ESCAHMO5tTQLIgsvILxfDjwRrkmAhEPUwgwEkDiXT0Fki
LhDEvIcbX1mj8jb6L4SdDZTAoL9C8Y7Mc4ej0rgzy92WQknPfIkbwVNm/WZvQ3YQ
wsS1MzVu1DMcnG3GWc+xudb5xYaZpxqAjYhXFcZBleE2ConRjdxwPbKx8s0Kjrpg
WbSga6qTwtAqoB/8hVwZUtrLiQAB2pC0J+GZKb13PFrw0Wb7EjyyyETMV9ny9hkC
J7vjRE9N7TRXkricYG7vged+GyR/LwSskFXfMSIHIC/s06vb/3J2BFGC2POILC0f
TluqGYPjqviV5pX32kvSwYr4ITl1iNpbHit2G77oahYAmcoQwa6XUqIc1RmiyzpV
XwoRiBET0dFLF0SEnmaHbZ2NzZi8z0JlysI83CoSqS7/ewvAj4odb4NJnMEPMDcd
dT3bEWrLOyB0TP10Z0nB/nwXy+/PFNSUQkRyy/SbtCAfO68112pgQPbEexqAffeP
gx5CuSxfXie+UO69xAyHTY7KwV/mWYO7dkonZwYsbSttSFN4knjI/qatJEdvkZV6
DZHVv6b9qMRhHKcuEJ7m1fFWslA0oTTaZrouVs5aU4ax7oDun0gbnMg+JSm1vCz7
ZInnAxgwScDhYMhYISAvXb6Sx53NQNT8sABWrmzw5Xi+FZi9DcS6xA0SsW9KLWBT
sdQbC+DqeWUOKabGgQCz1N8jMWZ4pYiFnWLtjYv1FQuEM5M9XV7WosoyFenu6DQf
SjGGz5vs5u3uKH+UYAxcIoln/frHOtLv+A90Sn2feNyeE4tqVApAOSLg8prJHhRD
+QlCOv4qT3IuY7Enooh9JPE3XflQ7FbvKr748cPn4mFKZ1RYB/AdNHlk9TcJ/Oqm
RwDgOSPf64b1oJQIsOb5z0US+K+70Xuhsc0JdjPO6tetfOGZRKfKQzmwdqxWf74x
0VZ4LLDw/jEjUtiTwyi2JRokXQoK98SUjzlWhMfvL1D8c30ssLdFssfqOR+asK2X
1uHLSHs1EZCgOp0hwG9enM/BluordWTkLMlHn/lGSB9NYlMLwfQXhT4x5gTN09uU
QxoGvh6p5lu0rVthzWsPlpYiTfBqMs7G+Bx9OsOXi50TPHbck7Ff7ZadsKEl7/7v
kAHE9vvxMSIm0kExCW3bOWfpM7SUKLCbirreY0dHeFRSctPEBED+r20i1Gb8AZIQ
qin9RcsJ7EzZHVICLDB9GTRkgqgAZgEOa9Uq9wu0DJdIqQDNN1872eeXepHK6zZf
2L2b6vLJcXAxxQ2TCN4acwEkZLvADQrtNd7dJwuB4ijmlcx/c5f5ByziNz3AgRaH
WU8xdKmmgIbGIoR7ygSolv/iCuZbi3qBUTk7Y9s5xpx9CaGS9sC/UT4hSEgeD/7N
6qHRMbXo6n/xNnNzxwXIlQ0L32NsYqZlYI2+6P7LYj0qdjBnkBPNdTX3EUwsNvXU
MXkefLqhDy5MXdXWiUnTEAH9IUZEyB09syF1IFGMS+CK9hPhM1YmRycoMEUPVS+P
Jygmvf8tydllMfjy5+xvm7p+gRMQlkywGaLMWpaP9xR5TT59yui/ak/av+Qm27EL
Zliy+h8WpaIq8nD0XRYLelsB+XttK34YesT0VzG2CMLeXF/kMpC/vtenFB4mJk15
ROhvU8cy9xoku64J2iMLVhTquvP8WXJSlybDlcE/tnUfsApZWs8g5AUX2BZCj2kV
LTXJuCtfoY6y1Ko9NgHodSGBJu6hBCU2y1x4ySPDzyw8ELcW9q9vVeW66PCVYahI
tg8Kt/xCYo8m7p6BzwRXTSiKkHg/vwWDztjmbryp048n1vd/4Wrtg4rfPMDGLOBW
8ECIXTlvMOYf8Yj1irhmzrU3JfmOVS02YAf0m9KrGk8JBBssEHX708ck3hVAiNnR
gLdGyehvlFdm2VLdDLmkW2NblBwmv3AeVG7Th+jF8fAqQ3ENkqBwMCCvO9pVU2pA
16/mp2Gcq6BcNH6jCy81UWhZvxfLoRyACHRMeO7gXQO1gD1UTC+7tBgmX/UgeUPv
STY3hI6wSHMP4IJt1pxDVLtV7MKAc106lJQnW7Oc3+6KXiHA7S8ytGmf9RE5cfd+
GMDG/mirHTd6sjEr8akavg2pcH2AY8MgtIOVh0dCfMupI9PbtHlQff6cDe6SuvYi
FTf+Lb7eB7IPhuN5GBt0XNYrhHTl2Z5niKKkSCdbRAhLZJgkJHZVrEPhg+rcrBGz
WwamFEwp4SQ3jWl03egvWn93l932t7bsM8iWtxNSwSUwj+0nK/e2OAuAzgJ6vYGC
+5sv2zXQ/t481tt1hBrbmArXetHrz7fHG6POMOchGTu+sXzkYvXu2UCJeZE9lKBH
JdcPskb6WO7Sx3wDPmFPzk3qGxaXu91k+8ibsrsIWUoWDdh63u0ItfZEcR8N+Yqe
BmCE4qaEW+ukJywGNN8JtxeJjDoy7ufGOEc0pc+EHoniKLKXuHWwQz8zarIag5UB
fs2RbMVkn00zW44SOywn9b5cptzzDcAc1AbJXZ9EBoJTct7zkOfMC57zCe12nHFd
WroHvqEw5iIhBWC0Zwxh0EMWpdh6ZWsnuaDp+AkG2cy+QuphJOOR+tOYc2/tAKpA
g4TIIQ2nizhTqo0YEEuh4gRMci2GMD0rlVeD2GAXynz0Kh0uq3RoVekpAj1HaS1U
Fe5iZeyd3lymDWmcTwUsnTFebdsnAD/0ISR0mWP9+Y6a+atsgQzzo38A1IZ0/m0k
k/kPdbYAo/3/LmTGURfz4SgS4TXGBMhZkpGyK+nq49xdy0TVldjT8BPBBGsgNDF9
UOHeoh6GZTwmuAyRpTUDTRzlXOy98JyidMVDZvjmVUIY/NEzBxXlWUjMbEy5R9nG
9a2ARKjkPKyt1Zu2uNfdho3k1mwTmEgUWh1R6KoWO357TAEK8qtDr9npRPMCYFE8
1aHkc5uHd+AMJbUS/2XWjz5X66oFqtOrnJFgR85cQep+RCnSI9L6/zZMc/SBD1YE
jMPOPJUGto4Pzc1f4Xya4dZIzcuMF0Rinv0GRK9tqK2ToWdtwok1R6zno/3sKcJO
79lJhLOtZ4ZOXap0SnyaBljiXwDIlCfCcMtFUyo5I7j9IKtxWdmLc3cUOLhYeqAP
613da0sDRQcvf660+f0EJzDFlBFqM1B8cCJKv/8K7dSBHf+NjW3C4dvuitgpnUU/
NWViAcnrfLeOOhyL4WAUjCIa0pHv0sDuoRcru+GEVDOv8xqJW8fYp3urBphLbfxx
cRQwG4TbkjJcuRHZes79tQdnSxcSOhtdHMF4piEbt6i/1GPs++Gp7z8bGGaBdO7F
r7m+OCthVtbMwsXm+HJBs6lzEL5//R9d1NYXtOpoFc6eweQxgliu3ymDfdJJmKt2
Dzmtq3iTMP+b/Yv5YdO6TxrTIT6GRN/vmCBozwgnq1VIAzHkEEDKhzaa+DAuLDgL
SHkEJJrQB9cpNC+GCMAQP9CZyCydUHYtkqFFFqQRrCccUpGI0MrY0ziqyXiQ5DMi
RMJbS7XkvzhLc6Gx8BGZN1EZKW1d55Yc6sMT0QQU0D49x8tIRKAofbikq/v6oe+W
iv4y4lx2tcsNbJMgZ2G+/123GhIRTlPfy6CXvyKNT+GEhf9afIM4Bzvx6ofwq8bg
lXRwZg3ehnDUx0xE+ablM9/QSmuk7kLrGQFRmOEum7qI0xhjXCRwXLWdxAwB2vbF
6GeGynmgF/dZfInvtwhyV7T3J5uYsdt7kpfe9N/Ij0SfMXmU2OzY+5P4FLOeLXwZ
EDQWcNpKBkqeWUTVhaHfWwt6wkSHhsA0Eq+Ysv0AH5+LXF80fEAQaPvgFfjimSBl
h+lUB4b9NjBVAAy20v10Hv3OL5LF5Fz//fNM2d5mePzQdy6YYRl/C54sgnHDv/Zs
CYe/Z+mcDN1rRnNXjPTwT3M4jUThQ+zUYn4TQJyzWByrgumZFpRKbYqeFIZtVqe2
PXCzCIm71kj8x8twflNdEAQ842fTbu56Hxlm6UHs6UmR+owe+hqzVdRX7vdpWake
lb6PrPjcClc+eho5G1NgpzBiKbGCdIAMWOPll2V60U4NtsiEu4YFFuc3sS16tQA9
4SW527T6gl0RRAErBmZ2/RcXgVjGaaqxMBpYZejVrf+dF+7lo7itUVr6jsxhAjtI
39E3tdM4CXyZDJsItU6w272xpj5vHiAVKhhC+KQyWQ8JBy9DDkfoKPY+r0sTX+Dq
qXeCriE1kHnM6DmKw6XJz2CzS/Cns83fcTRVM6bkugLc3OnGU3NoDbj0qyigK4Eo
u7PDuvX6bfZXXBtMwC9/D7Iedh7HpHrXHk9VScqKrkLkxaZr1eSg8wJ638ZbYfyk
UZtt0rP9Zxx3/AI1MD+FX9oK7ShWTiV8cTKBBmMjrQNs1HpNNCQBArGVKSGoB20/
Kf+/EeceibiYU9MM8q1FiG5JG+mXf9duwYqPV+jWY/2qboR6xGSYoinXSeubPAGF
YWyMZJrEqtn2e9TSky+Tpcp5gySseDcWtFLtncq3UAkwuhcqhks8w1bvDcgbWuAF
MzubUcxmTaxmum1W1KAKFfqgdpStW/N8lbsBW7xT2lEDa+2qDMn95vq4eh+dde72
TR3OYz7+3IFsVTHZlwt9rnZI+TN2nXOHeRIjHEVasqkXk5twNaUqA1rgh04QvbUu
7RRscHR/oAryKHVF6WL3GpyAsXUtYYKTe+EYpzb0cWZuzSFoJms0Ck+nWmIDTSvw
WL7tSfmAZAChxqTddcVEsdoLMSVC7gFFHYjvTyGRJ0JJEbZq7d7GbvflRIOT0uDn
YH625AAcFoNYNDk3Jk4G8Sc6DMPFMOPBhK3pYvuyZv0Nyi+maCl8DZ6JqAFdGGv1
jvchlPN7QQ9awvsQRKiYIgRfVoW4vpRNbQAS0iIDNQwrAS5NwglapwpP1VhbZQuw
HGmpQDEFHhqStEuR6EfF2Xd/WDxrStsW7gFS8XpcmRkchd04cMg29ZZjpJyLx6Z1
XYG8DSvXQYBkhncQWx++IezCxxWv9ses3G4utS/qPZD5iSfgdWEEboVlPmatl7w0
y/EO1LAm+4VjmG73SyF6y3MZ90fkOFrG2evDKiRYaDxtbwERgheX17LAxCP5gyv9
kX8sEzpLDN3MOUgieFJP0m+GktMgIVO2lrB3KDk4DbgR0mXf0AGXvSAk95EMx3qj
ByEJK99b0iZoHgYdZvi09nY9LL+r6cMQvPj4+NQEzNh8TGWoy+UW9/+VaZ6mXCKR
3P4Chs/HA1TWcYdHcyEqjeAN0/zJa6mkMZeEMwZzyN1aCX/SWwuYNgy+e3jO/IxB
51QCaM8oBTtSukHLjEq/Wkx4wz625yxeAGEkHi3g+8CdiC1KQk7tyB+6fxvGL6oY
O4hlBt8Ff5wRS3ms23OXl20PLvsTvAAivhgNzNkoQ4bLBPFqUwDEQmfGNepD1L3T
k6kL2hvU1BZJk+PA08k7Q7HBNhShngDG1j5XtWAaiW1f/3B8T6k/YZTTDS93T0jw
Tphbsxeh9uxjVSCUPWSMtfsoyMtOO2iOHFKwGKMz+BQyzuOw4dP5iJaSswQkWzrv
PlJ6chN5kHueS7ENACwVY0Ce0WbA0Y2QD9SOB2y83NPIr9Wb/MVb6oTXEtRb5ydx
EZt3LDJGrbVqd86yX9rJu28h/wlvI6q9oMNnd2AbDMxc0mku/BMg6UncjuwB7GnL
q1FHTVeCC+jAn3d8QrMnAxl1fLl+OpLsT945KxXCsqwuprQXjwOlTV3E23p+ohVf
EIthn3ORIu5Oxdlr/z4QO8fk7FuZswJ9feXhgvS9D1sjzN08UP2yHc2dWsRSmjmy
29x5qdcuDpDhVAxx927InukiJgEElcCPsFX5ZTW3CibMWKf8YXFIbI/vuojAUNpi
UB1+BmNk5AFzRK3Pr3aCmptJmlIcGhOthUEyLQgqel/Uvki6TZV4UePzTrDfkmKD
C/uDbJ6rWTe9UPk2/Lzzlu3AErtDz9CAmeKpsJZGzt3F/jh0LNzirsMtHfrmkTWA
1oiH8Bp5DsZrHwX4hA6cxj/uJezGz2bND9F7DAZGothiGgT0eEUJxRat94LFyqcx
wjuylzftR0E90Ipp//8xPEgdZo5RINnl4w9FWykfQTAK/INLvdKj8XjMXV/uoMEe
rwsiijIFjhzuGC25OuYYC88D4rJqHxNa1w5N8Wu9jqMWfNbNhGbO6foX3MAXmcZg
6f3B1hItWNzI0hue8mUkDFO/ec55XhPaqNmh6GBd7U+CRmKN6IiC6f/vNqRdF/9F
tZ4DSKC68vJ/kbDa8ntubqQa6LWkaHuDeAnNfpMN/YehY/rr4U+fMiF9JhLS8jIk
RUVHHc5/OFEQ67JuhQKWT30cf5z2R2rdNU0WDWtTslpz3wkElZUkXJQjS19TwrmF
rd6JdFUMjQ0t2wPmPhym0IqIA6WI4Zb5XmPxkbevV2kJaWaChhep11fMhbcFWdPv
jIkiDvdq4Uqkg6pXkqs9IRlQkcNVhS94faQPtd9KRYuVxRD1h6PzKEkBTrUIafIm
IXmIZdp0U0s0Z2pV4iPeUaY+ZBUDpDEDHGK7NwzIENFRCudb/MveKEidZAiqZ8df
nXslqaJNflbvfm90T6/HdX8eFAxpLaaj07dD4/nfZRJNkZ9XWbWr/x7S+kw9lSFc
JPOyujMXDAauQ6UZpBmQOO/sY8cGwCY5Ft5uBUJ3UiAYbyL8NrseXYjmWpKYfoTz
pTL8xTlxBkZCrvNy/7aRWfi/rN8tonvwSRf7m5MjJrgUPk6bJ90ksG5eoMnfy4IG
LaXGwY+g/gqCbwbl/haSCdFi0lTnOvAynS+m86pwu/3dst5STl3mr2r2zWiQVBwb
guunSZZM2d39n8hlVpBgGE2bvx20+Z8fGdr0LOkDPRDd3+GWQRmjtMOUtSIO/H2K
bZpwjtGFyIvNDuwTMN6uxvOl5xCTe/XH85foupUrPzFhps4zcqxQ/GzCLy/nFTsp
vv4wU/oKI6FCYUNl0tfOl4FfwEquE9LTyYajltHbQWCvB8oZuUqySiRS7y7XuLvC
8KRGSfRE2QE2/jrynUnT2YRXpXRFs9XNOtVvSFqsu4aIeEQMsggSbziLuKsnWWHW
/GGlvguTMpVw4pAz4uOXqNmS8YdWMxf9U744sfDgNz6N9urDsokYZ936ofIRhQN8
NbySqSNiHKo8vXwT15NgVBb3GgKUvf2mHGWOA3GDXwrLb5VyXH008KcsKiG1Eijp
a0pkaW+9pOonJM+FcKtD3w5bZ769rcqhVc1R85Lbuo3/x4aLaWXP/PZfF56gP7wM
/DgTnjRLmPIqCY9H1l3D5C7lHKu+725Wbw9N8S8f9RiALC0OfB5GoOEQCJ/iM3am
aIJ0KOvt/3TeDqT3OLm0fkvXPDUdmKE2/06pJvEBON5c/ieS/jeatJlrUb0UkKUy
/EN/ec6FJ3zvFnpYDxZAU9G2tNqQOXPpGpYTlV35K9x2lr0V/WN99WhE5QeYDPzx
vemBIg4obHRlUzdzoXa+QTCp1qbNup7TBQXpEKrKlyV6Ebt4JvIX3qLOZp3qYZig
2vnuAqC3V0D+twP9QbCOYBZ11v3h/GYdIuUO+OEAyJyadCSp6gLLhuCzKdVOVD7J
vAOy8/sqRuQg2tReYdGv698fIqa208+nLt1Bz8cLku+tvXY7yRaEoOAH86/NlutC
+tulfymsrY0dAUZr8rawX2t+dTCmlSZS6iCmHDmsqhYAQCa7PRk+idbYn5jWvSJt
oIw+P4K5/JaBYzs60pOZ6XQ5baIkGC7r9KNJn3A27F8nmon5NHGtOJjAMt8mViz8
DiWWcTWWwAbcvRaLaWlec/Lb4WM0Rj+P7zM90T8/7RgkmV5CBPbbtL0vOLtQn2fr
GRf+pIs1F6L9sUz+UXMYIWbnqeOpZeFvhBpRlR1n9ykhntSraDTGNlKxNUs8w23G
Zq4+Ls7yoi6tkHuN1AwnbA1LkMhDhznpB6873vEk6rY7dAVuJUiVaOx0EdnCPxPt
Z3j4xWBJstDwbJ9dwu6b5zcujO9g+41+ziLdlavQ1iUGDKI7iRuxrh4oDoRF6Aar
CyZWqMR/koyO3r6w3jHJgQMxMvlcfb8oS68f0dpSHNQgJSQRF1e6cKaskf6Va9CL
VHnFp4uhd2u7qTUqT1M0bzTIahcEA0xvgy4FOLqbLhtKg3/tsES7MyYtKXkx8NVp
EMX+N0c8LqbPpeaB9dSUVM4BJ36eUItZfg7thw9fLEnfAxb5gzlLuk+hQWAl2Sc3
617MVXVAcDdCnFMWhXy8W9gkfnqmCt5KPzGnhUzl86OqLjcj1vvkp5Mpv1/sEE0P
6rx0bylty97mNBZ3ABNILUElaNyb7PuSsmr9Mtv0+eidRZQpE1Psmdpq23uVATkM
i/5TEG0WUrra8zUHci4kk25LZNv/GWbL14/V9sMzFUaaDKOp6FO1j7YHILkFTHxS
cR4ZKghorcdHUAEc3Q/iZS0ycgVAKnBiths0ovJrc2GGyFoywQiBR8pjlJcRoQhu
8ZkdhC3y9a/ZcZnW+6mUvkmPUYEWCZlYYxt7602lyU+ykWVkBB0wMBcnqUn+vlf5
ieUeiND3M+MLPG8hLilcVbIDXMhvWLwWdUNISq19TUSV4BMOu+bn2zw1RSEsNlLz
PNO0M+v5UZrCnmpHEhEarvREdcBA+niTXcNnG3IvpcZaSrYPxkQ0bUvMTjvvns4F
mufU3cPkZqJ9xDuxUsO0iFle1cHyyNkTCy43Wnr3vr1J2zMW0Y++VMEpBcm79SUj
nGUSS9Mhvk6eTJybBOWUGMhmwwgLyDob+qGGD3C2OM/FYFbXK1thDiG+TJmTzqpw
HivYCCcNgD8mlk/xrkyuB2QVUZ/15KqpOfFow00JyjUDsj7unLKheKJ86aE2q+TC
VMkSZftlAMT+Rkg0Ov1vG8Y9niXMcfs/58dbiOkf4Ry9tFp/AGse/DGAf0TrkyTm
d1/SS3zMaLhVbAPKeiUsbq0kAg5uDnchIChx1NVGijrmj4tp5Fx/Lm4NbfoXVokH
FIfJHe2MTm4vqCwT8qxd2B+c1ci8DfIFZZ0MzbXU5vSTahnZZ5sSpnU8B/dDM+5j
HyJ0CauqpKLbwY+3L8PNSzlOBDaWoUjBcKbvo+mKfWdA7WHLO+aSgv/cUYw9BtNI
nFglw1OFe1NGGA/VCSXKqdvTE4QAff3groPuyk7+kif1ZyRMD758FCuoCfpHOwtk
PA+v2D0K+khK3UhOVE8AuC/0GRPJPMYwVmp9t14srwGMwHHz7Y3WvMDsVgqYaz3Y
4OSkJElr+5zL7fkpOnZQdqzYOhHzaxdtwvnesOg8NpKs/HHUvz+fO1Sf7DrXfKYa
mkn+Hkgzw6barRKWe+KMLIzunvR+PppZFS+H6dtMebd4lEsPqjE4YHSIqCTD+VP2
s2O1GQVLIVbdWbYQBZSGS5KaYpEEWF7G1UvVVSgILWRKVYfuq0crxV/js9rZ/aVJ
h5ZQYELbndAaUiVj3WuZ5V+u06ybYAErP/VFVNlDt8bijRCodFkcluYBRoHvumK0
rC9y3fKTK//oJnLcVlZxjUUQNQQ+EtWpaJMsM5z+mqAALucKYA3TapqXwQr3HYjM
NbhBejJRfDD4DhXdnYrD9BNpnUr7grDAyB3J6BNcsAXCOp7M8c5J31lSUS7TgWJw
B5KjdN79LtXyH33j2uu4zY1FjDx0PvqMrUgS22LQFDoDMt+Nt4B0u1JpcVjV0Sah
GYTe90SVAdREzhCRpCniIFKt0pLYtYao1FmtNDr6/ZoKBSHcs/xtWjJrQzLTy5gX
B9lMqivy1w4czUXOaUtbXRUAowkjs30lPjz0o39433hGkq8B8bpioh4MDN6BYXHd
wdjChnHCCeuwcYEJ82P/o7szTgZszkL5Y0X1jtnK69Q77DX+ivlL3Tdz7QazEv/n
vrvONaYWcJd2I69biALy6qP7p3CQJqtM63DUcaE8Cyl2F6gjbMiqlFEcLtyOCouF
Qq3V07l6SWXfMzL3XjUUTlxBHSr0h+lXacuWKa9fzOmvvsWUQaI+jWvdrIvqrOm5
tRlvfSce4rBYokxoGIJSGywm32ozS93vOCZPY2VX6f6WvyCybWe2PSg7S1P+PgAG
hc/8xCH0ttNzwo2/kc7IDSaziEYDCQCY1gezpk3kEsp45P6+E5aJvmUKIQ5T2S5N
geMs0ii4I8VopBmRDKhTqX+TSSZxdQbW1jGYapNci7HSLV/1ZHL0TiSyghFdGy08
NE8B6OdC8gCC+AWACYMxAJDQiXKrwWs7fjgxWicuLa7hJBXsv8kTDayUp1Q9+BWJ
v/8Tt52q0sDazRVwbcbVO51aCbFn/grTHjdFJ5lGpmW12ZjpnSKzJOQpzMYOaaQD
qlIcL6C2crdKX9GbFuzK8Idim+M3/rBRy1Vs/rr9FxvUjVkwyESngHq+HeBwUxE+
9I0vBRq9zo7RTAp1cQiEmpWWgJRIIVXaPnhxdIbNAXxk+M2Z0sDL9zypgfAhwlPI
j/q3VkWjBRMbA8GBr3XsXzY/qzpLeLpxYe75Boqw34P4E7rjuAuH5lZpUITgvHWP
dG7f6d0aEn9AVHG7+w8aD5E9tiwf9/M/zhqocKcHLYHIqBzDL+4KH1feH2WH1s3A
fLOL6TA8LeT8bcO8wO3uHlnyceTbx/oZXF+s1L0jq3IeTut7ZdX0vfzfuefXob4b
Htwp5Nlp20kavnHFSSmcHG487e0U9Bcn9L0lSMn3U+Bd57OwpUaFgM3CYEdSk9e8
n0GGN5QP6HqAi1NKOexNQZNGNFQUZZYTHkZJL8YPeC2kI6S6F8qKAb3/hrEIsYsh
TdfYYrdYjAxjLUFE+xKthIfDZ+47ZGIdErpd6cBmbe6YdAr/USQCbzmvWc7NmvzM
mCVug9a+LL9WEJ3Y6xkIZPCPGpeupC+U2OPVlc4ilcRgm3/PWPVtpcMkiq/BrOt7
eZGjBOo16k5jZmlxi3GTaal200fJdWxvI2eZYH8UI/NE/X4zGduzZnx//Xkef8d8
5EVbq80vZVisA0adIE96JoWbmfD0skpl+0IagHV43XLFUFoz4PUDO2Qug8XqTqDP
uppvapiEonmzbgxtuG7XinRkjOyXXPRPsG03TFldGCmGO1Yfde8XFx1lrUOL/EHP
UFEdEkB+/roBHtL9f9co56arXkXRIegHRvTwlOpP8Tzf0gO5a60gEvNBLPKlIefj
I4iTy21mveyQ4JjbP2wj+lIdtQvFjh5Ujz05zedvcxREX2wilDo/X3YTKmsA5EGX
I+w4XUaqoVzGjzGv2AdH7m/sqadPjQ7xGCLNxqS88w940tIa2l5k6NzHxYK/Tjt/
zMIORwkfPX9JgKx19H2gv1LqzljNeIx+J1Up5FFCLr4xC+XcHzequYokOicIsFph
R/HiTYqcP/3T4Z/Yob68AFZZYwDZdGHZEBDHlWDAFhjd4SmRTCJFECugVbGpQPq1
M8LtV8TpNDTDgCPSTnl7KMIHQQHFbA/qq+udesCjyvoenp6wb+WOazziDPEFIOSA
HbNr4HhRXD1+QW5CNS1JCfS37fBZFbpWcG5ULoyMi1aDU9bRDEZFC6ZV33U44Fso
G/n5yrbv6+zzdDV+J4HiwSE9ev3VbQymOOeiOtujeOEEGjKzJgNf2HTN0h5uW9v1
fi7Z53vinrT3t+ezlPtBL4tDCRZjexM4w/kJ5sbZ0aan77seW9RY2TQ1KOviMEs8
DwrcsQSttiaYpzDmboTww/OHpjMv9R1uwWAJO6edFkHoj/K8pVPEDe2mPqEyU5hN
qed3wwk5XVMtWsE3fYARckFmc4AAM98Kjt8fSXOMSlu8ERgBdHBRLdfspy7+ZrHv
EElACZe6w3Vr6hpmfspmzR4PiCq+ixYWeVuuHReNLxxB2we9R0GKJZg6N4bduzyJ
uFBkan2Q3ipr9Iw0h//2TDcfV90JGoRs0sCGJuwHU3O8/da2Ij1V/N8Ut5qz1HcY
sxuaG/CfHhFxwJOp38vTKNAKxQ042nWbiR5KeOErT0+xQsDN8GWJy2GW8dBx2SU1
Kqynom/9LdirYyWlOWg1rJOUyQIKIjVe2zBBTi+n6p5njPyJ2xH/zD9iNOsAZYAQ
KePSz3SqVbKK3q7qemIjxrjXMc3mleXHxAvzV2Gi7IB+4e1F02TIN0T7qgwqKYuN
SqM/+XnDydQcczo3FARArGBruBbbXGge91mgCIOwC2BA/qKfyEYhxIDcN5D8B1H2
MmUnHCfgKMKEfJCHLt2UUPpY1nyjlHrSbJswtuApv5lcQItJoHxkUbjvz8o2p2HT
euB9r7LuveCLhOyD/oEkSyqNNLqsErL8jneuOB7hJVZiy5K3LGKuW+DznAC8cmK+
01dLGa0DZ90B0Ht+OKEuVyKwIA2UKjZGEmRQ/I1cdlP7DGi9/xua2IIs+sj8JcaQ
FDfj+jd2DER8p9D5s65mxV8ftjALPs8319psduBTs2RSHhrj6tGlQr72UFGN20RB
fmCTG7LdO0PCfMY4hU2dFiuMY6ca9LYkb9cFiVMb2+39/G/I1DET3fTfkc1yZXaU
0vWcZ9PFQNwTbXswW1KxRwisiPL0xIf/xfFlsHTpyOki4MkThdQUYXtrYL5uEUVf
UTmv3qH/G1VqRFJ4h/kyubNQdgPO/KT1z0iBAcNLAMPwxYd3hsxbYJWJNUtkhQP6
cOmHnV4ylzuUmClIXVewOueebdtSmY/ivyMIKqtXBnAPlAdWD3EUIa80NCIJsLAM
L8gHjmAPyvYhZV62G+9QBRl+6OQXX1Kz1mVO4g/9MCy+jl/B9xpn6xePp24YqUkI
udW1mjmi2zGShxiUj6iE2V18bcujPUGVqIOWzopRTD/Yr0+x8jdFVKBhVcB1OPtB
QxBHgvzoMG8DCLCrF9fWzZRq5F57nd27eWdHAaK43J8wVc3ivmNkwvHHxSlDwD61
PPaReZeAm6wbwJJL1RM1LNgqgH5/ptg+TeKaLXyXR1WFKwx6KUN6IziFYByx45Ro
plOxN9sThwpVRg+Eo0HX2gCtdGiKvkzS3Rmha6tQTYeED+pX3PN62Y1gCJ21kMuR
GaNaAOegCjKXR26ex3AuwPgo3h72gYBejRWg2oq6b4ylckvaNlUoaeYN5tYCb4AV
vlTlReUydhn16pKcpMCoxgCQm+dbxFh+ixfchjcHlByCEzlAw1LtE7n4hyH1s3ib
Ld6cKk0t4O8CQ4CvKpdNUAjR+KGN7bbeBGyK7Xbe2678p2XoS2nSmb6JENBYPVWb
ufY110dLRaBkPZo1FokCdvuX3Fjka+/rU6OtIzKRTy+H9YktLaCHuo9EJpQML+SV
WAGGr+PeSrRWMTgHchzIdc6Bo2aHvE4LBOThH1U6ZbIxs5teH2AzVqPa2QseH2uh
pwwLLPe/pGXiKLODNHpErJ9AyoyWt3TboTm51y+RsRLbyiwGTGfe1yJSthJBGSdZ
lpeMTCiVVZuAhxnCjiwH8cK2dE58Sy6jIEfgjZJPwbq1fHyuppWxSwCTqDSAt8gS
SAJJSY9mbXwVmMkbjVuw32vQ48oK3LePpcUlaNgjQiwFBA2QVto2Kw06zV79ladE
RFEv7GdpgRVAeqRhGD4FztAryAcZ4QdpUFPxOzjIm6ztlDp+bjaX+vhEw9qpP5u+
GKzvgSXrG5OFk2BFK5EvDZ22ZyguJD8dqHii7ThnpeXycdJgWz2aSsEhfgQQ3DD+
Qg4yKbd9xYla42qFTRcgsW2TK7eWsyuZebGrcaRQ771wS8M+4H1FrAoyytsKOYym
SYFR2DXM2QRHeyhCkGnwYglNN3XALO2Ave/gC3AnrTeHVRYndoGgEvSiLAvzEwb2
GwTY7xotvYfnKXu7nPn4bItOVtpTOuwjb7IQpCKi1eTHYdtkd2fCwTw+RWGmyqvq
bMtBkUi3sYxRh0ePI5/okrNVmgPuwIDShUrPgzS/wOpKsL3md4w4fNPXcGWbqUgv
ZT68Xy7GvftzKAAdHq/hjX+mv4HVSIg7qVY+f+3XHxpQosLrywGDE16tesG3GA8L
YXSFIAKuJfY7hJBCnXH4hHfQQvSs7FPCHKwUwFxVdP5ySnBhNUS3qW28tqtYnaKT
ukICf9mH8ZSGaWrpyrPQepVLF9CKRy+SfJI6poIplpx+yOfrrbji0MWLs2s7jpwl
917ovGofKEPSrTsduKiyb1LxVQgSfK2jxkOYTaOdhbpDnrAiKpAy9yXTyeGn+Xpr
LV9gcQRAtZasqsUAygZ2XCsaO7DvcYimLgSM7kmYV4WuhBnJJyyWv4+DufBt7VCy
YYfK3SKXD7W1JRuR3KL+4JonnqSLrfPIOHYyY+gRnkiUVxXZ4CGvCqXD8FfjGlq6
h7veX6eAUldbw+j4BxmfjOfvwWlUL1S/WGheUam8lwZAFpG5p9PyI8yBD0mh9PbZ
dpLhdhows9JY2pTTGhTXR4sYo7J1PoC7M24IVGTOxTScbA/1wzVQYTp2cgDV/JBr
HGJZ2DTvwDR+fRp4tdmwnNWqsn6HMGn6EL+EPRX2Ops+k6/haUEElcSr36p4NFh2
POFsIBZq967atrWMmfIS5tdnIQ+BtVdAmODWPCP5BlJVRoJd2qnH61I8FN1B5vrj
30tkSiND+9XgUVcjN6/krdWf9Iylv8pqutoeFR2p15vBUqpJ8jgJS3nGAD6080J6
OamflWl5w01jdQ8uzSRWwHLg3mFLS1tLcPeDEYDU7DbXiqAYimUESuJOgX3XV8nK
bwMLDxsXhKwH39Pjuj+oDarlm4enTXPmKn9QQPUcBVbjVzrY1XmVRSpLxwqP4CaR
fd5u8cWhG2zGgrvK2cH36VVhOyI8f4bTcfYL9Dw/VceiaYp8ab8DjswebKUy1WZe
C1arFMfbmBWZ4q9GqIh0QTwgtQc/nkrv1Dlzk01DufCcQbh2ZyF8PrHc5iZCbZ0b
VRV7JityPawv7J1ab2t+7wvPJuDJVeNBrp2bFqZBQcl3nD6R7ew4ZHES6obL/5IO
0Qm0mt4FJMehn7IW6/gQTO6nWgTIjOTmuoDU9/GU5+E53/v1DQFiZ4q+3mmjbskb
B5a1wJPP95fB8Ww6qsS3am4Tq1zAQ7PoRZTRFisdg7qF0l6uOfGDztQqLszjncuy
4wa5sbce1qrqVurbVcyO6s4YXlTlDDr8dURPXBITpWVyIQt0GmnMyy1NsxuG6NKS
8lSxT8mQ5O4AK3nXfZcBCbMVE7wyZATIxSfsxyb2UJFGD9cnGWipUkViy6SO5VIT
FMFdwzFjtjgDx1hLx1zjYpbISorkiPLyCX9fLQb3HnD2aiyLNEnj7uUQLwmOl1Z7
qQjr7S6WZUXMEsavqU2q66i4ACKxw7jzUSWfdoHJYvqGqwRigyk5VhBmGXPBsZam
U4xrQzg6tZouq7jesEbzBfMwMxTePjB1zxDd7YUt90NpPTL8tKPwwuhkJ5028izG
5ZhUYekWgFS2g1izWSLPvtp7d2m+Ut7DkrSw0sLNFvn2X3g3pyCoqfeVe5a/zRKP
vCAl1z+9VsYJvVWGpNkpVum8pY621Jb4/+VsBktm1YkKqIxLOdvsHQ/MSQGMXSVa
mP2Za2TZ0D2Rf/dOm+abIO5mlHf/BTWvmvhdRRZKPhvf/kltVmNfmDQTJvO7M6AP
obtEhI7BLSvnGeo0TREwlQ5HqZJQDN+MZdXTuviYbQSjThp8n9wF88piTTLH1tXP
bluBaNFiufHEav7cjiXTUJgE/GO6T2WGxiwpwESjvfYRgnAWOY8AqVmwMbA9+Zwh
H+7vUpgs16Z7HrSV/mcyGw/6lWBl6zO0xIsr14F9sQ1I9BhvTr3pZTDsqg/sNmwp
pTlxm64xWJmoXj3Ppb8SpPFA0Gp8X0PTq5v1FNDbQnEfmPBd50AFAQUvXuXt1is+
3REMJB+dYjov+tFdTdPn5+BHeq+T3pGmAd2I3X4tmr3V2pkU0JX9v8/WACjYTueU
Z2O4cmM0Ak2Piio1tPUu3N1Ago0NeJAQ4NOGS7RYq1RHcFAQx57Lg07xafPyTADg
rSrpi7x2bd88/XEZeXuFVo+UUsGDYhnKTJqUQAqf+KK5/3n0o8NckX5xO2CL7c4t
jaAHpezXjo0J+YjT76rbCqxdrZBfwfq7tImOC+lXM4MImOq5ed83O6/AWROcqHUa
Uxbb76WcAGckWCYHQLX4517yn0ZVtFswr90Ld3nWrOPU2R96Gl7j2Et82Und/XWZ
aTeB/mc5XqJpA0m3WKcpOSs6FD2YXZ8Pty4iWJujGgnxVW+YqatadRWtuA1aXfbl
5Zlx4BqTdnSBzJ/TVLxqXbf0O4n859XIOFZZK09wv8E3CjbQtKUY4LmhbqzNCIaf
w2Re1fvbzSlrloYcgOK+g//7JtjR3uDNwuCsk8h1i4qubTBGV8alICOgROL1XNDT
ayBTqdt6qDprL9QrxKYLoFObVXmVmvmYDm3UH7ypeiemcCqUJg7UUA7cagcslKPO
XH0d0DiiCAIlOeQwyV52wG8ozsRUsiLerQeWliQ0aAdy/r0N2MJMRVbAI77GqZd+
FN8TfXSVP3VGrxUmEI2dp90I277wmXrl4Oe4yzSIBZylhKDQmeL6WaDc/iJS6K8d
AUZJsxAbnh0YpqjI3wkvauzf5l0SVWQqAnplXrbJL58NHLpF336h30ry2HBDmaTW
juGEx6MY8KET9Asz889yM7oUBZhLbRBFJ/S5bns/+OCBHqerax5IB9WRZzERh2ET
e5HO56tcnLn9j3RUsHogU2bgIgGmdiXYXuCIc/m6GmMRlJh6dpSbgWGuM5GMzDe9
DyVCmJr/t9rl6a5RBGkIQCj7UlM+pMk5ZXJR6oJ+2lbQihIub7wGsspQWjU0Ws3P
Pxu0Zn66Eh33FYNhCBtSZ8roPTbOe77+AgSC2B0tRWD3upALgtC+d4ju0tIoidwh
iTy12AihXKfxgaz7M5k86+NALXpE0ZFXOJn3qECickVnTH/WH92iXaPXQ/ux0Sk0
mKVEAK4Km6+AzyK2m2QUBOtV+gvh2g5hUIfRNDY0ajW3iriagTN3P4KQSheHjDPp
oMSdQ62XzOeL6QyTPH9GYO+Gs2gmQi+04cPKEQtRWnuoSUD8T+Ei/huKsauB9E7F
DVSVvrcy/ZMuAI8OlovGyOOEqMs6jsfrIX5HXuAlt3asJ7WVqPX4/88LzHep6FOI
yFwvg6pnTus0BUtHfIOlXsDVvlGOJXXR5IZwmO9GG7r0iPlx5izsujIl4S/rksgS
FZRDueBmqnh1bTiefv9TB7NfZ614n+DdpZCxb6tpWr55/7bzJQXXwqsSnz44dxaY
r4Wbkr7gHYvNq9YVIsSJ/JuVrl51ZMXFxMlFoSJyh6gTZ8uGS05dKPWd7NATmrzH
opP0yZHJ37t9zZk0CKNjKQSBjUqgiD7uO2x0BIGGmcE2kqBl5DLIE9WQyAPA1AtH
Ix+4d2A6q3kCWD7QiCw3MVbBgKRMI6qvJtOokdmA8Pq7vdyq8jexk3VC8AtdNgtY
jmpgg5w/H0xyYSm2lzGWeT1i5/oLGfD3+GWBuqPT1jovpZnz3BtAhRUfrqxEu5IE
S2PV7sgb4Dwqx6akTwjvq//OsZzrZwzBgtefx63ZWBozifSNY9P4V24MLhDt6wyC
973WV4ZrxiqLgr3iQSZXcKw/3gC4/JOzK7wVA9VH11/IwmVo+snx3M0MZDvbNkI2
G4sBuAye7aKf2JCHVcdhk8+QNQB+ge1opBnO8GIZlpSc6/zZin0kAAwQJJvya2lL
oV9xYiyIteoD4e4MozPWxPmPMK9oPXd1fRZ+NC+yIYI5ni+3LqkYni/gP2vWEF1A
z9dpYvm+ejJz7H0Ll0NUa5ouVdMgINOGledYR/0ao6phlQ4hqLy1nH1AcGoXi5ux
V6+PDPi4q4r1cwAJhlhQVdo0xVUbXG+zRR0JXau6Q4o557QaIj1WHpn7OZaqJJ8p
fMz4BCVRgDy2Uopm1d4q3u01U1vwp+/cPBFdkTz4leQh6qIKvMKxPGHBl0BGCtdd
l8bBJINexYEQYn2YGXzFMk58+bqnGCv+AancL4hYkBeE0MYRFsxVRNg6DoHQAfjF
7ml8dHRxV3zyayIIZwsXNo7vyZ85nOuTAIeuJYxRO99VvluSIgkBd/vwzjAhJk2A
22oB8W0rGCMGkPTgYQVC2AlVaD4K9mw7XRCACNjH4nKIEYLtRGnBwQoQz9iWqm6i
rhXnvMZ9yGsNLhSasbgGxRr5RQgYWxO/P1vBbwcjiluYc+B2vboqHXnjSEM00RHG
tD1+spt6PudV72A6ipMGnTrMoTbEkgGlbWbJLS8iyB6soJansmkZin8+LPk+IquZ
bxuRoSCbq4E0tI53oBAndZQL6xDRbSKYLSs4zdQ247pUi7o9YOnd0K11ANfnQo0k
pbdUo8Rd6xrM2a1w2jKxNmM4h9h8OnB9W1VvZhlgS2a51pmoqeQOel+0uIqhz23z
EEqmoGcE0f/Rz4enZdaZOqY39uLp1qmD7yfBr8wYdjTnN+SdR+3LrW51ehh6ci6f
cjPniMQjJTSDahTAejajdHfP89wskMKhQKxs9Mw8GrG5iduNv75huvvHB3Kv+j6+
PruwjaFYEnS//8YNbDRJqoLIEqkwsUsIgf7n/kdjEaoWDFfcVOVzzUz6FrPMEkcC
KE44dA+MnNLIO13HSGh2AYnfDeCpqbfx+StFy47LNUwXXMyl/ZaQ2WmJK0FmKZS5
CiDTUgfUBpFcqLvL+nqd/cPeUmwezIndNrYqn+DwHZZyPpWEX5afrEZd9Y97TYa7
9uJ8lqVBVcA8huEwETPg7w5Sgi76NUHPgOnBZqBGMdRzjVy0pCXkFWK133j0K7Gt
pc0tdnE1O7VntxyUwez88H8tqxKb/11jaksRIFJDBwzs0u53/Smu/0HAY8IBmfzK
tUOG5RZn7+Sz0uEMQlMG+8ifIhDoez02XQmRNem7d5WaCm8nLXOKvRNnGxloMril
0033ooPLCqTM1Vx/YPMA/VP1f7OPibFTbFVsKoyxCrTIDVv7pdSTGyDSYGaQhdVK
JP2A+DDerbOUjHCxGobwpVf05MtInHTeQX2K/CFtLMyvIlaSjShxYL7IulUzbrlf
Yeq9IW7z+ShQXDFXyemt+XWH4JJu180+pWE8+REv41Sh3S821Yo92hbPASunWNbt
5HgtYs/b9JaMJsgYwXN9P0bjBNR1zS6fGuxmoWLk2T+YwPn+bAOegT5+o600CJ/Z
VfDWPBD8H42QlUIWcjV7qHCk7umBiAaj8FS0EOh58u9kQYUiGadiXgidKrzLMVwF
NSZo6jhezQNMoZ7ecloohNn5oyxWG/cvwrmhTDIkMv+olA72Tq/UzSTRLwItLbRk
ul479j5Nh73ctRNWH3YQ3UqcYXMrKyG5OzIw1Xs+HkYhyf3JrilkETQzWsnX+7Yy
Ty47op35sA/WzXVwurkU71JC5bfCiJYyNbq/R+ZoRU3MvK2OF2hUyfOmfPe+BL5x
YjPs6dIlUxq9KoPJrXsB7d74h/5gtx6vQ7xwxlwYWX5EkxncA150yKQcPIO85HlV
U24tp/zVcdmaGhRzmRwEa6VxOnY1Ry1T+1C6xFUEqt5w+HRfy8PmL/Ym4+R3jpJF
RzK/JWOuk+RQhoSdjYeUxmCzG/aVfmfJPolCRdKX5KDh9+CmnkGBTtuhM2imd+Nj
Mnkju7IXWATTFq+/UzeKvsAo5LqfzbC3QEMEs93snPZWr9VBbhrdg0IAeiW2A+Ff
4Uyhx8yIWsHIoK0I1l2Lt9bYVIOAPYvMkwQOgeBdlW1sf9Gs6kvNG6pXQnt/uHv0
WznWekLTQxK/L9pGyBNHwnQG59kqYWnmFODGbIlSgwVkS8InK5nPibQ7Hc9HBSk1
LgVg7OBxLp1iEwVCNpQUniectarZL91ovmtNemQJEbV9LGjEEXUYczAinWp4MRz4
htYPFXtvde3kNla7xtnaJDqqfr8kRrz5j4Ulo7SyyEn4+R8Fjli0RaQHKS7D+pcf
msG//eHqUfid7Tr3kkBQ0HzRTeL1pQySTAAi/52fZ8oJlYNZecARLcU1lrWL8jbb
3T+XygglUk234xpjyql/BkZ86bKafGfMJXfm4sHD688uUerPoPBS9W320ehUcnB1
b8qKBp3xpcCUHDduJ9ovCxhaYY0NgwvAsjR/kpIRLzj/ObcZYOPV/sqYEKVcvSLT
6sNJg7EChr8HOCmeV0EptF763cpU6uhpC15sId0Uunlo8Dpqv+IdtQ9P8SXMmYfE
4vNv/LvMvFAl/GqTCaujUQyrkjEK7m+CZUoTie66qKDu8LQMZDqnYXCQNA49/bO+
u7m0pxHQ4PwoUF8e0GksohErH2mzxmIFvhrZb6zbBtOzdej0Ywvp9ONjgKLJrdvY
Wyd1WFhJjHSqDWXwx6lYgWQTyzPED4DfxbAgzSdIq3Pj/xsSXAhTbvQNrvh7yTBh
m5Tr+8JjiZ+hH1dWWzdyPpDgkiwmV/D1uk4QUeh/IjMkZzvEk5S1zxyxW/PKiKdq
OXIUWSr0jIGGhr6d2QW7SSMO9NVFxmqBQGe8KpJ8q8Fyus4EXMN1Q5xfWku0/Rmp
Z9HVOAg5mmuHTVv8PkxbXAsm0ghT5DDPlS8ufws5G49tzQpvbwEy/so7p0ia0rtM
ZLoHgBWIZnZ+81y9KPcORAmu/MZVtY0wIUKtS39tkO8LrfSu8xVZqLdx2kkZQARw
r8okRbbvoML4W51/QvXbK80LxBCWla+8Bi9tVeWwC9t+AZ1+idOEXkGR2GUb/Lx3
x9hPHk3e3cCbe7kjaV5kOWHFLlIrcLbZPt34rh8r7oDEAGy8jxXO14eHJciVsKTs
fqxTWhU8+p9No3LrHfs0BeDSeNo8yigMDeBjp0fLbWIkvV5RluAg7emGF+EEBNGh
n32xxFRfRHS8V9mAu0SeTx88LJdYjxG4BWfh0C8hQki7Z6Y5zZqSDZH+C6sTBPM7
1Of06HpmjF0PhEWozTX55sd1uiApmclPiVLvCYEnzUWKL4nWLQAdPnWMZaIlh/RU
Cb6ibjIt3DIdQf2w4sCWOMguDOq12SDTfmadWL7gE/oJyx5UxtdSDqF/EgNKAh0f
kKL7UeLIGYaby6q5x50QQIaD3/Wv287c+rIkh7oC6AZStjAuVykzKNK9jew0LXOv
7TIoNIs4OdPvOPyNxcf9kH7YxgBH0qGF36xpYsFVIO+Zi/NT3cLyUEe7blLQbduw
b5mbHFQL+Px0F/r5XfrG4ULh3BL3LdJZ6/DDxdtIeNfFMcshBJoy/9e8Lph/zQ0i
wlSAlCOVmeB2Y9BM3CsZQC8o29ApbaRIoQOKQx+yLYCQFYWUml0rCokbd3MFm8dF
/uRqgN6YVKlbOi0lenH78TqEGlbF99vPQpDiHcZWcvikzTtryWhq97aRQNIIkwWS
qxLBfjc/QWS5T2k/mpIucvMKU0Pf5Ud5GRRrs1WBuVXcWKXNVF/3TwkNis15uHxW
NqpNKXvtYOR8Vx32BWe+7RWMNBMZc4R/4B7qlRVnp4d5P9ccA1S1Q0B+Lkq2InPP
YS/DRua7QRKuWeDydbhwgQY7ETPy8NUcLp65tg9mzFDwXgRqCQ1GfKjAri980wlP
G5OYL4a/+/X2aqSYv0d38+Jsl6BwywrbbZjyVhGP/n7POxvXkG9yiIrt6uo2MpK1
jwj6EyXlfzsBWBIzwwTOc3mU6reWl/qqjK7Cq0kXvQLb5d9I6MgluS6hsROHBZmn
aKQyMXU2Xp7iL20I7RMIh68JwZb966t/zf8zsXlg3S9jkeof01xyKDenllYP4Se6
JMm1aQtGzturxwhcCnr44kbZvGBjpEHYhAYwAfrehNeNAV/+BZLDPkzpKU76MDtN
LHEjlLgH7WhXn8eH9dHy4SR1mzcGiJSQsaDa35Ig7qMgR7q8Fm3M/DlumraH0BB6
Zh6wF/l73TQ3sTlYv/Ml3m0duhsk3dq/9B8QWwOixkPdLZ0G4pNsyvlxzJVIgWOv
SssOL1kdUtxj/LB8VaabtS2Xoq3V6w5T7+c3aH9nNAPW6Xr5/D87bHhOVc7Dc93t
lweRyxgEO3dK+j+Fox5Ztn5g+rqbP0sBiGOAp9dn+BpkLgv6ZG3VfkjtGTBs1ukP
3rZe4QwbRS98eG/8l1yYL4LU0HbCoQHeR5WtWLjOFUEaRxJxWZcd7hJwiIowCMfm
GHRk5tYVhIKw6JUWydoZoMH8ZzXELBVz5urYbRXSg0HbhuVJXro/m6RtNPHSP0va
YdKfKGpR3tepZbYMZ8FjPIf9EL3i4Ichel8TEptC0/tj1xungmy38a2dj3NZwABc
ug9JErqq76lArC3S3XqO9bV9CZQOKSwrRDjUHv0Xs5tzVIQYBd2PsKo1fpRjSJXO
7Oen6fYc5XNvuCa4V8uxE66qJ0eeCisw5uWJAZSxbM7XEwE1KVR1XF9Syuswywgi
SYW5SEtCVWq+S3pCyTYU+cYIc8S0BKEkWw40NXl4JV/X6NWsawA2KirzhgUbRgwB
AS+TKazrcAtDbIZmI5YdlPvsugBTMI5INS8VkCGvtCiTP/A9/p8fouaSk8VOvcO1
220ua6m1b0xLB3zWr6ba1QspVbqgtvNBdKVA/+j7uVTLE/Z4+D2HchyfqLEHi2fX
2yCft3R2SgIJl74/v74ZoFwe1lg4L58PaArXV0TD8Qh475dLwAZq8t6g8RQcPhTe
sibrYojR+4vmgQDhBOspnLR6VdRs+8xfJv3ifoSulRp2roBXASlWhxfl1Yt3uLx3
DX+4N5ZeJt/7MzzvFHvPbE5Ytktmb7ElyE5LP+sMma+RabeZfISUahRs4F5FkV4F
ZN53tz95yaWt31gr7o304OAviXLzZCJPtZ+a/dT0eUBCCMp3Fma84RAW2CyOOWHl
vf9v/X8eqpVObhAS35VSpent8gH1fuX2V62ORevsVrreTqRYydSlWeARiJ/rZ94A
n3FZIjMQD55G/uLJRpTFBxxvlbX6YcD0DAOX1iVEXU1C8q/VIiIGBu12B65V1Gxo
DEc0sY/RYTlh88EA6lnak4AGA36sYU4UezVa5zvHDWTogO+0oglaGA2dRrDkBJy7
eaclj0/lalAWJ/zRo1DY0sDCzG0jI5JLwJAaVuGQr7M5o6vaKEDq2xmcSm4CmUNo
dOWld8bg3yXZaBLGWjeBN/C9Q7QX+rGZqOL8Cl5OcWnYTb0KXqEDyHXAisuHS9LQ
gYH3T9UqCRg8yogElVwvVeK4lCsh8yvhMnXKjMjYdKqffTBC+ZgwDh3mzJQNNmpY
wPeyi1sUDm7YoP4lekoUpInZXY9ly9KfIFkKBZhqyllzU2kTQ+GvkmyvIDggPgn9
wJVVozU7Mi9ppcamE0O77f0JE5OY/zCMa6MwJ5QFOs8KRNAIsoBOkBzkVHj6EEPB
hjm1wS7Kxl2bKa1+AHgCUlrg1AaF/jGy1V90XRhFnCC+AlVm0lw9IfrKhR9pg0fK
cZqijp4oUGiQXkszl85sLzF434zKoph5CPTrAnf5m/ZEadI5KCFNWnnNmZlvV8D5
dBqGIYnl2KKR/b4VebssXoeW2fGzAuabDsBUZbke/gw3WZ718b5VZ7LnWaFQ9xXJ
aooufgZxaJmLXxlFJ8L0IxLHzRyccfOPuSHdVkAYuzeSC6ud585OFMwGLJwtLB40
Jb+BLzoWgIXnH/N+bp/PBWNRV1EixIK6mmnU2krvcrcRMDoFpqvaA5cse4QZ0BH2
qZ2JotdLr47L8E/sx00ZqvDp1x0ODe/WUscs+keiH40iJRQGuNdG02jt4BSyHy+K
6m636uaG/cQY1hpt7L2hBDq4Mu1yistL+YCKgKnOITF273jbtc4m6r52ZBF10WbT
JhTaVpiKNbmsKiu8/zzQOh3w/s5zxIhd6LQgUDDNf/Supou+hbuvwUqurk5ivP9Y
bcaSE04x4xYXNY3ca6GWS979gxiGalFibSYKXSVifDsFdRmhrc/vgG+Y6jQfD5de
CsPKh46IwZ0odyH5r89aGZlBqR88mKN9DAtip5tyP7bOpuBPh0+eWrTb4gZoLZH2
2J5WQd2JwbNGGbhk+/BUDwCJA04zRlqwC0/1sHaQ2TtbyBudQOkQMkGYzxc14auo
0/NCKJLnPaQbsPd8JkDT73BJsO6iR8d6TW/Lr+GvgQ1uH3VzVZovELw+ehrXef4b
dxe7H5t5eMYFnah48vX1Vo4s/Gap+yyORIMREphL63sWvO3qEFFSBOcFWfqtsDxL
kfqAmM68L9ItSXEJHFrnJudRq4dcEv4j6qTLWpy1ADEZA+2H/d4ygcQMOF9H1SYe
OkA9xBy7f2Unb5P5H+TsYXuNwIgJ/8ajAqbbfVG7YXMhfnkHtWhn6Lf1A6xmthqp
y4SDANtghRXENjYzVb3c8cRgLhWwNrAY5zVQvjr6CdGC1dvQUekZmxDFCyYBo7m5
FfIIluVDDDdniXqKF0tH6JCOujGeedCnwZ+9Bo4RwYIbok1dZ+aUqTUUV34agRCL
WZBwGM0sK4BcXmX/lNOgObL4tJfW1vG0CUFjipcxXaLks3QSmzF8RdmvM2BKhuNj
sr28pvunHfOZaJSKkglfvRG9nkebpyNGF3GvpCwawewFFPT5Vr8MO6a/je3uZszl
uAxSPwgXF9PtRo7ZJuHg1I6sibwEzNvlXzKh4JVOr2LlL6Fzj5JgBCzQtl7Gg+GB
IbHLGeaetRtl2JYZjoLziobz6bLltrOmYf5r4tg3brpakbJfUvS8A0OecaY6SeLD
udnesIYdwAFWNxHs9uImVlnhkzThH7/y0yAYhYYai7MoEypWTqEaTrpZzbwh14nq
xE6Bc7zb9e4iHRAHzqJSDQbFuhdDVhmoq3z8k2ImwXgkhUyiIqwUoc0JUQgsJa+g
//JbQc1FXfn5LKQJPxhbuh5uzbpTveIyLB7Y4cAkG7hHdAUhIq5ZlYuutW9YO3v/
OIgALixpbj96EIzP48WMN2liZdgrGZz/64zShmkmSEWxAEfbEJpxPe5OvHMV0v2p
EM21LnLgwcZbc8xF29Vg1GpNj/yrbUjSIJ+VgTTIeKqQwt5U4DbMBvWR5MbdJyRR
Q6CRE2OPol8aDe5m9jhYqae1+yK+WRwV3pkxAHluRypg2M8LzuG0VFhVDI28+uLs
cVdHdfKHYamaKViUDKkDVCoA/l4x8hjGndKx681f+1QmzxPXuxpf/L/LmNOsW9nS
TQHS1yGgjHJW/S6sZoG9zkDe3ysv/kQYQSA7QMXEMiJk1amHc3Ay/DV48LCfjHDt
+paGogGIvSahT/9SpHbk5/ETixIgQstHQh6ZTNQBCFNM/pNwzl1XOQPVlnw0ISK9
bRZRsFgUAhNOFIdxobskMBqtFyWr1SLcZXj0g8lKwEsuQgs0fVeQKmxtDNhfmNto
Dgep9xBt1w7bI/GKILTNK6lKvCOM7KUT/1ztmjUjMRHBYYzmaVr7G1CMAT7XKZa3
KS8UCdLl1QxuL2zYUcpQ4MI1mbjKMCKZFL/2XTp30uEH8q6KCFZjoRqKTw/RkMQ5
gaf4LKUe4D9yY/GvmJ8XeWASe0fbXGeE5tcvfGS/PTaHzgV5bhSsnw0xN9ubprKO
pa1+lEpLIB02FpcJOt4zN+iHQ8m9E65FGUph1gN+yWUzmmdYInCANXyUiV88ElRn
MbSicjeJPDSrEZoKcQ2wqgqU5jyC3N1/HcSf6VyFOXMAW49UkLGH4T4Zmev7XUa9
Pk9mP3Nth6OHULug3xtGW+J0C1vHKMMLLSLIzULvgaaFpAfqp3en6kRevpXppNDO
p7xIMJAgh/aX0kTjqTay1+jEwazRxGXfKrOvm4VZx7mtXixfMEvQD+zMBn1X8Srw
RlJTtPRfYwT7okQT5+cjyNpl5CI6CeX2d4uToGedG1vavA2eC7d82qMy7rj8JGJ1
aTVN2ePHTzUO5vwcqns8b3Y498l4k9gf0DBvyncqjxX4LjGMlWXWR5+zrUppT/As
3XKH98ho1HF8Npiode1qA3++Pt9BQn6bluav4MUiteiJIBB+tItq21lyDqqQ9Vnp
MwLOMGGYIsX2LjMw5iSTWeBOMLzEuk2u+IT9GD0nVkHMMwIcbBe5RggZxboQzaLm
IHkRogXu2foMPx6hGa62E/QDX3USJxiWyaA82DLM7bUcpRI65SWXIo/ff6EBtKud
0ur5Auq9fGuttoVpzyP/Kjd3Cm0eZmWxWkp9IX7eAOmaiCV0soY5727ZMyn0Euno
HDdZPrkSXTlxNIYvHTJil7LiMfpFuc+DHn4TkMjzDYiQVzyyYXtMpq2LLcR70iqj
T/XZhe8arLNmaa/D23wAOS6Vifcad4mJK4zgl5qy7h+uDe1o09qN2ex1x0mDojaM
nP9v+hBceZiiGHuz5fq0I8zmzVQWwkssNVmQoqu7C9osso/B9KW6SSzEcSk9dElz
NpIdXy0ArMd2YiI31LswnLsKBXzwzSzLJQb72h7uweLs24TR+H7BxyjtzciPsFhN
libKYlYBJvGGgehkc52Zu84UzIY2LYQbB76983Y3jguZzqfbEHNzgmlLdaokrqT2
1Y6dxxITIQ2yVhbTbUPgZb+RYju3oJvaycQaCAMW2KF0O+dJxOhQ4bMhz67oRR6m
pOGa9A7X5kLGkoPX3upgWb9YGqDgVgwKkXrJY79pLRvHxvJc1rBXaU5eMzW3IqEC
xLfCNYtNTpq/Xj7h5rYPX8CaLEv1KslkshnDPD8h478OPijWfYiaWsHoes8Q2D6h
24st3Zlt7N2Gh+dz/ft5NZiD/pd0gyl7ZdLt0lhcXyLtEfOCHmLt8PdIhdgqqJg6
cdmVKy/Z9FUTG9sjYiuOnzQQV6Z0zSX3GPD2yf5/WHAVn5jV1RIDzfWktxFmFDfb
ygY8MYPW1AJC8bl5qaZpfin+QWucnyczKbEuNEcatqUKU4wPYpwgAthwtscLPfLi
Ce2JpT82IynOR0qWtwJYNewnU8QczjViOp6rpR92cyedoLJUtnsqTUGtEZ2D11od
XPhMXqWtmrZB+rT9LuXaVDOxsoQznmw1rmsLWDtTZ9bvUW2eGLMz8pOmC5y6B78I
/oWR0JWZmVDFku5QnKYshBv8iVDzEfmSEhkgvc4E2lcSAuqQXmB212kb5rhmz6b3
POd0lD7Ia4gl2AbVaTE845aa99XzZKIpv8p9w6jRLCv6jrSui0fZ4UplXDGqONko
BNgveM0+8jnKvAQYJduuv/mu6sgUkTF4XOAqsOrN9l/fgivD+4xirIVujG5w3MW+
eYoqUDCwLQ5iTDULdFAHad8tgNMjV15j2wLR4Ov9I8Cyp50GBz1oTwxdFh2zory4
i90RJk5phaLxedRd/9u9iOjizR0CEoUWmq0wv2gqMZoh0Fnn6cK2kIlXOGnNPe6W
lwMJS7k9+ElT1jrNzGy5qdjhqU/vYSvcMuOqp4/xCVrGL5uFx3UzJZP5rp0SSLhQ
OqofpIs7L+Z9tBpL/PT5ua/zmnNDznMfRTZM1DKvrFqHInk+MTDlCOxhFa0704Dx
xjaLJLtujjY+TLec7E3EcDLFLDKg8qXrHmeDDZR5OATcQLcwlNaDoaqEA19qGmLY
5GCDKAh5E1zZKxMAmW2XWHqVFDAab4VDLLpqBVntWUb6mMKvKkXvm8Exj+DTqARk
OqnpADihcZx1Zwk48z7RmCO6CdJ1T79tCeN6iiEGCU943UDYXeRoyHwDoe6wvh6S
VZzXg/AOFcAIio/UAzvX+OljA0F8E194y5df6b6twe5bsfSBxurFnd2NVfMi4fq4
vVWzfRDYKZzzlmfgmHTZ4LHiAUjF+Z31zdroGS4tdpQXv3keWPyTtsCq79WNbvw9
EtE5HEwHWUdPuHXk79ls1JlbNkcVMlbb05XZAhPLl2DRUDhcYkz9LY1owoHdYz/1
wWrkIg25rlYip8QUXxkjJHlytV27ih6SpXyBQposROd8VbRzzdB1Yhp9VwKyqL7K
3fCnVrHc6GqK9cIFYHtKM/P1SAaK8d9MhnTuH88uaA73iXulD2/AgrVuuLLwSQXb
hIY8hIRoDfHoHy3rRjkHdxbcjHHE2pB3CjHJgYOHJd40ODGrjnwLaP9ninfQNfU1
ZE/eslCl0OUHGzDA0Y1Amgty8jHH5MJ+fq8HuFMpPu2NiW+Upr2dVMDaQ/R23Mep
ZblkO2p/TFFF/y56ZCPLnQc2rhDJMXzy1o5lOCT9bDyB9IzEXGAiYOuNZvkaUJ7y
9eXTB6lxZ9W9qHZxb+BZtZH7SvUlXW4hoSUE7E4ujPmb8+bfOOEjVInyNRLYBs79
S5WIMuJGke0vR4dqHM18VeUSpzr6E01KIGg0jCf9m56hF4gMTVngdBEU/JlGyzWT
mVMgCp2uIkKtSb0PZ3UmNUdSUvrMjcbJ68vifgry5E47kOrpz4C7vV1t1ZJnaHF8
00rr5LBjkhP7r2ZWxgJFcwVVd2s3snNnxi5iGVZukfwrf/vSBAiJwjwjxp7VygzD
8R1KlENe/zEvlGClDjOoJ7f4vxH0qfzjMGP370dFwkRRyagJ4cZTtuMtaEzz7cYV
b6KWOHXNCov+JSh+XGrr2Sqcv9bI5/wFF8mtNBe+pi5Vz71/ntEbxx2i3FxjHN0A
yc2Zxb9Cg7c8hH0o75tIckNzpmHDbbX0azArY8XBGEW6qthTV204T3U7SIA7qxen
nqHIusOIm+oC70WgzvUSH7/2dertHEYFB124kYbyrn75D/3v/wEky/XnnbGHJyfW
D/vkMg3xQhG7vK56ZViwVvkhTVeqyABxlviglodqhNcnI8qU5P7J399XL2TWDG3G
y85bWiJatLHcJAoo762hfeJPQp4GSg1TsRDSDrVhgXsSGiOw8qDfvnS2wcfbypS2
BcS00wTendZVx2wqZ/GTfgu/MbNSYZKpeVpA0tPUF3u0KSd63RWDg+n5mF5PMW+7
PyEmvOX5lACSdk66h17k01AA6zRq4JtIAWZvekrrV7c6uN3qVnLFkxNYNhxVT61z
/12Rwk4r97+lfQXrVFF5Zp0jR9sNEeNTs9rAj+EOBfqiNQ6oIQH5u3JRDv0nlFAc
WQNp7M8LzdKNNo7mXHAxt0hz0F8g9WM6glMq7QSYuAmmwLM9wT4EMiaX71sItUTp
9gnt26WEs3R6T0FqudswV6Rp/zF3WeA6wPCCrQfXGFSB8cetMrDa5rtDsbDqDEkf
h/vEnh4uycvHyi49Ff3HZ6E/RLg53LqfSyOtl28h7kBVho1q8onLVEzzv6dr1YWm
WrIaG/+AaiN9BYY+Ju1Vjf0S4+OSpJ+i0jp/XSM7Vwuj6EXRnA6yACPeykbgNEBI
1hyl2hTlbX/JxaYQZmDkyyTgIuYkoaYDa2eiUKHoMeXRvE/WNNHBuJTZJMfCW+2t
ZgR5wH/S41pSD/LLOaagobZEiltg05aaR3UFF4CvR3VEg2rtbbqduzwehwV3/qvo
qyHno5Ov37CpRACqu66rd97zzppSh3iaryGotFp9tId/wz9kqjVSHeUTD6FX8W/p
P0M4hJM8y/qoRKcwgMwds3IjmtWUS1e5cnoiT6eL5DdM2ioBlj1y2ovc8PgDWnMQ
Wg7pOnUlCNLi5VeJCyEQCJImD67VISnAkv5131lOm9lXC1vV3c8H/uKY8K9n1F3j
wE224fbEL9pj7+OAjl7a1Sv+ZfFwXDy7+0XJMxCfHaiWetUJHPlRsLi7yVaT5pfE
7jfz5KLiZwv2azSQJg+MrM4HpMemTDo9WS/UOp1kDasd/7oFANe6CIPFia2XLWNB
AuSRbv4lqvJ/FodIi5vEf5El/bR4S23caRg4sTgNLt4p73kGo92bZqwLlPVHitEg
0GkYUKu1zXeiSLmaeKywS1OllXp51Xsu6yEu34+XLq8Kfv+FEUmOjEmqgeoAeYah
wGbVS7pUznRZkcebHHLvYsOmsBfCnh+0tqrbCCPzitLBsFPctVR2+wly9r05bsHA
bAK3uHmcK8DsWR6mvmpw9KkBN/h+LI48JOWuwrYkHNS10VR8t90J5wH82mEmVUJG
Fo14UlkNtYPNnaFPbNEw0FedrRX5nenzBl/pMtUqNq/IJkrOo50U2ytdFVKWHtAN
W7muf4WkJvHFFLgvDRPnaT5B+XA0vqTk9pPKXlG8VE5BvwGjc6GGPjoyOH7REONN
/qpkAbY+fZZsOxRRKRG1SVgm87lsQbRcrMxr1dOBBxoUE3JgYbux+yuXc7priFtw
8aVfLGKO3Yi4pq5NEuzJUi15Pnfh05ik+gH+Am5OJqw3J7Wotxl16244FbhR+Mop
zEd2+FBXosuL4oJQJ81nqLqNizNhjACMeusqwtRhqtkJtaSMrSxQp27FYhwfa6xo
O1uNjqJOcG8Iu/B1aYTRrEiRW+eQckU1Po+ygaVy9t00K2FcHKWUWqilgSHssgK9
NE0Sn7QlSdP1uwxryAnpSGP2i+13kVIdfUmmSrfrwEQkw0E6/IOcCxj/kOVAnjKB
DlrqBMUn74wZG9TSFsGHY+OivUXn3V6WPyk7jYJIb3tpha5D5FniKkodd9IwGvt2
mWcYY2FpLI+qz7QVKaAtMppPmPZf3OJcjh7DEOdhozcs7QxnbqhBnV+s8PRu+YEO
Afisq0+9AgKwMPRmoHJiGaVZgvcQPcRYmSxx5V0ig84MpBQJnjkl/g/ej73ts6wj
qg3AZJojQSL4uUHP1R1RiPFhln7BhNOs39rexMVAtBeld0f5DMFyJTISqdXQFK1e
Ti3aJmDoFVXujwk2uXGOL/AP1r3rEXzTK/HnGZeMRhEFhBbRHCqBKDq2PpbeWgxM
owon1P4xJ0OtQbEI4QqpUxVkGSPcXau9rRaUa8djHSRWaBcx5l/2C5W7vTBr3V4Z
7RRz8+4pnNeOzkc8lDc9v7BEpXpgTYhbCueV3+GeEdwtt+FveAMjJlbJRJ7A0zQe
mWL5VJmeUIUmbkBDs7W2RrnbrhjUcEpsUkq5apwaZ3Y+Jm0Xf6v7zEUe2gJIl+yj
3M6IUDIpxf17HlC0VazqYQqKwVyA4p2UvsB+2tnoBqXbr0zPnqvK0PckTWS2HKPn
eWo3GBfYiYJK7W/l1pE+gv83FedXiRzSuKNpQGdJHCtsRQziTdGo4L059vvNWE52
upYRhV3CCQDZl9RJd8ov2WEQ03txXlTxuAXoSH5FDYk06s+lr7/5618y9xQGVSZj
6Po5JPxZ6235J8dmzxZYr/+4cmNTnTQWu/IYlx29f+tXqdVizUxeLoLyzrWKjr5k
nZApT7DqZf2e7MXw0Kc014d3ED5mnpBhf0vGrWz5cfTon0DR1A3JS/qDLBlmVMoB
W/Zs4Zocb0rUuS6K5LVuy3S5FPIyWnR2v1Igg4FLqoAwXzhSB/igpc2ZSDrBf73W
gukBYVwwONd7X9wdcqeTDbSfmfarwpR7puecoMQ+spoy3AGjnopnv4PR3nTilSp2
tbNlnaNxjXkMngF1lhR+JNUT4pN8Bdj2pKFAj9qXWQMrZ2g7zWGpSc49KzuccaDG
ZD9gbRvXcCTFPVeu5DKTBTlunwWr+/N0qiUSbGRCH2nnaB0zhoNmryFQneurHEtC
aV7MWPUgX25XuN+gMRfkKXOEo+83oiC7lNwGkVia4gB4iSCS27rgdH19n4J5AplY
oyVinGYc9N2J+ucmrn3dg2nLgsfhiIQC+H273s/ExfGLiggFePm082R9G6ck3/VZ
cLYv4YVUyFXRZ4z33Yq3TC82SXF4/F3gDMVJUtwCJ7uW9t6LswwwjmNihiHHXKqW
cPDoTxDopjnELvAO2xlLACxp4b/xGMABcM2MpMX0Xf2gs9bGlwApwhZxG8Epm3qj
qdnyjO196qyy6wV6oZDszUIJcQzgIxtwl4sdfubFfybQlvLWCsY6yxPBJy5LK18d
01jPXbdAXFqkmVpREb4YS2OD0eaQ124aAhDrXboWg1tNy/8Fn8m9UEqsaT4ibYBi
t0ZWAypuERUg+cFbnOupeIZfHRwbXDBGK7d/SKdfSVXmOM9uVN7Psl0KoeqGqNcE
kc2YLtu3jcrxCAN9JlYIVORzf1csKCa+6PcTxSj8H71W6aZ2Vh2A6rQ9cVWdfT0f
s+Q1bbJN3HQVhVeQnsBpvw2jttaZPdyauepkoZSloW9yolgH23CKK7pa/2vIQsIV
4hroJi7r8bCKYCJDo6BfLOgJRip2dJCCWF9jjT5z7toutKvDQIiz9w9zS07iJ7uW
dDHAVPH0kUSsYekgG9V4acVlUjAhv3P7sk7V2TzMKtzuyUbaFa7Jvd0N2U1/1JJy
zHVeDoZk8ZFzsmvUA8ZvSYEF8jepZAppsb6vR0Y6C6jHq0m5qJiJOMV08t8RAd1t
oDHjU1df8sGUydST7BMVSJspO7HEarY4UtsFx6LcH/vXwPju//sjaOQgxLb3uCr0
PxVl4H2FIQxk34sNzbfz19EpxzyieY/JHhwpEZJ/KP5t2k8dG42xkqr73bATYbDt
lmQ69/w0dZsR7ZdQ3WpN5Nv4ZS8Qv0AkOXu7Yq8de+9kN5Xws9sihX+4MzJtypjD
QW1pcJzI2m7ey983OHDqssNPI/zpY6i0PFnFtRY8f64C376oVQKdFHbCNgbdn5ce
SiYiyvo0sPxhbjeerQgrxuzUixmAqcPtHXZLL2fCyIEhzQRZ/g7B1PFcZprIOqfF
XMaArQvgGzskIKYQv2isvo/Co7QvHZKpzOLkwAZ0KgSfvQxBfosdTHqIkygMepWQ
pMns3Ut2y1ik3R2ygAXOFgR1RSUCiKNN8UfmEEVcwujNiGSpOuDzW3GkOFi7xpXI
DyexVJXwvO6oo7yyxAohad4r5spuAJePV4Q1Jk3bzrYVXZRLP9nclizwTektPly0
tEXKI+YMcHgNsPvwoA9EzmwGyH3Z66yhL1LUg3STq32Nw5VjhQNMFbuF2X2X/lHV
V8/BWn8s2idna3poDIN4Vau1qgQHmdo4EzWReSAGFC/+O8vfBgbTbfPRf0kHDiDq
kQMhqV16zz2XTQ0Z+UtIRsSN6GxRgr/set9aP3yyxc3m+QUDCDQxrdTH91G5wAYv
QG2018FrpaaJo5BIhUXbDf50TXNizu7AucpjDj6CXXZ8Ff6U9xfwRIhjPP+FgTcw
cDDqj5Ag/hqbXJYGV24OVcKP0l87aZRa0x1Zm2e9nR+xJXvbfjGzFBFfwyio1Cq1
WjfAsPvZDD1Lw6W4ZNMz9f9a5nxiukiMUavrfkL74Lc0NLUq2Ep/wulP4N/aELAe
HyE8JHl4t2UCXOj8SJE76o8MGvJynUhVOkcFnrGuXIx3s6z6DhnVnEgLgNzACTVv
mvf0j8FFU3NMg4D/kDSAaRbG7Hh9u6YpLN+Vb70ZTdthJ6dI1G3olqfACPTkPpT2
qSDKqMn4q2WZpsFrx+KAjtYxC0aDUB5YDPqGQaq9BhhACot7rZK1WOIIyFqAG9x4
EyqOvepSa3Wu+TO1GV8V00ckjEg+xfyzHog1oBQ3nf8O886SNKk5mf+biOuTaW9l
ODTP0rB8I2lr6M0c1WErDC2yl/ImAOxTj6sXsBzaEgKaN71SUZKls7EXZ+gTRoda
LSmSqlmAILYTcj3DD8f6f8hzC8jokJGxIG8eGVKxx9fb1cXVa88/yAxX/GZ/HOnC
1vF0nr1PWjkMZGCwe49/YPQlpuyj2HdXaPhilAarSlUX6KNL8iOA8GNJhWT6sAP0
hmYG5M3AmuLXXmK1iQvaeWxb25q4QEmnWU5yBsVXH5mYQZAw+2Wr5XALG1OkzrtQ
4AxkCNLF8YA/54ELu6C1WepdzJjTPeT2Eed8DLQQB/rtkCVoqoUgubu9QOL1bdHQ
DC1ao3W9sWA4ltn+RsmBW3/K/onBxzKsxzcD6hdhRktGNuOFxxeN3EwnCdtVGIhK
21GxTkZhER79Y4XoiYzKPst/N78v3vOsOV4Oc0XvQlwOLrzRDGZCX7gUwYWxM8H2
7Qibb0m1R+Xh6x0KSvE/Xnuf+Z1UQhXXFXiIWIUS9u2hvfjJ1tHSVJTJiuSrFIy1
dnG/etYoLx3nS5f98TC16A478krMfVpGmG0Gq0Qpzk6hzxPB+qzEyePgJHhfZXXE
mzfVqnufAMGnkOrpZNzmiEJy45gSB6SB1mbSQMG+4dUjpmY0a2FQ6mptvRVRM0j2
ic5H6dc4ZlG8XBalUF6K1tcY1WFCrdZPME9QwTVdDuGxbG2vhDAqR1P72jimiPln
HKqXCZu2b0MKPUXAx2TN2i5ycumXwJCgKCNHvpjd40dYAT1DPHoBVdozpCd1Y4XP
5tGl/uCD/T7e++pAY9YQ6lJJm8L8yp9pQriuWd+EoiVdT1e4gTkfpRWpn8Ro/YgG
LSPZjNxUD6DMBNqiC1QjeNrTVK+8HKt39PI6P8beQ7ZnUtH40R9+99awWbtJmvMF
N0SF9ZIxqZc+EMgpSokILoz09bxqa+lfTdUO8elH2ebGc37GOdn4Wz6nZuxU6EAW
NRlxBhpxhcenhgjuW+1OVl2vlWnoT/S0fhCwqTGMa7ETev0I82sSlHgXOHy1P85G
uePaTkyuD3fKDH5aLwQVd3mR2BByvEDiJLTYlfZ1GF0cIY5IzrtKKaZQnlWdLIes
QEOr2fHZap2ok3k6K7xc36zMGGD8NOqLtIW0BxzKkvu8Pd3kG1f5KUgADe+j/qBD
iHjbkgRl1R/KZR+pseMh7mAc4MtU0G9Xu+RzxaoOCOusOtVuxz9m2DgufDuPArlY
u9YkuKaBxF8ZDp+QOOFr06QiotI/ZCR1hzWlmTlR9/0rfzsXwlxK6Y6nDdArAH9g
vhS+vkWK2ocpQJFiBJtl1MP76pAEt1Aqp/pW73t4UXxGWHn4HNNAFkbOMAj363u8
FSfEwo73dA6YAhYqhMqWWTFbzmigkLONR+IJC3DBMK1gKbnwBCVnU5GevREsrYEm
aht/WYwMXLw8KrRReqwEnyU7CsDbK6qcVYjsgaewcxUZ3K1y7+P3fgdEmOa1qduP
kP6WgqXgjuXmO8rXrErHcSW4Exj/RqtcRiVKwCyzzpR9rbDLa2g90CApl6+rzEdp
4pndo1HFNUSURvJn13bD93PMVYh/C6eTlzX4QbK4KHjkqF4aLYlGpOVA2ptOM5FB
qG9hlInDaeN3FXokcAq48u7r8mUJrmv9wRMJaoQ08kftTpse3Ug9xsNkWQI56H22
0ibUhz0KdHCdCWT/zvywJM3WVtxHv9+gsatlH1atGOthZZwqs7FkinjOl0e519ft
kCuKeMv6mLIm3D1y/wA9IXKvbA0mbCjuA9JS76eEpK/lDZIycWxpXWUCSp0wQuhR
vbq8baTEx+Ct+ld1PAoSxextw0njIdpfnO9DWZ8Q4AJ2g3cQYR5zDDoNPi/1P7Bo
RCxEBOV/ZmFVNAxRjn6fAEQcp1PT4mj5ZE6RmHv08Dk3/fJiYHkRHgo1Zqz3Q32t
+mfmqR0lw1m949wff9/6AnhNrpFUhO26tU8+dQc2SokLSnoOkAnsiOmWc/oKrkuS
QqbPgNzl8JnxCL2/CP17iFRYL9/JM8ouIMLO4bDItaWhDv7ypOg9cVq6ASRrWTZq
ksk002qCq3Nv9Jd7l7ViYyhRiRAF+DzMVyatlnctkVMj8xGAymq2Ln1FiRA4xXgN
/ztcM/qX/QQXjdbajxawh1+VElP4bDyEjfUs5wqLIyv4gbbVgTjJKDu+nHAVPVaJ
SPBm7X9KIpZTxfiV65dNpRoOiLne/8tlCx1rUzrGdouwvHZc9UzTWoT0z0z1ghkB
DRjVvcoBchuCpak6DS69xzLjzE7LFMUmn4hpf1lpOl+xBZ6wh5QE4BSJE7Sbq1Dh
FVbpmoNmTuogZYV7+v/T+vyGibdNOcfmv7wQW8KiSg+zg98aatKYeuLuiL8Q/4P0
/dKDrIcvbWb2gDo3peiZVNdz8fM++tCaajezUIK6n2ZI+Pk8igSUgVGY3rEmW2Cs
55YkI21PFAjKiOZ3OMvGSgr8tR7AfioDCdyU6URpahyYQWOj+pNL7qNHMmFx42yx
HVMng9HS+mf026Zrr4N8pEmf08RA7MhvDY57dHlamNv20SD90EuwFPn+AlDgkSRD
IysRGUv7gILSH4ChN+hS8JC3GRWN4KnnglSDIB15MuNjWDx0cKhmmHVn3YPIwcrD
1ZosJ2BNF7MXwaN4G2+Z1QwKF+7H3a+iJhgttHHh58eCjYX6MkGYhu0R1RdbXMFP
P/PvsymPOS7vIkQ0/TpdasXltpugZ4QoA4nUWHUvD55LgrbAjciov9uHCRMItEJ9
KKJKH1bf5Y8J48u/gvkg6e17Z+ucA++gaGz8mP/b03bkAYVn8DERurEZynRJDkj2
3aMoFVY6IKdfvLY7b8wYVyxQ5BA77nE3H2sflKseBAPlkFP+uYCeVgYF4OheiyjC
IqJJddvdIUZIDLF559gGaeTLncs3BdvYtC50PDX1iidm/3eRto252L3Ar5Qj4Gdh
NO6RKxkXAezBpeiPY9dcyBXdIVLssVGd1aOaR2DxDE4KKPRP5rTc5MNValsfQ/bg
AP8d4HziPD1cGnS376F36+QRprQLO0+0lPBli/oLdUg73k5ymuDlYhH9Ysx7V7GD
XwXoI92QAxXOX0HWVjIbnWUYIvzwIr+9hBAMA7LdM4X82FHFbKYDIoR8ejqywdpl
wCj6cIHfLY6DhohxvGBir13IBWdEJ1/JGd6IVKXfEbA7UE4iti73T9S7U8A52OcE
ORJiRodYX0ghweyv6fjxua9R9lplTbliFdTn/pfHKY3imy6NRL1WhBEVef5CZh5E
DFRDjcG2KgqX/C6y9RqtK8yaiVB7hRP4e6jTlF5WjTTAWIoQcxgL+a8yhLwcqCe2
xoB6W9UJg9p9sATcjs3q2Ng5QtoRy1ht14t0Ev5Csu8eEi19sWlKbBxgPbrkg35h
wTxeoVX/0PebNCsrDsFDRiraeOLYPXryPSXNHPJsLdp1qngrq8VxHlnu/RXKjoK7
ppYdHzUyRR2XLuBVhI1YNiw2nCoMJ+pB4KZ4x5XwYjBpufaJOAfQ1GVzLpq5f7ET
hJpxYBjSw9mlKRZYH77wL7KcQ0UHUmW2xhgZVd84DDCWPNzqYBIm7EtPLNFtd8mE
zxhQ3W/aGcSZX81f6dzcTThJ6IStlve9gVBK8FkWmzfX7qDn0eqnggntuv3uzxNq
HEcQcNu4qcibWREED9OVHMVjhh3TBbA6hRHlaVeQLYlIp686rrgBU8TG4H30Rk8V
TCQBTbC4s5NoVh1Ar/uyQp1eS7r8sVMlfIMZKLq0VWZI+eLNOjOsMWU58aG24mM2
h2ySfqGZrgS1Xj4Ej+ErkNlIWF7pZqZ/N153t/uuLdAKvQWtbqpkv9V6BlCjR+a5
P0/PFKoIiRo+dN3tWC1xsD2eIU+bw9N+z3THXxIiPOONlUxPcGB0kpWQPSUm0djH
gHbOQSYjjZL2HzFxvH+MHOPi62UBmGTY78SH1dXJDBmlURV3VSB+FD267FZ66ukD
9x0r7uZgUzebptmGtrFpSfSBjUVp0PrqQ5wU+6kH8A2piYCoZ0etxDtOre2py0K0
JPobptmLR2OrlxQ75p2v37OAO3Kwvz8woEOw6xTMf/TQXSAyxMyu2C0GVFggFKyp
OdH82AOCxCXI6n7PfXmqJPAEYDlaOMte/ffINufIy2HS++XmhbmeWw4473llQRD1
S/cuWXNkFYP9OPUuvY6myC5bXlCnGQAEWkm/2dLUcK+mkuoa19sxV1e3cmfFVkzF
n687KGdyxv7wnK4RqOUtkkRG3f+FpSxuzTfiIQow7eepDaVSezCDnPcRkNBWfeIh
gGqZjKhxvnpHA4XK6+f6F/e/m2DBgeUQwvlbRiVrmBzPww9DTuVdox0Yzxo1dr49
YKzAIfgr0YNzgGxwvJJ/lgtNEME42aEiS3UDAyn6vIAoJU+iDQGlW+TrxkYWB/lQ
wlO3DRbKlfQyV2lmJH3dWIMIwIVxDxDJpqODfXOHjjVZAqcjQHHayCUUjSsei/NE
XZNNsoe3doPSfm0qYTwaXqn77tfYnzEvg1ovo9/fWlklVXIlQGhr+DtLrC19BQrG
eVzHJs7/S5Zo0qp8InGguOLl0U4LyAavs9lUGhNL5lGc5wIVPyCXxkDJMYjnA1QX
N3acOUG+S2hVfhg7UmOT+WiN/SmuVRm6Q8qiNMz9Auq7R7glSeLnrPUniPwWikGM
wauV9wtQBQWLKxeoMwnzTA50TG6t03CLHS2BLRBnoORdQo8wMwU5xcbjRLJ3Lvyo
Yxnjfejr3Gp/Uh0Tt0Yp6dXAyW2+Ey0c9dSBlGRsvJ9FcCq0WykHim2c2GN98t3A
XWEksM7UXVZkPJtrt4ei2CimjwS8/nHekBJnuOT34xOqTTucZdEyIJNbIIaqyIu5
uggKXkHU5z0AOVkQZ+JJIZg6N/Pxm21IEhBgW4980vZKZtmVZPQy5NmQvxj4Ple9
wszVvUjpZWABjqUNmeJWtvuMMD6mYAifOsYcsc2CAzCGv5mvJ/AnUT45lYHDotBm
+Tym27Eh313c3DWIfvywWieGPgtV17epYPdWB09d+LpAzYT4wBxFl/42Qz9MGpBw
O64InupNBrv1GafhMXCL1bQUAjQ5eOWnkZGzaZa1NrPUVEdnFP3f5UJoLDwapKK+
abxf4A1B97HKkvCcIcybLxLpoi8xs2vfpIHxgrNE0sIh/INxI0j08fwcfJkFKNuq
H+yP+7N/IGIQanRpmxxwkJwU5TJx2eowSdRy9CQ/vNh6AhUXtchIzmrCQWJ8obyc
8KNyu5AQ3P0OxL3DJJhRVJZi8DLMo78znSBB6zOQz4INhjtWQ/y1c2aUEDirOUdS
boP5JH2owWVLwpsTcxoJL64/dkYTgk+07Gvvo+FH+qAB+b4fO0kqBXurmy5BdqrC
HWuh0EsFV//bGaHO7uT3lcb7+tn6v+o05VUdvDZfiaaXFyo+GqYT008PD9fhxc/c
O2jVMCQkxmvdO5GBJYU1dNGZGe6Ne8BrNqkat9HM3h3SudtSDM/DqkWr1NXQI96b
vNj1AxC9i0Y0bJzPxwJOPYRtEm5cNtCJWPQlh9k8705XhdMwyDpnVvytje+yX5zR
yPZV4XHoga7NouhgN9Qs/jKdSWCN0v8OqXcLGv6RQUiW0kjf4GsDyM39EPS2NGBm
0/0dL0yYuHK8xSbW2aoJehs+W15kZP3ka94b8kt15ghU6n23NM4Ojz8GpnM4quny
ENt52SavYrDMFNSOj5X8z+un+YHpS/2xQZ3J6ESClOguqntnJnYXv19jWtthRw7k
5QCq7PhHHec+5PR2irchqOdi+HqMQ/D8g7JWFp2gLz22219yK9i6UpY2AxgU2Mjt
MZW4P4z+NrI0TG7H4NhvQhYbkRSbLPvf2FPl15KxHLZ40gzTXWkLgekNicdIGBL2
1onID6XIM8E/pdAX8DjWIlxlCJspTMN48g8YDiZjMbZPKYbTqUrn6HFElFVdR42B
Yw5hGLZtcP5xXwo7e2cFLNq+xZWz9V4SD3faBobFI+DxaakVCbhoLiQG4awlKp3X
Nse0UPKBkPmq5OfjgRBbdH65GOcgUJzKKn2Fqy9oHU8lOvqyluVbgzQOj+3UMU0p
PuOFnQfCeU8afmbNY4Ucj9in3b76Whh9DYmgbh+8NAT+DDrjLoCK5Nog5FI+Tdz0
5r8SjonPn5FEDLJ85MT3JxpsW8i1+4ZmWN9Ulk3aJdNlF8eXI+z9a6sBMmuvkxEM
o3kiShUVLyTTonDQWr97GmE5/Df7IfeTwFDfqpXYbYp3G54UUily55s1OvhGAnGk
ZAXGVJNWjoIx2ySItID1DFu/xWHFgKEKCugvvQghCBdwiuxLINmSHhz/JhgYYFkh
PBD4gPrfa97CgILDkHcdmkENPDIQv6lIRnCBIrRyG8r6hOOmcL149YRspUgdqxNp
aEZ7dCsvGjybgVTAMWrOObEZNkzDTng0VvZ05V4Tg2rVFTAs3pe9AOyM27+P+kl/
eyBxNVX/QfcSTnnop3QWWuJRLsWUES/KQOLWj4g4VooKLjOJIKX1zvRgNREpZO8V
JXSDQFyqngTDFBuQe4A4xTYDYzbMlc+HUtwFY0O+xvsvsHGu0Ztnq7yDVq21pFtW
9BI5oK7Al51XyFKDRukz7BZp2QG3ymXz4NvVmKv9BGGq+YeBoi6iu9EnHaxxh8fs
RSpqT0hsC7GBT1ggb0mGP/aeN5gyjw/g1yYaDvRqFg/q4APEmYuPAEJaALWb4xz+
n43ipaRTxokx/ppDUxQ8PI7wcshDrzxqc+6O2MTxkl2KTRj2c58tO2cpfvk+/3VK
Xie43OVQNv6NfxrIhKo+Jb3SdCamePvE1sBLmixCp6hnYJZ9dZAlw+h/bqe4PFH9
K55wJK+6CqkjMYaXjErpDtBN1ww8wp3ziUkRgeqVoTueRcmzCGuUxT+k/wt5YhnA
DVejHiUfjMtp7lq0qp+EnIeor8nrnCDYKlD56lxDosVzwEfu8JfxobzSdsvMT/yn
9agl7X9JNUUde2gqoKPJYnu5lYrXKWsW0nF6dJS+qQiHhFGrDtIvbSSkn5q6a4vG
dLSeYo5R4NxG6HCEfx7s7ZxGRA3k56zNEGApsLrB2W+XdVR+IIMniMqJ/y1U672b
A5vaahmWOsiEgCRV4oW7YkAqc+oJHLkwbtS+oCFkNk5aqGrG/KdL3kErG4Z/QuR3
muHftRGtHhMmweY45IoIQy9WMtqrC/XiMx2Nb+emrpTEsl+7NA0czNCTjXsLcej9
klsJ5hoFCQmIzgVUZ4Ypzl5MohRVUKV7dQX71Le42N34FajiKC67RUu5lamniFxy
S4y7XxzOz5wBHD5VG70n+HxxkA1smQLn8e3VWgrZ3IWfUF2AB1fW1srEnKj8to/C
fixyxFIA+DrDHo3dQDfedCbvcDWMSuhq1ed27kLGpRux/3raEhcnB6ancFRa6Hjd
YIonvyDKkJn7sm/sad19SDi4Ae12aAZMR4xXYjhjqWy9J3g4ZPpqLSM+1G8gVyPe
eEvzX6yLqfSyWSaZakoGQ5y0Aw4TwmFGo9hMcQ7zLLtBE+d5KB4Cums/Zncodb9o
MN9EjRGDlvmdMkwtnTFU3aE1Fm/QXmThxVtqJPd5I6ZPrUDF+4H26eg9LBDr7vXf
vjOs+MH04IZ4su26kIO2piNCOkOw76QK0QQIlh8xvg5Z8FjkIs3l93MK0Cuzj50W
DkfVlx1QjhGjQUdQ+QtBKLTRinjfK5jSy4UbnZvlozA5wvj9LSrEJqzdM5+QvXym
fczozSH34eUoG4mqukzR1ER2n1e9Gr0sm17DjzizD3FUdTV7c7AaR8ukATMKnczT
5WqoYKFNNLq8qP+DMmwVuS18/1zRr4PuEO47aW2e0Wd8ZGQb/MPfp9huqe7+RVSL
tXmjLDd8hqfa/vgk56VkrG19WDDx75E5kxBoMrcsTaG+iRrH+La/6l9Ue+CFw094
nWOXoYNheCP0PLu/7NVXddzO9HDnDXFHvgsPaRfdaC8DVGXc5kaQMjeRQEMwODD1
fkeJ4F6C9snPiL0zejH6NFwRcul5iaggTM2kEz1DFwKdeJcCInvsa4i0IG1f7HYb
4ODLHnPck6Pj75xJ26b8y7OnexTNhkWq7VXdElcsLipOzqry0PbJ/sPAT54975rg
kn/+RhEFDzSw7u9MfNlpwpxG688kVGqKkoxHUyazlwlTLXt+VuwWLTLitKYf31eB
/9QuE3j7R3b4Sz4Vh9C//iI+g+pczqACBGAyL73dgk+ZDZaQ/zYcq5VVoL7sdNwW
69guXiav/TYqSfcPodVjd6Wtc1EGVN18uUZ32DODHOxLtKZZ9yhUd7iN8woeX/HN
Qq06cg+G60/o2xjxD4WYyRJnrow2bRumTe0Wjk6Z2Kw2tEvYVX3OuGiHhpqwnojf
pA583vazaDmQ8xVGan4KqkTRidMR/9TCHHZOlKFSZLuj9NGPeqJRzhWY8pOZ8lGE
s7H9Xgj3imsHL5qL+H6XFgq3PsJbcwarG/JkN36RnBuWRH8vDgBo7S4jZ/4UbDD8
odRAHUqMGduXo8QbK4Z5KFQ4reNcoGdmv3joZ7tKjAfYbF3twMEWmgHYZnc/BFG2
5m2mtmhY9tJfQLUgIQlJrXh+gUsxg1TPCGa47Zbg+vGdkkCP7zJ0OYLvu0K8lK/d
rNvQk0A/Wlmt1liPiQ7a9TLBc3K77xnGYrezj22aOvMXP9Udsv7QsD6ZnMIqLFKf
5+8LRqu3MlZGKBTYTUtzjcqgsgkzJ5OxlBPDtVDX3xbi9yLkoLgBCGWwvDwS/0jB
fKRjNZbM8wGuta4JDowTM6gQHT6LxlIkLF+LBwGMc/0bk4GvAods9NIHEmnHvnor
sRqX7nlaqe37iNiZCwibO5qvEY3UZABATx2Rm+ycsM9tHHHrr2zFBvPCEjQfd0T1
OGpDY6PF2cr8lsRF87gn4ZKmol2LbnMGnHocunwvovrGxoZz4d8NuDIxSByYGpx2
Rz5EeRCmWDSzUtrgyTiZF4cqEcmU5UNWJa/xiqX6HG4N4/N6NzUtoRx69Fr0uDif
NoYM2CeK1s496IgEduQHvUaHK06x0F+NSRt4sdrDwH0//Tw6B6Dd1mX68oWqry5i
evgXr7S43LPgeydW6bxrZzVQSIhkTTso/CUerIZPFgethp/4xQyWSot8hzqo+1dx
vQcjpt01omFT/VaLy2Yg+NmkVIeFH3wbyFLTUtQVrUvJcU2UDXIlv54a7NsVR3Yf
9QDEzI0o/GyB6e5x5pvgIaBw170aGhRv5XIZ+PmPWTThVSf9aWw0FfEAXh/9jHnz
2ppJXRc5ZTqktqfcZJdNyl4SSniz2u1YjX5Lc/12HbfMHMSw7R3QQ2ga1+vYAOLv
qc7qcp32hUWbnSJ491U0eKfk9hFfThDGu51b38iwf3w/edKnPErErOVWW8Qme7G8
iwyyQFiPDGRgqYl4vx/0Cv1DESktPze3lD3mt4vVevr116qVNV1JyeYBzz2ORgWy
YyL8IG7fhKaoEy8gm+LEhrxaQU99TAAv7ldS7x7ArZhaxW0C8WBCrrpuBZHIm0nj
yDTo0scPA0Mvkthrp5ZG1XNnJKP4cHMzmcXpmg0+6EJBWkLkfIjaHE/wHR7JS+H0
HOrB2GHQSXYXlBiZJT4CIz4oSo4cRbvWmQCqAOHyKVnoXTl88C1J26J1s5UXvY/n
/JSBNW0N5ZTwP/o9xta1xFxkIF5eeRlqJGPYEMLkMvEzjXesh0zvt+rbznyaKzt7
5MTDkLgydcSumgTd6GIaxyffZ3zva7u/r9n/dqM5poq6Na494qITTDVcuiloyqaI
MfkOGe9hJDMv7nXv/wFtg4Ccp4QKP8BQnOfGR0LDAqp0Da1uc4+FqjSBnXxdeaws
dIS3kp8SxcYWOj1qVNOhrqE72Ek3YtOMOb8do2YB/X1BTbCvHFE3CoXe495tSXej
u2rlWr2kWkdKYrjPrc8JIQ5AHds0G+JwLDd8q5PzIt6y+V61qW9LsaBDYzUupabG
SnJKteiUgLqQmDEf8jVmR9KcZaBM2WLoW2zoRhGDiL9s0Dyhh767POAAexRhGS0Y
4ewYBOOm3aOC+7PO4CEvXpMBx3u9IloTRqRpxS+WOxZbfoz9gQP0g4k6Z2Qqrkrb
7Up60Cf6QX5qFPvFdZ7xOGxSTU0tWykca6F5BN29/pX3/dPKWKSbPVf8v5Z4ECIj
l15MQG1mk+BB/p1eNXG5IwWypQWWXh+BPXtbCy9PP87HUedA6N2p+4uF0BcrSHC5
aC3ooiPeIe8yXhClgMq5WjalkMjdMBFOImFnGj53woYHYYx1Xw+8wPgTTLU6QRJN
Vo6Sy/LHpaONJskpnC0IhWsFNikDFqGmy5sQNiecb8JsD2dPTDf3io/KPkxfR+Rf
vhdT193GWiqm6On9v71CK+RybNLjF15AfF/n2oRSYEhZvp1myQeSX/d7FBC3c2P+
gUGckN7+wLnfrIyKsrb1BTBn8bA7w4SA6WNG7y5LKYoXCbPWV7r69NwGCNrWfR7y
E0nP7TldyJDHELnLHEu0AfQ6UhLqiidotjD3VqxU71yr/sP4egMV8WP4v4LMkLW4
Ze322oOtqMFznOZ3fTpzdh/eyKgRluUR2eANtWDRC79pai2EcRXW4DX7aFcgX+YS
GZPHdxLf/51zv+nt7ua0qEL0kmryXm59Zbm3UlZbcyZGo1HW9CEwsbJQE6yGR+De
L58j8nRAXQEF+eGvfvT9r9mkYmyv8TIp4c4s2cNwBVqh+KAZYYP0XzrJxvM/dQJP
y8F/1uhHAF5hHcgpIYH9EYDR9xR6VNPXKTD9+c6K6bWMUsiXa6RoLVI1JuX1d2WL
ncZZtG+WbtIy2MYxpZJfp6bETXsUgl/JK30xs4RRFuWzocMSoVeQMpUO1kW8ILNY
Kka2XOz33IRq5omBNzv3ot/91rQIYWPWrp5kVydNfxKzWmJeRLBNWvWfg/p3DoLv
83YGwGJ2OwULp+KxP9UNi9IO5uwdqA1BiIMiVIA0MC9E+MexmflisL7905h+Vx7u
keD+LODHQ+VBrM082dq4inkiGHdwSs3ZMHJojmarmGiQxgHXFW0Gq8LDU3qlquWg
TQgtJQeqUCQDqz+wdpASuhTtq1bNtnkdWQtH8wARlEVodxUUfG+v4i3+rwsN5k24
YdyMhH9bHpRgWVXFzyVmJ7K2nRmvjGPYvlhTitKX56xEbRMIUxLgZz1HqTJyQ0h6
P6YDBld3Hx9Jj5s4BztfB2BGFYPsU6kjyn3V9QSkKLBsIXHK/eYiSJdiX5jjshGw
pNJsGmkgWIjyFm1aOaB4uzaZzpVDJ6QGAFKF+wKVe7Pyev34OomWF2Qsvfow9jXA
LxV/IaD1PjVCdI6dA1E1Uw0YQ6Zgf89T4RcOlUegKx5asMn4wMgZpvHxICzbngzA
fEk/Vv29iaOwDPYBMLxotT1AB4VPDTUvCEL11Cq9qh42z0GCyMY2h2T6c4gC4Kfo
PJlAU1tk/ha8YTdPrZ/8sauNg2EGV+J7knap1dpukDKR+/iyNPC2WSZJc6I4ssvK
aNIYs42kQyi9sReQ2zopvu+myxLc33YtFsLi4HUT+nWOySHo6UYCx8yNdO+oM5v9
tb6Or8NeBL3qrczuIDL7U5L152ar7Gr32Zm2wLzFYGJwxCD3aZQUTcTVg8bqcSlm
xKja5f1nz9f1FT60tRKlGXiSBC+WO4K4mKR8LzVgWnAVbYmvw5m7vdeFXnQnw3vs
tGoCpoEEX7jC5mbwY1NZr088/hkZuHtLrUs9l83T3sDXdWAt5QS1xKg/6JLgq3lH
bST6l+12iOjxJAdEINm0cxgAfdi0k9SzmfUs8757hxfZd3B86TzFlWNpyaEfzWkh
XvhKSO7HrS7dJItkmMOV8eu+pqsmPUy7mnZdHIv0NWufmnhKvD9Uz2XC0LXLKofR
z1YFsaLUx9vK9uSrohjANllCYDxUargs/K81Qm9tEbdpR6wmxK9OXq4F/EeUu06Y
dQ+9/iegKfTYfo/e+0kcpBIhDUgImXf6CeW5mw1ZdCgVxdrVdVQGwOm81E/ky5fY
Ra3E6iRrz1Sxcozh6nCqKVb+ZifUBS+tyhPYWXUbgy3603j9dnwPJKk6ODrH2zW6
REzdwizfUV2dH/eTnO4aAhXwZ+iax4bsPUxA3Fno5EDv0SUdd63U4rKEczTEEemb
XU0bFeulQ8JjCnXvB7u/+o7TjLHJqva8+jj/U0UyIA5mwn5e/Xq9y/H2MXTlxCDQ
XuOY8NgaGVOceeLk6/mbqS35yHA7xULnPXkDXtdUtTgtJRVLZHiryqPyoCYdf9OR
Qirv6HT01VqM/aYtKMAq+WJzK6l0Yq0Mtpfh8+SDVzHCJ7mNWdHIztG8tTelCP/e
cUNUl7aqS5FVelVGZH2uQXZWpQV7Gpyb5nB1zXgDzjtF0fgKuLpPL0wgEAlBLhZg
4UWQgfxyu46cUVUtZ1VRTIW1KhOWHlAEysO7KOHAXgBxGVxwoj//tuRV0rE+o80h
mA0BBgc2y4vFDCs3CO4bFT3HrjrJcEweLYwFCDvtsKRb0zZ5oxVv+ksIGXj6/GK/
x2IPvZUNahbpDu7gXBfUf7FBOyOToQJvbjzDZqJ+BMenCcQgJ4XZipq/osdZD5eX
l+hNC2AwI+RBF7lbgzL0kWW8vDmRJv0dImJscTPXwavNtvt8p5vyE30Q+zdOrfld
WyOjjwy+Cxwa0BpgtuKtinXaj1sLNFhXqMhxdV3v1D61emT+mylIMseWOQkmogdR
4JkZP+y0wvyItmbWR7Z4Ue954sacznPRju4Ecjv67SM0gILe6kd64zzK+gauOeNS
Y6DmtSCCLDI48iD4buBa+ok5f3fkz+i64M/eKZVnVEtFcGwhys4b3Lvl5qR9cmJC
8G/vprD5IB1WG3mE32UGwgys8HermxuatjkE4XEveyFxYZFTfvwZRWFEQdO9uDQF
F+c0zhgCxbhj1IqMY1M73L6DoVI8PrlTxxzDZJ7+9PwEvtGhG3IcDGj5GyDebXMs
C1uGolZU5Oj+5bL4Je7vgO5EgK6TskKuU4+6uCWxgKa4Ge6t9dYrrJKjNWHfnufb
ACCw65MunfyFLyTRIFD4DUfyOgsuZLYOpA/5uXbGP3Ih7va2s9bidgplwPyER3yj
osLrXNDL8+s1qb67SsjQ6iH/5BB2vLmepO74PxmgkPiqqcU7lQ8Jr9WPBC3DBiZC
JB6k4uRKaUVwGm2H7YIK7Sqnl/JHoJmLfTR4/uAGsB55PFLCXCe4LepmuV8K76kY
/mnaFA8f8i30IxGWGBAcpbUVnL5JJn2VlQ4VjuafWIEj1ShkNpK5gWhYvuyN5y2L
PpvTvCopml7rmDAVVwurqR0bIGe7B983MfSm9r+N1l2CotMDX2YvQfmS34dcy2gn
T6OR+8QkJX6ICIL/y1YA+Thtai/brJjT+cTJXOC9UBN00iV1z51amXghuKMBUXPS
cYIq3nDRTN8N/lrHi5cFvFbJhi3SAIQY3XdKmX1QNVyvpJ1pt4JgCJb71F2Tz850
ugr4R0m4E4l8G03qQnz0IunNxJ3GKIeYXzGUDvUDU24lV5tM/ZVPGWYaZzW2QPU4
4PSVGHx/qwUNaed2F1gGkWXjL/hjCiYnByCGPP5jPw+yZTL2zJWzMcF7AzOKF/DO
F4lUSGUWdrmxKXQ+PCrHo7doWszR8jn4NUGfJfvZzhJDRQYisciDVxAgjBHSvwP7
HoKsO1QuqAfNbK17do7d59juqRY5kpo77TaboNDExcK97E6s5deiI5lUrBnqamCv
YBVTQ5MIaE5poX/ix46c5dnXKkxw+b/hvtR4T8+2ui8lXA7l3FU/oPXbz6a8fYq4
ojYZHiKFxIKrk7sKo53tLlHEdZ5FQvur6wAFJBjF5y5bQAG0HMzyrdfjv3W7PBeH
IF71r/ZxJ+pGhSihEt0xDCe0kve2nHgm5cNBA4JELWGM4eUfs2dHpI1dNbMcHJRT
s2LF048VfMdstC96cCRSQhtQ7M3tdQ8j4jiZmJ8Nun1FZF4WTbI3RBFmraHhfY/4
mWQwZ48YgAgN9uHSyXe8vsE6L6G4g6KC2Hv3uNDwXnbrE9Ygl4ZOf69VZLChJOcq
b5DJHDgC8DkMyMZXGjqzBA2QWFDcpZTaC41UPPzdhYEXXqhHd/X1t1eMU++CQu96
6gRB8aOYlMSdShdF7BUT7xAJIZspdm8gf9rTbOwmtiezxFsMvf7ro/VPxG1pq7Xu
GPwZizZVzT9I/r9YtZPUdyA/yC9kUaDlqmluZtaDVk69cCHrCGfW0BlPXqbtL50X
5Xxgs3+nHSvHWOw2+aHR4Niau60q08YJNF6Em721VWywIhK40xmYJu9Vj2h+/yuX
FM2gvtziCDwFBLkhfasA/od1Jl0ajsiRlGhx/Yx/rDD1kO/4vKxX9XblnC1wIXa0
zHzswcEYncM8LGWyFlhDxQX0WXkbHX2sgybMDp9XqZmE/aLAgs9eobpl5H6vqwPN
V1gs0oZZo0cBhKvtwW/aAAJIVxM4VCB7ke/w1MY2HBrWlXW0TIK+2ZA5I7aTI+Fw
KccRFBNzaLrx1N2R5/vHtqEFBqQv9x6Q/q1QK5WuusHZ1fNOJYWTA9oCgmfKvMaH
xf62n1qOB9qxSMYx7RMAqVBkUig7gsUzlJyfmzTl3UEQEE5UVEfik75+sIZ0V0Dt
yvejP8U7aWaTVsBk2E/Xi5qZowgOz5x43zzbrGdS2efgTrLE+acMgIgjI1AQp1sQ
FBDsH5DUrAifGmr1geNdtIB8tVbt+tDnHf1NpT3vfyChtfsMj4jHH1s0EeAFEBPE
Mhe3DJrZSfbNKeiL+133eOkKxgCSPY5vqUEm149kak8tdbqU6JOMmKOgfIfvxMak
D2m501POuYY3909IsWuWVUDgaYfClhayUKte/eNTpPdpqw3iv0mErx9uPE6UuDTG
Ks6MmeD0UOVROmA9V5nvBqSdj9sTduhjfQwfmNMj09fo6TTmBV7X6Q/PKGghx3Rh
jWMIrfny/0jNvB5vHK/fuvo719A+Afqs0gepsCrgwXwjc5q/8vm5bZcHFxrrNl1n
BYZfo//ucy27sEkyJ8Y7oN5PkHpVXZ0hAO7EMbFeRIBixhf3D/1wSrXlvYwJGW9q
5cycarQFuEjXJhtmpKQirQ+1eQQbzAklTtvDg8OUmIzpmSwLs2DzAd0ImRNdv/70
3Kb3UwL76MrCoVd1i0zqB9OHFmhPCwGWPijwiwehue0mOjUoYFbuHZK9pwmm4d/u
F4nEu9ucnft6RCtqy5qMtYBObM7yXHKvfFvFQaDLVQO61otPTvzIL4LYpRDamPkQ
xkbL6DOWoTMi/j0NFXX3n1hXFAvtHSuP72gGFbA+i4fJrg3DpIQju/gejhmfewwv
YjoCf7iyv/xy+8uJU6rKOc4WYuLc8QXzU0ffeCiril2LTgjt/yvMjCrhBdq7u3r0
wSfH9I+3GVA2/rB+URSy+ulD6tx5V3MI7/4Uhoji2b+n4JdsqesBcfi37bm4b/1/
svcTeseVBgYOmF4+dwynBXlJDk4SWdYZgaPmzDUHUwdSmrFSibDcbNnADY/Qb3Ml
fwx/hIRVKl297iXxnTqBKGeGBemhRjbEmGnPuHqwln4zaSBemWq2wtf9br7CULdH
clJPcNt8LuIlI+UrNLYVVS0t+iq6aGJf0hX81qRKsAr++mLKjGPCAUlWa2yXHaKq
xkTHmRi4fSeDpXtap4cNCLW8DwXRvfa8JxyhBG3rEfn+116NnyPP0sGwaQwqa+aO
WwmJfl1VQEZIZgeQQkO1a6m8vmED7mqi6OaOyaQ3kq9vid7CBYhIMtOU7geZcyYl
tTIeiJQ9F7hJJg6rhOggVdpei5oZGsyTPjAsNi6viXgkVRwuBL1wqBPQJiiGXjCm
lIW3/SB29Zv2NsQp2mSeYS1Vd+THRwEJN3Ac5qeAGxDpFb9XF3puLmpUxaoattkg
/WYWKqr1ifhyjbh3S6fQ657GWigk++ah8imRIMabs1ANyWabCBgQRxsW7Yy0+D1t
/XNQrbHdET8F4hnIw0cuT6Z4RViIxrnOG9qho2l7RFnr3+tEmnzIFE8zYi0KsRnv
n1cTLTgiOBnBwuCXfZiLCsgqf0YtS6Qgq6mpN1lMUl2WhzR3xn7cLf0dXyfGopuc
kNMh83nssrht+CKIoLDBQUO8BOqBa1tYv8TpNHUpNzztzEO1eMFzzeiYD7TyOcbm
ARhR+VPGMKYzdIm6pL9XjsuGW7NmAXDH4lLSEVAaZBSY6OwmT3ofHJWayC0/VQK6
eyACByVXroqpQAEK/qSfG7bj1UxP3F9Z2oiBWWFu4C7MXODIrbr+/npIrmqyIOj1
Ua4141Xon6Umhbd7gf7RwFjdcbWLX6ljYwdx4LqNwymaaRUWhyjKsY+t+h3qyGxl
EKycozdIu4Yg+iM3/gseKWwlF7++oWlZrLWtfHr0rJ/9/bhMacrOh3BXRJ8hpFVJ
ICXAJRV3QtDf0il5kOHBoxaAiPmw+dOZJgFtieDqKLCTA/vyfByOC5E00hsWXqN2
Y+s/3PFGBtJaig0EFrxB0yVbXtvOEljmXH40J2nnrURmx/QE2FUmk7Kz+36tAVxp
uclbXwAegRpHcMrduk4ME4hnUYXCpjlzx0zDsIBvZK7wyGww3uuugoqj/6d5jmsC
L6RfCG9KdYaf3Ys1rcqrQ0H59Hd+1TLatXPXTcf6tlgL/U0iXsYEyZvm9QN94VLl
uYz99/EbFQeoAqLcAA8M0lFStpktdHEgfIYTMq3duUT2hkixY0futpiMKsQnx+f8
JTyPqfR2SQLpcuWoUBwOxYngwjn84i6Y0sjzE+0cIuu0WbiLpdO0qa1Bi7Peiiw+
pHaTHWLdDiPfHX44E7YVN43rXFBCl3L8HPmqrzeJndQnNVGWoPaYx1tk5GAmI04H
IKJ/rThRG3aX453AXpVfdWazRHHu1j2JsyIRIvJ12qnYX/iWHEXTwUtXHbgCXIBf
73HFHWXIGSrE25tOuz3PbZ+5KrftgABGLpFJ7mxq5Q4arpDt1fj8M6p9SitQbTfO
GUFfWHrK+Pmrc2mLLvjOMgx8w6wJCI/8J/+/9S/TWhrKlkgyxIxO+yACaaNGrgY6
ibCI5coi2A+P2khyST3xPDSgsbNw95z45rM6YcdfD48NxdrLI7Z0lgjkhSIHnx5O
3GoGUZEiiEXdbC7g9hzFlUJLs+VWu3XJR31Kxj97luwdKJgAHTuh9CyPFdQh4V7T
JzuYCLRozoYkmWsb3jI5Pm1+Y0YEX+eQa4h1miRrku41zcXkPc946PJ7aiPdY+dP
m9pL2ua0b3kz3R68gjdXddGXEMRWQWHu6i1CSVmNRwbrEdivia26rsCZ5uDl01Pb
7Aa6fwYcGFCreafWpQtLR8/W1QCidVRwinVGQOaWZ53Usb71pUwDrXrc9kZfd1Zi
sXavIjt63NG2xhO0Jq1WWQEmzYHJgaldVSiRQ4BdKxyLsdYUlAH5C1/ujocOGLTM
70gLGAnnqnOtfqtrgTRY6RR0LlagrCgOuTyKVIjk9W4G+CZlvxUQVxikJQ4hIiEa
XxQxiyXarAmMqeU2eGT0ezd7js1h09fKutMwS8vC8Buf8oTa/vCaPgMNSYJSsXek
19q6XG1DZ3lBlEKgUG99hTguzU1VeoyY7B/2oi4LsveCYr5ImraRj4827vHDsWxn
i+sh1zkMJRv9f13igeRM8p/flJq3BF4C2UgX/4HQq/PGIuR1aYcGelpjGeHbUiM9
Sn0FRtESWBIXmZLnWMHKWrS5p/e4TZLmkF8KXUXyxjEkziTHV101as5k9mhIkz6P
gvhjEL3PajljY0Y3Qcjoqx9ZHrsU3bLCimp5rBz8+mSLwRKXsq8RE8NkjPtY3EEk
/T+YgYRQBmPBS+QuIJqzFigSOVBvCeguDqbHWQSejJzGTEYrgXWA0uEa2d0PFbKw
4EKUd9hgHrm/fBEO7na0EfnPJgs4p3Jv7EHf/0+MUCpavPImMHR+XMkJgiyFs+Fl
xF0NKtM7Yy1BBb5vC7MKKEOOtWjh+rcTDfDxWcyPn2AeRMfTlQPVCkH8nQtF1hvw
V07Bjxp5ia5jJ3Eqgg9pnBmbZtLT7k23TtK8CuskWAOOd6u938WydBFrsP4Q3CN2
zb5Ab919SgqvPv7mia7nyLYq4hYgRnowlMfzuX/ALHoOu0Luzh4NkDTXt1F8MYGW
PIQVqXQRDEA+rQMUWM26umWv7kmWBWOvqshfqwB3ZMYhXD4cKfY0xQ2+ON9mKkSi
btbwhucs4P5vqyAJ4tuHtPjufi7h648VRc4Pp9VuO+mlzsJXMeE8UIuav41QoW7N
Y2D3GCyLp1raCKb3vsoei4DiKuhlWI1HHWlPrkrhUlerb1Oyo/jAGc0Fi+z6vbet
3LMsC1QeWU1ERBZTf0enjneb6B3sxYZqGfnhGw4yJs3kBhmamvpI1w69Z7A5kurC
sActteG4VSbCwXu/Ndu7oOk70NGHhrxPkll8D1C9KTrPD/+KZzxZKsllTtitVPPM
r8cydE2ZlddMAbX7YSQwGbXuCHyChmNnPXPzSfaPs2lYnxzQauTn6GFYWkgzfemu
eu56GocVyPENbOtuIvYHl+PVlB1DlTzqvfi8Pp1AmcAMqE+DTLbxow26/+VOaMR3
FHkRolaF+SDfE120N23eFZRHMtcN+EkDNuVu9yA/2cduUQHCiJtmYqRMvJqSE5Tk
VniGfJF+Ch8rPRI075vDn78oKhspQUBrewlcQnii3VXLNQzPDf/PFLK6Q3E8aYK0
Q2XCzq5b1L6vRyxdedQWJTLBIkpOwaDrqFqxkUodLfY/mVhVSO+1856hk2h1+btx
qerYoTZuo/urycB2XUDbDTVZtS69Q055OvUha9HV3DCEJDySeZjFGK/P7rpXQ1GS
VmMNRBYTWaFROyTsjPyN400cBwZ5t8qwK7zSwVmEGh/iEs3SBDg4HPaH2u1NZDDP
rGWfCw9lFOeAjekW7EjLCB3PAxkT9eKG6rJ1iIAQXEBKqdwguOx64ET5kFnPyL6L
scS3fhxE59BrEWE51vJ7xR2m2nmOpghgxKbS5qTY5xu71pVhlzZUJqzGbZI2dPOi
F7lLjuu6tUOh2KdP751kCfC06n1/bkz2FGC7dClpw/aQPU4avTdPV9mAwpLjGKer
RTsRhgqponjnK2ckoCC/iAfLLEZQWVYhlitojxrG9pUvNQghvnwTilyysSwqMxC2
c4ZfvVHxfwH3V3iAhREyvl2LnU6Z7jJO3qTucuwsRNfF4cZ90KOzXD4FzOxV3z5o
imKFPkFVMUts21rs/fqhhnD4YW39pcbdaWs8k5PIOREqUY0r6I5664ZAqbpOhBlz
3VnIzecQkNVQZoOEYETKFpO+Cqa2ybEZ/+kxuljQg2r21S2DcFT+U53kgkJmi4TJ
KE6Hc4xZ0TZfP4jWJegSRHI6dsJpWGALTJZrKq13GrMIo9gLDQf3as3tCiKbF7D8
bvrYzan2atkGxH0Hvvs89xPhn3LdxXlgsDvPC0STtx0wLNY5h4LUi+jT4lMGSnKF
l21w+dBej9tcve2D+FBf83YU3hqxM0xcOIoqMIku6pBZvMGCoFPDhcd5YLd5PIl2
qGx6G9weaGAFdWgWTuSwAQhsBwDkT16MgsTy1DJWV3BWN+sXS8yu2c6bHpX35LPH
pYbvHBkewVZPkzQ8w2jWI2ggCqhCEphK0YES+rdpYxmTnaVvLSdo5IHH8ID3VyG+
0XSJfvk2t6ZLzcc4SGA2wTn3zQZGFYCrk5fQLaln4byqHPQnZnEkjvZ+nu7Wy1HF
JHmEODvFWEFvNEdXJDpVA3J2+D1dDfizDmrf8KygRgc6CDdKIykVr7uO2K+m6v4v
xwtjiAsSLJAspI6t7Zkcuj/6tvHEsxqDbMyvxeZmO4uUXJvYy2nRR3tosgdUCTMt
jx8D+Tm+j7Xmjm+WPtH0/4/qbvFG4e0Y2yuEwmrnIy0b9bl7LmC8OtjPGYR0+qHW
diCXf/fPnCIKZ1AaG7csJMNKTODF+uJ80vwb1g5D0u0tjDYrvywqmUhCdOXrdvBP
2IR7TXvSCltt+FTPm3qXdUMcj9ub3sWBf/7PdV/Swy9tREwCMVrgxpEkMbzTbPft
HSmzw8BnF/n1hyk+YzqhrBN1wdWnVNSNOZ6ryWsPmY9zoUrzyuDKvS3orFhWaZgb
1L0v1y8u3mFr27ou9OBV+piGCg3nMUywgc2MoY5/l6yNoPnPBz4urmyS6zThUwuI
TIk6uaxWHfIjmf0oleM7VeLS+yNHCfzG4O99sjDa1RUaJVVSz8oEHCH0f5Lu6WXI
snx7QZAvUDc1P6PaLZJAxzPhnORZCtdr4zls6K0MgAG5TgGveN/MwM5B8fjcWgts
K6WFmvcTTL51Lfy+Wz9li55y38QyNGqgpMpNW+9DX27nUdtcEnDXBF75X1bZuQas
R8C4qgDYdWWq6571j9hsR1B5+X79KpXdgO9z99bWKmmMjO69n6n/fgejTs1CcIad
y1WB6l/Lh3/llMYovkVJFBMnJtQOtevDel3JZohvXaypixWVygp6ea5qwC2X1F7I
Say33X/vdCkUOx70qlYVC30if1v9nwh8j5Q0e796241lOkAbu4i6KM/xDjBSYbs5
sNxHNBlpfKQKXz2+l+61GU0YfrNllVHU0WjQLFg0m0CySvLNFxWaNLdqVEMomgQs
xBlAcpoDFijwbSFEdykAy1cAvasFqKHTEP6Bs+9AbRtvJTJrdVUmOY4Dn/EaomJZ
cp73SCiPcZ9w27LhqHJqHfbo8poIdNo4KfnuaXiTBKOquUOX9l+HRpmp67feYprZ
NlEvIH5nVfREP+bMJbZwtb6pgn1AeMrVJVIQGVPAIzAC9KX+sWsfGLRPt4zfcP7w
nOW9KEZUMrRHBGbu3XGkJCkvGAHx26K4kor+AdP0Vd6HZxAwax3Rszl99B74VTd1
857TkYMKx7/QXdhh5FmlSLi+91/phOldRITLuzCXw3JZs/pM1XXNPVzGNOLPIP1o
1z9qKUUWj076/k7zBGnznz0gnKhGQsXXKHhmftM8Bc1DdHWW7bv8TikQCCWT8P9z
branKvv30Cp7dw3njDrEtXtmt5/NgB2k1cowRC5/ci2z6lSuEsnbi/p+0PViHFhg
BRP8JaWOpt/CpINFwqfmQ1F2KgX93o4l0hLL14OUrwAVMBw0har66pgDBx8iBYMa
hqliPlB4R/boCCUzMUHQkKrDway7Q4PQ5sj8hLl95fe3CRxTA7yhfxCysqnlBWk4
SipfdF3Y4SGre19z6AMFPbMGAFGtJNBcjbE2TNv4R429GGgR5DPJn8kwxEm5dlEx
0cHKZ7+AZCdof6hXp2R3Py0UAxGVNMDxmos+lONZ2wwOr2Qj8q8aCoN6xUOQWFkf
XFIRvxRfGYKkmRsC//Q/GQKwFfaVSvU6KMvekzepJbwjQAw2N39PN8DGwTA72ca6
fHQ/tkoPOFLuT/7e/D/0L0DWcu0gGtIFl/4wi9fy7YkepesvXh/zQQDYl13knJZp
hq42VQZWrU6A8WnbmTVp5pxZgtZ/aZVqdyPpelxtbPX6INFToAm9c58IlqoQ3C4B
of5bYIrzwUC+LjXo9UTJhZK6oh2ZxVS5I17FkbyL59+b5+6biO5xFgxN8ABL5krY
R4kYxUL5iA4rnUKt5yYaCO1qGP0tparlhilKUUFNZ3vlsd1S75e0ts1uvRAQ1HUp
+aGcaCIC8H874FeUfgmfGMlgKex+p1dqGZQhq6nZIYotd9JOJIn9pmuAO5ue+Ruy
GL+jHTni0kQPSNopJg+ru/8zFOsfCEZGk5plp1t35m3MAzwVN4UENbb/zdyZbIuX
7hjvHbaF6j5QzVFNIpHUwq8nQWiyjK8In8tDRMoHFsSnvwxFR5gti2ldafZ4RB4z
hCzqdevvAmkKePjtnTH+/InztVZmT0GDHpWhPStRgkY3gl7Sros2Ph7XwOWgdwFl
LVMqzvPvOPJthQyawjyW7pf6CHn3KoWWnpe7/zI8XDm8O8XGmnZuMPRK82ycP5KB
oUzuVfh7tYEy/UiZNXXRVKwizSDSGYLneI5Eyyql3RXEjZA6vW9OeMDg0L8LrS1I
kb3f8jDrn9/zi9fNee/yRgLGE3d48Ld18UY/AKDqk5x5YSj68BlrPWmCvun7rKvs
keVnyI2tjZnixGu0BX/XOYcPa8cDLkCF/MEmwxoP/6scAojrsA88VWL4g04V8VSt
iYH3SjeqAWztzG5JKTMmdTSE8qpdTAYUt2pIBuGLJ/yToF3iuFU7Sxg0ne33NdaG
mCxWq6DvJ0MV4aLMtsqWsRo/OUkStzE5lxEEnAcB+6nwlVx0FBY1BZ2wW/1VOOdM
oMo3cxUwOalJh+QZbNwt3+saoKph6L0WaD7xML4lcZwrixUoYsvdSfm+DTLF0qtG
EDEosRDQgoJKM8GNwYZ0x0xTLVubDfsvXCGsgKG8qxpjQP3uyn9KMp53Q7jINX/Y
kseQOyYGDpCmL6C8GTQKGDRkLjrVZzuWEuD4/OcPKndnYCR9Bvuqe56w/qBi+y8g
tromrYlFuk08in8iD6PLX3GPyE/0ESdm6R4kBBGYdNTbIjIGF6GHJ8B3Qh4s3wY4
zretf9o6rbae6b1jQokjjfIPirexwStxuu/hY3AcyluJGBqtajZNcvsjRIG7+ndx
zbMj+KTxGFYjhlN2GAngs62jyz8wwddSwlVSofS8cPnwAVX5/gE/IcQDz7+f+D89
CSj2I7Z7KlF0+rJxzJ0axnk7wehGYxw5Hcu1o7NFDp65lo1iFRiOLM+0+vpy+GTj
JWRMoCbELMovbfsNAZH5sFaaOMHUtSrzNOiN3efh6zn1fO33tBm5z+Yq0fwHS2Wy
AagfukEZ28lYaESCNfBvVtSq8MJKXhPcdxgIg8g+POUOBfwkExByAstTIPL2MaIe
kvZTrm3jRPV5cZdJ1Fupq4SCM15TTHmHi+re39DpLWBvhKlfuAt0faOdKIxU4mPX
cQ+KiZp7kB8xLSCI9/rqE6BgviIlUXR8b0OUUxkT3kQd9Cno9ie0/m7QtC5GFq5K
goqQGpSJPsu7YH1rvzWcvYPV+XCk27IoW1MZS+d1l1B2O/S7NCrGXqHSzStqtXtY
ekb0armF/7Px2x8pRm1vkr6aUiU0K1WhYWOYypYkHTvAT2p+Lw96hI6kabYAnI1m
VcX77HnuUgwOCtrSLV0oOXynNpQ3VgzxYDTHk/eVomgmkqjTno7JJSpycqzy8Bz8
228/YNvseGp2KNuMoOP8fs/m8+Ep7wXpCPzmTuTJ9OoVryf4Lhll2GWx74qvqsIv
Kv4Cgkb7DAg4dWBDqm8nbE0/MyptJkbhXktVAknb4vQ6BL0MJClopW8GVSwnYrOe
a9bz0L9Uw4caRSnJloXGKW0F8ka23dQXpjLvNyzoOEL11pbwkHPTo5QIKqxWVnzJ
h6MWTG/X34zqpBOzFfe+6vXtBpcK0w7JKqESTFdFXTLaImG8nezr6BVafKA8jyi+
trj2t6NkzQq7lFj4YIA6S+WtsA5oGyspS+wEm018K4BGXdtP+Up3yv+LxqI4ZH87
zQSXlYGxxfaCzvlaAccF+/YHcOQNNSDHFPMTzmtS57P/dtIKMfbtQaS5RktG5BYB
EdiokGrFg2oe8eD2Z7fGe/HVWcoc+CAdaXhEgkLeGOFZySmqCglFANTYKo1DsYRq
SKTXyqMLsdUN7XrPklJPOjsq4AA5ZQPvylTq9zyW94LWLWwmGiTf+b/Askd222Bc
BFVwKJWPdHTDavntrCFwsjy1XWzZIogVtBDCTuw2Gp4E4VQF1HTqE5xbCd3dV/kg
Tz/MuKQzmGeLRHrtlBnkYrMSSPoaM+piP5KOiWjRvFiFGm5OIDcjQipR72IZ5w11
sQrJVNs/33tuiSen5b2KD8/y2QcqR23YBxFq8NhnS4L7WoFxo6+/tQVxtsXOWEUG
SoD0HTI1pLoxSYcMXehUD30vbGmdT0tCjqepRRKPmRgrbxpoB+1AEeNU+OnmzJYR
QkhPDhj/nqPSPSWk9Gqq5v6eREreHqJ7fWl4UZvZDf9y69kvfvsljb5cLJIEn69M
zrzFDK+uY9wP8tYvBdeeW9OBw3Rsf6cXiQMBknxlkjaxrXbXJIw7rCw0RdvpyudT
W3HrHjsw3syUVgaEVyRzg0XMjq15eFMFMFhvL69WytzgJz3DJghpsggWNdLAVDta
VuQLAVhhERfPr69F5VSdWkICqXr7IG8d4h0uCpj82pySiO3QzHRLa/g44QkpfgH6
gbvzY48OJzHRugy53uC/CB/3S0pouJcpNxKlRRKKUDojmqieEJTyFOS0hRkwZtXJ
TrLoQkEqkTlbP/SM1FkmYinYxxVg5ncPB1wF6MgFz/P36uOKYZ+ov5onxL0k+CYY
aCQxSzmLuK+9wDB+edeAiJPLxqhEMDr4bIk0JDyn7agmEWvOQplBD8iC4La28y0H
0u3/rFKbd45iU6QNRMuD/n7Z/DqpgrThuS8VFu7ZYbfinJqCK2dO1h/KcFe5gwOO
RXs+yrCs4d42x6hho8nNUSJU1PF3BHlxlZISssjN6pWFsmD2Bb6G6gF9VgxWz/m6
6CUMWO3gKwqAuLZU5NkWIuWgj7B38JdEvMnZbPxJ4Sxo8nkkI3EGjlZXwSfJ+bzz
zgjtk/GweF3THuMOj2u4xpu29aO2ARIj6DoWIbYxaieZ/dxJIn3KQiOye2G5SL6v
5Ugf1qYOaNNRBjtJ3GD2ENgVhMsWO7FBdi2eJLJ1frNtg0ljv36XDjkm28dm9z3A
ZCGkRBMHmkhXRHukJT97Nfu0fvNlgyaYIjvqDYvs98p64zZlYFATCCUnZh5oYiBz
/ARXWC/X9J8Cq/uVv/j2tf2SpIJIu8NjeMbEHaN0kDLzKMdSZNsqJOWUR+U2Kga8
RhVcRufP2VMS4CIUqW+WU7sSl9SOWU1aOTRA8ws3WBdqhQL9nNwnLTs+PBNgDdoc
/u7kKb0bf4k1U0txgbwEseFC4HZZE8YKhonyy6a33PcJ/HfzO55FGbOsHmrDEgg9
uBvqaoapVq8Z6O06rufuXOy83eQy6SsTdJqQBwngYcVy5go/nyaCsj9e7gM93iqd
uuJ6s0R8NNJxilRybBxERqKi8Nmhu+WuLo3hNDdB+p6a0cRiLle3mKfCwFtdUGzT
Ncl+OtmDD/f4LSJTVkWOMH71jFuI9uf9xxAAR3mWVCMXSZ3BnjxD5s+RmVYUqruy
IwBT9jKab1/3niJR4Uds5Ibp9U/3KQnQsI32BVQMBiA/1vlIwP8tFggVeHqOHGCz
Pcw9QvinQ6pAVDX5Q4wMOtIVsb7VnXG4CjrebEi0sAlZB/NqnnLvQLekxYQU/BCD
gouvqlSLbdlxGJa77EIKenR2K9v5/X3FpLJfidnqUnygni1cO79Y+sfBWl1xxskh
rLiNcl/Q9RENWiogiJfp8iMC+Y/QPpL6xiJgY6ihG7xRatigW42fqFvPBdmswqO8
7aSa2jEdTCJVABKVwS9KQKySa14k8PwBlWTd1ozQnqUE0edUnh0NXZhr41x1sF2o
s5DcWsPX2pmt9iV4nfeLAGAjD/rmjq3c0xvQZj5aPJrYSOUOBWYbV3V8AnH+qkw7
tTzl85KO51Po4xySb72hkkYZ8IjVvQ0gjw2wcJGPUKfMV5MXH3intpIJE7FUhIep
xM1qubZ5O26O4/EKWhLCA0rE/mtTmjxRMYoWqdtMfoJpjidmlZinJ4Hw82YWG09p
wqX5RZQvo8cpWGQk++5uSURxmvhTkqC3Gv8gA4YT+vGJy18mWrhYmkN6IEiTsJRI
0rLLZBN7CoJ/O5fiqBtRvPkSxBXuAcCtickkmv9vimuXVLre3TGO7IfvSo1h2yld
udAS+GIpWKN+2sWMt/RyIxiYjVjaorp81BqIHh6j3ZHhvJMGLvkHXGTAh+10yfSz
gncf1c2ViffdUCRn7v65wLvk2bJl3Cr4Llnxl5ew6F0aJ5LUsjRNXchmSU23HrIW
rY7At6desi3bd1biw1tMsjUih4SIet8j9q87GTSa5OdJTUXqXlQvjknd4ijYdVOW
Va80hdkeM4/+SWhBch+KWgDLuLCQRZAlrqdW453c74Wzxoa2tfIhB4vMBxN4/jcQ
TYegDC/9JQEhL7oZ6bxLQQfkSg6acsOVz4oWEYDa/Ap68IByokYScvRMv56CqHUs
z7jyYpZvC1OTNbzP52Q67XQaAz1Puc5izRvficqgf/Anr/I8vhjdX6nbFTo4EfRl
nqnT7DyPAvyVSFhQubpp4UuX7mcRHUBhghWOjCvBY9UdpMv8O3NPK0g1DF35pven
vErEPPCQDW+Gihsa3x7kESIcw+Hx1A03k5WrI50DLm13RQ5LWo8QYtDzvUKtEViD
pGLhtgZcCcexm/eyJ6gvylz1XjPHeboZiOkIvh+Ekfmb/ZTkGRzEYiQOJ+V9n+6V
I7R73SLea0R83RrKnxOQ0FpeXqvSdTBxxloBsEMs97WcaclIlr4DA1eVMVUVvcP3
2H7/29clXlZa08vzqHVF1V6Oi5B7prloFipQkbO6HW1+Uo7mZNStEjXMfRyMxzhL
izh8yTx21sT6D9wjggPbQHn2J7jFxq2Z5qp66/0nYezg+nFDXI4GONA6J+opTJ4s
5oOcJWH+jJtCdH2hmBuTnXtXdG4v/dxdxuYNglhJFy7nGkd416xiSZzZcZFDosJH
VJjHIXrKWK5cZOAAQ4JKeCoUlCAueDkr0ul7MQpS24Nlsg29RCgBFAnJUnum3mMX
Nss4RFzTWgbAGRjMpjfI5u5+rHHo6/YnREInqFdvyx6rsML3YZ/7FMyWaQt0gOa6
Z6fZiF9EXOZTNu2PFGeMlccVqCK4m7ESkyPi1u+7BMBV2PbDosQh5fU3Tca6NzdZ
KMcaWKaIhtmKhbrIM1U1z0eFNtEeQrw/R7EXp1yNWcX/Tf5dDafchQrdvDkGRwGJ
PrjdmHPRL83xrO7jELegWWKIy8h2dD8L6tzQxyjAX3VEb6mOE6STwjgshH6rpUMo
+4TCnRVAMt/cI8ADcsYy1F/6VkaLwyNiHzAb8jr5ywNQrMx4JWqyMji1hjvgtjZs
lpq+LuriUqFRlSphOSNwTuh2PmyKOAWV98PaxlQKM5IIW2uqhJs6v6zRcQK3y9Vc
Xy4Ana4OyGh/yTNW4hMsN+LvQOxl2GBJAyg3J2YnWbsRUxdq9LiHCBpXHT99vtCQ
veMxHTd6X+lN4mwWui2SkrprcHs+64xQdtxPsY1BalCQPv14Is7v4D1OZWbZJrdU
69C7nQoXXpHA3le1eLTwgLoP4GmyZacHEsGI/ghBYjnrONBX/h9fabT+W8eg+mzR
ChjDuhBQSrqedk1rzoF34JZs+WyHBw0OAOgJ4DfHeVSdbhafqEmehWk6r3GMpS5D
XQvcsP851h8btM9NEpfmTRiWpibULd8fNv0HdduX2T2oozM+t/brUIuZelmT8hVI
dRyteW8IZ8l2ng5b6z80WAVb8bUwQBKVThdhfrhQIGc//Qw9X43kAn1lAXRZSYo7
PPuvs/U1UIkgQIkLYC80jmtYTFj5l6B2sSYSl8qv9fVoSfrHNtH9Mz4TuQ/HZoHb
OpGPkh0ppcPQCdw3cp+mTRn0ptooH6J0vFOn5ZcYbi5/dtYhV4ozo/eGiYXO+CqY
l28JIiRjowP947/udPYWlG1ITkBvI+hMFD/dOHJyA5ZTPqORvnwGTydV+CFeyJCN
8FHaquljWEfzTTU45JQUXEDjgcazKEP7dxEunKmHN2Y1Ng0ItLfO5dqHBTYPcsQQ
w0dR8PHQc2WGWDRmrEg5ZQzoisS9zWmwANJlMwKimLWF7FQzz5TmrDL8QTvU/PqZ
6Yql+Jj7LE7CaUb0rFccbhtbkxQUKY2FostT3HakhmHnJF5rKAxz3c+Ahrix7TuG
/8JMT3g/mv915WDKr3/2RChndn+7Vt2wtg2gpH2LZ0Nyc7EY3j6QONTDWOIgWivE
cNwVOm+1mPpdB3zeEsGiypf8WG34gvMcNnUGQ0LUtxyp1+7/Cdh1A3rOZDeY1N3d
GNZlE1M65ijHflvF4NiImHPUFoz3TYDWwX+Jt1U4rRfRFRXvaXGltx3otPNkYOw1
csp2PqTWNABq+fMDKBpE8bwMlm4Kv6WG0tWB5tVOV+5p/AHY83AKFGXhnOWb8wDP
dyLcTgCoEGEHtQFpkssN3YYWbX+LnXz3huNHi6SHE+ajwCfQrfqJrV/dCSIsqRYk
NTQWGzTcLvbbuAgZTlGTbKbW+19xiZ8r86M3vQ97bPIRnVPrqgTZ/fKEKEs6qayM
c+cPfSMh3VeZwcqBBTj7jaJOyff1YVyJQIH7ZfO7hRoTPFJ9ySjJmlqa9h3ob+Wt
1OJvHYNTAXDOs0HJvyX33BW3Pt3tWr6VQvoP5aAZ+KR4IYwvdpWQj+Cg3LmjuYP7
n/LOZsokFKwMse2T+emRVi5Xrcw/Dl79yuq5MZbJNla4hbFSO2pR8si3MY7qMEYI
Uh7+AoyfVRnRa9GTCjRG3nUoFL4Hp7tJVE7dpQA3kWHdBWRdJny0BwCeIOVQqB2v
x6eLFjjnOrMp5S8bujHRVb+JbPfyDpVx1Iwd5HS7yTiv2FQbojqx1Jnqo0iK7kif
UJCtRHL5sNokgA8rYJNcJWSzqQv1mhtRjr/tKtZrYEzX3hoacpi5IRi5mHaCBEDW
zaTfqaiMxDaDi6hoGS6F0H0wp9D22klb4zXhebKkC5Vuy1biXsogw04+c125InJX
WjJwCx0wcfboEg32hM6JdHTUXp0QhaSlTFG4cE/RbAZQZ+wDiKn7pHLCPHNiGUhr
nLfteR0V0t0EPNMkTF00pi/8YqqkD39DNspxqfQygbg6pBRvWEZZ3vhvQY6krC11
cnmBT3t6cClegb9O9hREZu1L2hV5XPLUXB29wkuwJ0y9gq6x7FPGYiT1PnqR2oEP
JRZW+EjLXUcxG3VxgOixT9E4mlGB7UVIhRTMgW5dLoklWIaglAPQVw14sMpGbixZ
XphZwxyy+kKXXtoP/+okG7vTCA4jHKuDGnafDG6jxUbDXUlP92bkNCh2upx8j2fH
NK+AKKcSOKHVEeYoAffJOeiVJuk3Ds9IsHklpLkzwS9DCxM+CRLvU7AsaKjRz7fj
a07WiQG6/FvNk71tA/2uPL0S4lrXe+S48fzpHUhhxxz3Syr61WuNcSR+fE1F2Fbf
j6DCNqlUIZnIfM5h4X4y7Rzf+DCQkQwk7dz4AUFQpB5HTTbj1gXz8XHeNBfdFION
gvkIJ5zCZNlrS8o42zkCg2zaD1KJZnMinLt7Qv0dqbx/buV+vBnpHjhQqwx79tzv
OuYwa9y9EqrDMyyzRle7Q18qht5LnjIupxXSBOPPn2IMmY2k1CL7esgK4eSb8wjx
CuxX5Flw/wMOrNoooIg07LgNQ1BC7f8TNAjyAIIXPSJlvwY2jnDVVdXSTyjjOiAo
sJiOwdI43hgOfQq4vUIaZvqG0IpL3MKvWjltGH7tGm1JbtBiOMjtcXgozyhTEWza
YpGvj6Q81adTXg0w+mRce3tp6YFlxr8WECJOZx0DDc6pIpgZpsaBiM53P9Tb88kR
V71bPqfOc7KyywmhEhq3VHUTYh+VRHaY11Lsx+kdtCcIA0XBahiwQMDxpq0ON1bu
6NiP0cKwL9d/oJpYd5zLPqlrjzuhDKcqm9p7DtekBi7IcrhySQ4+s2YpiwEmdkno
7NTlbhPwc5TM6MZnXNtq8YMHbfDIfe/vLXdxCerGANmnJ2sScqJqXZXEJiuy5HRr
KVh9eJqiS5m6IC5+CMQko3x2HZP591D8xRsL6cECJ9nDM6FAT1GM+0PjKJG/uQMr
6+SgYwy2ECE1AuhN+odJ5RZ4vsJcdgOeXrLtVHwMTnz5zVjMBzu2ot/drrg0OjE5
DdvUexa6BmuRtGeog2kLO1RvJd0c4DPJkeKpP7YEiCM5UF9XhCqvXoejEfr35+9o
wQCDWkrV9Plho/7adu2tjRCR+K4+hTfVfVlWqHy3hQHC1zkwYUplG3v616g1bIcY
2qbx+YStET1Nnpis2Z74ublivGIcylAoG5cJJours/+ydJDwDYQ/XtZ/6bTtg9ND
leMgYO40G/gwyTBq2P6WLiSDTLMOwgkFNdyuhBL42tEmKt6Aw7qpKlYkrfgEZ5jO
0vNKhr2lARptDTlsz566uyqxtOzmnfgW4uhhYSwHFeSg1GCJ1W3XkAREWo1BYfFx
vp3/WYoVpYbjC7EiU5kuUGtan82IUiBSeBIaE4MaHQKJJMAxpGwjjQGaznQt9351
NK0wHi9GICVnil63NRYtiXbFnNXIyO+aL9Z6RsjwcAxiFpQ/lIL3oW1f6DZrxXHN
2RYg8FPOReYb3ARuiSBr/DmtM5FWd3rZt2Aa9+6O3eTaY+q0qZI52XSu3gNn1Wkb
+tACz5g0t/+w0UoYohg3jVR6OSOvWKW81aifcLoQ1KptwxnNYsP3JFd5FfPwKkCQ
GMRHTlX90sVzEWQ2C3bKbfx7Dsk9BDdbkNGpp/1UiZyaaV5aJI2WUNhMjUl/C9L+
f1DP9HwWNqZfxrqrl9t7kSnrjjf9B72agMqyD80b+zPNdg8CiuCFX8RcC2ATVuC9
f8RjVZuRbt4niYpPhLrYoHknea2Zd2/dRrsdrjEf6GweSMyjdVJkNA7YVVrHryUc
WjznHqONBP+xzRAd0V/BsbMsdzcqGnPK2zHLs0RQBGd9VQKgPl76L5jEAuTzYhcG
kYZxJY5lTr+H1YtCs/rxbbjVjeSpHdbcWXhQIeO+PPRkyg/V4wqkCp4aL6hRo9wp
epxqGedlPmMmrS86miI/rJRZjVE0b3X45aDpeF27b7KdNPg1KpQXHRECt3jCHfMP
GVhLKqUV+ihPayeBnEq1W9vn2HvaaagWdPIJu943ers5Emkt4JGblwoWV/DMLCgw
vhcU4dti+1YyJDDlEz6u/cjib4iP3GPtFUYT2Hs2d1NhG7xm0UvIWEQG7mdnCkok
sX91Ijc//wQRMJqAr1kxn7eaJeUyZXs36i6YKgRqLLISMQ3MUn6K26X3iujt87mE
lqbb87wJ7yoWTsrNSuLWct2NHnPeXcmdj4rT8ktHbY7vv+OzHl7H+hTO60LgudMV
xQQFFGdfrBo1xUJjEtE4Tk9f/4dOt/TJ4OBarGnTUwFh6ZLX5xOXOue20/7xUccz
HY/QzUH8UW/fXyt9I5n3hSWQrPBYDX5GpN7AlWWgJruP8iX5B8pakmkT2ptd6dy1
nHh/txpzCJR/xw9HO1E/leWlsmX15fIZzZELZahlvMY08bovLRtJ+CGF8bfJIq4R
DPLjlU/l3x10ckmWIpINxbGXAN2WiP45UhFy6t2C1RBiBSns1Pb3vL/bT93v+ORZ
JnPpKePw88soiaGiV58rYxhuvsEtJM0BihnBkBYtj2gg5QLxjPIco0x9tG2LIXvt
aM5NB3CDlJ4J7YbUmasH9Q55HUCvFGf+bsDRJWgowfaVyrhEYCZTrT6DiBGenXkO
WkCBB7mdTfJ8TFvYPU8ff0Sb3hlhLQVjSxqp6yHz7sSLaQAPmsktxQu6Lok2GIhN
B0i4nmO3qufcN6qaZKSMBU/TOgXMq8fDl9Lv8tvXJp9umSpIYoQXXXAfEgCOkwdf
Q5Ttdk3cpEFiuAfm7m6ZMpgeUW7n7X99dGClbt8oQFC0JvEBDf6oclcolKzXBy5j
fsOMSNag7gutXcyfmiZWWPCT9cz7P/16TglMIec2G4XSL30KswwMmQTEf9cjmE/7
O33koBs7D4tiardFW/2NcxtZY88MMmIUdqBW6fx5rndoDeGINhzBXTT8sEuZFOSW
4UDTv0GkuX/RLe3ofuwsPH6CIL+4Uu502F4AoAdqLZNZ4XRw36pIhK8aLryy8utx
a+0GeTX8L6DbkQ1NfafvB1XiMAU5swqxw4Knnbb8wLyKzBlzbLozKZpUuFoQ/sbX
rwtCI1Wfh86f1lm5H9w04IoncUN9I1uiMmLoqnTZlCjXrGdLC6sy/4uml+pfVTQX
pYrr6tsj0GvF6/nABV6dfWf+hDNzznI0qH0GBJipDm6a1uAriTNOKOoCyKP1gZqE
BEoUZl1ra7nfY1THWDOGR6W7kJtUVNbtomZIG8ThwLKxmxlyrViSveZgGsfNabRU
Mbgga3zN4voKyE2ewjo0rKFW0JBpEOBMtLMcoDqY58HZX7SzckORKZ3+ZFhtjxkq
po9FmMeyooQqe16mbECy6KZ882bVwkYB3DG2x2Kux46hQRQW/yH0H2Ch6B7UtRQH
GrRLQr1+uChAM3+QYB8GAfIaTsOxk/cdyyP0sCaUyP+0hZRuHE7UP2gbZhZoiCYP
RRVSwx/H7Sw7rVzQOmzYMWbYsdBi9wGpWtVlTJp1ZONE0zeD3GAUjkidpT0dqbNu
sQaLQLB9gGpZ6nlov1P+mnNM2+2Z0fNYXQkXcu7jUviOZANnLjg4Lnxjyj/2PtIF
QeqJX4yBdrhDq0I6p/RxcDOun1k/WMx7FkJc8HfNnxhCS4ZdbwZcyrQk55rO7yyy
JXDT6SYDvu+fjhMtVySItrrZODzZ18AzrNYgMo3JkjBwfi2kxQ7GdRkKbhSciVbG
wd4ffVdd3WCLlz1O1WyqGnxzLKsgCaEZbm6kzs2IH1sa2lNKPMVUR17viHZkOtAC
Oe3NnyGO+V2L3QEHT0NE7hLfPhzjUVnDS0qlteV9xz/fQHD3PwWGekKN4lnE/LmY
c+ZnxQ5YahiA6qUdpaUqW9YP/FeAs8KTLPdbu4LjlMmlLPoS2LaZdDH1A8v2Odw3
bI0ol679diAQgnx0gcEkU/xsPmOrwqXC1q3oOefoGMBeBRA/hFLO4LYJgWflurIS
ECyhTXzb0lXblBesNBPn9WyiZN2OMKbfJibWCPo8mO7zLC090hFVhvhHqSjImHr1
4LjlcMyuYU+7uP4SQreqGYqFcYUDiJwVNdaDgDZniggrCtlLN35KOW6cR72pnrUn
4MxObU2JrqWmMN+9Ou1EFoC1V+FD05pALTMYrT3ipf0OdeT4SjRQoQTUZopQz1hq
zdEHc98rpeIJxdmDTJweqAPI00aWDZxWrpydwO6vOo8dQ5Qt80CX9eHT35rDgo7r
fo99orwt2J22z/mO9x7cQUVSZn73cnRVQ10e4J/Fr7+OSe+uOfaLIxlI8oo49nFJ
RKeyepHIr1AuYdoL0BLbWR1mAB98b54DJmI1ljyb3Le0ZTEB3kQscuqCo0qOxEp2
PL8/GCuqpRCJyAcbK17sX5AKbOqFL5O7jNLsJwJsrwVotr8I1dZTPN3dDkDDSh3I
bsNVkj6nvA8KodxKNNUU/KweaupaxQdBv4JUOb7PDTMrewCdafo91LK6+KbGUltS
IAfXwqYBmWH6ZhCS/SOEwluOw2ADAyj9tDasK/MyPxpAv6eqa7xo0bgi1rI1o3NU
z6h7we11/4EUaSi/sZwmszWF8fyukxqzn5Ak04hUDZL/382Np4l8XxHogXcCmIbm
GnXKFzRV2q1DA9YB+NYvEnTsNHXeIwqmiAHfMEqSGyoJIcCItPlaEwmN+2GUPBmv
p1Yx2wN00nMqu1Jnb/hO0D4dDyDd7Rb0M4TxLx+lMUrSopdtCX+rooo3qYeG7Nwe
DE9yqnv7B5ehqPf1uwkALP2OBd+JT+6+1CX5IhXOSoCI35hao3rpA/0NiCuyQyIZ
6nfccRcqdm2esN/MwdyEEKBMJytZ5D0/R74kjZLCljIOIGRLNERdumineC2CT4gr
4u6pk8oYq9kbOGw/QdvlitUkLopjN+M9GXrtmVuqKl97n7y/vYXh0To0Vn8pPdCi
ce6lIF93K4f1li3AvGnxPCVnW8xD6AALTfcyT/7Ua6hMRBdIbkRNvOtIn6RXUgRY
6wBQUPyFFylkZi1yWEFhQFVpPd5o8XiSdGhVy3Hc2kHj1Unq3ChYCrjNJzRA0gFi
dXVh54mIT3VcpE7g41hRByckL8ITTSUfHhpdXaY6skFxz4Twd4IyWQO8EUOSRl/m
/FbLstkIQnrPMbkL/2ONysSypfX4wFHvCsFd3kQFv75DJ9JtyaNGJVet3TWorBtv
ojVSL/VnhLDVhYJBNmYhan2wa2MGS91FXVne3s+/lUY8VMitkYxu1Byi7pq6gIxp
LhEKHJ9hpqabWjb9tu/T7Z5wPFIKhc6WItMTu/4HRzZQczLeepDNVB617xV3WJgo
P3NfMqavTJ87J+/zdPXUIhphIDBqThQk2BVQ7USN4HkXxhln9s2Z3sbiagPoNvXg
4Ip3YGxmM1cdlaoPewOJF3mB3Iq+atQyLjxyd90Ip9Av2ycR+ruyw+MU1PHTXeYy
mapo5DA36N3//ywBWJYKPnqw7hsEVtDAsSxs2tShQOO09BXOw5K8Wi1ClrDeyqNx
YCB4YUqME6rljY5DUt/UPHaMUYnopEKcBSHk0w5kXp91gsqM98tW81voMJyPixtz
yj2yJ2CGKZo7eyXgaUbTd7SzwEss38lIS2yRoVmqSmHY5nM05i2v3y34Z0Phzd+K
7Z5BHH/6/vw3pWvM5JqxAZmcGjZ/iFuAzbwpgELqbgsGZUSdU+hAl6sVE8QYzq7e
yrs9qTnwike2XJQB+yL7gzUzmVxNPZmZ+bD/aUhdBG8monWM0JXrAwoeIg4hQDg4
QY0xx7u6IpO/TICDdXnOMkLIb37gbXgrVzwDlzT4GW72Hw5Fqs80RCZj8TNzpidC
7702h7DCJjw8pwCZRiiNHhJlrz4U8Xr6BF61AVfIUoWZ/8LAGk7nIY4NwTc48DGZ
tA0XqIEQ7lVJrKZ/iI0qEhVgCKasBrSweQzW08AkD5UDXgGfbcf7oMe6/NxPajLU
YWuNKb4FPjtaTP5GeVZ4S9MYvzsh6HELOUT76ocrWf93Hh62UFGGsT+PiO4L0Q4z
JnltWLO0LzFxJh4GgAHcv15mEFUdqy8ckbehZ0Cee51E31p/NopxQGcAUr7SrDRG
EQVDzIipqhpPAfbU2nARGWNqZUmRhK008mAyNVBGfoemkGdeUGKRShmHsfm9s2HL
pBcxYW5dyOgixx2btEyL9LMSZSlIWEuvvjkv9k2yM7PcvGhn/MLjhaUIcysekPbv
a+ynf/5rbAdR8xqo2Xi89IINPXGCYz19GIXI0HvnAmxIODtDMre6GVwrMX7LdRER
xPUENlu+d19pDJURRH/1PdvSZBpGuQm7FqnWDvxL+QMI5h3WmbNWLrJ2GAKbDH2E
zLs7UmcE9pzRLMRJvwDSnyC6OGoO4epN+RFlKvL9Bp4WQ1AmfUaay0soG8p2BtVr
ySeih8k6ia6auAFl1Ucf+KQjbMpO+9WhKFLZVUHiBGhY7F25a/d03vmhDGw0gvk6
B2eIdU6/M7UE3sZbkrszCtONfYAnn97Zvz17eKAGP3tzqYSM5gnwVcICkK/oAR7s
L7Qokfu7Jiel2t8wuW+NO0ek5GawlH+//0Mh+xdYVxPrffCmzYi3+a4lE/Of9qDl
3+hKd9NuDR4brGs4K5OfXVcfgetrzdC3rwsqYOFbnissf5pUPyRJJdXPAc3UxiXV
epeFfTxyUPZ+b/Fo9EYhnZIqSJ6Gj0FKAyxSbquXdzhNAVUKlOn4z5jmyt6UGMMh
63zY3B1rgtQp6duvy9y7YkokSkfn7CQQAiIjjA6QxySJKHvoctSB+/qNbRPTzuqs
XTdJGGd5LDEgBUctgy2EsJCU9pOr8Z5vpWDC21KXdnp1Z6bgiBqI12R0v20NQfWo
FBui+2zET6ZeG5RMmzQBLCnWFwGUaApMdvzSDUpnC5PqrjU68qKra1cklDctRTdk
ASEvBjtZUTwaaV3G+ERPO6h4vRVAP5XRpJxI1EaxJzUZJJswrzh3NmrMARcgKTh6
hIuH9VccrD97rcThPuigNrUVM563NA+IVY6D8h6CT24YzAodjIwVVcuO2NfqG6BO
lhGKXKSPCBjQfKOV1vn9V4PdrjtIPrdoOSgKObYkPxG6fN/u/jW6sZk2WL/J9PLj
sZc0DbXf8MHFM7X7zyuOm7T5krm9vkSj4I1WHtMRN0w3yGYV+UjBZhDuFIUnDS/C
xM/CV+DV4f9b/VtmHeXifpckWqloaJiIAl/V1ZSBZ0jx03gWvKwD1pC8CORRRpJi
V1N0fCQAXc64yXrQ9gr5PKD473JbUxxi9T1GEYsM5Kmw3AOo0qe3j2jrzWKMQTW2
S7cSl62j1UdhHy270Fi1msGxRQ71RzSdS44lb7hAdwlzACjf79zRds4gQ40IFX4J
A6MvM4QKzjhvwfjmMtQbeGfADjkTmAJMPAW+O5ObPm15dSQPaeB79qQ0JRniTvSM
Gf0/0mm77yzQlykLF6+sdXdS/OKVoaY3rJ+ZAKb3XA/Br1mdNnZ0Tdw99+5XLs32
AdOACaMnD1DmP0snKq6+GPcvZ0oxvMZ6k+Ja27EVz0IATgWcjzxnb+wQSgGo3Gk1
XmAAz/OOiudjLxiqCIZ5WNtknPYI8aneMx0JeMi4LHRCvfYdaDpUGuyejeEGAUiZ
jDzL4j+iP7+QQNveI4lAJcSUVggM0UF662cIYDQCthFhAdJ0eIzHqNjYHnSFEbVf
cSPH/zPjoomRZyAqnBQj0qeigOxt1XaHWuXfGPwKPFvnjzSNsKjbYi3dWHLjySen
D8e8S717LTPF7ZMvBJpcT3Wm2qPX+/jNVZ2OpdPe+7Z88RcNzZkCFCafoic/ORTm
+XibvTj1GgECIVmoXhWmDBcspszUrVmPrghB5Q5HyhRYdRWkq/jguD0l24ob3jce
hCditNJ43bcv1VrCGLQjWzcu1Qu6QJr0u3zLXPCxi8JGLb80bUYNNe0pIW9ch3s9
wV8NbTNE1ny03+ukcmd4qdM5Vh0EWuDrV0RcIUEe4JLgeW4v29au72GXVEMcSrPq
WGFBNFPBq/WLqLlQ4zU6xET4/1KxqM7IrjPo/O4b9W1I4MC2uOBSGm0qTkQGkioG
O7lnQwuvaHMTidWOBWgJt7SREe2RMn49u46p0uP3wxchp+5/yHo5ZvthlFLIZk16
CiBrDhUaXbEDPtGcEkevUj1vbgLJi+f7K0bm+DgtcTc38A5wbdWF1UNk2Yhs7lPX
rxbY5SulUnXFpRs+64b0R67xZTTiTrKCA9pasvCCNwnEkIvLUW1CEMkr+C7Zvjb3
0vlhEx3yNdUTbC5k//Wxid7S8vxTwXmq0H9HC0D6lcS2yE1VjX/MEeWzQx6uJh9p
fKvCChwpICQ95hOAhkqupeYk7Qfeds/f+3EH5qH5/j/eLOR+JA9iF9rhI/2K0o0n
cHK4u4gQedoMSNHHREkQSIETYGBpY5Nc8kbrN/zoj5mB62/z5d1+jpjhybHB9ZWn
OdHrl7Mp9ZS2LH3bJXigtHM0hET6w+Suy/+6fZtI2BNW7xX8iATG1kLq7julsgiG
/Te+xQBFJ/3NGdIZ2oCf0ElpHz2gmck13f6kpyd/lcnh1kpLV1m279nElTCrxoRL
wsi0/rQQLGYM3bYfvjxZJ8bvh5VIp50R07kj++rRqGnaU0wvwQCybbDSszwcZMFf
1QNZm+xDRDfKHwbauyApDGIg6DhSY4b3BDgkMQU6tJJ+iy0RZx3WOQbWNj4zkMjq
Aw7f1U7C920bJ3ffgAlBORgB0J+HOwckz0x3sPp0fSY+/9Fk+3rWYy1NKBUUnTl7
JbPMsNOdIQkQxsBeVYvF5X2d2g980Rjfa1x0wO2bPFd6bk5u5T8rnTCnTHNoc+VX
rHobuInjzVkLHO6yqtHjB0m5jY5WyzVYB/X+C6lpmyUSZmQk/6xRB3FTC/fTZVpf
Yt88rs99rHr1uNcFOmbvdg0c0lQrSmSEmvRWY1czpJJgfGTPBxvpMIKBZ9BBnpzI
qNe+qpw/O5DhJWAAEN11noNSSC9LiS3KEeYzhsE9OPpgnLpDkDCcDTciTlDov6In
6GfUkLzVP+spQyoINSABl7DdXtRCUqo2tG+FOtNBB5IIcQxaKB/l3oFm3iEJQ9+I
zuZwDaTHZ/9pooIFLCdA7NJiscfAaT5z2a+2XB0m5MMX34R1bRtTyCOYX+y/bevz
74SYmtxtDOoWlOAaCu7h4HS2XMepFpgnpxY6wZpG9hMcVupE4nNw1NKV8XY/5q6+
RkaNYuBHFxlXte4NJuDL5FwIJnwopes47gQC7AbejRM1ikswBeJ2OoEDGdpAyNaw
snZsV+9C7v6BZ/oqe5PNGa7xuA3Vd4h7u1JXx0/UK//ST8hkxJkY51CJer5azVpx
giPYGkcb9+dtDWfVyCwj5zJPDB9CfczfybUPcOYf6QVcQ7P2RpSc7vz5lzmGZNva
BTmrrrUURV2qrUYYUr5fvgOkZFDDLWLXI+vOnXKvbNJB5c+I6y49+AqJfG7Bajed
xadyO9r6mj1Pmw8X+9txzED1Sy3LImpWyBSqhjHbRWZ2efQDolzbFKeX7WO49Ym+
B2CGTB3TAc9DRtxxmDI0NePemXF7eBvjEUPObfMG+fj53DjsmZJebTyddPKE+09r
2y3mYM7DCa9vHABaOMOvH1yLwWZY3dTPOtnHy4t9gEMFYPaVC6Aev6kR4a+P/mfL
tQXadvgRrWf0NqODshpmLquWZKH2E7Es7O7cfB8hON6KZrlEJQy6KEHubzr5/9qh
MhrNRYZLXStjzNx82fTZn46ZfBULzMG63cjwQFpzU1Ujf19X5YjNWLEW6UomrtOC
DCWxL7J9d54rh5OC4EB+TUi4ggrWrAxi6htHVzAYVFAT+Sdblyt37iXDQ2viZh+B
dDXexI6+CzyU/OKGyibJ2rxBV0AMxx9BEKwPSJTRgmAwQeX/gPbTF2Ffic+EvLuJ
o4aGdt4Bm/3AKJWzQjiw7svLEO+U9mFl3QJTl5t6AnFObBrcT8wBWAwDzIQ4mosa
iZz9Y80X7KHF4Ra0msuhiM4K22vRUEInc2OBhswZ5GuJbMcVIYdVlWBvkYQ9bVJp
I5Vq0Su0PnO239kD6igebnQCK5mXEM8FgFlnZvchg5PssSA9C9xHgnG5qcq4ETGA
aYwRKP4BMYBxkecsuBDv5SesXtGeZYF3BayovJJCDiIeLaryRyf5I8AzavnEWcXd
HCkwCDcQbaRWv2Vg/2m54IzRSImtiGyZAvhfoTkurns+2x9YFILGzPH4r+V5c5jd
bVbtxT9bKa8yvQNuRIe1E5zNtNJOHfa7QKhb00XdOLcb8QB9W2oItacD+69invBY
Q0+6flxqrE3XgFoYJ1WGsanAsvvO+CoPc1MvAOF0zdCI9Pqn6vAtcXrx2qQgCnP/
ghd970VB7dzWAhEPCd/7TlKH4lR8F/RMql60TJ1AvjMizSTSKLTG2jDHazdRN8W9
TUmDHBpSY+k4vOEw8aj4H7fLQUjt1gG+jiFWGFf9hQT0AilR6Cn6sOJXzZYEwLBw
A5rX35mzMyvJRbyFwh4kWgn+VFgVAVu28XxmP/wS0ZB0V4Ft7mnSPrfqAxqoWeSw
hDyflUMe9e/QIsCAiitbKt8KYEHNlbnwukPwM/GwEkqjfGbTBsPSTwJw+YtCd+wB
+uBgjvB/0fluySZbtr7i0HrN0efq9tBL+wGsqSbgeoZBr78+M5zk19MclYaY2X7N
t4w2QOHuvP7GnW1LNVYQXrb0E5oyOOvQ+aG7wwCpLIQnSxz6O0T4V6c7DNRMkd4W
F8qoTF1Wj/2VZEJzFlxZXWOb6kMdL7sh9qdyNM30EMAZF2qYRc0iXIo+4PWiKW+v
Jpl3L8/hebNDL+Dt3OOVszmP6Tyvh4Cyv36miWNSIWjV8NPUqp+CYLbDGHFBBzFt
WTk8p6qYw5IUrSopI3Fpw2Lg00LwZmz6ubENWdiEzLDFlJ+VAAvCW3c5MMen5mm/
3JUJkNFAVklKmGwDOy6sudo2ecGos7atzVRHIZX9C2zYKJYsO37j8fwsWZ5+F1iX
uSXJua3toHsTEAi5hEKY92x7UsYHOt5iLeHLNfOErxM3X1UffPfMlprZi4t0E7BP
UAGc2ag548I/LuFFjdpd1SObC8KOu5m0lrQ8/nGP+Rt0t69ylhBPsTi906bDIyWA
4gZN94v2bMqHo6RgQT/Ml0lB0qZh3UAImG20htdDk3Kc4gXuligngFpAuvhIWWhg
Yw6VIVdAV2EPRDrrfreZdu0wXwGlqc3SXZiPAg9Br4e1CW3NzUFCbPLcrQ1TVHME
FOqePp+e14rdcB+8JDArm3sxo9tw+0RPU+h9T4S9CPfICUL7LK74NVFvwDdmtYI/
gHqVln73ugtKQkkyqdVj9es4jpjxIZUvNuKX86XWY8I7Fg1gyFfQj3/H/waCVQH9
2gUywfIawGWoVzGpYrJC57L1UBFZ/VDzteM3LHTNuq8/56BGES70yH+tIdK11QY4
BcmyOU+trQnqaKiFH17uupBmKba0+ndXXCJcyFu+p5Hj5N/nd0oLs6XAZZiA5uyv
FOW0ugvudwMLt/y2Q6SoOUPgYtFEHbucrplk98mxXnk6wJhuTg1u9VwdQn40mmWx
57u27LhonzdCkL/DRNdgQccDUI7c9RZbzzj1x9OiDZf1Bd55SqFlnLl9GokrGyGs
g2jF70H4D1XcCZ+3Nib9IjrNn6a1kr1Ew0vFOrt2D1i2C/vt13Cj3z6OufFv9dds
levFjaTFIv0virxBBtVkhPBqlNnx4xUcQU0LJ7D8h2yJUQObE5Rx2d4ZWBxiJh/b
ueQ14V51+8Fs3pAaUrxyZG/p4/5h1Mc/huj0oXg3cZ3UfSvU20kdxLC7paQrU7k0
HSsZ+SL7bsOGGQaJNJjqTkb26kALm/8KqCUdSg8Mx45pPhQ1QXACg2mv2eSNfNXE
3xUbaTer8KA2VwQdeqjGInuJ2Xk4250L+73cf5LQoe74hZlZBHXUT87FyPAosJYp
6VstZDgrccX9HxI6D7YT+olck64LCkmF4tB7UAv6JS6eIGW5u9I1QOXOvWGg704J
88fXJJ5Kt+M2S6PraJGdG0FCzvRWUGHeQSkH8c1dy13NkLImOPfBG6mWaLgnfla0
siYM8Qf7GJ9IDU5yObfKuzgNwcaTxv3QMDRSjRej4ywJFVHtpeWEJtJLkvPtgyNf
TwOfgbt+xwgEBqTsBlKePKNiERu+LBqj+R/TSj+sBybIYmKTc5YzKpu3LuxboOi3
K5CL8uDXZbD3ZUGIH2iAeCtJKCW9hedojXQw4kJ11KN3So5SEtWrkVTBJzvrtAyu
fY1WuJaSNaVO6SK+aKNqtuW8dodL06x/f7ViRZejHxBECA3DVrMF0rwGQHQcblEu
U7nZpFoxqlLhqxx81sDt6E0CghBidjFhnRyQ5RoaDbaTw+XwdxC/nAuhJ3gzScwv
3Yvxl83MI6yiwt/WVOUW8uaR53DIiQ2EWmrHzMHoLqmWCfrznBCMSzCusgFChtIK
EjRJwG2CD3IJ7p0+ED4pIMHJjucUp19wmZJ7Q4+lb+LUVnrq10gxjDRMHKwexZ8d
oV90gDWp0kAv7TepghFVU/p4aUUaf2ZIk0AdN8QfFO7kMXpeIS2oBONsnoalKQFG
16ushQdUyGdcHU4trqsvwMOONi0xOu64DSAgHYlvQS/Yn9ITpBQJtDy2GcPtbifp
XpS73KXMGUWxVQi40oD1fW1fHK8/R3ZVDfu3l8rZgGvex/Cuu6qXMgsrSl2YMpdP
qxgCY0u6pgpEAjguuMi299I5gKCxAXn0i47qWyTa4nmWxEYu4Y/grasinepjNOz3
oHqHVir/iubJDY/ul38D64lpfw4WR/L8TkLY3/UpcF8aCUqvwNPiC9NF0EBc9g96
KemjiMXg/lDXEEphA58jT7tLqfjDTDN/3OCG0rSv/Kqyz5JbJ+Zpd4tFWiQJmDD4
PN9XWT7uAxwS2Frv4oSwYsPbZXhsMkZ95M+BhPQKV3fZ+PQYqe37vMmpDnfU7BCx
L3oEEbhuCgnuIDyEN3g022mM5fphh223jbyUqVLTZO+bh2TMao3W+kOe5PvitGC0
/0hSEVFueR7PGlWEiqiRoeAs9LgUcjiKCjGHgAV3Cilg3topn/syQAEBjAk5/oqa
F6xDdyx+j3iCcX0yCYLRlqmT9gwgvWLOyCabl7xTIrUk+bQFVEnItzWK3kA8PRAU
fOmbte5pO2Nr7xc29v4CFPvUmBgaNuO2HmwgvKFJ71Gq93lKm/lgw4bX2k16+iBW
gpIio7deY0Q9ujodyW0qFZA39618fj84Fn4zMJu9bJlWppz8EcN47sBJrz6B/Tcu
+MtwHpIy2XOA/aSWK7UNcdcfU4oA30NdigbU4qKa+iP0DF/DK5pbKmq7D4YXsAA2
lbEuhJwrSrYkJG4WgcBSFCgnZQSuFudT4zRl0B7OFdR9Sh2YjvluSQF3dRJi3h+Z
qBgbu9xp0kImgdvnASEHFAur/9RBb+m2jnqMc1o+eLJec67sAQNdYIWQVch+LjRY
FV+lDTyCCqJB1blzu4mlh22RrWDXKiwnX2iV/mjvnOLCPpxmvPwUOjnJAAXYJgFC
dYK9/pvc0Y5J0sco7Uf4yLUlupROfgZp1mU3b9Co4ou61iO6IMkzVZXbKdf2SyMk
+MIIfKXX+TtMKpvC9T8VVh6tWLB66FCtCKWK2JjS1MRsdb66PlTsRytbRXq2cwjV
N94oXH1U+GwQfjti6x0iblMXN/nZwMI5NeNE8hjno8TAZg3Q7IdAXGS4Z0fGdk48
eraceN/5lNruDEtf4JZ7QosDYwqNbH+RpSsP0j3rbtDo6t6E2w49QLM+JZo2FJ6K
Wd3N3mGzdcdvjDJEZZOBl5U4S9ozM0RtXkOR8DrI+46lKcjt4D4ouIgU+CtOC9De
w5ksNyH4R37rVrcAUxovxZjX8xvoCM3W0XjKIMft++/hoyJVUixW3syXozJkxT03
IdAaI1cuBXnx656PKnGfrRpwaVtfoX8cQQWpyryjAa3bqoPUEZRi+8wxxKP6QBt8
ssu973rcAUwTXrRSrriDh6Mxjmve5Q9ORGhYR76P92C3Ec1AtNOS/eRBk86sE5Iy
ffuQhiI2m6TAj4O+B0raeBfyt2bmo4JlA4yn2fvx1k5IpJZdIsNHvoIleqgk5yS6
bFcGXNazhQUzuu7xWLOylADLKRoMwj8DlRQKj71zLpEstj+Xb7xxJ1KLzHBWQm6/
/HOUCSny5Am/0UJYNxEpuEGrpQ/Czlrp/gFja15vzs7PEdVK01FhitxNe1h+vhIZ
boJ+sHJtolrrnqioQ0TOfOdBdxrje1K449jEj75yAkayWMMM9+dpLAnQ4oCnsG2F
/6FDvzCTiM0w9gQwU3IHizzI7TNECeEzJBe4FyD2I6vfkGVWDRfVL7M2omhJ/Tra
jATy81xB/nUtPRFJzZo2v5oeGLN1qj/Ks2QayMXxckddzLGX0Tt0H+wcQ2lWumIv
UcePWLiB4Stn7p88iOc8QkGYUMGDuA2femXpQS3ejhjME2JDqOFUO8I7VImusZhZ
kUYqf+Q1ZkYUF+Bqn6Qi6b7ozdTctuN/2Z5MYkxZt8l9PLlCSfxj31h+3jFH5DfG
SWChiHEikfHODye5LJC8HyTUtb8qBM+bhc3RMdoS5V0hVoQiacfFYSt9/OaD5guv
t9a+Z2AAZOgQqlp+cZIlNgsDw/3qkVgvbnXOTTBcyBX2fg9US9APpUF4aC9pGN7S
xVAZ+L/ebleVn3AGTflLLd2ergfXh7CtUsqkjd4MVzJCdgsclIx1864qUbZZqKlu
tl8d6MChIFUN75FRrzXerCOGdlJ5R53BhE9YRiYu+gOj/gAo9CHOxZ7tzkPLUCFn
YMdhwiwesxXEylXsMi9/ddmiHwzzDklPTH4Re0x9g1XKP1ZkDsHcimdxerhhI/dr
kAimZuDq+mpC0U3B3SoERyBlFFIwrdN0hZ2evv1k+dkOFtlhO8gvaPkNNuv5Z7gn
2DYpa460q8SMeAQsk3jsQj3LYP6pNe7WcmlxbxV0xLlhPGrJk95iyRhrTl99pkjZ
rGWh5lqVT6nq8+oHAOaF2p/jS0I4z/7ZnbfJYJOf1GvbmAvQBtHi4aPYzci/1HVy
13ktdarrWT4HVmZDzhdFqGCzuNfjUGJFZtmNvvHx70t9vx6gxt4CIZUKc/UCdjey
bSde9jUajio39K6yZfPxcs5P16rd7jF41bUvSbQiEO6JC04u67cjW/dIoCSlAtbJ
EKQ/0gxqGLaYEUp//4LeTP2CrnB2ZJv0bkp/jEX46+r+wJ+KxQ+T1sDuozyFPv9L
s8pYLdkXXQL05arBUPqzUwiYdQZgyjx+tL+DUKWgFYa7lqIr5pGpaL7DFEbW41bF
fukgTTWWQYHb9jlcwXnOnRoWCtjCkg0I2HE+JPJaFG7GZR4tXqtFHQD8yoENecD4
2Y102l9FkcENn4Ec/wMwNWB3E2clWbBuYIKiIRR/vNx1/peyexIqi+FWzKzXcC3x
3JZnKAIMPQWFt8HN94AgpOc68JOim3Cl3GTfRvMX4IguZjvAGjn3+JW12CvjJbqD
eLRqtwYc9V0AWGd5gSDVplrbqLnHTl5W1LJZ67nNTg5Mw/kYcffgOa9BHS6grK4H
tTpPT5LHdAGxketPUmyPnAMbZ8u4vR3OpecRwg6fe31HEK7IBdnZzYQ9HPz4m9KR
bd8g2/aLmkBsxYwMenBM5hsl5gotHB5Yk+WdsPpZ9Teg6GfQh6ehvOPFmPStg0EW
Tf7knrN3Sd59qvMotSXbjgEodkZAtHfMwNWQ5WonptRcDuAknMGiVPZY4TJObzwN
SbDTJVUBq0P3Em1BunAzfUccN8s25qOgRid9s7NEovtzRf/VoD3qFaOIhk/N3zEi
2xvl68KJAzuYyTEov1H29tIz0n5TJKQzbEcEt4Ib7E+UVo9MeVxoletAtcc4qMJG
mhEGnUvBCP7VZ89Rm9D1i1hZ+3VgHYtmV2iDB4jC4cfE1OT+ZSoRiInQKUJ5FxLZ
3aPF4dkEBVPpnLKJi+FhWkG/Z/4tLCr3FHwqdwlVG6xcnzSMRexcjAYBo2Y//BPV
8lTgE6wdHNGnXeY3y66FkBOp7MlGt34SYMQVR8BQ8vLjFpM5bHX+k/q19TWCNEyl
oKU+RgGQLkBd8Qe929CJZTE1JXfo/YFoxxR8jnlKFcJmy0MsY6bMnrT3aGcdlPDt
gR217NxKZbROFiJW5hnkYYtnHx3R8rHItKEbujnjArV/KZ+SDVmEbabQmLmOzUWW
OzVV/kMTY8NAg9xQfI/WTbw0ZwJN4pHwYBIDw5PbLHgMTnrl3SG6LeD11IqV3Lg6
rzOMqF6GGSQkZh47APJ0aTJmI6EDEQWxJcFdiVRjA78Gr/GcfH959TZa7lBqkxqE
ozTrz20qqGwoJon2Prte5LvqJMKdW7jQbCvDHr2BjEL/SNduB6bZ+OLdxigiZG5G
fGXLjc0WIoninHyGtpO3KGZZAaK1a1STUbuQhBeCEaHZQgs+ciGNZXR6GDzX1UBr
lww6z7hzTQhdP1LfEHUsQZh8YfjHbTlpbpvrGQNVVOtwAwDr2kED5K9K6gVbtiHz
Dw7B5sYcXCuzDNTPdfJQTCusWsy+PwZztTtOEoI1OVq9HuF7oNtSDQp64snEuJ9n
ZEBV1sk9OlhUB+ypA1XPkU1dllyMlPbNE6swLflOAzDjgsW/huLaj0488tPi1ape
UMFBG9B1xF05W/FEb91VEReuvKP5HxmUgTAIOrNPfhvtUwkbuKS8SsZRpNUkmOOq
3AqAa4FgkOIrT6Qk2n068abjpU9+wTaMWqU58MEDITaVIkiZznvoU783hWD6Rd1D
mcpg+0RsrfwAr/YEhPBtC2mDf32e/cWfmujfBzkFMChSTIdvFtPH69fJvsaAnMIW
lUGyNpQansmpFHlLvdE91zFxqGkPBcOFtolthtCcCjyhVTuXcjvzI1g06VDOCsns
8fPS9oxrhNUoauxVs7gK1YoyO9ciVnkZcj8EX9WyBbgCcqX6Os0BmInZAUoNesq6
cUlRGCdOutFFScY7apq0BS9srKc0c4v2y5Tu0CPDo6ngVTYC3E4IprUSHIcwg9I6
gVmOBkq9Sxt4ArBK6J0KZ1elNyKBcoR//Q4JbriEQFzRbBKjTFG1ctyfcmvYUuUy
TtV3q417ymF3yBoNaq42AYTnnBybN9Lnf6fz/8LYhTichHEFoqW480AOvU0N02Yi
xnxk1gW7VvV0m47GOXOSCHNqLdCPOHYNSSyTnk1cD2aeEgzwfz9snNY+idhoZHXI
PS5PaSZOk5xWD+rqx8v5LBBKqyqSbTRbIKVyJ2EXi4cGZYgwptdTpRaNaAMfpPcp
6Ip27ZemxwBRYZPP7fVIv2Ll5VQZFVNmklpJUrccYPWgj8128YQTIQwtZfCtkWry
a5YBWUz6SYm9HpEIprZeowMM8UuyGSLA+sFFC1tfDsbrIYn5Aw3gx75qGsAVOPuz
bZlO3Y/3bD/QD56nj9yvJ1ZzBQfzfB3CuZ1xZ2ajp9auSo10DPJVxioU5+aG3PuK
UYPNChFkKqSuRiji06vHniZ2iWAW7mIYnhbkBMlyOBw4sFMoL6lx7l49GtK6SShg
8z3B1D+zwv6hwyIGYTyE3LTptvdkKlbqyp6CYQv4RZaA8odjfUWAluq6k5/4gegs
+YcCZn3xp6tK66RjWfaZPlTGOo0WbKEDb2/t6C5ibaDzXUMBNpgKOGBsu4I5hnwq
p3xCD0UPdm0MIVt+X96cLXVKFBo2rAOmWgxVt+kLYEBvLSQQfBNmaXl15gWA3lis
F6he5DKMTSire2S7yQ+e5dbAY0Sy5tOhpvLN35g3T+W4bT4pMlFLJkRfwkerLFDt
FhYmm86rg5N9RXFGBVAu41GyVjBdOpmDjj3/qsnKIpBZmple2/rP2TCkvWzVbXQt
eOIbKWBoLrU8KRfs4XhuI4kbVssxh1M9WvbnvYhgrJQqo2E00uhmNaeLD5LPkXLs
W9ht1dtJHTTAZ4GuaIe91ZzBvxodMMUilBP+lZUS6TGK7S0g+B+BYh8un+vBHwF9
wmA9Nc7S6xdeX7vzgip/kxgIUjYzA6/J01ZawmFwYwM+FcKr0VHoROlxdA/r1qVA
I+CV/MwCUjM0p6lOYmwUQuZydrVBv30luFpdtobDLGQRPXZXmhosc6+PYvjOcFh+
++YPzAVvQSe96Pv5soVj0lKH6fPvzfy0xw/e8QS/iJGrwd9+0f29RfibQj4r6cQT
t73N66LjppHHYie6GzV2pjMatiHtZmSbJ3Vo15/CFstKR7tv1gQiSQSKAVi866m6
rVrvm2E9yOph5muv+a4rlEBRvl7DZvBmIKvNJVTEV3MCgAkg3pR5/lzt7MWugh8F
W6oxfzEClU6DJTJXeFpRy4kVnoXuezS/6TGIc2cEdoZ0KjqKgWCGzytsaPkQrGN6
DBMzSLviC8aeF+xLc9h38duWBPRkazoN0JqP8AJKWi+jT14F6jItyJ3mmHstzcAW
RWM9kcqa1TbuMFPTa6I0C2PfwfZ2lqA4rsRAMEHPKhpjo2k7e5YyvPEXUl0ZmD7R
XBAxxm9iO6YKn9/bLWfe1KfMkYwc4Z9DxplOGMNZd2+ft5LaMt2pfffbxWchh2qi
HB/Gk37DVjXNBh1lP5bN56O+AYMVX+nN4RVfDJDo4XpStt0+ehfc5LXJnTSh1Uwh
CQOrdHiqLYWXZ1Tg3BgeI1VADFn0vANIOKtYuhUidWVit8MzJfUbROEf/MkceZT/
/RU74rfViqwa+FA9yn+jcrDvx96uaQBwyICXVcaBOxG/7TrOWbSzwrhEohwID7c1
jaayELTKNkzwYD9USx4KeKDhVC2e2JMDRQOLLCIB0L1UY47HQBI5Ko4N8O/3HvQO
+Gpumr9Oj+kfdS7dtX6r2YZjlAKgebzgC6ZEefi8rFoR51H46nm+QbLYJtTIGPeB
/t9zfRq4NgYEwily3HT65D0t7UoXmJsNDruVsFzGrbStQE8l8tP22ir8XCRJOg+j
PNZ0hejQ3fcyYz6Er6pXUtT5ekL3KmFtGSUTZeNJ2qAkuS39S8/J/nQc+LgelRXY
mgXR1qTFPpoEwoOLtEYV9AHTVcxQQANc2/Nf2UC7x2Ae/MXyOT50nIvSEQNH/BAs
JpOCo/vUoXiXbkQZ7Sozw+a7AvCUyKzsfapxutk4ZPply5wwbRHyaUFYOj9vBhDb
TmLSpnt7aTH1wujaTimmV3kHryelg6L1VYZfrvUcVfvhuuumZv7f11iGoT/q0ExL
KItkknwteGDPWLfEbyOIQva8GeLFByHw3CPjjdgScIQeBydeqFZeTfGQjx328vUo
m5PCXvwDZkM9L0S83+IFSxp0EtbotH6qWSg5URCzCVjG7bfI/Q30xtmzwXR6w/CO
CM/vwNQgNPfZ5GjzXWdBMraQHNJcgvSpOU/72frBJmuGMkknxzQpW7ZkS2ibSJYQ
+30Yymyr/bccNxzU4I6l1w/t+oEU1AFBE0nGLogJeNuvi5p40dt2cGk4TpIuszV+
V0FEmnirDlbppBNqYQH4zvIKcNDhU8zQ01Xak0xWTRfyDQJYo4lqP70ndYJm9T25
hUONbSVdmOnJjuvnd+qrNb/ZxTOQzHcbnn1AOmBivWWmc1WzEVzMNL9vj5srCwrz
3evrP3RCpfwXh816b7T3XP5GJnvMb+taEZrtxfNwHUAjy91RPBgs9HgqcptjQ2fR
xEFxxoFFvQjGcNkSaDUfNXOlRskgvfMdSGVy6MnfYzMfNpkbLSWORArN96OGmagr
GQWsuY8owoKG7NvZMG6X3aMWIKZrW8Zrd5qYvrxRmhul/hsXhfH4YM2GeQhcpNHY
mvnA6CSOFraIaAD792xS7UGoyklqz1q6APnct+Pzx8QcBWJ94uVPffq02ASVnJ1w
MzjUWorJra6yA91hzRYT9QZoX6d3iNQ1C1zpu1ca5nGDGP4Xb+k7mN5ma7giq6pR
UGcSMeiAy1mOveqm3DTk57vTtVUaUvKFb7edEZc9G2BpsWUIh3R0Rpo+CsSOHjD/
EHKtTZw/WlF9l8G3apaCYdUz0INS7LzbpuncMQjz1FJ8ha1CrUkmrxTRlY5NW4TL
502tccddTRScDNuJ8FkXBe9+EYCnl4dGhNAzDR9m2z4CLrzVBMTnuB4LthqRNyTj
K++qCpENTCLGD+92g6h3DdgFM8riY88K0t79g7hMVumEK5AboTyXbgMTK0R6lFD0
oLtNBc930w+C7QMQpgDqCWhKh22wZnQTBy224ank6CtT9mS5iCmp+fYeBnNPkzaQ
h3032K4eErjJHHttPdFyNKqcW6K0IVevIp1rK8X1/1F2U36EsqexQXAWVhq+GNiN
nlrJDmj01My2v6OO5eLycnnxKTWbyYc8GnkAtbvGSdk1To9ECBWK+BTJ+9YzlhUx
AE+braNpMrpj0YrczXmchwZMq+TQHdKiiVCcY7clp9ifM/7B8Z8O04nmv1PKvfos
tzGM3IWbZ4qkbexUeoYxfmQeQjKF9ejjNHpzwv8p3uCa/YdxirgtKe/eJ+mcbsga
fJD8ek1HkJVTrePwv0koTe9Dhc+zV2KZzCYZIeQD/Dsj4DtfkkGkPIAEU1JBh0r5
XfmnxX9G54G5+C1lc77c3LEfPjCZ5OIh1t+g0mZn6np3mNAx2P1w+7sZBe7zjHyU
urV6WYDBD2Y+erSoG86hcVIg2csM758YaQr9TI0WVRev2vPxVz4G8Cp+H8vOV941
ejuLZ+S+6KeFA5gAZrXxY+L1uHB1cSH9x85q8qbBIFMMe05eUL41RTpxOWWYYmgb
jrc1GfdwPy0Axjl4yJK1d6SxHQBV5jnpnEATfGeeY+3xC25GoXvsDAl8NRoSxl+t
zB5pPeNhegsgCPzEncd2jRf+IPgqO2RoGT4b/9QrVvR2wL6UiAyal3ULNsQCfkVh
mhI8zky4BkeyTzjZnnH937EIq2e1zZjIdMB6qWUPLSnDuq+7qTCax+Ffxs83/UYn
5Kp04A8EyMOSLfhO9MnX0O+wTCUPxNyuQolfx1bhIVW1zj2fG7HE6VrimFspMfIy
LK8i9aQ/YrQHMOdKBgkP7Em1hOZsNTBG3brOI2Xh3/EZ8Zl+iJS1ZZqsjlr6PQVH
F1GD0cBr542GX964ElKTXr/hcb48rLU6lAiW9n0SrpVehKS2cBx/YCh0a+rrshBq
pVfvbdyW6Haoiq87DD0qkwemHf3JdtDqsgLZ7mGdYmQi+g+9uWPyO9vJCADy84zT
b7FAHV5rrPNd+Q52dhFT1u3QbnsyhVm6m+gJ8U4ObzMUqTOEYWQc6XYuAE7usDnM
2r4tuvzBjvNJ2vVQN0FrhVtzGkP8pk/FqwYimE8/02s5NldlFpM6tOh3dls4NvNo
sumxPN5pOW3w3sd6+8hZ87YOSExtn4YGti0ZkJp1gtCxRCA38BZ4OnVy85O5m8r/
/YDICjLmBU4hDZfm/Kwua4qj8zNoEj/P3EQvnFdZ0EiaDZ8BWRuRW3SHtzXT+lH3
OWkaq36LnCc03Vk3Myjx+qQM7df2AyueWW8Hcy8m+OExtfJikFXFvEuzyXUJ19J8
Gy5G4HGuyl9CAxzl+dSOQNeBYYWfI2Dbdne+hOo2yeuEWmGMxVjaBimIyiukerYY
+Ja8Vw6d5HFVlVGltLHQ1NdEn58ZnKQXnC+wkoZk4YtW8o6a6txTczL8DntBaPK4
fiIoGc+vNXmx2I+nv0h9auOFZL5IrFIJwkajRe5dg1hKYUw3AFgkmdN+OQlZirOM
asd96HAjyVK8L8kvT81DVMZfbemL9LgAh3eoyDzQm8MPQSUpU7owC2FuqDITzx2m
UZKuOuwKQM4SQdk5azAXqsvWPQjx9KtxP4yUToTXyARHuczfAln0AR8SNsfOUCgE
TOscThYxWPgo64qFOiCWSL7gCaG7JdcpFk6VB/w0qpAgLgLwjIrpOl6so4afR2LH
2B7PPad7fENMhCWXkuAK1XwlvRlJFpgGhhb3Y/u4/bSEmiUyEZLLEbjXhMFl+3iZ
Y77J6smKmhC3thwGGoGiQvI/s3yk3t2rxbKPCaP2jYAihdA3v+GL58uisJ4rmb56
x8afQCpAppBMWev6bIvq09PZ7t8tSp5MvkjbYZSOa60/ypcACJUvGcjFn4PZma9R
hij5cICL62e/pOwJlTWpnlgbsNbFI37BlgjH12hsJ6L0nYZiY3GZnemAHotTcITR
MKtEFv2KMG5Vq/DuZHy5FDgstMnWD+DU8sWHWuwHk7C6/k7WQw6d+CyA/GQ/SeG7
32iI8Wif3PI9qNomM2XYzC7wpdIYma1ThoDAW8k7t9eWO3V8MXcnyDclvTNWRGJl
pweDxucq/yc9xS/kSNWFnJ3x6ILxj/IOviyj+KYtLtmKTd1Z4UfSdyqTWVB6r8+A
THYwAoTnu9+VJVvJ9RAHg+2qUJryH5qs5JyWaxX3UXPY9D6UhaOZ/iSQq7lM3VdO
Z9S31a6kGYnqofCjUlErR6L0k8zzLY346zA3p4/m4Jg5OHyKBt3coH58KFnkLqhi
eClL3MI4cf7M+yFf46Yq8K6G9ShlBWml1flmb5F+ZgHRs20BBVmwgak0BVSSm/KG
nmYD57sO3q/+Mmye5LiAVXSYQq245IRgDnBRY5FmsaZHYca3+OaaDNTqoOb0qjzc
jgd0bg5PEY92dXCi4qI90r8IxkmUtfjxONna/k5nMdpLYdzAns0JYd6BOcidtRmL
O9Z4IC5maf8vInc0p4oSdwgOL7mUjuR6mkTDqtUfp5tEAGw+Z0lvM9zLxG29Cggh
cRSECTWbEyEPEm2C/yhWC17WHSylJxZI9p8WmPc7/ZVkefYCmc8PeQAggsHEbfxF
I5XMCvLftOC/M8ThrGtlwZ4o2xeImjgKXZo4qHMSSEmV/Mg8s7WDfLCb+6uExliN
/zz6UjGHKpSpTQStoWF5dNKNnG4/wbvlFg/pEIvi+BKD9vd0virSx2/uJk66pzBF
IaopeXdiZTcP/9BxdE/Ch/gZToad9HLA+kk64vROyanQLURVr8AMjfajzho9gBkp
Qxhvi6zSgilPZbGEex7cN1mYf61hroRqojDhOVEnJoCJ6NuKlsJReky9v1Pi7kUM
p0aTiqHoO15LFeij4NuAn2Njez6MM89rrGcJnZcYsO73fa4iXLooxFVYy+mJfY2q
wN+6hlw2JceQJZfV1z3fRpjdvaQJ5hIjhAu3k0kb7RlxDk4H+HBlXzzeIAOmKkKu
sWU9njxzLKSIdwz2dhpKQxOxQCEpK6BvFJIi3y73kyq7uqTrqE64kRs7QRB6pTsU
GPwtHVAFYJv2RRhlV59hJX8XqLyhYYjOV5YgQ30RkZgOD0CDI8/GcE6uXnCYiKe1
n87p5klUhBoHYqwgdjKTweCCZSMCpOhbT1k+4gxO7BmeBsTdGS99+M4JdIRFD2hn
+4Tp0aRirTYa1KLIcfZjXCVUibp629Ri0/FqeReU01c3txPy8kDjdIdJAV2w0pju
uHXVjzxqsliHMeweKxLCqkp4VwUqm1usmkv6zFCJwCOndUQXfd1aJh3AR5Mrfk1Y
Eex4DCexdna9OBNchT90QVkSptwc9+g2ZazrUz9q0HH5Ft34PgBWTVQxHfGQN5XS
f1f54Gv5rSkCNwbqE1CI8PLzDhWb/K7AEYC6XHsZEDVxcsIjVy6E+zYxw0sKf/AK
lUY/a3X1fq7HNMELpwLe/1d4d4uirXAH4LwWjzumpBdXZp+cKGuNELz3K4w3Nyot
AVnvOuuKGj3ncXQphSy/845+tiOMi/KpdivOJ4iXmGuS5wAxIz7DtxrRZlu2Tp5Z
hdLnrizuf3cxFQh149eUMck2DtMO2HmkuPtPHdeHmv1kjpH8gH5W91B/pd/QhsRA
8jNGyIEyKMGftFcDgJZsxMTDEKVZQ6pTMj/oZEnoauqPsNQJV8OzMak0C6mvU1Sk
Zj+q4oZ3e7Z0MMJZsgGjWsj8NfbW0CGgAK/sNmlJhpWkUfgD+rtx9brODgz300F3
EV4Vy/XZQVAertdrdaR9VQ2uDoJZVc3dT4JbcpJTLyeLdk5jZqz3rrO29Py0Cpmr
j2AqLHgF0Y8cxX+bKs24MWLzbG63pWXfVmFCZL6kNSLRdw8Db3PQKIGRDEgz8y3A
P6s2RVtgva9DYRrgO/lzh+1d4Q9mMX2U1LBy+bVaUtQWEdoY5qDh52jdM5pFIwp4
nTt8A+1/sZDDcw3RN7g2HLDsXE+HozZ41AQOBj5TTzAJZQhTbwH6EsIvs63tLye7
tWFxtlgLVg68W0rl8ePlZPGlxfnGX7kBMXfcVGgkgyHfiFgW1cmQAVYLWmmo4wMo
S/f+uxqh2oXh9jG7NlX4W900w+SKneKGrrn6JjnBC+NwkSN7SugLhJECJkFgWm6J
uwKhahz2cuiNVD4s/zePny11WntOKYiwePnJ1/c4+rOJ4NdgJSil2K+nejX3Q0ch
3OJvRxtc/7CZoyusEW/8CGSFAvehjQuD79YAl181nyzOmT6mlPDTMiGGPnNnHihY
qBBO759RFMc1f75lyTsh3ulLi1ueK+pBQGYa23sGCafCyIvamIuafutl5FD17RoN
stkxMTmDRlzgZMPqcRYNamNq+MU+BOcW7Uh7moAju+8O6AvTlKTwFWHOynTryw6m
GY3xtpDBr2z+i9jy99PtwFUJoXon4qWU+0vkIp+s7ZhAu5PV0cL2+tweppiCvimU
JoVsAcnYmipXEzx+hNrT1Ic74xOCjYUdWBwI9sl8AukHGjrPXXxIBILuvw0hhFUW
ezQ6B0SR6w4Q80ZCDtwdOJR+MTpwRncXpoR14K0axvTirRPj3tN6yGoe3uAVhJs/
8T2XrgfCRlN2tGLIWmF7/6jC5ad6ykR3aFz2HIIDAtWRrbnUnlpLA84djZsPPApO
8YypVNd6+ge4do+Yehg3hk1uL6PyKcArCKj1Ji4oO1mMFBaRoWox8xLJgloNvJib
OV4EcZpYqDE8pLtcwfzzPkluhhFrqXHhfm8W9tpvxh6rZKUJzx+SOB9myLfC+77W
+PTb0jtdVrJOvXi0hOz12449K/0oRKyWIOWIkSNcQnSM/W1rd7kXXqwOpFxYDcph
NPJ+WaxyBZTBb/wiv4g02qLXVelyNFWEioy7AKLdxtTYD6JbivWHPq5gZc41fcPH
IX2qJJrxCI0JIXzqjqwLwfpTkfJqhGbYmmMFI+CjGInle4oKULF42xF2O+ksSYOV
ZgPi08wg2SuvLs3+uCdlUr1m+juEZbtdaj3KDCvEnNCa+omb+ASqT+dkoCqswCuP
7GFjwF24Qyh4f5T9v2n6UyftZF1hC3fxlZpBZMk430au+QGI9DXMfk8a1wtj70cM
aGUXYzFk6nEWzptrDTr825C1vfFMe0cFTDEIIAXm5QCUN+v+O0V55lrILLsovA5P
eI3Eqd+bvpeMiICp3d98igBI2h9lcdGisG1c3rzEK4P5zO07JViS4u+SvnoHkG+m
CLxlP+aNFVFndfQwu6AzCSAWxz1QESndw9qEFobDFs8osRt5IysO1AwY67RoKCEd
TPT0svZrTt2gG2omdeSVzHFU3b1Kehx4tue0U+UgQT7t/XWLpUQ8cZt7Kz0KksPM
g3UnuG8YFg8wCjZTJ43/y9rI4x0GcYgBrVkndq0/j26HZ7mjgHqekv7Dic6koglI
ML4btYtIIsVfXQ64a5rfZLlqquHXogTfaS7tckbKDFEQN89brye04NxRfYNNH9oO
vPjuxG1ubqkRkpmTDFmllcoLAcxDBCrdcNz+0KZ3V0doDUe6R5R3rTOKKtjv6/RX
yEnBd49vi9oOa7H0Tc24GgIsTRxl+6Z2/CTqwjVoWN9QqigYLSSV9h0BeYG4y1MO
MoaiyPOjmNVCsFOr3HfBNslmCUl40s0qz/2dJq4e9+qzfBxUcROhZb8/f+WLAxM5
NShx0i3xXSQWIz46O7pNpEhV+HOcuPWMNdpmftbH6QA8kUdLgR7bEAJLRpErp5w/
3dHZZeKAx0bXaRxHXs1ZzZUKfUYWnH2fHQYyV6xjiXUwmJDn+BUcAQFF/FfxJWIJ
JWUMaIVCYEk3+nTfbNLYyeJoJXASqqms+l941nWqRMCyIwfuB9onNY72/9Se/hkX
x2584Kcw1zPmRFKpB/2ZEu+qTpA066xGHfZcY2nzxNPLDmwNPXNWQauuCLU1vYc+
9AsfDKZqiizcOdC6noI5ai+CBrR/9bDICDeeBSdfkoClEgsIscMSrCbz4T+bjXKp
ofSrjCm8k5mZpps6wX09FnQOsYZNyXVkJTBm/Hg8Qs1kewXQ9tqT1321GlYPneUN
MfQvEhdgbWzCIwK8Wt5nRsoku+UaAchf5l1MQJr2B3Hd1fe6aYIU7VfKjB9z4vcE
dWF5t3ttU5ffhwWPSLNU3yHw7mjNY+srgc84VImHF51unCpY6sbmZUl/hT3j3pLz
iS6MF8NcVLc4JEa8wkGOPZZx7ywKQ7AmLC+xxmq4LOZAe8fOcd6IUITblKeHoRcH
egckRBuyBaP3MMCLJ9VMmsYxDiE6rQF/ogrPyRGwPMI4Pbyabgp/qwet2M8c6zrp
xzbMcI30Y8Av2gCnXCdqn6PGuqwHMA0dnUO5o922CG7JNQS7RwCyThKW2ImJiKbb
9IB+zZDv+Q41vaCH285dwZjPK/WpyeURGg7bzgLTIKj52k6Kn72n47wqLItOy6lv
9k0YuUSk6It8wLnYkgSCKP/HS07aRr0YQXWi2Xkw695s41pVeXGm4Wq+BxbruQiK
cbekiTvUPUgZSBXpoPyu3huxnv8L5mGOJWJpNgtQJbz5NsjmtkSmT2+waPPUz3Zp
lzCv5hMqToF8r+KaoIvQ8cwCl/n3NQLAlW6qp0tvAPYZLDCXgiifAqRtkvG4slbd
Bf1LFeMZY57d6Eg/XCgjtlJT5Rb1xnFp7qmLbTdR6OuEXka2uWd9MQzFmlrAEsUW
HM0IZ6SotBI3wubmAeAqexU8YSXPHMEwEBZMD07V2ZmGAnbMsPpfv3ldVhDTm2vD
tTfdDEC8HrDIbnNDO8eLv9cicpAxIdjOz5Keo37oBUVquVYehFZgtAhmg+JDwHJN
egoeXKsVVcyukuKpGNvO9/SUDKkkNQVZZoBETm2NjDxNMM/c6g3I5CpxKpTPTZ1a
vG+MLqht8JTUyRnjBMX9n5hT6mTbxqG0g2X9gUfuYUT+DCJTz1cswSxfVlEzAKii
51WQG33CJ/sSv4dTkJ/PDq3oX4gr35O4EBJZo1tK7JL5gDEFpcHvx/vRu6lN0jw7
v2Yvcm/jJBazvyC+ELZUTchL+viZf9KN6+mq581lJ9U7/PTZQTCoS706pQTSstD8
y8x8b4T24oKwBMMvD+ZP9XVJOQawCrUKy1Zffd51wPQBMs8efzMjXyC6QObgRUpj
fCbOJ4pddx49B+HBKe/03VXgTBppfxKp6tBYu4jlKP4TGvp6C1F6bbWg5CwzBZ4Y
yhoLx5H90Qvg0iaf8+YFauVbipP0HC6lqtTQ41fMSEV+hGKU3XpK0wzVwlTDgrZg
X9OQiceKhzl6tXRWaXkdY0SlXSBzzMP7HzHApYt/y2xTF2F0rb/0IMDg5KBIJMl9
u8X1IIBUE8/+HNUEblmwi6yovbKFv44nvRfxz2EMNK7W8aE9jqK89hMrLAYnaaJJ
pf6mJa+FutXu8m7FdqSR9xLYHW/EFv2+Zubfipno9cenkdBf1Hc90U5v28zF9Xb2
kOauPdkrPZ94j7QPBD5HR2JwwKe1+mIrNQ9qzmWSJtStnyUub+9IEESWRbfLDbEt
aR30Z/vLnjBsH08nmNoHA+Munfd7/zXP+8NKvIfB/7ckTCP+YeTJRYjeKQptphXJ
MX0B0zzUcqiwVcL8EYb+xW4g4mZhgQEpUp6vPITWeiOFQa5caPLjeEaEPfILMCA4
IVacI3zXCwSqNGESuYB921sDtRqWFKAVJbhfLMMYDycN6EvTljdUsURlTm0dwmS/
jonndhozVtZ/FSarQzqUFJEFqnsiRGVe+uVxsJt0jcAAVMr7SPPBF7BZ1Q6SO7Jc
HwNFCgYBCUgifevYQmu6oRG56PCBJSRNmOmU4e+1My9iLHzDbrj9kEq8SYSjfQQJ
fxXpCgHyzV9BgmNc0CmyiBDNbq47fBcA8J+ymq0tB0hd6hmTtyJAftFtVDLRgwuC
yIWzS3fdvJqUL+4FfotBcP6WimRp/Y+GLyF1hc45/+9JRDS2qu/lfDzuDPpAg4Ox
nnowv84GowhyFJBJ+Gmg5QUsqnNePAMpMUvT+0G1DNgNBmmQtgZkwW+V18ZFUXku
ZJypp4/ygFknw4JMlv8v1hKZFNznbdWVMPU2ffjzXQTxDanhVKw+KuCBsexwCH5i
hapQ6bcADrWEpgebK5lWPbZdVmSCrFFxAS5hmj97P93Ag8P7Y+2uwjlSJyo3iXUI
3CrePSo0dJPF0c7oxRWcSsmxiqd8GYH7n/P6Lo6Ep9CoUDTq0H1EIp45XLrQnQ+I
tMG3zrVViGCRfJzusXOhALhXWrImg+HYUoOZaPlasRjvSvOxT4U/Fd/enmE54/Jp
fDFujL/mk8RMoq1rZDsAeThRW/SnfG2LqTpZx28mIAuGejXZT7MXnpt0HQYxW8L+
R4ycBC0hr9oNsOPKS5Or4s8BNCNIGmxIJh0zJBR7oRXp2llSbWQHp8C/97wLUxeX
SlEIOglj2mHQWUuuv/gTQesF/Q9M0CQ8MreDzn2DEcx5dUKoJJiV3Ts4/V1p7ctu
ldWU/l+rvJXOBndkmVNo+485wWpJ4yZwA14C4hXf6l2lV51Q36NXiI/FquZTT7+G
CTy/Q3WQlFuL6QQ/26nZUn1DAGYyosb90LzDuHm/kbs7citaVmgEwTJKHUJPdbLJ
Nh7Vh9mhZjOnvI986TsJySfmWWbvWYeMHcJrkplhdHTljJ/M+KlYCabXK+HdnMXd
sC9T43KdasNyw4uiDh0x6f7pJ1jkshMful9pZMC1+YdX78f2XzPHR0bihgUaw8ki
LPt5zj17JZ2BNI20l9OWApiFg9HhC/xvnvbKfaWcLKUaQKoutNuiEZ3OgD9lozmA
adcbaZXeLk6PKlVVEGjC1OyO1YKXhFV1rcDu5sWwxWmq28YgtdgkH+zRmeGIAiq0
yjf/+qYMSFOnWwyfuTFRCq1vzKRLaUOXHc7zkO8jMa1shk6RZ54mjjFJwwpKwVsN
nk0IJFrbqTcWg6mHMKVNfJ75n38Js/BL2AWCLl0wKMfejVHQ7QO6leOJVblaI+C6
Fw14xsIMfy+WrYem8fI+ekMRNEfthmqGA0gT2Y5wMHkKewzUAv3y8DLn9xG+H7Ck
ONqaelON9ocmqRiqBxqoy/b4hZQ64xnPE4+Nl1RcbbGfjz+aFvksintLpqp25N0F
Vl5GsUhgNCBinmAMRsMmy2xes1GO71ajYpoG09bjce4tn49aBvgPEll4mS0KvB1f
G9hl3d7IFKQ7YdWybvAlkvYH02AMAW+R2XlHQlgmfFKovC+jC4hkwoGUsslYX0yD
xltKuJgnlZadfwP5Q7LZZr9yvxArdHQFnR2u3WAxMi+jRICbbB8CfF6wrDoa7JG2
tOX4+y+X16BkyOsbOYjVFCzfTBILRWdE+jt9uelQvqKbEl+foRoTSW+FEy5IMsg1
1e9XXNDEMJuit3Cx6NcuFMmK2ljpR4C+PZ6sRDBPfwpNPB7lBj3wMnoyPCsjAfmf
zKxTtgjwIxbqpFo8YQ5NfiAdSe+zRibT9KnJaouZdY77S4V4Es/tyeeIvH7rTrSj
8gFeM0piuu7hOJxLftyib6egJGCXOe17GDmYIsUZpv4Y09YL6DaINUsRjSPgwPv8
rj5S7Wi4sq/vkyYO3m3dXb5KRWg+IWifNq7e5oPxZ9EmkC19vLW/I/Nf6q4ygiK0
IL7vR30qE2os821YjuS8LXYPqpmXbdqQ7lKRLxYsmRMauprD9/3xxH7gM+Yy5DVu
Qn9W1lf9xUkgwVO0yEVFNOY12qtSUVr46mgZuSAuu279mROEk3gqP27wp1ggGgtW
r/Gsi544F1n/zedEP0h/Uq4v+/teXkytnoENDJQQg84smyofmcx9MAv0fH337CSO
91cdrgcR/MVCkQ/4j5iLFvNO6o+E5csbQVqYwdS8rzBH88J4TWgVoefrStDCb5pF
GkylkyEBWnez5CWmUO/w5+iqfMHVpCTiwByCkbY045QTBCRmXp0ZxQiNH5PpZVfq
e7f3NhI/aG/5ygfn9JU2gmBy6X2U9pNBVvsER7xfgYVvndAGbafisqnjLsu3pMaW
nxdgSOQECgWJwftkNdAgJo+ZyuGl4ejXhW7I5BQ2QzhKsULSnmeJaCY/5n9en444
p15s3otBtDv3fGNqvcBGYOXFE3g/wj+e3V8gu8IX0OCcxL8iXKD7FTRQ1kWHFXFb
sVrMAAEYVm6K5UMHeJqp476GHFLCWKJfTZHIv7Dr5XXM8pESSUdF/0ifSbUzbDAG
e56A7KMimBkkShV6nTubX1VaAZvQ4u8KQY06wFa1Dyp+dgdoMp5Ye02xASRCr6/x
SP1NDjvs+m9twKH+l7fOrkAcXFkA87uzT5VrcIWxgh441ouQcpuOW/zp2y5yYfpQ
pXICLfhsG0bElQVIPAt5Xt+Bkoq4GenG/oz1oLOtUEJ7pf6CeZOfrrKW3eLf+JLY
/rBrszrxBVHd/pe74rH/Uv3iE1zQjjGCufvOh91s0M5CHYNMetVPfVetfW9uXtC6
1jHT/Wx6qwgiuwL3GPY2UALXv1rfHAsJJxeTkQWP7xVlXgxLU66XykekxKTEVlr3
GpuURlBZqh+dALFyB7GI7RZMzT91MFPHYtRCbcSrepNiLjujxPqQ4GoY4jDEL7pR
9HYALyi+LMci98H11mOsQMbm+JRYwnUG6+zTEKklo8UVlaXorn6cQ97WTwSr93mi
Lpgj5lu2ciX7vFVcxhAbRTsJoy/s1NzRF+PpwF8L1uL4N65NdtfL207oS1GFy2QX
uuQqSGuQG6r4g3wQZzVMzi4YEd+J1T99HXmleEoyr1e4AvRYgG13Nx1v+vbx0DT+
51SNONpRWeul4jRGeE5xEhAOIz49syig7zAmGXP1EzG8r+2nikjhONRl9OWLzes9
ec1aTjGHvxNYWUmmgWLGsqTbc1j8r7/LBaB5QN0NNtzV7kpRcHaaNcxkNa+WP03k
P2Oy20Wu5Akyd/AjLCQM/He/kX9w9JB9DQ7qjJDXAm4efoAT6M/IyWKXXVLDI44q
8kpryMw638lQ8fqUdjiWN9SIMWjkWlYfnxJPVoeMt0/2P7ldfdr9hi1E79Z4bKqr
Z6xumcfGDYUoIOj9m7YPAa+vytiiDA+o655qnuwiAF7FqIYEb397WCSYq5MHuAHC
rSTjeYeMPqIpE4arF5hkBrfFUuTyucbUpJS8UQ+rVwUl7JP0MLRajzKJTmNPngqa
1p+sFgthyDMCo1FupENJnRINgjx+4zx1XxLT7SXcirDB4tT+r1M1LEkc5eCs+hAw
Vjlx/33kS+HbhkvPImtlblFsp3jxjBbocem5pblfRwcOsEz2I3V1JeaeMrj6HcUB
i4aG+TWNlNUxNBQK6C6UMmZHo56iz5Rz4hNTm34ly+XkyWgptPz1OSwzTc+mFwEV
V+gjFBl2duUXeab9pK3t7vGMIDy11zKc3eTQwTETsyDEbAaVZTWbDX4S/lj9CC7R
r9d7MJnVrKcYSpIDSHOcR6kRA8kN/51FnlL2NMyq+MTK4Xrb+BYg45zAtwcfYltO
717eK86iVAg7Gp3dzrJD305zovcg3oDUHbmDPcG5u2gQplVxKE1X716vHUQ3+gEy
9gnCTkGt+rYo36UJSAUCUt0d/ROQV8ZCBDcDHzCpjWEwM7NpCkfNj4DV2nNVGxRe
NUBo7PF+Aro7jGqsg5GA/SoCIc+n+qcGIoDSq8VhV6xwzH9GfSLFTYu0ERWh/niR
qCrthhTgvskh3KpOQ97tql9MI7U95aUYxkTgqLWfKcyZidg4D/Z5msumXe6MCJYS
QdmeLaW76HuHbpAUMdBw0i67wjfYLx+kLdzQ6TNaWzqIX6BjSbQvxYh5kW2tMyeo
siINk4qINng0g3wCuVu/pcWT8Jk0Q+l5z/vwkXvfqvRGDlobCm9MAJ6TbAfh6Qwn
+PkSchDz+k9yKfirdzHo6Pi4b28VLkygZxLZ6G0Hi2b4GXpMNwTVmJSWsGN8ha//
RJT9PoizBqlqQU6JTccZDjFmr3v1oyg6qYRcdvpfg2CltMn0YnmEi9YRpI05PQpv
nsxQ15nz16vxKsrDwz7JzOB7DBi/pjpeZpDt6/Gl5Dj1m8UbNGGlGTMJrXMiQrNz
YJwvDjjCLOsAFAVqE1o3WeOalkReW1hNo+0k/VFIvDzqiGcyo56aUMhsCcAOsVSi
gOOhvui+MDr2cbbT+2gRA+6SfHjfBe9zju/Vd1K4unp01qVxcmaVubeu5baaHUs0
ZUi7C3Ts08YsZxJz/CAxp7e0RIIaWaZEK3pLWj1OFGFNeAnkai1eu2apTkgantrN
TFq3RG477bJ1FRvnOMC6n5SHke/cPAK5S+onuKHKOV6S7ZWADUi0sMwpTuj48PiG
rQm3TOFxn2rbCmOnbS79PtDkDlx9FPIkrY17qVhYLxtwQJtPsxdmnkpXKHV/kfxa
Nn1bsy60c4XJY34A5f12kIg7vTkdc4D2M+L1N8uTTHh6bMimt4h+Ii8DDQ9ODAh3
51IU10THl4v72zOwIvCwHGvbVuFxnbCjGReMvtRMP0PSPitguOFHEFL0jRT4fVdZ
iOEPrTTt33BgPAUjQhDSgc01mxEcTePx+rqTVLOSJj9lu4CMswh8v7Jvs0eSm6Fz
ZX1MF/jKOL2T68hR1Qu814HDqtRuCE+Df3Bdp7xU4TClOq8ivwfm2zIdGP1rgbPC
Jzo/+zwdn+rWvmkUGflZ2GdSVUJHX0edtV2k8okP8u6hyh9fnw91GI/lbf/QoSfK
k9Ryz9DEraokiV9b7IZBbd/p6BAffz/pTYgVauWUpyOFI18zEmnzfpOMTVOoKoOH
vNzWlSJKSt1ZwALnLKWDnlmBAvMSx7anXU5jC4rDvdwF5f1yhJWEUgx754ntX0QU
oyeXSr62Fl5HX31pqxnDMHmZHKb87QG1vtTPOKXYDSfOgEEd56iAUSex400eebPk
NsBmaR6Uqh1JszOrUwqzzNDtDCbl8t2Piu0KmAxUSMeqtD2qXYJHD0BxuDe+iRKx
wmNbpIgUqsBst34G+z8Dg6dWCNQ2o3wia+N8bH0JhxoTqcSLWecsjdqKFCbfcMaC
5Itqq0u3IA5VDTY1zb+LCWnHux/F0i2fp2fJ+6XZxEJ2ZO8D67nrv9WjYd2Ke0fb
tABxhRjMzTukDvmkpPB+x4iePYo0ykNoeoYHWcjwwizcu60msgHzluXw9YW0vdiv
i22Ox/jwlGPrbyZneeggKwOJeskouodLq3h/rPU2tNpIwYPT+c/WIvakUFEDGVQC
TWKdaEgfPL4oQdLIWRH3KXEIKL0SoLb0h6py4oDpY3WekJPzTMRiinEYgyr6ICDg
GHn9VxVHPSsNIAfnrHAgepkbGgAcjkXns3ivjtd0Geb3i3Vbwbdk9e/gt+TDitiK
WRS1YlUF8kvzFg8o3JoyxE3kX2GOkq0zyfVWN3B81eW5KFwEBur6HNnWBfp2hLYu
8Xs1v8t3HxI0CoyKaxrtdhX+sp+xJFFZRv5GEDZ9Z1F1vHV92MihWDf1baWWa5Br
K11fP55S84z2hMdIjjVkUMrGmvtspFsybVcRnwmhwggDUZWndWjBkbx9pmJPuNDN
8PfD/u2fpd70QehcFl6ZZb4dJha8rNfYX1ERfbu/EMh95m6UpW8pHeY96imKPaAl
qguw8eMXHHs+oUc6cjUGE3STNFlbECOJktGbU9ICcoK4panZywF8PiXAlQs9JwUC
GFGjoEXQryj3ke1lsN2zrDJ6pWJiVMa7KgDD6BHZ16fxZXY8zuYApA9xui4vfcud
DKt7s+B5rVhdwNssg91q9GlByty17ELIM379Vwad87qNUMggGX3fDx5Fl4Bf85Ob
sIbGWByKyQyFvUzxDlN6uJdUhrEccUSyBQU8g6K9Q3fkG6PUBkb+8vui+Z9ltH2Z
HDqC9fl1/nNFmaaq8tmwWNyl51j38pBql73dCA4Pq+UeGRc6fBnopELYzpqq5ZOn
CIAAQhXDP7lqQ3W7Raa34ZMs7T8L4BXxLetHTJrG+mk+oRwWWt9gTPuk/J/tsR+m
pXIBuLmEAnjWFdRsgvUoySMi5oK75FRY8SbsU+cMaGwhuKVEpsC9rFr7NxCDlQFn
zjmMxgEfDrt58cKRqoteyc1/BVBwb1/GBfdt1MzUzamNbyn9GClaFx4nSjPgKr6G
2wS+jUIrCCnSPCfPUr89trzgZTj/exedNqTC6q+95mP4xCqCOMlWfRCZQYn/vCQl
9ZZ5X4m72P1bCqMc3ZLlw8QSbPnKjdSXuxYD+lZUepnoCHsNwNcyNDcwPcQrnvQG
fQtQzEMFAtyoMQ3z/woz0HAEnCkAz0wuMYHyswXQpB4RZVvSKNpOTBehetet+Nci
fDEk2/lK1P04ucGu33zANnDMu+J9LpsVexzgC4K/1OvXDOxLi2S9vgPKMqRChtdD
3ONhJmhdKjUTfxXpnKXIUgohOVP5PVb9jmSGh8z6kaquFaEncdmSkY0nyipfF52e
TJ/WX9vy1t7744uXzxkXzNALKmVISDSCP8XuggsiNgwgLmei84mOr3xxTKWTJVzp
xGCIoJ954iYzbHHmG81BPn3kgBG/3Fdn6iSRg0+snXg8vRdA/TFY6Qd7YLkaCLXf
vBgny1pP9RmIM1q8UpLzuokJ28CsmVc0InBlbOchRugEcmet9Iv4E7w7VA52qkvP
MHXhPeMIoFghkeY1/tGLUEHXC5h5v+t7tIX+0BAJAseHsD7sMJtxtFBu2azFRrlO
KiaIoG5QTO4AaxLWd13FaSiHcKduQ13aqJJps56gHWN93EVMkg6rXKDnldP6kjMP
EWvJlAugeYpIm7ac4zz6Kll8w4WDsXLCtfLwOvR/uHuB5rC/rxO7yiqqo1Z8NMbg
yM0WXjt94fhlspFbpzpeZswf01DOBJbvBsoZphthx+BNL8ncCA3ouvbqArmN/4X/
1cvZORLdZ12cgjiNifSUZtp6sT/pLCx+/beo1IMC3H/lH6Xy0sSEKdHB5Djm0U+x
2xgcyj2u8ftVRkpWtuZSrHvDRQRUg9s7vyvcYy4zXjr4JysywuWzFJqjZkldbMa+
2uGbaipwfTe44VuLYOfrI6PQtibYj2eJzuep1RtO/64L2lMXlrLc0G0LuVGunebg
lbThhjxnif6ZMZ3KIa0f0MlNUYTM/CQnnUEBSC6oTvnBPlw0OPqSFE2bJyvfdf5F
i5utN9ZHiOh87I8wNFKFZ+NA3nCNDzexvMDXtCyZT5/2Opiw5cMcMqCvg0u6S884
hs6IKjvyPPBWiL9ZJRqhF7bfYwcjtDr2QIG+dS4Khwf51rf+jJvaoYKt2IZaFAQj
dxDDutcTZIMohpmvLCe3mmtd3ONIOzp645P3Eh74MGdDWYT+445LF2IGIjvgMqJY
en0E72AWt0NYSoddnbx+CnOr2agWfrjbSGHL/1+dWiAYcuF4bRk5SJ/tz6vRZwfh
CSbMMKEfixUrhfmH97PVT6g/NTUeh1hc7MCSYZsiW+myVWbK1kkwEPJHeWCZFcrJ
bk0r2Nv6PDmuufkAo2HaoL/VGQzQNmPpDDzh8+ELa49Y/Mu9cpkrIttruuhu/z41
HAdBOnFAC2jrEgZOo42pI2EIbjR5bDZ4lcVvRdhnLOkaUFWtKSc8y8ClON8nOyAs
xUakupFIaLOKA2H0sjb072NSvBV5jDxpuR89LLWbrts+nkdYKkQMmAzcAx6GuOQG
OgMU83wrKpsuP8LnpKQ0ywvpvEkD76KW5LzGGchexdjfI19yXNP++S/Mrha3i1lw
wyQyVCi0EhZ6cOTIfsFkHHlSIk7RGHkU0terufRPnx8z278pm5NGGKreJ7QeaRRx
9yVq6p+253h7cOAgvcioDhZ7HCY3vhUN91FMSrKSkEMRpmM50eLoL0oujS+uNw0U
O2C2/rzjx0iLwTG8a5ODzUDFErXwJweaNgGf7r4nQnP90TAjE9DYmXEk1jhfBWIm
lP+q0fBKN7PHjXgnSi9f1gK5Hc5zxVsIIHjIWOjMbl8xMURq55CQ2oL0ZOPCsYfr
Aq43EFS54/3+TFGAEdl1+5rhUVlOKZtXPK5LX3/EGNePdtP4YZdWQrdbuD43EpMp
w8yu70fhHxJcCEZ7HJHfRuqQHKwbGXu4a3/vfzbSKATUE/4ZB6OQUR8xxHBucGCc
tY8/WfO8DscNivDiJoTu0cshMG5bTmnsj1011k2c0gfSlJcGIQehrQnKRr3dutQY
ADfULLshinkzmHhnrI0z2TO1i/qrfww/m9TpIfi/3blP1XVWB5/iSbgyd98eJGkN
O03S79/aRg6x1koHgZOEvXce5THSC7qmXxSrzs1dazhir00dQwwv1SQ0gRkNuAdl
1rEfy0fmtVQZpfKGTtZ2w8G81jMrrl9TV+HufRpuNhLaO+B6PidJxMqP7qUW+tmm
XPrtZUJNlImx32yYq0Xek0BaMg9uZwQ90qdoyDLYRoVpN0UOCynBg0z9tK5jcG/p
saOs4Zp71/t9Wzk0GKuo8sz/m9TRkbXIX/cUOWJRXbas2riu5/n87GzRoT8DoUdl
KJEAEpUKNnPCjtCRrnufMozjt+AMm+bkKERVwqAcHxyYKDiGjzfQ+SfHXMgkZ6hF
P/yOyU/DhVu6vJIftRAcoa/klFJA9kFpclmuA2YliRtsQIK/pATfN2JkA5wEboLq
glQBp7899S+xhvcNlJeXPiqtsbdRjyXVmkOAjnM/x7xaSWGpQYo4av/9t5h4q+xo
EwsJgaNkWWNrZdbh+Lc0RTJnWaqE5HyyYaHNd/90KFZqk2XSyXHfVlCPuWp1ZGYY
msVBXKtpDv0DgMqKAFbqFjA/dn5ltyFTeOMP8sKI3c2LOJHcpR/8Dia/Fg9ZYUNH
obN2o24kvVz4efoZVpAgYYP1OdrKL2U0k8Q5KFuKtbzThMxqPtAemLfbq61JO7xH
jp0FjztzjhjeFgIvRP0sXYfVHitxG76CbHmUkGpJRuqZFDlsXDulZrdQcTZ0tkUR
u4Y9x2u4oRNjMQvTduuZ85Z0q9XLPFcirUBu+ibkKQm3FF5bp4H9vOsybtG0tngR
oLhzFdOT/TDThRGMag9sh0QpzXCTT+H5j4xqcp906ejcDbBp+C5hCgMy9wjnjJlg
hJ4te6klxXWkBt3gQ6ezCquzM3IHyQkh+z/l3mIKSMHboMWMH/2vqNT8b4REuAHV
3se2bnq2pcwqCTWDqKVJJNoTi1fOP8U9qDd3/BrabWGHvW6TUAr8Egw1mG9eSEum
ehl3QK2at/h9RcBhnrHMnMH9iS5KomgTx3qDROIFJPAcgJJHExmM1axIIvKWPbzz
Mw4CnUEWJ8BPPQjgjuT1McO0VgFsNp55SDwMZjyRvvs1Q7RmLRbkb0ZaLYghf6WS
wlHFN3mJot+4mY5QjeLFDrxzjq5FuIzf4TD7pn5qqGG8tWkgd/mI4/XWmM2IUs+C
dV6Gu/AASDHVn5oAYMm5oUrPXWcnejEe8pdf4+WV2iMXXtxU86A9TGhjCltRSD+s
MBxpSRPqjxq//NYta2ridmPv/UMLYym3Hd+qCMuNZkz+GIwrGXNz55444OtSodHX
ZIAAsI8iCwtdsnSvaxsef5Krr7UJvqsS00CFulAMUDfjcmPO0462WYaif9D2MUOM
asU18Wo3N38nCq7HKi7f1Kap7TBwFGPYG0+pVcQ6lNlW23sXmXxYfevwhihaVmGl
hqhpJss3nbdETB5ld0+QUy4+nHHNE+fvPs+ReMn8EmJqSMY9s5nOQc1Cmx4m9Ttl
fgKn2oevMsXACvyp0xRjiS0d5ACqznUCnaMvD+jg3fddCaI8yGtel3WbbSY7pBvO
N+xP35UGU5ACm6FOCe3S2Janyra7Zye9JpCxcKuOLw95x/7T+ISDaqxX0Klgj6kG
uJ1YC5YKxvHL4baW9lXMZDbZDjXw736h0jO1RgRJ21kRW06pqxdd5Rf7rr1CMePx
9aiQ6cVWUQyf9fc1ewKpzm6IZQhaXKgyWJ8dYgH97mjdFxU4xtRJNQbElKrl7py+
ky5LswbPvQ3NhjNRjox9l+NOERatKpEucbfbD2eb8XxkaBjpcaj3z4uPCk7OQjdG
LKJrHjmCWDO+jrJEeDyni3XjAoFIPhnPFGD4nu6IdVov/y88wOgjZZrzC9gfncLa
T0UDd2wgt3rDMapimez/wbhL+iXrljKdh0Yp2APKAoUEPcgXqO04qgJ9PcoNudo6
KQrv9NT7+Tj4fmCF64TMyQbx1BhEhhvR8Et/rQAjX+KedoFuV0JQw27pruyhayGi
CFX2tJhcK+hLzM5c5BdzFrbahw/hTHeHmpygLQTS57zf80ztBbramYRBnDZer63/
q/LToT3HdA0cm7NY0fuEENAmatzuOn+H0uPmHxO5OV5Kg+urQDCFkY1fDl5Km5HG
+TVGiB03pBKMsL4X6mdw/6gDdJShUMCACvALiUZGbGsaA4OWUwMocte8piVhqCTb
psRceSX5xNmMP2wH2NTaDj6KVeqkDrTYrprPs6MbtlVDdOVQgaMwD8nM83YDfH+N
Tr+8ilW4INPut628vj5eYgjY/uLXyHrFHtj+mGY1BUHse1+PLKMuC9yEwZOcOpBB
IpuV93JPRAKajmhA5LaFfLmD5DGsVDdbOb/jtKda4k95IwRaXZ5TWUHNd589R3dT
s8DVzLDXFfBrzoVHycdvUGOpcPybRU+rN5cWHr44j9sVzmySCD6TsRhm4ZQx4MI2
4+fvbm3l9heuhb1Sr0tB+tbCn7n6BOAjnLr5MNZEjeK0TGlU92OeE2zPvWiDVBQV
CzVo/l+psLoRf/YypK7XdYJIe36nwwUpHKvYJH2ourjSc2+ykg84U0g14XpVVYMK
G7YwgZ8tmpGwBMz1igiBtnEV0rhLzn+ZN8IC5PmVfFnTgQbIa9czi2tCGUrYUQiQ
+E3+gf1p321P7bGD0UwqbWmuZOppLt4oRN2zsNd3EHnxLbxtXP9SFwOK1GB4CG0e
27wJrg5njzWk8jNGz76Us6nvguO+tPk7gBSs+ocr2TaXeFVJRj8O2S62++NQ6ngX
gyganvW5kWMv9EABgJ0maxPmmWoW4cNJq9l7Mnf6cuDQoafpszIhW6dMJbAU8aPB
wi/woTC8quS5yUwTn8rhlNw087JvVBkeKXGV5hB7L+Vn/1qsoYN3ca3BdgI4KgwI
Fc2GbZ7VDuA76IWx8y85LweQaTYk9mDm8nJ8tbv3TLJCQONsVCPEHIHepurjJFVd
D8c20b8B+ia8mpaCw6oTHvOsL/W7y6WhuOlsz8wxVGGLJwsbE/AZtPNb2zRs1+Di
RFewW8CULJ9pdlJ6Cs+0p3r9+Lz1vbUwGqL7Ri0GtvN1irCfTDCTM5/MknRo34la
KA19thJKy7hhOyloDtFVxk3R2cy5k88hKZuyQih9jec39wIsAux11RHCv28OsmC3
XN+Z/3Pu0AEy+k9mf07FgGFNDxr53/91wY1lQzGdXo4vyIJk+d3cI/3WJxiy7bvC
bTN8gFzKpuJna2drPSqxe/AXTW/Oi8NDbOG3cz8LWkxGpKFSlGKQAONxXlgGe5/X
qBLTuwagTwIBsmwot+x8/uBr05jqS+YwRaFovKE7x+jDiM5TcquQc9DwEzqzPxZ5
9bCJ65rbJ6Txfu1+DRkPqbD8Hm+FPsTVz2gQsaHvUSMX6pOBSPHDb2YPSZ5AaLyc
b+Rf7uyjSQ4KtDaruyW0iT/rgxp65ezzSfzJrfjEnIvwSS/YnqzXQswW6AQw/Iel
fqeF1PRKtA+79uQmQVGg4f8w/TjKcFJA1V4ZdK11gf3IjdbQWJrKP9RxP+X2UY1r
/8hHE4ebeXcYji7hviykgEFq1b5dhEbfvMSgkPcnGa3dCbHhlNh5exc/oj0U0nuQ
x6A+EC00XESQ9KbHcDJBddkka/qtuW859CvKzNJFu0za4B4V124byQ/ZiT/5qSg9
Lqvq54ArBw/9w2ycj+IkIM4rDD2xiMWinJ0a06t5hFo/xJMGPtXg8twTqEDW/h+r
XO0tgeS5UPk5yHTebUxD9j+f4JcIZxN70NlO0kcmrY5gcWA2K8cNG3t8byPWhAz8
1Ma5fdU13byV2hreIfhvnJfRIZ4/Eli05isMxx4rinFTE7DIRM8Go83wDbZe0wbe
MX21Gp//4dR5pr102BujUI4zR20schMWfGo3wW6OAzTLHUzl+t9toJBwe1/+dvnZ
1xcoE7HvxjCwOiZrqEvqE90F2CODkI9oVae4QTaPiVlqqHtuT2zTJuyl4opjRs0G
AQ37nqcUwaPs4ZUUnmcXbuUWWqkEN/+pwYCgLtJGolNqn1TE7dQbwa8Gp6S/bvV8
lobZHbmZTk5ux7q//SZB7Sob8vPsXZGB9wJQDhJDpXLyWeE9dAvxuDrCirjj8b8k
yEeER3uh4CPNdOVL8gv889sj1UWKLrYVwvlwBQd83EaK2uEKd02JnMcirT6gOaWL
MVWVX9t2/HWVJQQ5M+fPJ+L3EZNkQRSlTmtAE+22nLwDYjeVnFnIQyPimuEj8+ia
iXggqviOJzJRjnydBQHq8duBJpBfSEXIcdRQXR1pL9Eu7JMirkVxuoidwH0q7H7v
MN30FwfuuRVw3q+wnBRyI7e0lKaEWjgH8BD8r9XBfdMHJsNzwTjOgXeJmyKgI3B2
t43dPWiAmGZ+wG2xx5tXQDNJfaH4mldA1YYxIDiFTy8pX6yjCLmjqOhnwM+GR1Y0
WSD7ZLmVpgBvtmL/88uAp5YKWUwaIB+zjsAFP/C5mmk1vooXnftdgbwQUl/H52l3
4pJybV2WyH0fqZ6rJY4S5LbCBF0nPzfX668gDooGju0NmbzJWx+qIJAGrrGErIbI
IeY0nOjzoB5vNfKD+1kS2wBT3Zsg5qTm1Aw7Ls0TIDq/C6Vo2j+yZvE8EZAWwex1
ujccRSEv9U/eAj/6dT2layr/zQRUEBWwLiIPyNmmxOj2CKLxljmhojNPPP+qDwiH
UGmKdr0O8Gd/solhAKrjRkLbNnzV+DYHG8WEV2J3nScMGeRS0RvCFg2yV0sXLg0+
3P2YaZ5IIVu9gxKMTULH1mjZD5SMQ5mpXOAPIn67vhivaeWZnTG5Z5DSvqvp5t1H
rtpmRlmyqsLfLKqMiY0dU7/Zg6BXaA20QtnIVCRxQ7s+DWVt9QQGWEM0lRDWvdYA
4BCrM7ETVQiWhcaRvPeKwVgIW8txbWSlAg+u7SE30zmzffyfM01TXlolK0DW/wNu
zPNxmbKS6PD4hUMa/GcwuQjx0qXuM6EJ530DF7uip0M9OI7fN6psg0bOfM+Vcyu/
TSnck4uKAM4X3ijxtL5LFd5JacCjM8y+6lJ2bb68Qw53DjokZ/DrAYP2hDZlAGuw
eTcKFce2gFWAMOhnqglJa6K0xp060NLoLxVA8gnFyTo39pKrSsza6Z7lnxVkOXYR
NJIhDly82iREmcZ8ASNq5mnwzI48wF3j4esHPhTNndOtZ9tokajVg90R0OIpg4sS
tJfL+FnZ41cg6/8pDKjddGKplvNhwDo3ftZX5J2Z54MTcNuUmccjzwgKgMa6ZLbS
VdoVOodq3e1asRpS/jRgpRIKOi26ZltRydUuzMuPwsB8PZem4f8HOp4KYxtGRCrZ
ltDMT6RxO1Wx6m+oEAPQZmE0truTyCHlkKpiV93S+PC95vGs5b/vhuK1gu1A3Go2
KGXwbiTgSOoGW0Ju8BxCCZ6HHNd37eTZyXXEeGl6qFaRtrJUiux/kLFl6GZ1sGUv
+/TqV14mnzA5H63S/sJ1cxTqtuKKPkn+cMHo6J7meU6ir0jag8eXKEx3bXtyhwpB
jE4uhfDVAtUdrJl/RjpSiUKXJCHygNaSOZgFIvIEf68bI3c+bKmeIGS+RthRIRlJ
ehdX1ZO8Ci/wLpqSz4kfPXSWcX5M9R7jfhbP+KolDZ/gKOgGox/H9P6hA0xia4il
KbFNgLxy28Q7Vr4mz4zUD4o1vdOz2wRTzLm35iz7Z5XStyIS1Zl7sW1hUAEv3Hjz
VCHXqScEeM7YSuAzu6iBI2kVt/+K0OtH+yICoH/S6lf21C4svgH6LyeJcM3vBxtR
cKdN7owmoEaSY+pNHNS50yHspItqZPTUFe6/f1VQNoijuKtva1k3NY0KB0rPfDtG
5ROhEklnNT6VHIzAjOJiq1CFOEmmm1ive5Sz3oHcNjAc91XaM3aSFVV3xl6w4Z6J
qo4PgMHQJDf48gp3G4jEGBbCUGY0stDgdhd0N8lKLF2ftDXSl2YdN4sm2XQ9BGjf
nx8JKbfDpWs5E8Z6qr0wf9oXasKB4U/tIEwfG13GYCLs3p9KWov1VysQ4//tYPKt
4u4Qq6LKNPdXb70vX8fHAV7RnfAXUHSMsJSn+9diZ+2mXi8JRmMpawmzKRMbYMOG
V35claWhgB8MmbKn7u8VW2J2ABP+z80HCPfX2zXGF0hjkPj7XpCWFSgYZpnrLqQw
7BPGTsGezGv6w/CIJp9tQ/xi5JS7tALsK+DDQ0WtQF7R2rURP6I+sNDvyAg2uAL1
Hlu0tlwyePozU+DW0UOQwuPFd+XTiwaxpZcWFNqiDpoJKtjOLMCSV0ETiG+egdMh
fcdthnvUfm8O7275O6zvLnuWOZ9x+S2lSO87TPaTgdwkrC1EouJLiQwL33v0LJCp
zbLIhogj2Ygg67BCJLgWq71ysE2C0POO68KzgvbqFYUIJWQarodJYasCeh1vbytk
Kf4AM2P05jsn4NKhqis5yRTq8+IuL+iZAQKQ8oSiIIBiIVtZGIolxr8RS1pxFhHN
NpB6zh3D7KDfcED32peQeRBVorRwSTkC+a5SUmV+ydlxUyacQFb2L+rgU4X11xjX
zy7j1tvJLIzXqpyyshIbdwDWcIAHYcok7Vvdab1Uj59qFDoHuKgxFwPYItnA/iGi
GNV5dsJ3GTcKuK4Qyyymh5guUTYAB1kQyLLGrJGJrIcefjjedLjd7qHOWsuMEH1p
Q8Vcmgl5vQkwsB1QswMylOHDClIR2PTrhuAgWCCuOu0/y4UD/nUuSb8EYsrJ6TuL
AdgS8ZYWYLL66AmkqwYSdKITwMe4yVaZlOpqkNDGsfE9uZX5BoM97D4PuOQ+lfRU
+gd/wGwvTTQfkJf8GBiH2i+7VlwrfM1njFoOpzI+IVQiYOsb8lFnBCcGgffE444s
bgKb4jCX9XnDww9buAVQ0O6gx5cRd8H5A5j/kVZWwLNeKwtPbwVXtgVGcsDyzkeY
Hy73KFWjPi36o3Y9M64SKzikhQ3uZon7ftuy/Hz4OFO3DTCQDuUZ011cgrZfLWkC
aFn+vQ8dCrJDiGgVdXUwjzG/vZTbDKePb/hKFmEOYe7soN6V5nBZViU1DCf56bBM
9ETwz3XiXeXbtVFA0RAerUlDqojacynZKEUpYTZ0O0OVprs/Bku3RYcCWc6eaXiq
779/pelhsSjL1Rhr2mKHp3VvLVJcNkLe6ymWmK9IQzunFLQ2KqWuKJC0UA1CWDXG
T4mPe/x6PlNl0ZlkKbbG+LrNv4e+c7owVPWPtSUYh63Zdv5RxjW/2CylkoOOOvRt
OaUbHGOi75hfIOX24SPNK/XrDteyWAeTebuVT/bHhA1tJcmQjiYViLuC1y0sXpDX
ox1eXwdj2qoIJ5/n7HNrhD5Nl/x34gJ9KePOTpHSoPu4KZcF0b9m5ek+BbIRfcLK
NNIiFIEi17Kp/OrlZgHUaIFl/ojBuSj+AkYOp1BXv2pLpXusJNVdAvzfsCG6vJ/T
RrEbX5LtCnXMUyd02zQQ3nPJYL/sJcAVjLXRG0MtFIr2FUVmevrUKNCc1xJTIKp7
oV916ddh5Qzuh4xZ4K6TR/NKMsPXz5TVy8EsbaACMTciQtiz5W2IqnsZfr/b42tJ
CFlLobTI01B7niTaYPZbI77Ub4qvFeChledo105/RB6ltTMueeiGJpYvI4zRpbNM
G/Wsru0IeTDXygcVEiofRHpOBejNcVyLQ0kbdBL9MxzhmkIaMSZi2vVOovWLkcr7
oLaztgx4CA+YiEXy+rAbqkhaj9y77CFdylHZ6RZj8Fe88D6NSbu4nugcUhfMxwzk
RH4kAtFbU+LVWgrvmwE3t2wIMVK8uQN6D0jyyupu7HBfXcTlcmc2715KMDCcPdVV
h7v37vsjg7/h8bcXAQI9vSmMk+werNRxcCdOC1HY94paUOwUc1q6RoZZZulIj9cj
3aqlT0Qg/f9VlkO8oTyFpg2uxcxqFB69PqdSkC5zAbQyCAjYixQD3wEb4+ee+81w
EbkcQcnAkxUSVoeMQR6jrcWVtP0zrZzFMr5CXXIwjJJhHXSEOEMrnbByrsxGnn7g
NR0ro6F94Dhu0bz3tdBGJnqSs7d6noA9fFiG+OyBfmyAd3KwPsx2prT5ENbPGwhC
b6eh46wSoGzGNMXCBhzX7opTNHoyhf/Ze/He0iaBwDJiLwaMWPwEm/1y2ZAV3GNz
96qfXzPtppybmYhsWl3Hv5t0IPj0pftmCrXY2bq94h3fRbcLLrvTPhF2ZsrDauNB
ZroiSoZbRXJpsmBLltzDH+xRZQovcqLxIhykp1YDO/1AZmcpCe8IEss7pLKwhhzP
t8KpenJxItbHiMqpPu2q/r3XgCq3H89O8eZpPdeDVVHVEf3l+CRN8jQJY+tGZmk/
4yNig82/Ul2BJetf2JsFmMYhGrizBxkYuCa9xszk+mydxAO8MbVL3/wqTUcTUr/r
ofNaKdadlcNCTmgMQyA7Gm7wec7CfBvN5+UEbirywq6RgeCWiFkeWKYyIxlfchEp
XCoiVfnrGWM2J1v3+5fDEgkTFz9H+l0R/pGqa3H4cUy7VYZX7i3hWX3NvaCRSc8o
Bqtf16FdmINsJVw4PdMHngsgL/WEWLkal24MZZGTchg32bBIi6iOS7R3v3seGoyD
sV2tBLmKc7DxXDw0YFde2pRB8xGzjOEeSZ7rGeZgCbM7PjPXQo3xf6enOEnLPz7X
C+gbZfHik9mwpyGekl9y8FHAZllKjbYnQhCK+UMBMuhUQrYF6a9cDEYzBe7bNolm
j2FLZKZLbwt/YxwIkBs9P46W0Gj+BaLG1yLdl8QnnUYg0PgG1a5RQgLETBpvjeGO
v9uXpcOCZSToT9DJH75BNshOFPZYcyVRaNTq87iXIo4d3yPg4xfWw1sKOl8w7aQI
EI6h+gAihoK5W4Otxf9sV1ZProuRg30ZF8bJBbZjuvz9q8a7e2i0Iqmb60YDpbwD
8xW6iNJbi3WubnWhrUkzaElRH07nIKJ8UPjP0Z+eOi2hwcdzZ7zyfjxlksz0cJa5
YrVbIWb2nd3hzioaZZdY8pHD4ufAozE4e4r3nQ4sVgPbALiPrIIi1dZpsrS1jNmb
Rqu+N3liVAnAenipYbL1Cs72nDR1HxXMsF06KyBCEjfXcTgKNr2Jbw7wC9OkvmQL
tCUYyQP4JiGAzo+5KNpAJQN5+pVVLsnOJRziTPG9YlGtC6tRTk6fJUdQLAOmU1ne
qkCcO+Oonjk8V/YkoFpzr5FfVDmP76ik081V+uhP09Y9bkGFgkVMrzJ71uZbcyAn
ZzfuMlcIfAleDGgHlzXvXJ/X7t1Z8la8UfFfZr71znHd1j3aweoaAwrAM6F61oUP
yh1u0ZPJ/LphLCzc+FWxRoL4pWKjHPSQpxrAvaml8RWCosWcUrVO6MiwlmHYsIEE
ugiAxKmUfeGFW5Tww729RxmC3k0KR5f+4bFTRvyfgW7YqR4DimROgHBw/fnVIKSx
rGoOVILwXQ5cfj4GL9lIFZrq/2kOvqWkGhXUcHYTVI87YQBYydxwyX+4vi+FMROC
iH4c0a5mo0u0QN+t4z4iHdNlvYVruBBWzRFBBA0gpgccfUj831pqjdFid9EGtZwt
uZa9P9MKojr4xu2eS9LCthoJRxFbHQmZ+/Y7NQ1tguiJxVQhXbQQtqs3P5Z8OIvH
1Qrb2oXa3arsxu/8chPKtVcCpt10pigSRETAUY4v6bphgONvwI5MGqyKwGRb05vf
lDAyEpaAMASnZAiNpvFrCV0Vv0HrSLhy8tW+uW8r91G/6BYhCyJxh6cMAfB0QI7W
gLD6UgaWafhF76pVhnSACimKEaoXvb3f2e7P8vzinSK+vEhIINy3ZokyRkGkdSgI
Iw8SNFSs4Qp0QSj3+Z3PxkPAb1Dz/iXxu/c2LXsROQ4rAkEjXlczkb3HCRVv0t+e
cQKy4eutK1AoLtq+Lw6bjrL15fMFo5OYz24gqKdT0UQuvqaz63TWeOrR7+lq7lnp
eqd1NFsMs6jRJN5syrJ3JnmBbUf5ld9C74a16RXrkqpD/WTo7/nyp/JS3xqEpjOw
ChyRL7+nab6diYWNM5kEkr7Ecz+qQX4Ps25W6mTV5lQXyouzmnWklOXboRvvHWUY
dQRTV8C5ZY8POEQLzyamrnnZuOl1uy7bliYjIjmP1H/Raf+rk5kgyoVM2dAZfwnu
WbHjWPeJ6mV3QYdL2KOU0ySP5jp8IRqqX8gbPYOhMUT5CsFyDaDkbk+eHxixzGOA
ZaoNbBzMdFUexwHigeD/WVn/Q64d9l7cQ+QtVPhL96CBubPvs8HjhDQvzlql83H5
ubDBCGw4nLwObIUr0v22Ce/OTZBRsM7Cj3UINlmyraTo/799VDKnGXfDdIYCqYG8
XzTHBk9ZjQFpcGYAtenMw/FSy5gTA9m2kqQtGBFWjpBRrCn5EK0ICEeCJm3J1A+d
Ylh/H87GnpMX5Trmx6kHyqBvkam5+r6DEjMtiLn1CoFC8EH7//OmUUsH8xk8KiM8
867YiLuVl5spEqp34yqkQk+1wJtQv3Jdd3iocZCu0RTrJEcYiK7hSDBYDxWpEqC2
ikTMLgYjLB7TJ5P5v3J775r0fnWdH/EpmTYjbsrg6YurZwidqe7NWHY/8QW13eys
r7wCXof8ojiOuOzwLPqaB0hsZvEiBlcZl174K+x9MuL7ihWL6V0ANTUmoM4wMFer
FboIgAqqxI78qm7LUhIK+C9BPYLXeYbvsPWS2dFS1VJbzcFD3Z4y4ynBtD/SXNwY
i3Dlb56ECwy7AN4NTUAcFBfl5mmirf907znqx5hiijD4CvVghBs169imOyvaTjo3
TCg8tU0ZynH4KbVlO2u3yJuTiR9FPUfhMkrVy1mqp4xWcw4Noks3SwWID8SNYLC8
Zu1EPwjjMgsZx9PITix8FUSvrKtKapNYUqNLMUJ4tjBstjSrGAln56iwApTOEUYL
EjNMRiE/hRq03DKiIh9UFBYZRw6FuSNpH9mymkDWzMqokKB8fWoDL3W6ATx8x9EM
YWni4tJdfQ5DkQnZJVTDqFuB2ZAlMiWcr+e5qlkdshzTB3JLGY7y4+dST0p9cwDi
WortSieE4CA26fnCjwlIXNf++Uyw6L2gKYvXptbQj9MUo1OT3NthFtRQgzxgdy8/
VHaQl7/HIdjY5lDByWXtE/vX6T0pkW9sglJ2G2pRQF0f8Ti84TNAbjBMtM5QQ0UN
TrnCXEhE4IIn85cTSP1nYX42PC4iqQJwXGuAAni6j7MHKV3GZQZeESDpPpPCSxZI
4Sey34yqt/tjpL4wa9nXI6gznqCPtwZkiV8K/ua8tf0+o+UI5kU/A3f7ukRobn/x
SopsM90WvAo73Pi+jO8NWEK+h7hA/RVtgfbOYeWhRhEkUYNcK+b9WoyMV6Js/AMq
tWnQ3aq6IfM4iB7YW+S5/d5h+ZO9GhYjf/RhjrUhlOO6o/zDgY3kshxUj59OfHya
MrvrcW04fdQNyuVJ2/b6URxgqctOIFcHblhqCZpb1iMk5WFq7Th3B/erkIFPJjtp
hdljt4G/PG2kuOYOy1lFHGattaGXHISLcLgyTQ80R0sjNyItH0XxOik/EYIqXr2+
Af4AU+1t6dY1fOUcssUrZGRAmwzWJirnzAwCbMGZSgwejkI+FhZttjApzUSihIqp
u8z1dDBFjGqYEhifbDTquYNDjfOSadCI+Ut4vn+MvySUIQZ+gQUgHAGKGIxdriVe
cjRlFQSgYA5Sp/3R3Fa1x78GOvQcbyi8uJ7RuhzkdregR42ZNUrfhs/M7yUuYwKH
rqAg072og7x8XeR+TWge8CTPi70/Gu247eynZa9JNQEPglFYtmbvUFwUuC7cN6eU
LtJk/FjuxgUzKzqUJ0R5UDI49qgaeSmgMHRTVwmIxNKvfdnrNEquc9h2duR8xMqx
+phuhy+ttWGhxl2ZahuDNsRyHY8ZnqR1rEnYWUoNUFr2UlVpYRqyEZOmYDRaAz+R
o21Wmi9NzJnpLUCF0tTSXtJ07lqMUTPzsIs9gCXxxTD+LRTF2IKLSFRMphJVt48k
O4kQWnjcqFNvUNAWb/IG9XWivCPTMXeqrsxrSN+oBI4r32MdCaWZzYyolDzsjoPk
nkPV8UA2PYuffb7EGUjsSzdjyjXo66cTBx97yX7qY0bgzqwu1vRa39NaDvThsLJK
78xmxbeYq9wkKc9a96pVy9bhlsqKthW0AIX5U0oucOx9TSAQHVb4zo7c8QKUcICs
rOqdFotjWMsZtch3rH1dvJEUTc1mve8WTxAbfyk9r/N7YpjxEGJ/F7aIaiYbtft0
SjktTKXPAKgdGGNi/3kko8yCb1Ny/oK6QpkxGuh98lg4SvRAQTs2AvobI7qcb1Gj
eGIdXDNU/J0kJ0HjhCIxmUi6vxnFf95XULBb7cBkWL9OzcviOnG7YksCus7jEuI9
gkZFyiLGoI1ylYbAIwffX6InzX7B5ASC8qgykaahQauD7aIr47t/nSlxziJIm2Pb
OdD+HhvRDnhUBvRPSiHHIZv5z/6VSce3oGVCB9HsebFZ3Odttn5/jUI/aS6Te7RY
u1UBQwuShMsc6bp9VEW9vntZlp7g3/QnqJoUspNVHVLn/xN0dg5gYy+Wr0/R63Ge
v65ajESuMD63QMSbjR7wvY304A4MGBEB7ZK1Jxvk7XJ4x+7Cw+5plJWEfF+qpb0R
DErgf9JWuU1bqJMoNskUcS4/zO3TPwdAhf78t+H11TjaVMcg5OpxDlUWkl8rGssW
TvvdzSXz+0vCF3ufhyVzhmLVgAFEWzaqIWuE53fxCmlmH2q0H/DxVp7GHGVHuFeJ
luEajKEYNxwmFFa9++93e03OWGHN/AAaRCG8oBTsVxSicThu+ES5q9Mwni9mUxZ1
gdWUojAvadZDD9xJ16Se4ksSEnknzlOnCa7g/eiL6b9+Xvj62c8ORqgT9MKoc8Kh
69W5SgnRC8MTcJ5g+tHvy4RTsv8ccQ6VTKRcgHZ3M4gg0INhNR/DtkZSdLmi1MzG
CwBzM+dQUyPsnv6MdoLxWYF2TRif2z6eE4izX3c0COKVsN3UP7MGb+eW9YvGLF5U
l40REXw/2tsF9oKqRMjng0hEkBJsLa/rVH455axwZOjsZKYH3O1zZjOhVXns3paO
97ct4VDZAHTwBGPfVrrCfY/v/nSQ2y1Fn463mB5uVj5KCLHhZlEtJUFlwbTW7bBM
hQcpyMS/204HEavJznlb2maYdlW0rehEO8+MYRgQRvR44ZjUt0gllT6XC1zBnM12
Xp7DQL/FZJlGF0kzrSTBRamXjDciRuJWEz/Rij3BW9azSWRDajAZziGcx3Fg9shu
lYzYuSuYfkEHkrcdmR2ZnCpzMX5Cu+nF+R/jqCkPT+Vzxgrx/J0YoP4eaVNvj06w
AtMOzU1U9b8f15KnELSqJct9ecHxmDady6T4h/jCFmZ6tPK4qWrhhkJJ4Mxk6KRV
FPos5oCqfID4bdePRF754lILmR8AHeMfuuPElff3qYFXwt3DIfDFoIAMUiDSlPyz
xNz4f0jdXIt8NH/DqDL/8AMWgGY75QMn9rRycTeSI+uacDD1dF3zb/4YYwPO4Aje
uhce/uhK1+hYS5ZEwp17eoVrcIkbMXggtdHgxS6+1Ki5vWkYuBW5sSd+xjHxRBFd
k2VPL+A4AMdK/QpOR0l1Oqo/ZFZPmhuOkyGr5zXWe0PheJTlAeRPNAC5cJYf4tJ3
eTtCycA029tYXpT5fWtXqMdA/9gBajnfyOM7X+YEYxftSqgEZEnS8Zdevy5KEpQU
4+CX7lFMh7kgI1F4Z5L4V2yozwS2eqOgN/XdBmfhOGHvFPZr7F0wm0GC/Oomg8pM
F92FHwCgcdCuVf/NKmxJtTh33r6fnt5kEYjEfzVGvlQAqgJiEYLNwcfU/XwQgQ56
lhWm2HGwAgNLkPMEry0cLJlQtOakPEoT/Tyb4LATaS2i0GnAZkHtB3KfmVNCMBd+
1LqG83fqb/YtUzN2ISPtbbT3HM55sJp4KG0OkOgdw4x25sHeKBn78zVzl4sDimG/
Z2p95B0buWTg411v6Kc35cYZFXOdlxyEVlBilvANhv2QCk8HKs2oupZv95R7MCqS
qQKvMITVBTR+4/17M74hp0ewVkxC/UjXIauh8ZPn5Sae7ylddr1f0kid9CIWyRR0
IsyJdQ48iQ4NkLaVTVOtFkN5bEmldqPfUwIiazwvHJSz/IhVzSJfwoM18F2knIeH
0ipkOGcdKjoxev51RQqc1kSMXJQcsch5FVw2UhY69QwAYGir/nIQuhyxwwTPf4b9
T5BYC5M+edlWtYfcUPo0ezQmb7cgBBNfr+e66DPv2gWGimEW6TLagMM4dB9T2Bzf
65pEEkNExQDkzRshw0ox66P8ohJva0rTeCBgUqH4kymiHHe608DP0BeaUEkz9F4j
iGeKzNfLDS1Pudndwu4DlqzO59DLPlplvkLScPkW0r63FdG47d078H9HfC2/Uc2C
zch3lipfXa2qeljOIWGZimB72IBKAYhPdhqK5uV+Kw1MKcKt+130XBFgTARkp6cM
S6cd4TZbZqZ4P0Kx9g7TGuWFErjliMcfhTPFoyxDGP6RNQ2C6jXJB7jAoK2AlFqs
JWGcjQVBlAeCcTq6zyzokYoZYlLSP7Z2uiUaoqvpEbbleNPHhonCGHlxhdWgDFT+
YqdJdKZjozH6C2wRV6YJj+cKO1ExM9uFX6/e5elniugmGI/ENr537lox21JzAWxs
crkNCRrLNCDL/qwn0Eiv5sKz31gA7Y2A+MOaCv+wNjFTHc7N8r3b6koxOW2ZoacQ
bgQw+dYgSS31HlOmIrBjJzrq/US3YouYHCcQGI39IVQIV+uErOHA66eNiaWnGFSB
/3OB79WMO97zQ8anMWYLOB8bNbpgJfKK23unZuO4PcWhMNR99bK9zgEjodC8ILc5
eLo2NP78/dCs61MtgEMuKqaewQX5SPgstEf/QO2CG8wn0/OdB67V7Idupra8NLXz
UXszsmHWS5ijj70/nvsd1YdH7WpEX82dM8x92/ysbKFbqjxcVPeo18x6m8f6pjgT
PKudAV1L9Mk6YcKX0lB7CCrAY6zOn/jC/HBBn690cmv/FnczshackTzlh/JZwH1X
UflE5DknR+zgHdCwUGZNPc+SnNqfoAmsCGZNj1IDkV984T+Fheq7MQeYnzO6IlYX
5X3EmC0NxbZ9GPvBAKgKtBHQgH+m2DS6xr6KNNVBQMfATRDsjdCYJzkdwcr+fAeE
OklAKiApfMu0gJ9s68rC/7FqrO6/XNZwam4Tz3XSmmEZrgZLTqZrI0eTxrQqSjXa
j/UhvZK53MoIpy/1xTn61AAtVRrQLlxMXcoRm+3Dx2JR0s7uX9e+WgEK4VHzOG8g
oE5jexDEWAZ0KikaVN9QdKswE6lK0jo85Ta16HkT3+N8Gi5PNNHMn/+i2DExraaj
NSqM0nu+M/kpEqzYLo8tsefHJd+fYWToBxh47YdeB6E3w05zWsQBfYtz8j+D5MBM
DSCvilWo4TJUO2+Cmv5y4/LSUiK+G7h+7SqN12lGzMwpAsxECv5wco4Bo9cOLxga
FOqB+2tOw4nqEQ/BxeLvWKBM6cRyS/Wrji1P1OPc7XXBbiremVYDJRbDkSgQ0HfZ
mYlKxNcI1DL0Zd5QYtqb0QzJ4R8z0Ouj/nJtXQVTGGbGx5YYW3tlqsBUrlCVcZI9
5k3ty3d/oT9RUMFUJ68JGfCabLKiNx4lxgd4wBCM7M9IHL8qxwqx6S0Q5VaUqNZj
4GVDXwBj3JIVUgnbegyHdJbd8XCYlg4kuBjN2j4GSJhgf8DM1RWyMXIkT+B/Vxe1
NU68Q8rA2EZH2T56ItuvO/S6zQrqGH0RcI1cJXYV1ZaFs8or/IcL7XujpUOjBYeq
fganJHjIqCzMy0ksjq+sfm/FhH+JoXXWH5yEQstd3kkrGochYDbXKUTNYaNBVo3o
ia4vLJiwIeUoAiDxzxla7rDSwqk8oaJ+WX/oYFpje/wIWGlO//YQaDUzE0G7JMWa
DYuYNjcQ1w+kXUajUxFqsL9J6QK9liN4ycQZtwKick41sWrk4Gu6HUBpZsGsbO/o
/UmGkFHHf44NqagIgGcbbwxoOjpa3CMmzcQDTAA5wniw0KwfgXrOaASE4kci7/g6
IduP72XMAPM5H2WyIgnP1yqYdlbUeVY28ag9ljSs/cj7FooX2FBGc7WRhiTMvDab
Zu3AT7yyzeY9VNkQeKBA+5G/EN7+VbqJivVw/0U/ZGZWaVb7KEhsUpBgX95i6glo
MgAcnVYgOxB/GGdG0bQ7EFdQxrd2PQJJ7SGac/K9+/YxW9/sIzu3Rg7dMgCXV5w4
T68eevEAtd73UvNn2H3maUa0My3RTZgyyK/NLIDdW1XZvd10rjBOeFGhtXjznaPZ
8HFLDa4BCoavHQVmTcc6XEsF2pGlyJ7dY2awt6P1bpVo4dx1NAylNVl8CofQlTnn
B2clbIuMaL/7npOQAY8iSCd+B7pSv5q9HjsDeAsl3dz86sd80y1NtmiGd31IYdcg
Hxj5ucFSC4bYpMby2waIzQ7x1k6GoMQZJIPtEXcrJxtYBLSgIkIw133L32XwEFWX
f+4UZgzdFNA2dJBqpa8q0e8n6Api/RGZbsxOrqDTryDL/mKKOHoOWyxBQhM8ps1F
5jPXXqh5YbVfnRS/W1iIxuqtEOwQHZ24kP/F7LArDXCnBgeE/XI5rZtv/uvJi4JZ
G6fnRsMRLJ26ziygUioMwGU5Cco3krNCUMyR41oAJ2Pg2nNk0tMQftZTavR+7Lx8
xQsF0dlxwZ+zmr7p3Gd0FguDW6wGV8B12KNze+PSuEYmCT7w8iCs2jOXH6KeOCtY
yZceD3lfHIW4u5kfz48A44YxmtwQrBMkASpUBi9shLenSdhHxK9GO7CDb7S3OzR7
jppkXOnkAbViPvlJpX98CDo0NkZ0OiZdL/Nz/DOTkWvbKEUKVztkply86w5IiAzZ
zPB+fS11XsXr/yDMKLLr92Mj2bMEIoSj9yE1CWdqG44smbKpBlFP2k3mFriwcvGe
RGORENJvRh/EX5zlU4FUFa5epXr/2b7ZwWalzVKwUOpmohY/clIBPfao2hrDVTNZ
PTCySxqJF6a7FCzYFI4QAEUYdMDt8GKBCbej4gdZN5ZkCfE1YSMM6qRBTqBLUvw2
jlZl5eE6FC5KkW+TJJZHEKNY6I+YAtHjr6RZEzGcns3OqwpLdMgDOwXoLrq7/xAg
/bG65jNOIhMRe3nwFNS6qkbHj+WS9bJ4YzPw3YiHo/BsSVTiUMcejdTYH6ndUSr7
IM+PkUp26scsbKA2ZvDnr6mgNRAyocCMmJ/k+FwG1dwjIZOvpXrgOFxsqGXNnAOy
JLiDQw0vu7ZEvFkTf6kQYvWrJRU98qWEwOEEa8mNLQgHZrTSBp43tash3Zvs+iZy
MYVHe/YqVQCKpV5Ejhc9GvlhjN6AmTZyeMvGU8TSRkq4QQovQFIABYK8NWzLgVkf
DWC1EHfBsH2rcYiVb62dxmhQQlHkBP6S+5MXQEpHqA54jeDPV/VL0eYxDz+aMoWo
yHfqj48PhGHPFwyrhxkRKs4wyJyZUzM+YPKLKDcpAwxwMlj6Qdm5ryZYMZADwYzh
FA341i6N80mmpEhVb5bL9OaCZGfPHIrFbeX+Rg8ax5sC9cOIzu/g/6jcWOArSzj+
gTxNaArEjEUKwIHKAOJdFam//YMBmuB9eruSjbR/N1CuzaEeNgx+JnjpyKJz4YCE
acJ3Dx9FtlCGXEGtrfKve9oeGNYW83tLfpp8/Q6uJwZjnf9vr8vlWZwx3HTrQAAF
Oe1nT6OXsQbk8dYkZT9IIRI+GptZ1nvzUWNrVE0whwMjL7dTtxpt30Tgu2KufSui
ZoMZqbX3SfzsgyjfN8mqXs/zvabfmF57OEAY6DeD/MCGvalXplyKV4X4MmSIG8g8
y/8ZylpXYKyq714rmYD5i1bJQHOB43lPR9y0gOt1buRLit20ILR2KGcNmwWzDSBy
aHJgm9vuGkG5IHJLfQAqfC/lCev5LJwmfeRYqz9AhwAR48/AXLgX0k5wffSnjpWW
MluFLDEjzqgtcvQhmenXigpVOvHsv9MLf209DfNvw0+jOGlCdoVDQyjZ5Icr3vAk
ThY/5znF85V9hoKgZfi+YkSr92+e43RiqrU+2USgJLGxRsGSXbC5FH4GP3EX3HfV
3EGUdgIsn9Er0cKCm5M2bBwJe1Q/k1yUE7lv4iOvRSQjwgaSDdUD1+9g/PuootYe
pClAKHVoTLfryTtbVCTNtTW3NaPqKR+DaN3/G8mFuUC6cLmokeaIJoK4y0QSSZTK
9xEZDBepsriIGxxQOh6dSiEjKERKwak1uqScBbJTiqapQglp3kT6+MYfgevEa8ZH
sCeo+VG5rwYYZkhQD4j5jzwglQPj+0VEk+BzkGFBqfZSbdouJUXeshXXREzVwbgN
ocD5lqa4eJmbcGcDi9yDfPRpzyY85hVZsHl9GJVhbSGRVISIiPHH0lnLwLE7g1OH
BIZQyUbbyX1TlLBwaGt/rs8V5fsgesV8R3dtkEFhnFebUWoBgBpz10+6mk6MbrWx
chl+zYzwFmee1mwdPfseSDdBajfQ50hAJWKQ14qMN9ImXsJlHkiA9gjbY+6tH3gb
0QF2GKWGuVVlgXqjJ8cXJFhfp3wnpppXBdGJ15HV/OQDR7L7xanyD5ERqyNgon/B
7FeD7vrYE/yD1cfJaDqKMeWgAIfxnuVrBdH4VbrI4hVSKJz9lHcQMvff4YP5zFDl
2fLtl4o0Zp3k7fgFtqP4b/wbocUMgjofnNEBHP7LhoXc1k0kfpWQiFrpOHtniGBr
2iygNjL1k0ku3ri57XyYaeoaNBHWqv6WBq1Up6B5hnKUUmwCF+46EHGEyZhGXAbU
/uIQWNkNdwCf3R/hzc48RE17PTE83/TkkRxd8HNwFc6uKHaNQds54pm9r1YEvojs
virmkb5hyYZ9yrqzxN17bLLI2TSa3bkTa89993HrCXNRq9F4HRMzhakbp4klU6ld
LYqj1GsqbfGkFrE2/z348uzLRZHNFAEszHFg82UOP8z84R3hbNNahsVEQp56Zv+L
LQzPT6c/E//uv8hRh7Qna+NESypp7E4NlfBU3ulaC7SDlUcIlLwbQGObqt4+pjp/
8Mg8M77nViONNQ5EG4ARiLETQjgex3rSArLJfTSkCFu1S6q8ShN/VBwsYy2U1geT
EHplLjkuRl0sarmzTdnelxzuJFjuVyvLA7jHf4EfvzlrHXJqV2wE6Y+qRdvk4XMT
kOuhIQvXalNoXDfIiZ+/D+yCG1NeXXKOKNORQ7aDC/LlXM93Z7UYcUlCuobVg8Ai
mvHfmaUiAofBPBsaMhB7itm0EQ7f0L0yQsa5FwOdU92X3TZA+TX6AwPAQalWlR6U
2+DYwbD//67jf9N9ZPIYpqyPDd7N498L/41VF/a2h6T8MzTnP0m/v1j8YcmkrRpS
z5c81YTraZUMvVNsq7xGUHW1NCxVIxlQrzAafYrBTM624igKjoGkAYX5KGoQ0ABX
ngQFMjJo6ljL6pX8CPrp2hERuQJDoRB7nEQtu1vkBy//qleeiq3Y9DX0Ph/uK12q
4quQPWuKwS5qM4S3Vl+85pE6dTr4AAmtbx8J9UOKxhO+rASB7rThsb9kOrA5lK5M
KCsNqgPJ8qCCCTNr6Kx3JoKp8L1cWpIVWD3WS/DoAMjl3Hju2WShYzqjaj065SPv
+McfDHT8pvPl6B+T13SNMYW/eRAbN1QXpPuE2ai5FMAAWT1nmfiXWeml+geTX20V
Smb6puUKMsscnX1hQSAL8Y8nV+q5nJQ/sL+NQvAFGkT/vr9Wlgc60pdYzVcmRuCz
4l2bV4knQ7iEet/Wy0TGwUrEOvgc7O5tYKbASo1myaZI0Xz7bdSTlouSll6SpQSs
YcZLRT71ROsCXD7Bp/7FdgRC3v2pvSUEe37vlJ1hf2bF2gpeBripd44Huk16J6jN
CEuE/AoAIYRawcudRbwma3HucDB2yOO75ke7iHJdOBFUCy7MZ3/3qZoK+Xno02Ey
9qx9mdYsdPUzTDtQj390V2ly7IfZEfeui/6mOFEP32yez6+EPC2D83wfI3Vd/yTR
p3Usku+b+BWrJWp43hyVCVxhrw+av/DTdPUlSPjjWrs2NQeZhQpG6Ck5qWMZLgmN
DDuInnQAgSXPKpWUFQ1SWDKRDit+ySarL6n4dSWteTnswQ3rTq0MsSP+7hprJELW
h3pg4qubWfNB6wAc5no3b+6VjQbwDtwo4lXycS0TuAsMtidklB2DSb4CxXUWUl1c
SjrQZn84ZcbzGtC2+7IAKT6guqM3CsxWYiXqY7fyUr8daZL7jhVZqSPoYXTDvW4y
AYZ1ZgSkxthxWLIVAnYsm70eCIP9wHV9Lj3mjOuOK5DAFCh9jtDDAZLR1cOqppzO
V+cRIlIiYXqc1VYRFt3YfOGVhW9cKq4R1x8uCkU0J1XFwjcqPVh074WsOHteOlsC
NcQQ9jpw1SAqY+cuQTr6VmoSQnVyexWe5wBRajElTOLee5em+Dm7typgu6JtmTTG
vdd8CkqhnYbb367tWwBj5SosfWxSYjRmlYP2e5bUShNO6loCN8/NYAxl1w9HVwse
er1KsrxUJ8XFVE7vzfuq+tgIyxNHRy/3O4oTkA9YrYMVSyNe0JQAUm+3C3OAZW7q
CuDO8rSHik9c7dKNZEwqXKS1avhTfnoRXiWEbHz0ou1svooPz7alHKzO0O+qNvif
zy2qCqpUkgpB+ZddPsWPKXOa5itlCklMhICZE2B76DovPwp9/65foplvIvC3SKCY
MxsxULi6iwzQ0z3N1xTFc/EgjW4BNGi6MP1FtDWK4yrc/0vGHvy1wZsQrtykABwY
MPkS4HsdxRXqkZDxSknAi5g56E+L7eTPgkFVUCAgvxBkDrF3fqhmxzA4u+jeXBFE
rL334T0+OI7yFXttpiBvLnzOdkhQcnBqJO8/k7mXFj6Goeu5p6jcyCoY8yUTPcHw
nW6pAsuvSXr1JOEktBjQIc/H2N3p0T9r7wqL2IhuRE6KL2pqTOsk0wrM22AYsr31
GPZyp7kAMuxO2HapyFyrKHDrQ5W6kBJE7wKZ92EjubYQ01HGnD93uejGGF8EosAM
0tcUTD0udkiU6DMyExRYTgXLc66CMrj5I09eZnjJNCyP8i0SgbAL60SYVA5mTNhP
XnC5xyQQMF3V7675axA2wD8fh768BlSFj1DH5FUr0pD6VkMVtQPBj5JQDfFdNS4h
ya4IT2wJNLjyyx6FlvWYrJHnt/y9p+DAqxfWDo1zbdJX04Q81BVSjBwrO26/2UfM
xIdOg0RQylmvxzw2y8I1+CP2xF2/Z3M/w4DttMZVYupumFQnIAGrSxgqeZ7Be2+n
50L78g9mM7aDlL78WQ0u8DqI8qxUhYIto6fHM0DXfi+eBRp9o+DX0glY+mM70Vt3
Kg6ICCuthRBmpfQ71HCFy6Drrm8nbfvrVKQZ6NYWDKmftmH/LXbV3PgsEKhWIOoG
s75tMZR56HHx9iHJKYMBOjMvD6owWtZ01Vs1WqUJnTuYCYpViZB2dTyDF4PwaOxs
un3ddQeRVIpC1LmfMJMOSVLFTy0/Cp1umdMaxYbbN4L5eIlYF1U2z9al77kUSIGZ
x/SojUVXlyq6/I2h95iJ6xxS9inhc8EO02LTCRwv90PWykHUb68QWvYejWalsRBR
1kDwV/dDboGh+cMovmZ5kGNLrVeL43pY3cdfX0lhfSLlx/lRF4mO4qhhFVFSE+RN
MceGRlkofb8unEc1RvEnd6+VBIPDeLeNnBpObskUc+PbmN2j0XtiNJx+X+241jk7
UpbiMOCkgFEaxsOj5n0KH7a9FRKDWZ3BqDoXB4BfmIPVcGs0QNgSc3bwdLpnZHq7
j715BIFttZjEn9DUycazLcbwWezzO6BcKR0SgupdI7bO6a8rq45iIsNeshyO4hQb
O939lBNLY6DbBkPlkt7GKjb95Y6xMTtrwz/iXpHd7iMPULvIgf5/ZVBq+zOU1qp8
YTbtJxM/NNjjbv7+U6RsvXl8JWQlev2hL1Ah6B4acF9gLByu+kQ8O8JxQTun5XMl
OyEC9bpeIk/LZH9FdK0KCRq7rkE5cncJldUmaICKtcvZP2fdN7jK7KKYVAeuh5lC
Z1MQSDR6liv76FCunEzuW0Y2aEeRvBZ0zhdvmBzFVs+u0U4e+y6BGNO629LL2aH0
FUSVeuVTzGvewzkqVeTyjKgIyJv53Q/PKSsiRCAE5JRRk0aO3U5qzesoq1LHmN7D
540nGHTAEfX4MQzV10l1UEXMx1yhMXFgbaiNEtHXNt/+NCcZXNuaH+VyFnXRJAHX
Xfh247w6ihGUQPngRHY+6oY5OmQTj5RlRmX1pxgVkMJraxverOoFOS9rT4RfmStl
s7d52UeXKOOidkQzU7FB98vQpWbTg5OQImoLQMNBFQHf3QrVn41MSB0g3bmR54Ro
1TUfQ/iT+xoLi/QroJ1gALyYCjDXwiUzhs5ZzFXKgENLHlth4aEpDu/rGQcWFKEp
80MdcmzcVWviXDNud4fSPFiAVGfzbhCalC6KQLrt863YvY/wZGMlYox8CaoGmcH5
ubN9Dv1gcdC2+ZFP7QGvbqny9OhjpUYqGGgvomLlDzmzNUPUhPQ++zYJOCRj7YOq
DQvDZElZIyJ2JQ4kkjASfEcqZ1ywWNIGSN+rYvCXdF9suSlSoGHBdfh6s+ijhD4R
uyCs2uXbUCofRySCwB0gaYAsx2BciT5x5Av37/0NgTY6Lkf45qglchC4EZtEsKWk
YVbswTqT00SYKIc/NpFJyp4OXEYLqn5DCWWro7C/sRptlUb+h1xpzFgMaClhPbwM
ZU4ZSMR7T5zJ18VMZ4VSwI/Rjsuz5mw8S9etw55cUG9JNZu9z4HkbNA/7E+S4DDF
BEqnVqjSHoGjhW22aUN49kQoCU0XnMEF/ph1NFwGU9rARC5/3anYhpjHMoK4gX05
yLfq9jeTjC1LBfry7ZM/4qLMXtiDyHtzVVOtzg0R3nMXnOEmVuDDTjwm3debGGio
1kYNdvma4KlXpqXFivDnNb1dqr+6qXXmmCG8cn8ltXqD4tpzj9eJVVTsAfWBLYdY
MhRkJQTsVBwdfBvfaaedMNLobb2Fi6eT4vEF2lx6lvlwHlP2e/wFMvsbabz4yK64
8FAFDv1iHgGAlg+ILsgTRb57xDasbCjDwE6SYePTfXzVjW4tJ5G5+WOeoCK+kWsB
u3ty0CYPMYi/pugQql7ARiSyD3Tn+/idxJllr59kGr40MTma/NeA/IvZVf4i5mEu
ZrKla9471QWTB1nY/8KJ6uerQosmgD7WvAElVLOLssyZUkEWPUebeNF1Fej8fuAj
rOkWKFVGQwrokVTEbV29kDj4rmDJ5MpNUiQyHWLGsKQhnyb682OfplOngM2y/KkV
coOJoNiig4T1UXhW964MnM806W7rUD6ljaH+bqSDau0JKK+tXjXuvfjLpdlW0xyk
bNwLvFERks2wSlE2GbXy0cBYJGiaIZEtu/IDGpdCa29FDp/Br4iG1n1IP0YHMuGw
5G6g6skh+bGIM20UKQrV08pVqhdXLGnzskB81EValuXJ5XDDhsZiYDJFjLFFBykg
l13bDs/jqa87U8iy/SFN0m6rV1EwDXNItCvtKj3fCDeSr8/aCvkXRJI7vqfrOh7N
uwbVGvoncHI8C6p3LWxdsb+D3f4KcRFjA2wSeKNiI3GS/P5SgAimUy202BsmFEcb
vFt/WnUQA8EB7pY0vitBfyparPA5lKly1J1waJr7VKdOfejkLuD3gPy9umpekx7G
KEeRNH37Azvm1ox8GmfD5+aunb7RJGU+kHThOvdRwsIJ9LNgKFUGVD05cUWcBRVf
3Ol4UMQ65veewNBLvdmWXGr9LeZI4n3uHPwRbZ0rKRXGMgKUQbKDRrEWtOG36N2i
xIqqwNGQ+bNGu/VFlqOgldqXAKy+NscvmxAgQ6xNg2XO5CesMZOR1aGSmb1tconp
h2QcIwthdA2EVQshICw4mKQ74EK2IMsgNOEzzYHSWyLyD/71gvXTvnYHpit2XBt7
JYODdAy3JrC2AOYPKFywUvxlgn30k3GGXBAXnCcH1x5mpDqqzXdLpOMZyjqE0Y91
19TE400WCED33hQ9Osers4S8qOtIQra4O9t4XpQqwXy7qkBGrBC+gOdk3336V/2S
q9woNfPnLhwrEhZizUWuW9JbZUOJHjWkBQGoPQegKUSIFg3R7R0wL0ZGeH0bJhWX
T+UrIHMzpB6V3H1nHbRQksCmjgdAhETm4yCPLHXkiCITIfdUG1GgqkmCkVmR7bwU
kH40ReXXf+22oJiDm32u096WeqviRKxwoloHJvwdMQLsDtDr/pqsQ0fiY1nFBX1q
Wr6PtJeek6XzG6xtEKGAmxVeiKJyOan6dHy0m3AwAcEYDFeO10irRFvMTnzWxEls
MJTUaFMC8rvjWY2mTCgLhA9+dUYWD0JQ8+k2+EZLfkgnJkOgGRtDwFHEfMy5vZy7
6NLM3BO8X4ssh2tFsVK+v7nxXIqMoxE250DvrHnt0PRQDIv7UPEhcflBbiHCNEg0
4ztxubN4/TEPYQ7/3AtIezFfcDewfUwsNqFcMBf+p2hu+YAenCLqWQAAS2O5mOxA
90wH1rV+J2vGmGIP1j4ZD/iqYDz9YCJGDv299a/Go8jCiuxacV9W0K26mrfIK7ev
3i291JcMVV6dqSbK+2G2GAHZmlzwj59IDl56d/4+qoNOhflFMNIQoo0bmyj6lJA5
dvmGZHHcZGPaN+UgI6rzrmBwye5/Pedn+FW1rIfuOFu8Ia26YxBqATwde5E/OgaH
uMvDvytv3kHoOaL1hryp3XWiDhN7b/nAxQPFKXO438rPYcSF7EWKbiXd9NzgQzBR
KXkx3r/HtZkC+KGbaGNo4v8/kNQ9HmdqEaFvri1U8c5QhDSjkjamgrLlVKkb8Sj7
Ax0CXyhlp3BuhOWkBIu1xUhl+ha78W8Sjbsb/Mm6wkRtf5/TrfwIBcpHR/7A0Jdy
0HqchoVvMwva/QnQ9qkTLw5j9C3E+EufVJuT7PleYSL9BobzRnNX6+fbSL3ULbII
1XpDgfcBujW+1t5JccIOxM70wdRFNa1HmCeY2SKcbjC1BhOxuTyDAwGNABFqcFtP
Mu7kamNjf5IJ2NqMUiVY4g7vcag1H6UFIyK7RoqPhU9QGEGqc7WB5XXGCM82VbQO
t+XvlVuVkftwYESmUbV4zOugX17lc3wIzc5HuvDZ9gt6AYnV6g3SGSMwTue8YwXE
gQASSVxZVZjoIS719P0JLetCIHjlzVeP8olTsXcJ6PsFPBQkhU81/F5j7GHgWIhb
rvjd7j9cy77nivo6hZixrAWrBrZE5QBDUiGEpF01iuaSoqWjnkB0np1Cg5ebNuNB
cqGpjsBslFE5JwMJAA3PcMaIQeVeaQjT/1wojz6D2UHS1Nu7wr2G/mgr+RACcK/G
5/Sougnjy6QFXp1i7nLREvn/YRuhjb7xwyqRMF4oX2UCrWdwVG9gNNBchKBYVBPA
xEkH8N7/JObm7PqLoY5AtzlSRbzbY59H9MHIonNigfO8TiKwi0KWo7KyO2yDaiB9
a1T655lsmr0FgzRCK07ifuC6tpdT7LYkZYeMAaC5iaGnPQlx7jxNptcxKFQErT4K
DXtxy1zyEvht9tDNCzCKj0aFEo2Tiik9QsonmjTYmz2s/CNgW8dYcqk1+Wk/35fa
Ux1CFvgAfeo4opQvo15A+CtE898Iv7t40sCoBZu3VoAOW57wMKK7XgEL0giEek/f
aArUWqfpipmVxQyZIqwLSwyGsPgh5Sxa4t8v6Rxl74iNhbU6jIM0UR9ACRsXLpLC
pmaRURQl/mqBOxa30CdDNAX8ly4m6e6SR8ZezcqvMTF9LRSCwIzBFYZP6SbQwkE/
XqjpFMknmlfKkgRXNotvpIDl/q8XPz0/TtE7L52WosH1c4Oxkk/GOmTuKIvXxlbh
PJMXbTDBmLbKealMHySocvzrhPVCCmyPJFlM4MPNSIXNSwr0Kw+x/sSdMaWAi6IL
w33HD0mEocp+WzBYR3XH9fmQB+makqxTq/GVuQotI9uPFex0Z5SNedyDsKK8AwNB
PUE1KsEyCIYhNlcpwhGgmG8cNQE7b+EKn70H8tLklmRA9CudSEY6bpsb8GxPwp/Z
RSfThKsO+FQA7h7evsxFMbchLyMQXU5qRmPW4nCAeGZcmHSrZcs2dTsTiFzyQQVm
3raCC99vu671o8z7J4L9n7rcxjgDyMC2031XkEskYk/ADMO67e15E7NODgP55HXK
TzBiYHxd7yk75yWZ3xUx6uW4TzBQEhvfkgCbHJA3V3qraSaJoWoQi+yZxzYPMihj
e2MLpnWkQgWtwKdGBTR2YZ8aM8Tk/+FLEuZpApjsT8SVKNzK/pyzyS9p0fL3DyZi
tV929QssMXhjW3kY1NhAFSdznv+tBIdzeCgURjLPY6TN7Zymz4RWHvXYqDyvyhfN
pC9P2QSKdIOSnUBPxs6anIX83XEUcMkMfl+Vk+qKG7OByL8NG6ps/bAoBXD19bQ1
irnjy7nrq99cps1UULDZZx04v6/JEoqDcKjzIsThMuwiJokOJtO+MjdKL7vwAtyA
R5GJNVirWkHPXzDawipe/3C5D6N9X5/4pXSpdgRmHvOgOdShFc+Z6G8K0k/Or0oZ
DvHCkBpZy/JAxcIL5YH3ISR60T59eJHc0/6wErXOE/qF1n81hFCuDI2m8aijuejD
gRL5KMqywQ5ov/g9IBNKcloPtiLfY7c9QjdY7wEn+p6qrfLw2698U+NZMNHWiRgw
dj5jRCUpWmCRWzKWQXlWNe5mpJwF/8XW8Qbl0+3THgXe5mZacLA1m99DLeFVP/yl
lZNbh1hwgWV00q2TWAINehB6NMizCgtAJ6N6JOw/dA4QiioisDAF3A78okQGCEsN
qdBTBCqBF7gPaKjaBXiQUw3bycMY09YwakDcF5+A9G5vn89CZhmSkd6IALDKXEV8
OyiXnJaANHPgJHuozXFCaVwPhHEzXpWCAqG4t2OU6eY+CjWcnHan1I1Es/CzwJOn
pXpn8o/xBlaa6a01+kFqZOr/n5/cNbD0hTmqNx8lJD+0WD2AeGVyN3U2NTLtl3Y3
IURzMCeQ+8H2wob+85s04JWUhBhK3S2mqAk2Be0YY6q8ztyl6aAceBblPgXEJabO
0XzEfamtB0xZy1ZY3qV/n18y2ZLjgYD0pyksWUGfVkPjI7W8txLiWNkONtDOVSH+
HQp1w0SDKicVNIhUxsj60p1UU8wh8v9VSC2Rvixj2w5gpPgveRj0hf9xuOpNHRMj
joAjdnLwyxtMNJd3NSQtbl9ZqC8c3BDmTAAPtRnrz39aKzxtqFRGFyltHtz3OFbE
viKEclMCbRkSgog+ft6fbJycGj7GgLvg51rdAk1+KTNmmPZEGTygRMHeSS3JdJoa
Xk8M8SIGHojoTGx3Q8ss3hZLiCP21p5kjsygR2H6hCVhN105RE7ZbfibnD3EzT5z
VkQdb6djamGyoU6neICKsH8cegUn89JZkEQtJzTwGuXtCaitj77w60I4p4xSlkTA
+xsgIIAyKEtkxKzM7ntb2BniwtPTTXxSw4AUJMEzbyt2vS6zszMD6CwIzbQNB6jA
9OwD3yA8Amf+FWuEUbG+8xcb6b7bskyMLO268AL71juS6GvCkG5wNoX/KMw71giF
15SxzeThUeSC1nPg2w9BeM9Og/SheZHriXeUDZP68LDuVtpmh6uHCNKDMy3Ze14k
dynGMUqnaDg6MEAyLsq6L0VeUbxc++GdaHOHy3P3F0WQ0u+BRys+bm2LQE6lbN+Z
q+fb+DsHnIuDHvIMlx8jtASWW2JwjwnJ1U90HHUiWsPsjhn46PzkeiLvIGbBF7j5
BTahtFAGoyYHqjeB0F8Yae9AXpVtcUvnfQ9X77Z3PEy2JvcP2o9FGMkzT65n7Gem
32E8p0Svbj5lHW1JS5KOec+Xv/ageH39OXmST6wQZgmBrHE38Kv/rawRugVmPW9g
x1xKEOTHZ26Ksmr8Dyg2pEgjaES50YZ7pkZz8sS9yaPLBPVF/fJ+TO9JTzcLlQ8q
4L3afQxB6fch05+p8QgKSUgBQ3isIUKL07jySIkWPup4/OBg8fLg/cS+TvJhfSvy
+Cah7WJvZD1b36ZpBdGuj16v1sYAWUKSJq89DjpT5DDFSS5KAkpfh7ikHtY8KhYP
1MmWOGZe95D0BcRWmGN34lmzLS5gQqAU9AMDGImMTDYDyddAPUM9rvCDnSFizCwl
zuTh1LTlHo0ZE21l1cLA2eUxQjIinGub++xaNd5z2zcW+L52OHU9Wu1G5a5y0Rjp
ot9iYOVC6TneCfNCN7rexuo5RFDI5Wi8nEw1oKmj0lebE0jwV3Uow4uTcLJGkxbM
epHTGIFsiqzqUT2uSviQNwvTI2XB/e1MNOUF6xYETRwiQz78Cl31jvh/3smiImVJ
FQgJVR9Fnfc/uOE+T1OFO/J8NMhDbFNwPH0LDBEWfgV38G28TgqZMQccCoIfYW8E
sRC+Pn436UnEdmAz9+4DjL6mQHfIohrl8eaarI6ATSCaG/pIejHjJXCKg0G3Oa24
1Gv3CwnGvC5HOPj/AcHmGYIF5JeS+lKYC/9NxX8xCxTpll8HUsJErwFgeXcEOo3y
UeAyRtNvinwm5sxbupkkaGlvhDSvY2YbiCmZtyLUDqBVJGmfNnvXbTbkO/EMi/1t
4XPm462DIKsmghwM9QNJQBij6rt6sOdIKmODT6+2L9rVyzstcfCPcKeG54uoMp3I
/3Q5Q8+DknFH4utEhNYWXWH29WMbHWA4cUIBUifh/xjP0pgZnlosPdMIlSoQHzJC
00MHCHsvkFM7DPptOdnjFzRqg3zIvLioCfPnj0kn+7y1rUFXsph10upwKBLKANjU
RgLR80aFzPkPVZzXq4/TOSKbOzgYZwN1oHDIPOo8Y9yZce1VOZMevx9w/zFxyc9/
X3LIobQ2FGHPfXLhRVS8RsQ5yCiDrCyXUzB2V5hIZVBujsvqYyC3tsvvdvyi2Nkf
yJsubEsCyK+vHMLHlv177+X4HKBnW/o1vPQKTkJReas//Fb7lxGbgYFl9vLaF/hQ
3Q7WwgGHN2lzE66BT9Ncvu6gFgg5jbJ+qFV4ZoiluMntuzw40CRpZ42kT/3Ck+Hn
y+Wc+vT0s74XKJ7WcXOXTb+NJgnn4Yp8yWGsPFeg1zDCQbeDtjEg97zJIBbBxLaQ
KfHyeoMHE5jrDaFTIltQxVA1JdMkw4/nXCWEQOyT6NmEQcrYecvxwNbeyaCzyPV2
XqNVUlR5g8IaSMHwgixYaxuNRqfC4RZlcYCbxSb3D7Zdnh08WUF8uKWWWBU3w269
I9aIRDnch/8o4DjNx9t6+Tf/YlCqgpzUgz3JZ6c5aR/PaFQMceHUdexoE9gI90xv
1/JRGm2ifn1yah8hYzRlfq2xUreUJWXm1/8B0DjIBcYRMHaR6m3cCO9VEHGhwSGA
AbSkI3byQHXzOIUQL7cSizer/5vzxZ/PG+LWEsK37eWGQb5tUR0SkZvOYskMwScz
vMAu+y2deyvHmFCOU2mOndJNuYtH9BRnmGBBxRCOj9MHti86RdW3fdIJu+olv7YA
A9Yslnd/n4THyqClYeF3cQpaXjMq1uos8sh5wwlP5NGODtl38GXmHc3Rp/c95rfl
oud+MgQZbZ6ll4Uya9+SQtBoqoSH4X8noiWTlXIc3lmUGQtYQl4238pjDkEbrcid
f95EgZY2G5FMdjIEb+IGn1E2Q04aPUmQdcPEcORA9PRgWmQ5YmsKxm9DYR0iI7UD
D9R+PwiNMhh5KWrKaAyw/XjrPvf4gqEpbvHk9ovWUcpzxeyy0q8jhX73K9yi7Aeo
Lutsdt0rB5sMSx56fSGGmMrgAKCAck4Wblbg17Cs5Cn+6HTVQcDjLvLMsPWvjeey
XLOtIscuprE6V4smeCkngzMzxKE2ndtg7CQfeVJ/Y3vYBRVoWnyegA5dAfDVQ1cE
KtU2BsySzqKGe1dG7zaM+mUt4WSYGYMSWbtC2LqDW/Hkb0+VLb9/TrDbrZqVOJAX
jHC4NCJyHXVJ5t6z6rHKHjyIUfwaAScPjyMYtCVP8JEjareVvQnpy/AICoYGp04L
Eocjpp90/smf2Zlv7YIB8xmNN7Q0Og8mDeBF8bfg2NyQsuvCdg5VMi25+1zYVbGH
gkgfe1ikEkWX6Hr14Ny9Fqhmcq+T8D0IMB3FYETguKnGqRZ5w8oK5lkX4NPXHcnL
K4t1Q8CO7Ki2tmkzHR2e7VUBPHwVJdWpU3YxGbS7TctDc6JM+ubt0NVVHjzzvKoE
QC08FXvqrqz1kM9vh8K93puj6hEL5T96cCVb2ip1kFjDhfGlxrkOl67MaUN8UH2X
t0wHnhjYPzlfWHjZdnknyda/mzMMO5Ni7uBO/kY/WzlfRXOL4gBdS3c9a8HuacNA
MsQAmz612/Vlic8N7bv5GpoQWoKbFKLC5UEFZAraqmVuJqpFeR1zc5M9okxowAwb
DP5KUaLQHWGHt4hyLVKUrj3hrhIFZKeoXJPX1/qgALFUXdBxRbMwAu2/FY3evtZ6
2xC/mWBRel5W7ntLtMJor8v4lU7LkTmP5bQskfkl8NoMp863vnmLWlVXzuer/ytZ
gI6r3OczmBf791LVInOGVer5CsPItEWirlyqQzY2XMFAccDlWxuUNPh+XRh9mFic
wgM4JIHFh1OZlqofpjg1yCsbSkiiUZZ0elUBS5qaqCvAPGECF0QIVLGunPq33Cw8
rwMilWCSf+LztDxkZ4UqPuhJUTH7QxRb6Dk3rcnGvPPCSzyJns+8yIC+eHvKT0Zy
AhOvr3huwSNbjobolbbWTM/fnhAwW1JYuSQ46vOA5tRLMaz5GIo6kvQEKwlLTNy5
wGqOx9mib/plSW5ZFyhinB0Q9i9bTw/r+mYvhIZY3NWmp3kWnsP3vYY2PgJIG46u
JQQcqlu3vNZHpFyomWjUTMYjW8aqkd55FQKVtb5mtLbR3oRXYOv1a/IVvFSfUWpH
uPVSj8G9nCDoXx9nu/OzUAB2w9YzL8ij9NliHN71k7qUmo0rSae31aErvkR9Zq9f
9Z8NUFFGQxr+pqivMaEq2sJ4+EUU/JVSMuekEIQn9FqekwZVjo0KdlB5P+3CsDOX
ThjFSiW6AZhUc41HLZWcNN/qvKmSBR3m9bivgZHe2tMbZACmG2filB6XhfWVsNq2
NGUoCqSauQluX9TA0UPuYagqnF3fF/3SYEhe7E0S82j6ZNt45ZdFOq0gOCv8HUx4
1gcpA1Mm7nQpYqF0nOwHV+Kyux3vTh0jypveYLHxX89iOv/r3w8MISPYIkXdePrm
iMgohxoC752a+LSF5LmHAiG7mqOg6rLOfQ3wM+AhGhoa8qUhwpVcGPkuEGF5JERC
MpCbaTOy/Zb0NyHgXf2CgvVXkjAW2GwDlcmlEVyNWjxVKMhKmAM8e9KBk7yU3qpl
ZehaEI3UwrUdta4PutGbPlNsZaDaR4CUry4pgZwy2Vc3J/IX1LSx9SQPHdU0AG3b
aXcJ6KCpFwBQVFGLNHPE5z9gz8bObn0gpmujD//T2HQXCkxcXKRxs47+zfm9aAQI
D0clU2/OjhD//fQsLJIEFa03duw043jRcwAvIgvD4+0LH+ZoYe7LyJAtNWiLNmvn
OKqtDJ0ExdqtrfwRR/ul37JD6swoOiD56uDLmzwvUiXD9v3D6AXRb5Od1blaWmC3
ygT2ywesBEdCXFac0TM9RzhOjuzXBUn4jwoBtOUFRxE6ORdY/dzI3/DXssmxbqHm
eLVcsKsNuZEYdKWQNBsEzp7XE/HbRCa6bR3KAJX/iRkp09ctAtkoQhjwwca553PY
b2OxDVTLavlqi3OxVE+oA/PquRN1pzWg0I39ISyOR9Z+bfgjzQoCUGqr6DI6tOK5
Hg9n1dlwpOHJu2KnRo7DxSpFBy7LIBo3j75OG4IZCZuBgUs9qG7xd3c8Ttk5GDkl
8fjnZba/dX/rPtGwg//P2zmealF6Mo5tbX+yDDzasq6lZHNdK8uHHhLKtRvokOAV
vbwMDrtBJryLLdqgXVwY9hcVb7SEjQY/eAqvLoJcNVmqhUnrTg7+iXQzqLjLn/4W
96P+H9qDXjrz1FSHHgxbp3TiHrmYepjHo4Baj03eKjiloBDX/TpyicgE9qGalQ/s
xAp0RGY6KIrT7BH5uuj0oVGks6I6BtqGWJxz5ss6za+jm3r4ygz705dG9WYTj2Z6
IoOWwZcB7gHiATuucwlPccZ18KGfjoN8t3q7kJ8wD5oRgJML+mPPXAJAdl/84972
6K7VknW2TVLH5DI1u9TS5GsSMm6vs87LV51igSz0Oma1tribN7j9P7DsolHMrr2X
BhCV+7SuvJNt7zbwkI/UNyMkozy7zUcQP8Nt3U2U1ZxqEG5ygygZvyLqWtfTDrQH
SGQPpY/6cRaidlyUwHQQbmsaN3Qr6MffOzo24FI3RBemWTtEeQUvObZMReY2OsSN
JEolQg3KL4O1uZUAfHvumPnCwBdQD5L2NJLDucfktGIKjsA2fxkBdB+wgX5wDCCZ
JHpMbrSXfDvDMl4hIOoQ7HBOe4qcqQTK2nuJt7GkvjF2cZht+FtFqj4hr8R6IaxV
UPwX3G6VZMz/nkqrviUBTqRBs/p82rfUmbVzFi6JSAkpcviqFDxmMsFakeD3JaPU
56LtEsj2LEwmjq/o69jjIxMX0xIIizNJJ51uf0vTTYf4Ujx/og85nZe1LpujgTO7
2Uz0DzgxH/dWSp5FDCttZHpFwvu/5qHmKYKbwXmeTL9rh2CJ3Ftl9EHFH4R/j1R7
WBI4J3KNjlmbzhqvaeFTULkLBXltOs8tLF4eZsanj9VBo38WFgZ6GwQeLVdRDxtI
1T4o/L2GPj7gly+Ml+jobezQT3miRJXvyGPa60EQtLqGqqhw7YHLs1wWEnuYZ/Y8
dnfWKThEOOJ4kjylwYlEiK1KdXkvB+YavwRzRTttCOsoroEYIy63w5HaAR8vi4A9
2YK6T4Wpb8wKQyCMJt7fil/9K4T3RMjHx7/uAEIiYZoVuUn1vftqylIetBm3z0QP
S5yHJZd8kdkGkwOR/XzK//o6bntgwQeOxV1+1Y7X5BuD+vOktC/KZDY4ZiT/2YXc
22vfAq/7nEOOstKdyEmnVIHsZJZPub6FZh51i4EhDPqytWEpuFoCoZV/S1VLgdDL
ir24m1gduKwpqJ7CoVHKZ45sRkss9+ZwJJtXIpTOyXQx3RcFXT3E34UPFhTHca0m
iNHgfj0kZu0xPOVqf1JmynNYAaNPRdETJrY5UYUtt99HeBLleLIx9vCr0xl+LQlH
jtX+hFxku4GdnfsojXiZys4dAhipJMED10okatJzWSFQ7Fbbr4wC+OFRKRHT8dMx
64EMZdZifzW0E6XLPPvhTcWxjGrVi2DgCvdURySemj2HQswC7o8+DFhxjgrO0x+W
wUynMcF0oqJlUSWgQD+r4XWbSO9aNYO5utvo16xMsroqSX34Gdwwcp6z2Def7Z9J
LXQCvjW0KL+yVE4hJqAi+DkkjUobqC82IkrbMfwFqLR1uSK8gF/LaXlwP6uk2fHP
w4szXhCU4oaF2jgZYIJKByWRcDmBoZ8OzbY7cGdEKZ7V+XXGrr0D+zriKhljGnVd
nDAoO1AbuQ+iYMU43K/modeYgRmilGD1VC6QEkMVRLndI71SSG5Cwv4V6UbvvrS1
K8pY1YuBHlGMFUFF/hm0jvI8U3YMSGEozDSe91xaMH5w+oxaeZC6Z5mBlFMZb5wM
MRT0DtQZv9cqTGCloYKS2r2I16HEz4xPQ1hEhMU8/VuOMoaFoiMTM9gyR+xBTO6i
7bs/yi6lSfpmp/NxvI58RZJe+Aln4urmUK8W5EviAK4TTrWOUqhUPmGpbwtuy2Ax
oF/jFL+nWe+m5KsGZ7yxepROER835vINuy1Qo9Q82nTttUdj4u6zBQdbbHnYE7n2
kzuBsxdFN+rRlwH3kB4I93xjQtCKAZvH+mttjJBXO3xywy/ogpgQmd0gauiOvg9S
YpEzp8ZP5gJgQlckbr4W7cMqA27Uzm8+IVj73uvddAVUptMv5B0flr42b/cWQU/Y
IicRUq27IztVqOX9N7x57HwRytCnxbdf+0u6+yPoGrBQFhd1pEYgCwoY2yEDd8gs
h6dzYRfNLUG/S5BDehTgDUlqsL0LJAo8llr25E+IF57H9inLVWdxeg1fEUIkmEiH
ymaUbTJxMEx5y+nBQDctCPAQsxm2NPQ/Aluhjp+TIaQ7X0pEpsk7ybEE+dV7xBWL
x0iP/RXTjuHWWzcDCtzZY6pEs4lNqe1hSDNK/2UqRztTj56vHzWI4oy1PPY4pgld
ZDrMslrOoBvXaKLBq+o8i6uRIDw4wffslrWbrrrG1ttElXMWxswV4VnjIfoVOluK
Zlgo2bXyMpYuht213FhvU7vTh7G38t73Mqf1NmQ8K9bzxgRjckv+0EtXY5+W8JDX
+AadkY3KIQmBdb4XCsVN/NzpVGB+4mesUOI5kBYK/1xe0sB043aTooe+Gl/TbiWn
GY4CIXeg4GMIzP/c7S4BMirSmXtqR8q+6m1LVKZNdmsiSgHEdhpYWuwFrQSHcmxb
fYHKUFuOJaJm+Rx2tyLdHBU/Lh6gEOrpHW7UKQBy95eORnkF6pEcBuLIEo1AoSG3
IwyZIBmcR2FhT8DFjUbuVgiLHiV0N5j5FBPwLqIuzZ79fDUf30zau/wIrFPNuZKE
P53JtExMgWq4Rbr8fz1zEoZkyRcX9m9iOzY2xR6GLS0Mbg0RmPSkL1yWPWh8Sqam
FPsAZzp/8OsphbxTKEVh17nSkmMcXowJuU292nvitfnuG8vHV5DDXJfgaVx+Kx15
t5+Yu2eN5e8wtMpijeLD4GwA4mKDbhQzlVvUONxmR14xN0lqvEiIHnwfWvFFrmXC
o8ZGQDRC2bpLdOxPwN7MGio645dXPwc8vtTJwk+uokSk1JJjaWjWdCFuoNtmEtVk
/EphkCD/irHY0foWmFc0ikdAX3ARvBNMSaSkNN6/nxzEMhu021rHh7ygmERCwjkK
3LfM+vvfZI0vsWfPU+dQQxP35AJCdFMqDn+9/ieT3BzCtrVHldP2HMwJYQBACSDx
RQ3vUigwKxojUN+N3AGCuQ8S39skQyTB7YRzEAEoK2FuYOEiMgkJTAcJMqNVXW2v
KKpeIM2dh87vuBXAydWgfkCmeZlHJd5qMjaUyVx3RSEmcCaHz6oknplc11wspfZb
WmQnvkfRrtzu7TMi5KY30CR3vXd0PBUIzqd7fezaqAacVI7Wh6VTEUjoI8sAy0IA
95gfSuK7UX7l7U/VEWuq2w/KdFKI9to5gkRpz6SfmeewUg362pl8DQ5OITqnvsCt
nzbonTjPDw6bw/sLnbn0sx4ReWcQJj+5fP649hSQrcLuySiTPN8LfjA5+pEF79MG
aiO8PcEU27hl/h0mKPupMtVPxEISPS3OxYltPIG1d9cMkwUdl4IhIP/buxsjN4fK
jvNLOfxyYq8f4AKlkXuyiqRXRF3szWR2yzSQ0awpBHDXo9YRMdtPMIO5nGNIHWJh
t5MZW5eqQ7FwlQn5Z3WYmgdCa4BcnQbw2kubyhrk6hhjEUzCSZYI4+zjE5hBw2x1
10srAkRfe8NIcVecArnfqvTk1lohDE2cB6nmaQpv0tLxGUw/Ga4ak/slPjikmVCM
w6TlTOC34PRB2ioGDxBkzU38+uSTkmY7DwhG6ZTXM/0AzpQyp73Gi12/JLTaJePq
pXBx0NZniWXtqTWxjg66GLft9TSXXCM0ZoUkUIRrKVG9KirbDoTXSaTVO34F5Ke9
RotJ9ezGRn8vKt7BPgcmG1mc8BBsqTrfslkDh2pcCnlJM7M0Ap9aqxlhD2plAvhX
UFIDdwnYRJYqnjDGrQQ3Q86dGfwh0Sk1yWRcQgW9W8oPkjf6fNnBdojySe66i3ip
oLov0w3OIE2vp9pTjbuTdqvLRwXqZ8Ww2XhaeIc2AdyCb3FPpEZ6KTpd/mT7fBTK
Ge5WXXKDc8xx2j5teV7/jNPlpdplOvxqKuFIBF4Xzyq4JFszFINZH8UMnxkje/nc
9VXGAD2k6sSDaH06Hevg8Wo+/wG4NgTqgO0yIljghpMmXKMTpbHoPhdUItWfOU1+
hpZD80WU/rVbfCXvHQhPt4oZiFv4ygp8xo61fBQ1y6H4pS0LgH6ekonbyWh/o0L2
dPQIWuqK1LBmgSmfAEnyHEZusUmjZ/B+TwVYos7uzS177ahDQM8EIyW3B1aF5ZPf
PDK5yevw28QVDo4GipZz1R8lVFL3N6WuacrWOnz7giJltWC6UXFyv0hrmjUqTGoW
Vwds8+VPNZ0HvX2IC67BCRQ6s7zsGGCjejCNiH2qFMsSHAzRjVnXwKIu2I/pRI60
Rtv889GFb1ta7toF0MhH/spGDdAidVjTC8/8ZII3AUhk9r43K4DmGqzaavU41XzO
FVdd8mwGF9BJ7b4UoqlFRNUVluG/CXzdFyOUeBajpufpUHyNxMt0ZUcdmx9YVcUs
CBHpH9ZSRLNTm8W48iKVyOwgR36xc23oRzJckWUQZAI+66ljhJsvM/9RGN9vHYZJ
Cj4bqWLPo+zS4jBk8c+NMyu+I04dg4lQayvG1dUWYrc9pyJkE3Wi5vbmB3TxvPMV
N7N5KrnuzwHmcVoKdjdMo/1HaLLVgtrRcCJNp7zF6WlxByllFHb3e4Mq2oufu1up
BMk0ebXtXgzsyOZYDn5jXULTjABdBOhf+ihNUGP+l7XO84jCd+btmxLaVip/BpiP
2lBBNytWmYFSstboGFPvPljMKC9aMs/MfZJ/tKTHT62NyXAXZ2XTHcMxn0c8A5PV
k3QP+XjNM8EM8lj4qJxPd4CjY7NvGAXuUerhKdD/i3eCYQUr7xyDhvLCRqTIMivw
aoJvE5yn0VWt2VhYtHRBCTy8zLSb7xbrxYL9IqX15KqnTGRGPpEcVrIODWyXiS5t
q+Bb5FzIKT4vYLt2/VHe+Wvrq38ay22esFvk7HgKrmYkJGAeSp7KPuTXUZEWLJoQ
QKpGSMHx3cn3s9B0y/I/opmfYuOH/Fa/OGknYbl5OlMWZDjL+KD0NxIwgQQHTPJO
nJk8QLZE2//lc2OySUPlO1mDfxdInR9iFYLWbTtS+3qJ2f9i0/CHAyNEa7yP2lEv
9ivdAb1b/vhkz4dG0tqWYFc+/pjTA1VSHSJp/CRzZxH3AiqEwGdJMVW1OkIpCohO
LMbV+jB4hoEwFVeOR15L1R9g90n4nqVV1yIPjtXlu4J9lJGDOnIIeVWE4mUM5C0X
RcsRgvbItaVLyXrV+Ngv5o3Ncs5jMyO1E9PoCv68bxKlxubuVDYXUJmiQI5OtYCd
YRQvd6bfAYhk8Tuc4/wDFotyrULI3B9O7KVhye/+vXukCoxXEAQRGGC7bmIAhSgb
ET7O0BRBhs8VcCFCjlZYL+fMdkYiEfKSWwCsr60FCiBal9CLS8RzCS2Wku7KRLiv
Hk+CdMVnw35h3AKJjW6qmd4+11+eLcFD28dJhQa90s373VHAqnB8sdj6j/KP9Z5U
VBpvv2RbRynE6BiSC+9ji2yQw7HrThGBk2PWB83VFxgNlcPIlU3vlls6qcPvIj76
d5coDJbVvfczRZ9j65u/tkcTlEaXnLNl/ZIkFE2hNgepFsfKT/IF1S141IpsYYdu
jhbtifb+0YIzRikacfZqQt+3QgPFCgkd8bfUowyo1ASsAVUu8s4H4cmnZIHxMLd8
5bxrvuH0k4V8eKUcn3BpKyOC6KRNK08gCZOW1ONjDWB2AxwOdUqpd6PwAi8jETvp
pYPeBOwNhYn8BxKtrTf3IHr1Rov5Xe53yFJrktm6gLEU444mMkhMctXChEPG8o9h
hx9HBaygx666BYMQCHWQ6kIVfrE79CzJ7BDHTSttpMQpc2uicKhWLPzPnTeylQ/F
TrBUiDO7IDdmW6YurcG6RGZxNcml9v4TBT7cUh43u8ic8Pt2Roz8Bh01mU3lEZWJ
COTb/O1TUuvcxGr5ikROsKYjWjbkX6A5+OZRNBSvmzvoHPBPkGWejrG5VMCOEpVP
bqwzoa8vHqfQT+dNdOnW6Uzup7d5ynDfo/rOP7U90OYQKYHA4bKLwSTb1hxxa+W/
0raGaKFGA5r5oC8G8YS2x0tXTC0ufgcx6LC8S+D5eiYzs3ckjVwlN7Ttpbz3GmVR
k6tbZg5qbaYlDKEcvT04gY/el5sHtptCP+v3hrjHBA7UsvRezCr7Za1gBWVcfqly
DfkiBcUwrAtB8HHLoqda366Ow8M4zylE/wCaiP3tcNjxEmGxItU0zw1hwrPI5jNO
Ipohcn9TKB3xR6U2CrCaH/Ehx8ppFwHJQBk1I/1uhYPSnqXgoD96uvyiND350+QO
OCXaeXnTPUJ8u27bPtMbwgmj2K0hG17FT3+qprFPsGHM02BtlDONa8sfd/vWFrOo
BJNlgUu81z/myFZt6MYV8ZwpRBD9OVlLd+MH5vMobVf4T9xEtnuiAFjPQKFJaNLy
/Iwp5jtpMCLwGIGgJWZuhd0YePnvnZvziqlUBiGGrgIUaGzFKXxHRejHUdyVYb/q
s40xyj95Nxhc+nG0AAisLdeF1ufR+aT2CGNg/MI6/KJNJxHxI9BI/QsArpRIqQ2b
tnvh5B3EO0qCPBawAQxyN1Zrm18xUA2b5T4gVHvOOrMls9myzlzxLRXI3CCkgGpe
6uoITEjWlye6eDRU+P6Pz4kEPXB9AKywOdxOPE7I/tEJmUr7kOrKAHQmKJgH1kmB
kZbmSe8oH0QCrXmsDiKCZ1JexIqqq5JSaPQ+GyQyKjnour+DwZNMgMtnEbhkwazi
uGy/cHuu5u+3IHSffhVte1xaugMBov4WvcHxYcB5WNbhyxcXu9EaE4KjwzmDhT2q
bnJOVHS5taMW6mDJFwzRwX1vpUQnO3H0Sj3eYrS5FCNocYnrGV/r1Vdr1OX8xqd2
jixUtHgNOCom1lWMultztsFJkr7JAQwl723LNXVGYERH+Xmtn3T57ZDJ5MjWdctt
n+0zeFbGmbaeyuF0I6Dsg+THGXSvLwhTFBOY98kKcs3hn6cJ1TQhgy0QFPVQMJH+
4Iz2t/ZsveFLsF63wWgWH26Gs03QzuR4s/Gub/9/c7wpPfylbzY75qv5C3yjmaTW
wtvX8eFSRwBg41xYMM+fK+6v1n3Qc3ZdesbSekUNGYFUj04GMff6qCImh0210kZF
wOaxoJ7CCfqyJdMDVH2VD8a6OO1FBL5/1dmIfiFCJ+CUmbnNIpTneVIlnII9r45K
o+sCtHfA4cXi9SgupxkMajU1GRb+Gp/rcZ2XBr2dtlsCwZpAb0ANgB8aR9Yi0XoG
JXw42izj2zNnPwOs0X+SNbG/uv+ZPwJ7HwWxr/RdepQczlj/A9fZznFiqRjF8SNL
U6Vxl7HToyVAjFY1Q0M5NRJco2ONwzKs9Bm3ECI2TFrK5czTUYgS/PQ3mcDl7K01
1uwl0EO+Gs3UyNewzRc/zR8bVXqspL/c+LsRKuiQ758U1YXis5jATSVQU7rac8Z4
gMX0rhhbGFY9XsuGlVjK/ZsxfAfX3pV+XHML58EYVCUcnmyBPz+Bowdf3T6Fwqkj
eHH5so3dJJuaMqubP5WAszVlYKgqhRtdlXVhms4ZSoCToq+UHTSH0SsJrRQMo+3s
wT44mIYJVmSbteKNNadrEMed6oqSA7K2wsA5iUa4oT+QuQXqR1B3LqvWRsB00AAT
FhtmtlWplZ2DvKTonWWeVL6FhiK98F3MdsXg/doesdh37UEzqHpeTrdAeWvUHI/w
QIdPans8iwJsZruk1rUzgzgz5lqww9vDUjJmj4YdBD3aCkx0yT/XY6Im2pLYZD5H
g4PBoPZpJDWiG38EsrxsNEk+T2w9VvXab5IJ8U9lo6IpUcP7CS+CvAJc1zZgmTsn
+N0xruPimw7fhwoj/kpR37OQuw6Yn94z/ielq2F0kwfIxAbU2KL5YlaTUXu4lgRP
1B3zjIqQ0hQ1fmb904gekTw7b1Hv579r6gA85zXXHex3qsgA+smFVyj5jG22cVjG
BKkkHKCumywSifMKiESumSL7VIePHFwWofjXoijSx7UHcVOZtyPuj9IrPfER/PD1
AlPZGePcDxlOX4Vqg9ayksOcxegNkt1KvE092Lmo21bUFXD7N+u9R5wBYK1EdB4J
8d9bjO25leLdwQN4rokzWpm8MwPKONVbYs16XkWWb9GcN2pOzvSUDG5b+zHVR1qW
ynJTIK6p0ylwwzwStw7oQgdkdLXhf9JwNDcUKZVKejO5DKUvmZeyo5qqJtkHivs5
St9UJvGywFBQbqPb8l4iuEb1J2vqltCfCBpnFG1ct6zLn/5fBmL+XkATJzNLOJi/
fd0xZm0VKAoAq08PiPVQVVlKeoXHNsmLGZ2Y2Hkm0285EHCwKpxpS8zTT0/YG3Wb
VI9IsdLxKuzYNZLK6qqJ17GOF9rmnZ0RT8UDo0CgqWXkK9JvDGIf+cYCkonVb/Mb
uLuAYxXDmSK7nNPcTkxkmI+w+VP5I9LQzDfHSnz7X9Eq0W4/FZTfgAIMC2GZHk4T
DLy15wycMxCWw+Cde1Ywbye3tFBCFokySUJsnAB8QVC9W+Am01SZxaJ+QZoM0etl
4jpQmKClvSJAazHQwc3smwnuetQqpVBjzS77gn9PpGX5J6hADzNs2bqvnxmK4QuA
79ZF8Jzd6xczUkWF4eV2s7QWhr7IUW2MbENZ3yPTJPv9X+cqFsqI+F8DrZCUiRQ/
tph3JUXZLPtVeBBaHreolA2VD617WhyvHR4MvMwwz9DiLwQJQUA6awmmOiQuuDyN
e7VGZui14MTN+4JzcAcq95iY7bmDQECMtnhJbFn205w41gBIiNsOI4h48FGVy8QV
T8WjRM5tyii0BaLvWNdRbeB/Aax+hT08H3D6v0bAklr9RwOyyzrKDTRgAX/+s91o
3trb9djvpWSkctowDe9LTZGkt6eCTT7uWYK3mqx/SOi97WdnS06hr5bBbiXNZCyF
iJ3ZZmSekYYIzdqHkPFhoNhUxncbkkav13xFiKikDjJU1VuOWoX4iFF28+nchR17
HC0KpXqWCbfPVWUFHxcBInx7KpZ5IA8yw+yVr5eu0xx6ykmLHN7DgXFokQygBYBZ
zGPQK0RmBxG93kwfAlnuBRaFRbY5vBU5NGNYA/+y1OnEAgK+5QFv5tEfX+Zgv/nn
H9oJjpQB6WWhm/IL7Sf5vk9OcMKRhAQcOCEb5UVn/4GhnQSrp8vadMuMNn+aouXV
MF4x7dcXqAbmyEt0jHnn/r0cBo8Vm4ansEOtsdL1YRlqLGBya4c6O108aAsDb+A5
ENjNgd3JKLTw+iTy5F5SNzDvAztvV3dVOSp3vG7Jl8S/EW47J5XzpGrczGrMOXse
dTkUAIdZgX3/mNtUZJM9Rr/ffvMhwpRhOYlTElPi1PWTf+6KKs0ogofmWYTBbcSg
EXZrDNX9OBUESE6Dkljg3QwNiZ0PznJz7z+wC3+fVC5Ih6vp1PMN4/XBbe5dHQWq
IwMOHJ1lQBqQ5sCHVnLPyIZzj1xAAdqoKrhfa7sPXOBO2HP1emPecMtSxkvG4PmM
2+yMvPUXC1XiyCUv5dZmNd3FXleBzLuWkMm/JuJJFLqLhApdDk1x50tpLNUoQO+J
3oZ2Gx/cZkHpXavPB2y/Y4aSOOcZQ1tpD3jx/P1NMP7Wd0iJpv8M0sZloJvQVnzT
aYZpOYjFMoLxyxYqkA0hQIZkOHMfmC+ZaiUekpsd8vhPQ4yw6vwFcgpNBC63ReZz
xqiyVXedTgPhHW5FnOGTGDwEcRSl5x8RPhVjbM6u6OX9KjeRUujwXCRmZvOsobb4
nZS7e7/NwgRDamW05o9LdpWiykCqvSRiPL5zl0y8egYMK1H/zpn14qvJcjvK2GXP
aMY/547TX6D6sfJVmCwPzM1jN7ajo77LrpGQaD7rhkmWJW0OE+j3POpDbiGEtBMK
eygUJDwI7rcTQtfQVQSMuhxoivL1R1CqEcmIA1aaNzuqFsq1dTp2C3WrssvE76Z7
o/1j+dC28/s1T2MsrjjRCs6G4ItHc100SWcsJCn+ouMciTkGVLPGHDkp90XkG6w+
VXIBNqqYjIAaoPQS0Qv5wRaOKdX+666AkF5Ly6MBmeet8M+GPSAuhh6acphAVFSg
uwCCNe3hzvr51NXSecWcg2D4IBld3NVwf/N2Hjs+We42bMShvNfGyvJ6P5D9yIEK
5Y2C/IHTQXWHwhl/ze97lGbzJ9fQvIfQTXa97FwPBfWU5si9jNRUWZywWEgxpqMG
UBjhSyUlxX91ucMQ0dGXy/FGmmYqIDs/unSpknLZsAvwI3kkWnQta8cVr1Fc6Yr6
fIwLe2+mz3xndBWNBvr4DFXCzZwbqRffZKGthBMiTqBBuxJkI7p1F0ZZ1+2acTTq
aiGWrJvk7L3tmwKtFZDNaXHdqjnQlCS2doBsdAZ3oLGEovSgoEu8klylPExGNLw+
L8n1hiAWlYqY6dmuawMUlHAitIOmTKtx8DxMMcdzr+CDFCftyH9rK4w0m7pBdEhi
BBLusgQmYjUxp4NkZzhciNGxmQ5ha7zRSD0J+Iu12oorgP2XZtKXFZjJ6L2gss+S
NwwbXcycK374ZsRQRgQXGxPLj09aQLnbgQI8/3TSlBKr+Bm/iOYidp79SjSEw38w
BqmPd6bjZJNvjkbsdO7uS296elH31F8Nn/q+qi84WpXlCXfMXTd0DcKdNwLn2urp
Ur7lwnxQMMAPjZ+IRIn7aiiQqJHy75/8/NIQ8ajvNhAS2bqNbVtadE8Hn+AxInru
hNinugePlcT2GFMu5HCA84phAJFSaFmyYCmTCdEhu95CvIc23PQbhpSoPyqY+1u1
zlKMZNqW4JZy1gmaPmgXD2GMIddIY8E0ql8sDtm9Sh+MRTsj4C6iF7enOQSIk6FK
zX+SZyykwc1NSUcea3wfIli6um7Mw8g/GdJIOt/mPc/oUr0KdST41agZOgh3zRLQ
JtBHwjfBXP+R4SI4+U2slXjUeMd9vFYzAjQRt4+sZoSzeoD7tGBF7VSrkU24qFmv
2dfPUfnOxtXyh9PLOP0JGRLPTMxx04Ab+mXzYBpUZaI9Aedl7FUmx45dw5NGVcVV
O6SpgLkAQnWB57fhj9YiTkbzJlIogNYxaXzslKzZW5t/dq1qe9+tFOqTVsDaAWCf
fgEUfZXziCsy6dGibeNLgoUTlgZS1aL+KdihgouHejx41+VV0OozBFXegfT7PUJT
Q2dsdM41vg6i5rImzAn3T5o7g11flRSaMzOXMv6dPVICXSm3AuqpfPPYTR/vc8ll
yXkcHN95yDUI56oODMRBgP4Tgj0H+jTEMYcwZeSelBGQoZrQ29lKDPULXG90rcj2
iB1d2e4VJ8jP0njtff1qh7hxnUn1hNgneaBnxHHEj0JZMc1qQ0McL7nzi3wID6+p
gDeuWwVn5LbIN+2EJxz8TqROz2+ldqPtxqfjmKNQj6maH6k4q8waSqiTu8UtYbVm
NctpLwpDUPx9+iGr3GYDKc640Kf429JoJGicf3bSbtpc9b9xOMrRziJOLEzLNqsl
SgWVIUmN5SbUwKxEaQvNcwP8bFJZ1S2qQBvEtwBViB7gAD3NfOsDlGl5w1tZ+e1h
N3fTGWXYearzWILQNbx1JNylf2pZe+rALhCAqrP3kiqyIP0JX75D/j7ud9hTO9Cr
TOPpB/z2wEAU57uIrdiSzgetyLN/aQYdutuV9JUt4l6Bospcg5eJ4YOWv8IPgz4E
lkbtrvFtKKd/t75t+J15HGRG2apRehWNG3LtTgsyZkKFeOlofcN/44+eRsB/kRNS
zKeyE6OKuZpcyj6yQafAv1t8s9QQQhloV5Jb7CV4Y2xhyNFTn54+Lwlt0r4jmCdl
rEh7joLlTIFwRrMeyh7OMrCgO025l9vm09ryf6XG2Ao4TudMa2ee0RCsK4pQFV59
ePyom0ulO/RlI+1xnxsR1nbQcGacNz46b1ik+hIHVTTrILTvWbEGPJEJ0KSHW51p
Tlch2AzeAJrWMqveZpkyn3G+gfeSZ2+/4zVIXiILVNXZDQUdz4FOoM701XyhdiGJ
HyZ7BMco61FOFrZ7f8AAEETQ4QStSXP+Xg2av83jGEn7Q9oQm/ntL67Px/E+FsbG
0TTpezpaIRGyBdWgXgeHHX2CYuyiTi/W35PNFLWRimUD7GILlCnIAQxXgiajyA8J
jhHzFWYkJ9lc5yD3JelVRk3xacrUW079gGS9xETUA/CFROzTyjpmTihP6pTmcl4u
z9X5cJ6ckIyf1w6JuZbPMOX6MugH6D2WJZYPWB6Xaf+GVQWG57aHTnuOzOjHxNOv
KWJhR2OC+v7XdLfau8k0GJqqUOT8kXS5XKlTqatX4wWLUPTqmhp/tfxPQtBShAJl
JY0arK0VMl1U7D83Px9uvPX3js2DheCfrqStlrxtW2+cT23IlDzxkNNKrAy7bK2Y
UvwPKxlHP60DsNMTQE93ESqsFnijjTRXPHg1st3EqbqDpw6vHvZEdKTWSerDkLdo
noF3asjFkVHwa/SIYoo0Y0dPWWouC/07S6XvHu5zVeaNV11dRmtt0NljgYaVkxII
BMxE+2L52ei9YaZwvmMev4jlx1S4tvosfY0bGWALVslzsP0Xo186+VrKUq9xGZu6
pHfP58XJ+y2dsNb8fD44S6Rj7Rg+Ya0akgJgXRIZ0UeL6M8wKOfw48Vcu9vqUbaX
m/hxQQyFvUZxAqAfgHJkvp+y2v5qicgeL+q/b9DV3h0FDO47BUb6v5KHnd+nc/yE
70bKzkgWaqItRbptJaQjua3Voi53YO6n8dGmYDHeWb87pAObbieEK/ztFi4lrbF8
S8v3gme9FzuuRwm/+AhlorOlwX5t5MWNu1e1UUVm9INHsNPmR5wZEzovASejdHoO
fWrROBgcTRuP12GlVpR0NVI+3GlodlL6wn96xtsiyysYNhilOz86Y/bf2wVjHOsL
CWEADcffiiCmiM2ks6Wq3TwQxLJHut9XEt2GAHA//EXdznyNksMdmPqqoOX1pCgZ
h6fB58sEnwowZ2NfDgamPuwr0KiszATHgqMb76dSWbYlmp0oglJA4Qsi0kyMyiZA
6Wvlgbsq6G/CeRmLtYaj+Y7iOUF3X9QHdOQG9m4PtSan5+tO9/bSSRIY921bH9mk
FgdWewjkcEwT73DXsH8CsDu9/GsBWAsQ+ZdwElaXi4WSLMosf2onutQwVRCXAB2b
pB/V8WBxJJt8RNcajXXnBKJUR8Uond5ye/1QxiDpA8QFNmXrgDEipBmO05ZbzaVc
BJKudMNKrsgEeyGN7wgs+q1+yYhXapEVi9gSuwcXUo80ZCT8olHCVFpkZT4aEO9b
sLKDJM3bk3eiZM8Veb+ifzFkITepS098rmBz83xkLw0zW5A2/fEdhLBv4spP6Vad
wHpzAD8/YuMHDTTK4DApngBUdsp8qSzP8isbNBOIvZUg7g1iubq+X6ZqjU0zT3+p
5gqTfCdMfliccrgcJciG4TeqsYA/QqulNzpAoxtvJhFLTRfV/7BEPctdT2Ua6mEp
neRbjB8fzyoRWC3qbN/zaT7VQh1B9DwhM784XtzhUPUWM+moOsr0+wsKlPoOyrPv
zRbFktuT28eJNYYeIo8RhLPsTyKUdZX+3V3QlTK1fa+JtPjJ56LpfnR8Qii1ECzc
9lVGtuj1pD+T3h9U+opstUs4uXmMocGLtDGQ2jrmEmdtOySfmi5mSrZKqGImwcxg
YI6jSi1YI10Cen2SkjbCnDP8BYWMApIsPsNavrTJrzIm52z4mgDNvAe4MBlAn9E1
I4mNPMTQqRRW9NftVaqQR+v3v4qixDYj8dt6WGnmSd9FTffElzFaSesV0rPuO5KF
rwojQB6/LIIAoSWUSzdJrkK33JipYkR57Um3fSGmD1QnbcoDKlEzSdMMKX3szDD2
wxGGL71mB6fCjoaPy2r1zOsx1YCkPT7Blu32/mW+tjSsfDIpt/TLef5Q5D1tvTiw
o61J4FyrVPNf+kMZHjSegbYJRtEr7pzY1XfOJjeJ6JYjsP9PHpQiwIAOj3NZlCVK
kQbk+Z6JT9vCJkG9LJDu/1eCSoWVx1Zvuw8BfUnSBvcRbFriIBElYY8Hp2pAJBOE
Mor3pqme5VxsVv8HYxyrGA5NsvYr6qtkh7xZTQ9GCC3n/887MIcxyy+4exeXuj1P
61kDp8uLUPSCu26WcoupufmWgFSvhfQYBrPvPz6KZeAr6ek7imBRV4UMktJHoLrk
TOKz7HuyLFYRGx/8jXWwn4/319iM3+VxgmkA9ubvPaXrF3cBI6wX/qR48tfZdUkK
JiCGKOV2KQ9uMGABEfdtzyqe5HabsfzfM22bgrWsT/Kobz1E4aawrcJ7ousxOTW9
fcND7wCxPhlsj9P0GbhQQHWVuBi61yb9m/BMFf8habxUsiKFCGj24kkG9dbcoMl1
w8XQ/y3hcEtkc+elhEI+J5Z7vK83jNUchI3AHy6DrEBwojNU6H98VcmRFqkwXOV5
Ww6vV7VSXQ+A2fiRzwoxHHzBycnWP2c2R9/zGiBUK5o5J8IMGPxG/43joV7a176k
9qDtWDXSBmm3evCD5OJEEg7/KZrJCqwt6U5mwWQbsElK1wP7uQEYM2mClZWECQs/
8HUW86NKPEMJ5OsGQfRGx5+ZOLdX5E9cVh3k4cuwgGxW9sZVSlbKPJgFaVLMG1MK
+3YKhu40ymf0EBMae5i2RYELWfEsccTak8V3oqzN64O2CRmJWnp9fHOUvS5PUPEY
hiHy7KMWNmHhsVXydX04em7S0SkdcDjnVkdiC3TtPnQEG8ApkKxbQ20O2KaEoJc4
fjea0ez47Hy09cp7VtV0A9PNaIBWo4MukQvE81wDD5Wp2A0Lg4TPgZAmwGeca572
nfbhvgFyaoxiyCdN9PBj/jXMGhh7K5eIecNrnjm5tWlm5PJ9PiMQsoCywnDLX7cQ
2nrplVfCbgiYNOVQupcnzajpfVRP4ZB1ZS+P+UibDmJf2QJNWktjWgrrGA+e1WWC
7ZhMReg3pMrjN7UL4t6SCuKRZGsquXgacB74Yb0koMzPo/8fVHqpQRBmJfVFwJbA
NI9oj28fPicI/41Uz4sSC3pAm21AVLlGa9qPn13cTMUXqq3VoGxFzCTeG1aYnkFR
7yraNqq5tJXzzHMznbIdZfepFn8e4Hh6syo/MvrL3NjqBrIw26W2SGFU+WTuE39y
88OOoI0GSnQhJrDPs4QWIbdme3j4bqpf5dX08Pj0G5oV2gYvaX0kXJu9hC//eegz
r+mnoibTrDBW6PSdzQvNPSrltNTABrpmD5d329N3TkHOf0u4aCQkkZSgHusNETpJ
eF1NBvacsbo4oWveacr3qfL5iEj+VOFrNK5/mITQL7QViF4u/91Wzs/HkfWPvsmw
CMLrAG1gV0UvTcduTGVD87K7+mgDKw6WMswZZJvYpSNBmXz+1EYk2It6nR+R0x8N
pb6m2NyMr9fL3Zd11iglVwyku7j/wJym8ktcAxH15e/UAyZEvGJ7bejenfuD0ZaS
7Z2GOlxjCOtPVY0BF5D0cBxycKd7SMTyylOHyKNZPVd3gEgcvvJadxvGs4QaPdtr
MGfxT9a082CqAiZXm7enEDWehmWnf13MM5CN4tpsuzyPiuOLhMTx3Zawn/iz900u
Q41jRbv6uucXcMjmX8kNjumaPQq91dCj0T7mHov7S1NB4A4w27bzSg6we6TMZaYh
Pv3vjyY9WeEUDngQnHJgwMO82bJy8rD9hw6ZgeVyvzhD5jlFh2GgxHwZfSrYS5nk
COS7b1bJQSNS9gsn6p3n00REMP5YtDPrY1J7mjxvK+E+vCszplKLi/NI1QaDpA+n
5nnlBEaDB8aR683IL0hl0nxeclTvY8RkReX5APD4hgg5vTylV17tBvMCbZqNbJc3
2JcLADmdsJ+4rBmjlBE+6ViNrZayGTrCo7kLNvrNR98FzUODQ6fdCZt3T58CbJ7K
zsV/pouqdAvpQmk9ZaAdRrpbmutJ/TVZqPqf3fyt6xD9cVS7Z6f9Is4x1SwurVsj
XZUr1a0kHYp5E9fN9K8ZWcfmOxeZKTj3ibFcvu1W9ZHUOalAtsrHo16hDGEnlL62
I/OJjg3THINSu+8RwTjwqkX7BFOobLlmWfiNWRsILPMcCZ5TamlHpb2u8nRQi7Ru
pH0L13V7m3EDvGadRT893tD/53nptTwmKFN8Ha7nBJEQPzgN31BG57+BaGmkMkgX
nRZtTITBvK1NFJnc0WbjSbb2oT+v4WSOZjlt6wDJOVaiQdmqD4LDf/20CYRaObb9
5Rjs/t3XdDsDg/K9lgX92UfsaYaTRl2DmZL/BhXKmtfsVgpKkjpAxWnzQMABUuyk
meQjJZdQkWRdflPt9Ev2r6p1qFTE5Zrg2I47baOzldUSlOa7uF/LI7AGqwIMgRkZ
MOQZakmMyPnSL4dJHlxeYdYbdrK39+X3c+L/tzDdrbq/ZdrlQ1pjAGPkqgC6jqY+
b5ZF1/YEMN1zfoKIg4OfD7oc9CVhJA4PVRP0Lkbl0xHJ9Urzfrpy8zhEUnhefSlO
a8ghHGxdoW8078rxeaZ9Eg7dp9UQyzjx4qkgxdNTpPGfpF0pInIEBAo7fDAi+msz
HdyBC5HaqD7+c+EPt627jNj7AMpYVoZsCH+wXxqGAj1N4fjTCczaOdQlX3awUrdQ
SgbHBHuBCeyyCLioft6b0ZqlWYHEzciGEZ8PhfJGWY+yVt6cjFut+q2PdNWX4n4t
Q0S8DwxbYmVygUn2UMUdlLm0uj8YKitSIRxbf9+CKmteETydvk8Gm3lHfpwj5QYU
O1uqZkLQk8Yp05YBWXrN8Bxi00+b5ma7Aj+K6h+FQBlm2PRi/ez+h6irR8lXZh7K
EAiLnUqCTMADrkkNoWm60fZLhBwIquCotiTmXmKlPeIpR15xls89T7yDiqQeEZPP
2hrjtpbtiYu9OniBYOdh1GbQvUXeLwGNMRr8HTWrRsp8I3pXU2H6nKuApW7WWTDZ
wuKpyMfyaqYPb292/o8+FLIYRtp6LqCe0JJFZEWp0rvmZtO761iTMZ4SbnOx3aef
enaUrGWWfGG6fCBaFVT8ZFVZ15RHtchAgGfeqIAsuBX1KeA9r7itSV5rcCPcT2iV
yXxlR7fnUXP/VcsEvrkqsU0n0UHssJ/ow62ENqFHIsilwfXepMmgX+2hX3CFolaW
ZbKImp8SeaO3DD7kLujYeMTidac6klXazCFs8wHLCXqYjkhkv7wc/bN6lKdPLfBW
+M+gT8B8PEK79OkzqxR0qgFBqVdWO+wGGvBBO7AIbW7CfGKRtYqZ79BqXJOK40mZ
WZcC2XcCN+HzjsSFU+4qKcPn0/cw7sm6QbQ7Mfa8Q/ni9nTqwftHSfpDI7iSQpy2
u7Ol5Z6qheHJj751Fo42dvtg1boE0ne6xWGkfUoa51phlqqUbkgG7P6XMTa9KCAW
rY1+eKMobIgzPnmoZD6jANsWY5m/qqARkhueeaDrQb7i/X609vOUXP+KIXYD7lwX
8K16X2gls8XNkHMj4pO929RU6T/2fTiSad98syHhWPNlaQBzKnEf/843AmjF++83
74hl4HhSuzDdJ6uhjjYL8i3QqBmCzRhsfY2qSAJyCodvE0YzmP1+LG3ugYhEZRA7
MDTY4/YA+dqt4GHoeIcVHjx+KJoSDW6rN9qTIM2+kdqR+kN86ztFjOXx2qMrMwfC
D7C4bjeY8MaG3/92php0YcXdwFCzZjoNU8UMN43/7TYvmcANyj46ZxryhpPjjc57
+57ihg2z6TcE4NUux2Ovn+mnGFCUh2KKBfZWGFR42z7bEQ/ubGPPpClnLQLxNQQP
s8vquw7pi92QnxvnC+tSlb6+OgVlH1uzBw2gB4r2/expVw+sBSda2DTHi8lgQxVw
rh4QJq+Z1u8t95/CuHG2mU0DaTj0gZvM4x6NII2TE+b5RbY3/dUCaZIP2wnWNPPU
te1aUZn+LyajDdrqd3A0vYbk5kFryuEs73NNubaafnM9tPZaj/wv+tZ9LRN7Ewzg
gAi20QN30D7cmWwVsnUwKm76IDgPt5B5zB4DRVXLqR8AABhD1s8sisAuduv0vv6H
Pw0hYcpsDO7Tcgxz3yx87lJLdE3r1Xx5ViLRBSRUV291qyRXUdz95byxi44/QKPM
2WidVCPJmNPGPfn7n6httCSi+QaE6PAkdQOb6H/hKGSoxLrKD1ZE5w8RxuJbZjLI
99yDw51eXuw/MhQlLxMmnb1s5KNujzAxsRERB4el1w5xea+pi60duHc4Ru2iacLj
9x4AnJ7C+N451lN7jDfhDkC+e5vaqpXK7K+IWp6JM3msnB5do7zClRtG6Ulw2eqz
Fot6n/WSV8Xn79SmHtIjx8F/mi7/ldTHjrRe4hPFnYqjFJQZq26cEeh77LhBC5cb
VnDrkHmKccVCooifrCw7JJQJJ/AoYmtocbzPVZ1Yc0F/X+5QO4276OV7il0Fz7AC
FBPhGnUQ1fob3zh3E3aZ3Eo8S5Of6QlvgVMCJa9S3GoF02bpuqWECoJlLPtlQCTq
Oh/L3wiVaz/9BjXcOG7k9hgAWtJudj0O+eghlI9i0pKpTf0Mysbpi4Qr11f7n4LW
m6mX6qnBdicWWn4c95ER+TQtc4xE9lknIFg5sLzNpHSTaWMwxXWwhRg29Z1ROQB7
7aUTtWBXSvtYnE2bIP/RCik66/HpEVGE/BhrHYiyPQ4aj1FDesiP9QmMT1K/y2Vo
CULzHbBR/Y1dVRarkw28RfKdsJietSHvcLtxeFosRiI6xXNRrAJGRnpuWIWlCCUv
ivP7pboFTcDy2S/uvsyiOoWTe59k+ED56B5h1ZLHj/EalXzsQQkwHIc5qpzmsw0W
ToDRoh7cMKHVeuKgErtXvhueDXRiY8WncC5/zXq/D1nBzM2mBdnS2+TpfJGFE3+A
FyFLSzS+o/ijVGkOZtUFRlUAIiZJQ+6y++eXlGaZ667Fo590sDh8x9nZ1Q4Gk4S/
57QDCW09Ercz0luubSgdTUS1Hk2LEokJezQBYFu0fKMij7DFbQ4zZw7krWYJ3Iwz
mmpMrmKbsQlWtlDBbl0TtZHmqwlESd/mp/WwdoKgxLicNES+c3BAv2G2Wza6pbCK
PnZh2BJ99PW30E++PkM7BQc9bc6NNVhJ87ie/1pkEqSjEWo79cC7Crr970/68bk6
tru/hg5ES5yxB7lzAO6fVe8T4nuReSe34UatHFV1bnbXfFjqr/+MCK8foXGuxt2a
UUJx9tg70lVFFMl+5OWtbLeO1P55IP85g9u6M+m4fIT8+cMUolwZj39Iid4st+Z7
ZBG6r9NlLrPX2gR9I0PeXLjvfa8vCcyHN3PqXKjywjOQEn/aivbsxZd/pDh1V5uR
/VvAqrjKytUrXbQQhy1COt5f4shH+ALmuRQDx0wEZhbaFrxOfsVANNYIZ2DlB9nd
ZirAXnu7ovi6hY3ioGe8W108LxELMWYb9tGKf6xydnVOgzuo9mb4ssa9bdDUVLnR
97O8JMqQPxfenUqlsbymHnHVZx7Lg8pZyHE03UCQYflKzPJ5hsVP7WnPzZ7D4kir
MbHv5FzK0oLGCUZ8A1IqvUhmJtey8KTVLpkERrpvp/eqW8RMjbd1MLw5I7VmlaD8
zu07YAwy/1a2vhoFTghMfhpxzdlk7vtp8kHsB2SlH0irLci61fHzpmWIZ3qF8sJb
OeRLtf8nEu6Nhc5GgmClaXOOlo1ahVbgzbxKRfP1YZG1fYLxDLLmwsflyRdj1dSY
ttaE/0kz1jBoJBAY6ICd6C5PIzmZQiHcgoO5/WRg1gRPKMy9rSI84lRVs7iEr3ji
DEAdts+8E3rLYVb+wEFyeIf59roZBOH+RiONcT35+9jWmRQCdO4FDlItGLNuna6i
VzwKI71XY9jVnhqx4Vv+u/OXGCPo9A0j2urz/bUVpRJDPT5uwS8ipJ6EtWr0SjVc
xJgnIj0cREC5yw8GehUL62nc4LpjoVfiklsf5veiee3Gv6N2grnVOeBRIetrE9mz
rMUbH6DYV5HdlBzbr/TACH4ouvCqL/djWvDWQWo2BKAAC1cFWQx9qyqMj8f3RjlJ
k0rguHxELn96C2l9SOl/rNSTJv2CxaghNq8qnKevlXMp8gJdX3PqAW0JaxN0VNmF
zS/95L+Hix5tbaHewgeg0wfGss/sySTOqOdkWE2aI6e5Rgq0BA2kBZ1jZA06l9uV
clFVnKdHL5SZ/CoQPpBP+3safxjcmnTX+uZ8g5Qs/kRrLM1UjLx/67yFr0Ks62sM
fa1AA1bdNvjWNhrsXTVpBox+gH2jLb6iyjcdKcUY++QXXD0HMHHszcsUky2/CsYz
YLyBDwuNWZSqu0MZrTE6Z/Cp+Xk2TZgcz4nslwNhzmwlpcm/zyrm+qneCOeo7o8k
BgVruPb0dtRDuxNVH0gkHgvIIA9g236/80zHC/YKgIhKeJ8BaaZ0tRMz+kafMQUu
JysO6CUPNMmluFDt14I1z/JLd5oYLabdTtVqolfbCqR4tERehboHDiYrLzG/rAWS
GF9JIBuAd2B9mD92WJMZSSi2piLw5ibIfg9IS8N7ktpGdlJ2tJJVgz+7XUDzIhai
HQGxo6c8eefdUknygVxNq3VA07aepZ19oM9rsf2BzjCKF7Q3MWz8qr3AZADcYHYA
ui3UhyL5mmi3h+lSU8UBcA9dk6sGtbnVpRgCx2XNIxM0imERJwoCeT2p3HG421Ds
h4dRgceV3hHTE+c+nFkqyYf0hb1kESpOmns8sAHyfNjUNpfeK9i6ehqLNC5e6rli
JMLUfn7QbQP5AonCPsJQTszkmCqO5YAYDoOwlrGKVF5WsGmTsphWSgB4nepWoSi0
6mh5sCSacC7A1uMIzoQvgldTPYNmVkIGw/JrOd3jMoUosr3WGKSUiyZhX/lxKIsT
CNAtYAL5Xq1IFbPabdn0/T1ECLwiNJcWVPK4ZNR7cY32/N0cRVoMN0X3QX3AifnA
AB/Q8OzFfW4PsCOwWypGxEsQKHwtyIJvddTAEfJ6qPO/zSh0pwsKC8B7dOjBX8f1
XD2UShxRWUOBgdvcntbPPwI+DUg+GSo+xfS7wfL7sVaChPkhbRmeLb+R5qOUlb/K
JqCkN0KGoYEmmXOc+K5vJ9254C9Iyy7z4aI0ruGDkJYyzXHXd77AByuIeV4AEy2W
a0PbGRzwu9TljjjS9Sfh9l/3cSiiziqzkuOgireV7Ir33ihbS47jikPLFELV0gCh
OwCIUU+uFAW9oOvJoMGNDGPQPP30pgUIn3igT+In17UfZeLwYBgW+/Qjn6peNp85
XkZtgFlQd3SgI4bgs8dYIqjWoZ01zv32E6Mn0OEioLHQjXkSG/bfMMaH0XudNotK
6lVmSNN8KfaINuIDwnYb2rkA50C51eXSqCtq2WzM+vg3UpS/ONiAyQ9NrUe3WuD8
THt6nB+m0xqux0XTnAS3F/VOG7fhPB9joZPALukQ8NNhkEArYuIfsy1/VD6Brl/w
Jbd0Dz8/O/ftFODMv+rEhilwXNRVROJ2Z/Ij4GhyKs/g66ERCcQjuNAWPw3DeFKh
7g2LM7cw8YE/m7tDWc/pPXG0NtEdkhRvX53Zju1FB+AiBxB884xURX8av8wLapEn
4Adz6Z6jGF1nZu4V6YqEnUWudsn2WX/tu+KwqyBKZ/ElZCXmX7K8z8QYC0QQNAKe
hQHnRbzKBL4hefnTnMqyrNQYzLkWQwGDUmNddILAlPQU+1hjr+FQVID2n2MRxPVu
FE9EmGzkTZ+FNgMfPKSOwCuGabwyR/lXAIqGT7JNDIS6CwTMIgDqRcmgGRq+jic8
tLNJEvVy9BCTCPfIaqZpYrbVFR4am+0L1HRiyzZQpFn89az76gk66SM6bZhB7R40
3r2gEjPeD29DkRcVBQRCIXICA0oEkK0POdzLSkzD49pkj/urepDG7uJL8OQnz03n
FSysEIIdcIWV1rVFE3W4z0fBS2fjAGKwfl9tjN1589PnkUE1y6qjTH2MgljM9Dc3
zHWftwDATuN3w1A8vtDVMqxETD235oUUaAvqyq9kE7IJVUaTxejbvzvYI3AhPgmc
ld7jbgYyPXoE7yOV7/qm6/wHIlmSJ61JM59qj4UM+3z5oS5UhbZop3EeXwfGupxy
5L1esBbDAFQgpZetZM1vWj8Nk0T/upq/O6uDU1pj4bGcc77TqsG/HjMsN/lKL+P/
GbX39RFw1MLkn/+UE4BjpkEQjSDzkuVIa2guyWep/6dgdV6D/r5Ih8saxbzgYVXx
6myuxIt6tOqlgOBTgIk9PohXBf9+srU++rkHZeDkl9jT7bvzLX9D4mHlS7kyIy1a
QTcRbzUnrdB92jZhbUTXvCRv1r456hrMGLFeOe9lZor/hB3+L+bSFqIh+BSE5y/d
0ol8HJWXaQn4u9pubI9K20yyaqtBYTN00uruXNoU4ZpbspuVswh1vDf3MX+vdi92
1gddbmYbiF88nF+VvFJFct/tKQ6hi04SejvWovXz2zQY2zWCMAEpZgOMMG0y6EzQ
U99j/j0p1//h0kDSPm1oufge3AcQWZ8Ql+H9mnYZNhwjgN7khgbvx/THaxo0if1v
Jgqq3PxYvPPB8lD7JKMYpuh4xmYaCwdLb/5rHuMtwyDL59jVd0zqFA6ipEZlSTET
B3UUNN1uTnSkpFxSdqk2EHau9hyQbT+BEFy3R0lejTqQhsc/pltAZTTW6YDmgiiV
vLgluGXJIUMUQZyC4HzG83nU3go6whi8Nm46faqnOQtwj/gDiEUOzQjE6nltvkUk
wE9t3vQvRabwC8ZK83jbQ59uhULyWjRAhETzGiGeFoRE74T393mztQu2LRMZC5KB
YQV2yE9clQCkjf9cMqO24i1tWVOI4uy6cIjqaIDmGEPqkDQMCcfrqS3P4e8qe9dI
z4xoAMc+cgnefCFBPJCC2L3WcHZEMVmtp1HDw6GjKpchVVbbcitL1PrFgOf/wYMA
M+B60Z4Ds9oNz2cKQJxfFr5BfC7tHp6dmrEgyAhPrhYOm3sJHQB3u1dCoMGYlodT
Nql6L4rhuU638yA+nFRCb+h5cIMRaxNECuS72dD1I5bz/J/w/aE9z6geJv3ictWy
AqQ60Nb2xDxzRa0wGoCKjmtgLHbqc9hiXzWC3EFbSQ34DVxBjzRhNMWFN92VHzBI
8Z3zY1KMuAJvvBc2KgaFLlVlePTAw5EelOARqLhrbEFr2/iEtpGXGjWSS06lgfFW
kDdJg5UosdyqARP/+uf5Zm0znm06Mr8x+MrPhESyKdFm3PWwAMdPtIKiLb0vVlqU
4grOwY3th8u5tj7ErMYUNjHxF8HQexVq/CNMW277BAk/jC4Vt23QRCyosCcnHLEX
910hjQaiBpRBP8gxsigCFoFcZeL7xuLZ54jvK8N9XDgRySIgahhSmKlxDc6j5fR/
33EOo+gK6dCik+XCW+5hn8ksinAvIGDHdyRMX1e4WkEPCe4a0Or28LEc2G4VQTL3
+eiGLg3o3Yb7HXd68yAwliojUIJtZ0ClaZsgKZkQb9/T0arBGJqIMTNNcnoRBHbG
wrBAoahtUgpeJBtVdjEwxayQildsPkp8mljRSmsllBvcKg49dDY0h7MiCnwNKY+E
CEQs8WBML+nGIcsyStnPezRoV1TxFEnAimSehE5elBphwCrJ5025ghSh/7VH9V5n
fy4VHa/dMM2S/Hmg1fXkNrsKGUKoWXrgTKdjQtA8wDepwKnITCRWBaQ6tIvB+N0p
gYamLvHRacU57jHbMOaoeCJssiFkjQvUbTlXMu3dOhYTcazL8CXQHk1UG/hiW6ig
4Ke0kxayLUa3bw5EYOo+MADHqxvwmsY0BNzEjzh60Qqv0J/RsjgvlalNDkUsli4p
I0jeDAo2T3i6e8Pb5hxXCTA+wDjySctPnYoAYk4R11+m3O31mQAQZP7/C5+JjH92
GUn+HETefAbb2N+AQVkO5I6iyDCbSw3qhdjYTvE0hS2sl8tPeIiV7cOR/ErLmQZa
h9zq6B2CZPrC/vhOmUGvRkORNGRIitBsEq6TDoYE+zLJXoBHtALFptt8+I90YQDX
kImgiiirzKs13HfALpFONIOsPq8kBVk6d3CA203Lq6MuA7spmQuVKBdDD79K5ww7
c+lOvkZ+Wxy9fli39t2TULj7C1VjiGIVs08M+8P05FBjoJKsXM07ZcoDDOO6tnN+
dnNabZhEZRkTgJxLyYGjzPP6uaxNeUxOVpT8Zhml4x4rMkro6jkg3a6WPjiRsDBB
c1wpGAGeZ9P+aaU1IXsF8RufXG9vlA8iu9H/9isBvybzW0KNJ+iNIXSvJivNzYOT
46IZBFRLiC4TnDXPJxcEir1dZYMOyRb/20I/VM5qHUh1QMuBAL20CillLV3K7O6i
RejysKvEEzHD1Xf0Q0zL8oxzfeoiKfSwF2bAmzTo0Gd3jQHHTOthXah/yYUeyeVR
M8IOKTjnBBb2yXu23jfESJLSiHMtEVrhxaJvZjk5q+e7t9UkjALfbLlUtnUWLd6T
XiollRJWLcI6ixh8msRcoiczqhFmEmg6BOjsjFbLbUIjVpZK/hnnkddQYFF+yUDR
v25EBWcUb4z81Kpzqi5VbUz3tGLgjl8I74gY3nT7OlD9RG4AeTogCY8kcjnEIT4t
r2VQukkE1RsgYz+SOegwbjtjtUypjy/N5cmMWp07R4csa+548twC5gHbgCdWad7e
PJ9xAhuw/N4OnLBy8//HagCV/4zvO+kihibURzi+u9U8VhNuWj0in7uY9zfQaOfF
p1fe+KajmBr7XSfd73LV9hRDzTf9aw5VQj6JG9zYdt+s4d5NdZSgsyF5TKKImiOB
1hFi/Bf9cuxjs/upo+Ody7QZtJ6azSH9Obfb90gq+n1bGa37JuPsAWyv0yxUEyN3
/THtcaCR2/90GH0LvKTl9O/+bje8/59Zt1tyqaqc1BhkKHN/ghJdZfL1FLvX3EYP
T2CY7iXaboKjfAXXYkvOELeoct7rsMA2TibrD7LUldMgvrCKud7Ci3KrHbHG/Pb5
+fM3UD1OkAaLD5/ZELR5zjy1ZcIhEu1KVfcbsefuEi+RTYpwIGsjEELNnBbI4er2
qjjSeiT66amLsDB3iXuzPwt0+7R9IyKDpPtQn/aDPZaQLWnxNod2hDIDJw5mDoYe
JbAiTBcwIc/asYzwhFLDY/yyKIInD6MgZaBYfzx1bWTAHAUUs04SsC+AMPa02gvQ
wdrdQElHlgbWQ2cYYIRRHn+FSmiaSQX+nC9/wE5JVle4ZSNycnrdc0oH31/V7bZD
TplAlf+TzskzvD9vJu5nDWuw4ir/n0VG0IwAIf0FLxVGjeJUNv9It8aQhuwSKFUJ
/v0pbldlmr2odR4bTx676R6iidpAnovi+6IuR6s+pwXW9HsBjCxr9zGxetX7iRN2
jrj4Mu63WfpJIlf208RoIAVJtqsXrCrkrTVPbytj5IvUDTo9GUo8vvf0tqBRWvbd
5+JVrbsrvWsfD/2pqSj2KHhgsksthUA5SsaGuYPK/z2WONyFbsLgrZGR2akeJMsz
uJ/+GL5FJquuEj/V0wWCO3EiRVJw9dXu9rYIan4OKLwbYO6clnh93JKn16e1XzWo
3qjtrFlfT9uFarcx1YgCVpvWLMNy5gjVo+rOUjkgRLykK2JGnBrxB0CW9y0/CPIA
MKHdi2gOCBYcrBJhirGPdtbL2mCwJ8XYvNHWcQu7tLT2lHg3WcTdzOZs4tqYkJA2
oQnzuIB4T/ZbpMnn99nm7CVL42Og3FtoqvN/RMeBu7YjuzwjIEDkxiiysWDlFb36
84n0TPATrl65RrCwU2PwNKbZkFALHGNBeyfPDZJ7pBYCTdZekd0q7o/8m5PBE/eN
0Lr6+SvpgpZaCxmmwO4xUyQbOFfglo7sFRGRva/YjSZEF28Wxl0irjG2CFCQBbhD
jPbFoOcFjkths0+wb+Au02uybJQGSJKzejShOBmUu1oXi8wlIuxJTgbRPUTE0wyb
u7JrM3/+touzXhNJqZ815gI9GAxSbkCCgMdAZCwAoUrR3hzN3ISDeT8t9YwiFsIR
BJy3RijXXALJ3QtIQIE8T8D7IKsI22csbOGv7rk2cV7dmgjLMU5qfCWMwcn+2Vmt
DWXBLGom+p3FCXhgvekDguz7hkoxU6gT4fbUsROVDX95rjCBacMeLPvQSTP1HuxO
o024BRZyzAmjoI88Fy2Sj5V/zZIEFWaOxYXV4MxST7ZVEz455mUsLwEGDGCaOyRM
/MXHqGYK27qW5UXrcdq9JjR8KBDRUZILZIfY23wa8dCM/6YgrX2x7z2xYKYNdeWf
jsg5gsBggU7d9AXn1ZoxwyG9yxZ2jtelfgdZSp2lrpI0PMM0EkJy7+2P0UIqQfOv
5lCqAk6A64CfdWmSGQy2o8B8QjBfp7ifjyjWRxITcr2bKL91/OP2qURbdQOZZTxb
oy7G1088Sp1d2mLylSf01UISS9vYPA9bMeMUtdvcrH3LQaKOveEZ22BF4wphB5tl
4kaAfvT0fP1ZimrCBPWZYmob+fZb1SDf8khl37iLpAvoHf1ZxNWofq1+qyvvpIN0
P416n0P6wUScFYa96McQzTpiL3yiyC6rdxyhVh9IMqDCbZEhttW1Pz3+KK98o7/W
bT2gNGBQnZSqpr/vvMUavM49FU2AqtNrP7xxi7KAes8rjnBeyu5w3NQbWKUoELAe
3p2oYPXv761zPKLQ8/bmwvPTsu4CKZww6rjDit6MEXv4J33rsgNscNo2EkrS9tCF
9X9Z8kH5NJIfypGugRI2M+L2VJvi5aB6Jp55oCY70RkvZ9VJWwoPdQsFkexxpXC+
iJ+P1p7fTv9f+FZrEkr4ZwYPXRwIHPktFkx4Isi+I5VlHl85v/ezRXJyHKbyFAQK
P2PrSbwRFdiu+ZBubtw3yq5YpJe9+NkqIYWZ8HR2edJ3zDPf2bCudqZ28oAqzCB2
hX+WGA3/HGYs45T+7v7dRSPgDGPQ3iwfFk/WEzxz26yfRoG02FnMbMn3rz+MLpkM
A36wZR9n7nfqFNL6BNHJYZyZuolY2UllVl3BAFbZLQhxptkvq+mb+8NvhmBqKz8+
ZUK+6+zhs1Act+5aREbj4Uu9CksXEsLukNwTFR1Yjad/NSMWv30WI/3WOV/sbC+B
nW1nX9Ai6Uwx+rWZP9lrdKS53lGqVZT1bzbdLhYM5/ghyuRZ4DyHa2eza08hBFSF
/pcXTYKTuXk2em2W9zwCmXnwANm1XVqZ7DHkrdqRpHYpzH0BD0FYnTbgZdUKWIjn
xyqjuUzxm2AGKEMtohfcs7ztnB7pHq+fLXVeky6zmwtb1EpZrP3kkU4hfPMqIJmO
nQoOXEvrO2nyDQuVr1JRIK3g7MW1+oX9WF4ZTqvhh2JJDMjmULWPoU9UE/NNM4M3
3YsMOl2m2chDfBS/bcmbS2rnbIYtqLEEIdypVlP8viSfZGE67bkx4qt8RSLtxuIw
qoOb/VH3w+FquCjp7HCx1/A7Y1ctQiog8nRJWxn57tf14K8+HKWko6s0cJ+eKee3
4L6PcP9LvYXjmYAb+yux29hZzXFlISq5CxkRmLnsAOCt4dIuH1UUxoHz2HTi8/pF
rfX+dQHHFbxdu3PCMrnpmAOPE49aN7Ab1Ax4Vg+JcQ+r/uVHo+4OWcWt0wagMH90
Z70T8JVrAYJ4qD5e2RBHLQNYJJd8gMZCQaSGBNoQsVN2ZFY9YxYSNPIH7qQc76rq
oWl3pjratPcyHxHz5cat+lbs8a/txiRwonH6f5pOYarpaRtUHfQS42r38MUyFgpm
5runfUAXv4gl0W8HFg9DZQanci1ViI2eZhurSzbrbu0v+Jam2OYXhs9fmhOUMEI7
JZCWkVbvEI4gXFzn8/KabLw6MEjZ1DkhrXRVIrzjZhI35il5jn0J2nuQMS0ZkyLe
CZrSui3bsh6Lfnwcq62f5Sumyp2xLJKQS85H0VCSNhZLiQoq4IJ3eS18XAyda2om
IE5JY6YAdzc9Hs6Ob4vRM4h5q49G3YhAFVdE78RZtc+Q168KLDk5fzwEmIMeiGrc
7jFax5eRNLXnP/3gvUWF9+i2cHW/xBle96XwHNtDxeB8mtbsqgxSV08AfwK7nvNJ
u6iScITWRUaXW6QKPyEdAF2UrTxGbJCy9ogsNZEE0EpAOhd5plSAen/sGBpDeK84
OhLZ4d/+S+eNnerx2VQZn9yoKGH9BTFjGnL7B4CzDT1YY3w1/6YYi3oQzaiI9FD+
sYqzdsVZz8Hbwbbr3Xn5q8w/GhrYkEI2KdczMxLj8e1WLDxgE6m3FlBYYz6LH8cA
TcUATdF4iBnNQRge0bCOAfAoC0z9b3rmfrpUNeevmZwbFTFfYgKZFnxbJhAWFOa9
Z3EchlHtbgsj5Zq8tbCoJexCJhShtY+8ySWk/5C/0KC59/Xmd/QfCeVUCu6/z22C
vsPW9WKopaNHD6cHlqcEKu6Pjav2ZRQMEdohNp3RuFeaCiMwwfaupBTLGnQRiBHi
g1BwE9TLSQh2ZIjXS4VhJdn5gpWOoQWt/AfqxVCz5gyQfctlZpYJufBXk9BSHAB2
4BAjRoHbuKn3bd3MkXYP3oHVYIyuM1jEzQ0TSW8+nKl5mcwraM3R1pPYJD1LJ5XU
ciLGpNB/SRQfc43EFrI8XpGeo//1qplwMqE/AJbcOuXiqXPaUt53X0y09qwrkjle
acVEZlj3xVm9hpEg950PCcRzkiLrLROzly7oRZhSqIkV/5sJB4XosPb6DT3HWTBV
nXYv4B9uuP9CH8aKOl6C2SYG+LqjfAkLTc0Ug9kkeFqtzVdwmpPbJ8yIhwkeHQgE
05sNH/12M4buWO0Ku9sJcQ89NC168kVt+VhsGG34CrqyNki+Q1mdzG2ed3zdybnR
MtQC57rxT45kNS18/wzDHlkO3RNZysoGo+I8o3wQ6LvZ2F06t9Xi0AYiUivvakkG
sA5OrdIMFm713ZUDpZRCfYH3ruAlx/cqx2JvG/PGPhDoPlF3ghg4xsOM/+Gyo13r
jdBr8R16Tk0+T+GUOrXwIFxtCy2tbj3UTfqBbVd/+6jaqtFAPdVy1E3bg0lgMEJS
75WYiRPqzMNK5GkMOXHaddYpDi2+l4lYuqs8PEN/nvXkjHaIL/lzNP19n/ZzB5OV
na7ScUT6WQWRFTDD/xBo1kEKm3Nw8l7a1o5e1Aa+8J5I28XUQmnFegdRvoTJVyfF
tnU0wYNbSE3y8F8AxtcAtm2s0NfVdu0nA+6hvqMyBXlZVdaxYd8scPlDg68trwFf
0XvkIQVxHGyvBUbAJcpnSlG5DMIaRRGWbxRs3xnZW1RKcKyBLLHVOZDE5XlJlUix
wih6wBdkuIwkVieyCMg1Xbm90DecZjtjOQLgfKNytwxzPbD3+huUuqpK3slbeHcI
Avyj4ivBKw8EJCGxWDlnA/Ldgg76fBT1zaVwBspKENd+VOr/ZDg1LiH84FR8uVyu
eaH7ZrWW1U9z3Di6ByIUaESy1ALTUBPmLMd7rqC4tEsa+27VS2immyh5njlXOZmw
YmbDKi0qZztZgS36A81wMq4WPyAuyvpH9Oq39CTY3NyyItTvGr4NPQ+CAfyrjVVU
EH7n7Z+SY2Y+F+U0z3l1eFXQMhEOW9MVdEC1dEylIAtnyTIXgbx2G5Cv9jbXTaix
WP8OMGJm18pQYAZK5w8/C5qKP6bj+W7Yxi8UwPicK5qLBsNBx4rbsOZm3XPBE8ae
9qsZNVB7RoKvvaG437gVjgv1PPIJPzWh85770cahYTWwrhrd8fIICQiEWTwL5JH2
7m5TkXjnNhnFiV0J/lJrTjCl2rCCVQP71V8WsokO+ze0IW80Uk1OD0ZuNCO0+Lmo
bHNkuSlOpSkpnkyd9+JjQVXkJrJd7SWa7uTLnu6Gl+lxwcW+Lnn+BuJjLIKbiH5l
SX9Ti1cOzae+087HiwDawJqUociW7crtoyRMMAhdTe6QNfuVxFwb2yP5Ty/FB+/W
NNxoF1Cd21FWn3/mTAFG5hs6BKtW4Xd4wvU041HBQArSFiRtMSbnPRJFidTEaXo6
0z0ImL6wTZHh8R2ErG56rIZ9q4niqXywfEGjPkpRr7rlyPyKo4yV2BFwJnH6I2gx
2D6Bxx3wXVdLPLymZBtzEJ9E8b9xPVId2U31HjBUm5gjZpvkkXEz3JnYnYYXbWqo
r4RNCmwHtLEnyc+aKxsDvinfB8YaLbSOId1dHK3LtIEBcQ2kiWxNysUiCGjfc/QV
vWIrAk1ZTcwpeHQxAl2grXskFonmQi2Zo3DFi/aJnX4oHCDhoUcufetWdMYChcC4
RMHwZnV+1V9/mccFQo1C1tMJjBpxOKVXyoW98qcxpOZnr+1dLt8xYs8k9gPhlz0D
JF6Z2/hz1+M4lL3YUg2diZ8kY1jehAWOvTt7y/gKzxg5x3WHZG2z+7cz4InkOC7l
abbE5JNiaryrzN6zPHeTl3gU6CfY9MgJwc+/9tc8MQcjms8qtN2Jokb5qmVbA3LK
ZCsvew1vk7rlJIIH1KpLdlh3mrYUqqSjmYtTIQ1JVEi10QMYyRidtFj8/sciz0zM
SFEL9pR0aIekHbxaFPVwNmgznKMcPssUGVdJT4VjQsVHma/9MVaNIP2/QdCyidil
A6xqTMu0ZZZQQyJkYUTUGRaTON0NhAfGuVmX48cvjumBJPZ87o3X6op1oVMcCFxu
hGVh2XXsRl5izY2GNkSelgQNin+6VgNc1xkSSgF/t4dql93gbMxGJvxavWtfC96o
H9QtwjiJxzigRYwTqTTwW6w7BeaM4GWFY1kyMdRX/EOY0rHJukD6oy8uPNKl+QhZ
tORc2u3npsTCPRTQoyuVJgR7+TRjSojM3G5YTWAqp0aKIxikE4avwbmRftcLXXMd
iI6g7PFK8sIWcdgKqVOe9AwlPusZ/crk41D4cxBisXQZoqcQdDl5NxtepCkhFvaX
Y71/DZwnvALMI+NWM05Kvq7I4BrVNLW2a8zFq/XCsGoIiLLd5lPmeXsSbR81AsKD
9PwvEksqrORy9FmDCutoNY086C7l6Tp799C/cpL3E9chD9YpjDkcajc2gh4hWmXT
mU/dSIwS5rHF6r3BzWxQVZ411VNqo8PU/hFZCa9dn6PjsC4TsBl1SoG4AyJmjqaU
DlrA7LuVLiIlxU1SC1ObQQSNY7j5z8S9HaLDpXu48mqx3bEgPjvH/axI84vPjXGE
MjR1qDEokECzkOJlFLwiKgkVWw/DMY1HgPWv46XyK7gAiPSHu42uS4pBFF2K6dD9
nIymhOYeFcvo1t9EcFddMJ5ZGBU3z4/h5LTzsp7p2akwAlrmTRmJ9zJiRiX+C/1y
+e/l7Fm5KWgF6R4udeMPGw6DWAqe73a9tdjeqbYi2VZLev2AQm3vqhbSANdg4lVk
VTZrONl0wk0zKKYxlCle7uy6wQDnvu/Rcrmch/ncPDEA5y9eyEMbU+MEXzY2Ajaq
l9QuNEAyaFo9J6R/c4q0ucQxyEexpa5lPTV6m+Kb5OpP/HtZ6EfDgNHfnMKcL+HZ
UAPoAafyq9M0fcxHu9bbMuKmQlGVjv36YNjCQDyfMWtEIhQPeszSNqbT/iJNriFJ
xcDgF8uDXpi10JHP4DXGDUMYY9H8kW6zodu8ox/FZnCR6SR0fYEullt3G3RX2die
mNjjW7XzgzM0O+IT+oMoGWsnM0dJkxKHmJpL3oskJghCaOhXQR7dP2DQ/wENFiaN
il9WhQOWsPhNC5OJTmXVNTG3apM/IH4hcJ2Uu9HkBNJeFCreFd1MwvXTm2GonyIF
xNyCNtFxkZtyFQuGot3sDXOs+QYMNWedpQHLiGh/9Fvw1deeyKy/SbOmIReMFCSm
3eo1iLKubw4if9ycMK+uIzK8b4xR81cMkqlh6RPox0bkB/Sq1lGqaY06wE79dTxh
yt20YvkA+dHF9iSJvvL/KGhDTILXdLpCe+JSmNaEtteg3NOGbQqdiynzSRi+Tioj
reDhJ3cmkwEBuBi/KxMpmb9WMAH6Opzn4zSyf2aLveLP1iF8KEtq/E0l8MSsFWYc
SXF25km10fRyG9/yYope6vd2OqTVTXcz7cZgmQtCJWLnS3AaWG46iOVKOPRO9owM
8ZwVibzok7rzoovccNmPY/ZaiP/OBEQeOh1l2Yd4MydycdQOU4qjh97hpHnjvs95
paJj6bcHUrgsXEZgChEwVIubqpxKCqKpYq/SKDTWVlKHCzWLwY+cFQmrWMK3Vtp9
PeM9+yp2/gE9b+mEOs0JO0GlNM1Io6KJJxs18UjbAT8rYUHHr/uLra9oaSB9LusC
OrdLwYKBm4GQ10LmkaxNTPpHWFRxqX624HorUs/pEpUK06I1u+LTwtzheLAygTwR
reG53EMZESoqiyU9JbXwKN79o6+2ORfGtOtpxzu/OAy7UpC/xTwk6gJWmln6w++A
2gfVJzsqK7U1t5PtHH9uY7WPJqoITw5gOYc5d8Y3yjulwWD5PI8wLY5IbFC8GXux
oPooKaqLeB0I1JR0XCWzE/N1ZApKBzYQsgnu/YQnzH0jfR1Zv5rCXyEahsLcvvUB
1GlgldlfrYLchtxhwGPtxSRM6v5aoH9m5yQ/q0khXCcndn9r/BR2QD8xa6eCB8W7
WIJmPcUdXnqhwIV0RWuBZ5oz2QC29ijZwQCAjYDsbKEtGPTplzOLo/VSWjYXUQu6
4/5v1obWRlAKg8IboEmVXfn+rAhB7mXOY6Hzj4imz6FThFuqaiJMMzQ2dHgTrDzt
47XMotT24foebEPVa+xMKl1GCxMMeGbQpJFgvKwjgkggm/PB+/HoO/J2TVYVPzed
RA41O0tYyhva2yIQM6qDwBdYeXV7Rv3ShwfSYKWYAZOAvQkpjWnFivg7U6J1Vx7H
jkIUnwMmJpNRPf405Rt8mPkLT56I9IkGP5eQnLjiUGpSLo2Q996dgN5V6jLAGhgy
KHWqWmsb/Dj/HGY1LItcsZvnfS1a/LytXRC8t94LlBmOn2T/BVA8Lg3W00mbOi5N
xvOoNlaHYNWPkuWQMNDqNrqH2CroNteHpz98+CBYoO7cYa1X1+JHN7tq6I0DVZAR
mSYrLeiDcmdAO3tC+IFpRg5O/SOH+mO3L0JK38+RRvEai5TsBegvA+MWYxv1GYi8
IUqN9+U7VuEbeTiFZTzr0uDv327tQ9d7JVUyftCUJ8D20L/EifVfro0rgABpXD44
8jJWKuTarws50NYDkvv9nJilD02I+9n7xk2OCnOfv0b/9GpbISNy3RPzHl8Ii2HP
py5OlqX2zr6MCkf891pce71rygnkvOzX56jhAbksbRvLW5a+SgGW6zbN4bg1of5Q
DhVqvD5BO6BUCMCgWuBs/1kMscwESZAUoRtrZqCGNDjxo4MJhlqEmBc6vVIclqBP
6oCEW1z9IE0a/ZMgAZRa0fVG6JtmwTjT2ULQutVAmf3DsFqy1utNBz1hwxK1ILOx
Lq9TaR+gZZKAvaOBf/jYiDuRIfDmZ1y/dRnuPYUYJN4s+Hve3EwL94suHVntGyNZ
/FMByuKeb/xbpWtJ9lBxarfjEBnawI0o4yD+eKyUhC2KEWTus5apUL6GX3dHtH5C
S5qoP9yLJ3sdNkTGUNC6EzEPo1vR41RLtA+J4j/2nB06myQqkYxtjObaw2sxiaIz
wGS96r4zMFGWh6BAo0P9w5/0YUEazvbUi2RBMnW2e22XfSgbVW80kgxOCCEj+8VQ
Jc6jvO6UVbv7HpTNT8DlxbQi0cI6iDqa5h709JlnZzo3DrEaFc+EtpB9koM1NgE9
MkWawnL8tytggWe/StL2JVmV4Zzf1B9ORXlzQP5Vhr7NKEK9qSc8VddVYEVhb7hy
D3hNHhcgaWSN/EvMoLSn+cNq/cIvtao613seTNoIiwT982uNy7zX2t3yttOa8OGH
T8oRRMO9Oqqol0wvJ7nEELdBqZYcxCkoxQGknTvC3n23+ofCVhczlj1ArII9T3GG
ArYHfjJKlQQ+m397EusowiFwO/3rwlFsnLW6lfLXeGRJ6GdFo8WTJ7SBbpOy97Dl
MHqSbPan5RNZaARmZF5Xy4q8Q7oc9egQLJIQwUwJlbQSh/tlriWRTTm/YUCOOF83
uBi2s8zZXIUG/x1lWeAM9xVX+WRWHLTIeVLdYn2Tfm+g8ljDpHfwZhbqSqu92z9s
b4PqjAjttwbEZIxckLMBdreBwcLDIWZWb1v9DA8o+c/G9XH1zdAulw5saXPuoU5W
57fErHn0K8tBu4ENwg4R391PwYIUo+LHGqdfbFCbVR73AypOauw3yEFupDhZVZ9r
UQhfrsdrXULhGRO4PrTtMKn3hhzMHKPl9FmdS3MXsvv7OtHoWELxvZ9ZHa2FrHXR
UK6a2/du5BLsSCFwPTLsVL8TCBdvSGYmzONEgaNR7H0t+Rpn8HJLAc/6hGFOg/XT
Rxjhbzt5vf6B38Idpqz9I03Qj7cez9pxUdQcXmw8diw+rAxw3zEYsHEy/41RhpM0
NhNl6aTMw9JPEeEeRlNQ9UFBUFHmRj6Yx5SN7tXw6x2gqcggMLkytmtS6GdDaGkh
EonzHJLPr0Esrpe0Eos3529smOqsnrdqg/eeUONW4Zaumrj37P6ClgC3Qr3WLJJt
OiAthcctnOKX7E6xoK8n4PVgyph72YMUnQ9/Fl15+kw6bhZxEUEKOVQvSTAV/Aya
CfSxnrfF3FWgrmGlE3LtIh5E7J6ApBdBc1layHpSAl6WmYvY8UAfdDD9vZfoidv5
2G9iyoltqfJH1KzF+XK71ONolPgoKMq/i1Mrs2ltwxfAcx3nRa3nbjqRJAAeX7QR
xieYaDD8PlbF2TOq7VjBUL6TbZoHJpXgPWbG/CkbK+tFyovUJzhi61wZqMzU4cYx
ER8J3+c1sUdLwxMplvTX3b+QTDUNzOiTX9WIu5YZ2n+WWfWw5yFMYCqrgbK3xnGV
32YYnX0vPR4naTHrVzN0O/zEcvmzPpDdamiw5XOItqv/TeLoKZY3CIp97oMwPE/6
Ecb1tZMlFHfIPmbBFgksANf4nT5egnF5W4bqM+FhzpwHKrAno53rofwHyA3jMiP1
x77zoJcZeYqduFMP/ZZcUTW4a2/C750I8CdacW3a5zEkflgrtgTwPT7OdMaLxawp
DLRnKPQRurCwlATt15OGSTtx9YXrfcR9ze6ZpZ+psvsvO9bCyXu0koSgMoayfuYq
BdChhetyFzDr4GN0AHKWRB904Q+TIy5iqep4wKUdJqq0k6mAsSiWtsogC7lyhAH/
aJZnW/EO8sUqeYt1AbHonotO50I9Bu//nJVPoMy9UoTp5KZ4eUdjaVJp10CsviE2
O6Go3i8eUloWG7T3qDegLwf3ZK8Bx6BOgKUeLLDKhKD2Bt6Gc5fSNRkvduXsrx2r
uEfi1/NSgVeZ7tTL2mUUmFvIczLLDlNvzEEO96N0xp6qIzgIPZ6R8f3GY12raUXb
yEg7iq2xAHRxjceo6g6jSre4V6UGZL/JtZj403WbZyVZFuGvUWsTNzpkVs2GE65v
643Keo37rXlN8LFC2wC96jmhDAF0ATk+/JfrAGmqnCrxV/F4GmmGa3/YilD5vCOy
SMF8c0NCd0SG5JkicvbUzcoPm1vQOCCR0eN14SbRLi/YhS0lcGXp+NRRaOFotk+n
iTUWy0eod8C9VwJD/VIQXtzwoU9nt9rKHzrxwq4uskZQWuSP9KyJJiFqquAZs5VS
LnGB5p0HucEPlKfksinzSxExaKe3v+5g/P3lbN8ZGE4yiXkSLTdg5PdmmDnEvjcv
nsI7DeF3cy6/9sQA5veDbh46S1uuZlNlPLq69GKzUGMPaQSAuY7ycTLObF8f15sh
HfSeqycZ12X/wIu/X4c7vjuX298Igzgxe5A6aCEZJeGkntDSLuSj03IcFl45mAVK
HKtNJo6iVBvV0nqqmyh7LtlDHxNjpiuFG302TZ/OX2SN15pqaQZNrxck+Eilso7l
eZowEgtqqbWrNrh3UAbBVPb5faelyZKBevQVmQGKP3NLeG1iYVeuU6Sc7BnuSGWr
LNWTbfaBVdNHOq7ecqe6u7vF4erX9Dl3PMd+QhlahZUsMsAmPa1bOc0i++OUrImm
Im2W/vm4GJHTviIo6dQzk61EvB5DTuMuT3UQbUllm0OYA/azChDTwrQYJNZ9JfQ4
2GNrAtWBMx+1nFdVGoLZ0rPgvoMg8GiVOu3YNA7Z0P/iGJ92ys9ZjDsZKns02Ptd
Hd874d50Fuslhj7H9CxX8Zjw8YIWeuvibl+0c5+YUy7x8rnqkwJ3FAVyHXY9UHKu
kW1T0V0A/cg2FTZ4xFrd8ga8oCQO4GcJK4390kg6YT/aUX+ATwtpeUNVubsUdo0D
pnD7M+FlRBUgjm6eJnKqqTt+ArYvOfwMrXQMCA3NUFKwg9svdzdMxpeHdARoEG3L
CwFMPwzCyW+NB79/+DSyJ2J7hxaXvTEmXQFMWns0Ai7+JV340KjmsP2CpXu5ALIj
una/bY0HgRl5lsOLYvPhZDu63/Z2dRWPjX8fttkp4Z8RK/TIr65JX4C9yp4zKY1s
ZkZktXtomXwg+Ak1ypKJhYBTEqQaM8YNBOP65fidcPxAtxGee1RlcUQc6tKeVmgp
rxvXh1JESjDZxw8NLbTreG0dIKE/4suvbNSAish4I7mifQMPgtZVd49vdAmqtEdd
37eQCDgWwTZh3dr9j+HTVoADY8Z/ZwcZDaIoERdbgW+wxvYokRLr6fzh8viKUgN5
EWi+PN/UpJVB0eWvbglAH8hAmD/R6R8zFZTWtgZPmmEeVj7DVopagjMfo89HiKsM
YkBr0pkpnTBBnOG28pvY4c/fqt8JOt5q16JvOWRotSkdG8clhM6PkGqzGWuXqld7
GDNHgOer6gwA3TqCo+YSVMRFeyku6h/j9DQjNix9qbGwCEh2/nH+RcuOmYQ3CuBd
mR+79NHxPrDuCzQllm6ijw64K/etJ/R3c8/cxzjFiJYdOJQgUdDIG/bowA2RvvSR
xitxNH9oVEq8L/HJehBx8hYnDRHl8yfb1wU3VvWrBSPwy992HjJFTZYojaEYR1yj
5DfYKlHj4u2KvZxaHTvCzyy/u9kH+sK1CfILUvKxFy/jy6+3OPamENs3e+3NLfnv
4+YzGKbzakjVSKoLevg54JGjymN+qttqEFHj70eeq424OvJyUOP1asnfNMpYaZWK
WoR9fsVzYZn11sAVvAS11D9jOD37erGZrRGCkaGTYGJV7QMF0tIRc3Ke/N519vA7
cOhfBDI0fPENGK02zg3yMrOU7XEHBuCu531jm67ldXtH/2ZcVeYDPZYdDtJ6GfC+
HXEBqe8C6hvaap+8G7E/1Eo7lazRjy9fV5cqj7FpGKRMSvDc0BSsYk3TkYEirmSC
CBrMz9Kp0GVyKp9UTRxyxcupUW2+V22iNIBUDhprTxi7HDMDFIogWCyVlQo/yWU8
kvcPQ7wHUbPPfPI0qQC5UpARoxfYjEkTCej4b66u9slGl2PLijw1kLjlBLqfNlMK
BPTZRTYjoW6ddhWg3n7zPJDrP9O2BdpGBo6SWNf6NgX39xdmymqgbgdkR0FueQGm
55mZf8+77ox/Syy4rgZTR+7yqlxnoAVqDYH0zFzF54EfLWFJUglq5euWiF//K4qD
MqhKhiNAi7EnIMbM/7dStKf2WY3fGTWWsMqQw+ClnIcWvKm3jJOdQbjozRq3+Yrf
9e+ZRFeoBm+pfpMkM/tDO2j1CVBgg+ZyxkcJrTz76V6QcPnWMqmitOERVr8MmlFo
UjYHXYeUBjq+8rFs9zfivYK2qCxP3oHo1gIgos09HUeNUQ+iWdkXYZZyaBQJUDWy
pQ2VKKkXMq2lszg3nmhaN6F2aw+aBHEL1GbMuyAI1JdaXmFnTDaMt4Ga4nMkGaUK
MNupueP48yARJFOIbykqD1w7mn5GSuS+8RvFMmVsJ/LR7c9QS/cxty3k+9pbkX2A
bwj38k7CwmhFGImDca5KjSP4I2nBXXZuXrM+vnBP7PDdmwJKH1YwGzIDtHA2D78S
fTAnzzEBGOq8tzQI5WoP/p6evCfaPCJCsiesMGY/u5ZNc6Q987GUegu2p67zIaJV
GZn1lGxaQfViTMR8tH1nasclWz8udsbvDreh11DtTMyEAyVJ7OwRZf8VrpDSour0
5UdqgTY89GQ/SDjZtvAiF+SWnTrvbwFpL9C1I3kIorc5sDlTpaXDTVoDhJg5Tr1P
TkXWxhkHuwEJIdMGXvlniZiaFHxb9PdfnfIvbwz1zOFQG1qJtcF2neybuMjHXBH5
vjcPTrjhcEHb/muU18V+Zejab0CtHSJY1NEW6jcui6OOFhBuygItrIvA89wzc1dR
OUac3yB8cn8SYF4DNU0Omk/WQMcdM58PheoU0dv9yl2+nCW1fyhPYRscy4Q+L3rx
SctlMfkQFO9N2V1VaujOEBwcCuTJsoKracQsJcOVH6EIRtrX3AnSc56UPAU9m22M
wIkUNlfAeAVvOfEf3r8qCq+Bx4mIjyqNqXZb37v8MgiT05L/9AumtDcFoprbxIv6
+P8Xj/CpyTE3koXEbRgSU+JFchgp+LNQf0QHwUl9l/u2PbGNDqCLYCITEEglurd7
pSuXCGMdomPqNNG8A9YgJxbJLPCMovygUF4t7TR8k/bj/pJ4sPPKHMiSiw0yDWEG
UaR/4+hLS9DZ1a5Ne0Uxd9iIjKmSJMt6bBQMvva2X++aObyZky+6GU8xZ3s3JKaj
K29q8CTqGUyJYSQDUa2mTI+r4r4TkmdAkyJcOhq5q9KlwbwVEiq//EKHnfLGNbcG
pIk8/AqYzV0Jv2f9kcfWXP8PQFK0RP4fH6HZXfkDuZCSXYitGQ27Ws/hOgzvvTJx
gVDJjTXSizRi4RBwIjuHsJpcyCFRhx0xO0tIl4nsHe5DiQxwK/zPFiWSC8e3j+A3
lvT493ww/jx+W7YZtFZ0p0+tqBY30sGDEEAjCBoiASPyVM51NnZLOgoF2AUfiNUZ
HBePNdh7IUJDHbNF4T1rODC4WkD42hY08jr6Ul9HUjLZJYaT6SGTJ77wlolfronn
IIRMoF7k/r7mhuk+01FV0vasT+C9FfkKpFKzuUD2swnufBBJ+1a+vkrCYbmF4BfW
uKZTWgnUAAn2F2d1eD9SutH4z++t03ZsfQWCwxMUoQzAUjpzl5dZtjABJOg6ytn+
LfFria8tEepFABd3yZg8djiFbsz32FL58PTLRhBSsi2Qyudt9b4myYoMBymQ3bxU
CVLAPeMJOrmoONbXr6+bt7rDbrryZkMia/+14AIRMkoSPWN0t1c+KcpM8cdIQjQG
v6sybtBV3UMtFIvCl2KGP0dsOtLVumMy0Qt/MwbtXCwbEwUCdLkFTSC+HDA9MMf6
+8OeIiBCdd3ahYRa84SJJlWcOw7GjdKkxazpzWotbeyIGS8/AfnUmptIpzH/wSUV
TDFBAA/xIoz2CpAmoTPe7QOHT0jqozVbu7e5D6SZZDGfu2wR1JH7KzeH2Wddq7S7
v/kVovSf26RpLt33ZcJbRb+Qz2vpn6kcD8bH/HEv30bHxMnHgyPwYsh8/UcKZiJR
bGgK3TJNqvCPW5FpSypY8qlCYemtrLelR3ON8MOtIjjuI9XlPGcL6KFLxJ4ATBz+
rs72NS9LAAUGrHjsiwb9Zv47rHDnNOwM3PpWdDnt3EspvzlIPMgo5FrNUpUQa9kM
L8q4HFsLofmr6oK/S5btBYOu6gvJg2Q4GmHtmFp1TC4aePU2CsrTXYvoYgI8vfkN
H5tfRJK19BfSprtCRxMT9SAwW0et9R8bdOGQbHyIyqKxc1qLsOK6qjImjvN+6oWX
4Buj37s0T2BP1RpsTP6tUg6cNyANzBP00Sv+zCDKQi0PbCD+BHgIDE4KiSEKKOBL
bRueizIYWuo35vzMAZSi14LYfgMMa0treoW5qgVC8LAZjG8Kwk/3eDTluuabku0s
w5swh8Bp6X0A3JgRyfl9UkC3IOmO4QASDM7a0eTg3kd0FZDkKfPIvv3kDIlohZc9
dy5nZcMNbufAiWA1ie7PDNUotxKz8KB4Pp9lbcVCMDOle3zhUR+cQsQ7N3w9mDqL
vYNwwC7hKvBvhKkgFoFB9IoUxWEBxxPcVsnO571DvDOAN8s/4jtBadZf5lW3oMCZ
nhjTY/5/sqQ0ZH5V1n31DiYkQbUbsW+u56gOY7tVc0e2dFP6ti+FXMs8PGJ0zhfR
zgK77YkZy1UU7x3QqDZpKPwmru5xP6dvASIpyckjjnpRgxAOJLJBQG+9zec8M414
lik+cEG7DN481Ua9VC44oWU3JER+ofq4G9bbYobnh4dfH2IjlOGmysR1yOb/A6bk
lSnCArwEpoGtfEwZ7lynr5JLv35sl3KolX1Bqq9b1SFp33ZMXCiMmNAGshcuGN5l
80naQpsmoD73yPooPudpbsVvq28lWMbbbQWxJ16Gy7+qHhVNHWRBWd4kbPOZ3gF6
qC+d/P7oM64rc7NU3aCakTYeeY1rJvAZiOwsZcO/2c52gV9aSXhRNqZ3NcTYaJ8b
2Va17uqHY+EtzGAD5U+Vj1jsiRoLY9BJruDjA/RUMRGCdmHZWi39q1vsb0DVEttj
69uD27MyZ40e7KLMIyj0RYINk2P8pkXgFaYvwkjOTFPlt8pQxrH0g8rDuuVVkSEV
oa0oLnqvNHqjKKbm4cK7NdPp86pA2KB37Qnq921wuGlvHsPSzWpGnLES4/XCZ+PV
G38cufOdVMHK1OtDjgT27vGpojJ7qhRrhjg4F0QwiJu9Esz45mRiIZif2G8HETJT
DDrX09hCwFztJHEISrXHCs+NEQT7JCzH83LAtfhjg5NYd5rtWHfWak4FtfIrgIgN
oHYB5BOnwO4IyQ0uSb1n13FnYZGQJczneJn6o6uJi3Royy555krBiYlKNhYJ2gzx
GSnBlufLwlWrhDQ5lOn996WpNVlsy0LvS9/fAvHvZsJTxUSPQKDP4PoWTQsMI6tA
0hVwfuFLQduLO25ObthHOgKqSwGBR282mpmannJ0nWUlK7aP1ODTKriVB7am/LAv
VFp6ojZFQ3lmdHdgsERKk/zuA5Bvs4ozs6lPcux16c0ZCX7QCJA7r10S1QGYthTu
20Q1uglTw81qeatHiNcaDAFIAs77wDU76bE4xdbmmb7FkhZuJyCdy4YcyhfZpqaj
M9b9rFdZUX/PsfE0+MZkW6V2a0tWvayPVwd+8tg/MVIV5APLNShFHQ7vPOs16/R0
ueERyTPT9E544D87NWrgBAhBfdHkLrKYgp6uvzoD3m7nZSUluLa8rJgMCJ7dSvCW
6DCHhuqL+1hNriGpSE/zQkz7k4vhYELPSwrulq/MREC/7YIHT1qwxeITd5bO5a2p
KYo4FAu6CxZFfzVa9ZfH0HSwrM8WXfUQGWOQBRQpUMxbRIa1GgIWYh9wEcO1MXlT
+OXoQbSuaumG76grSc7cNPQAE5VqAH46mhohtuzg+oDH+8zvw3cya6E2yXRUnm0e
BnXitNmsExrNOQngAISO9frxOTQM38+LRvb92iHdRT/PiJb9OrYUHcu/BstkAgt1
C3xmpFXiJK4OipND1H/gD50C9Caa6smldhXLGvRrQsEc5YZfm8odzARnJJKGnOz3
0AQyFuj3iFKhcI5pK+VPgicw53vESzJKwv5PNJHVJO5pHrbbZ3lyQYiZGGLS78jY
1UOBxki51xbm2fRpJ1oz7cpUKeCgQJVfu4SYhcEe0o8liKNtly6bcVFhPvsknywv
Tb87y0SCJ7jMCh1UdrJzIDLqoEyH8AHFJgOnbX9fn4GNbiqRNL07IkqS1PtzJMIn
xEFPfSWm8Br3Aq5SoyvbI7vzmfsRoUJlMEfbbzSq2OicpPlYPHvt8dml6EcZF+oP
qaUrnIPuUm9MAb6Fa3tRT7wXX7FRp9wcOHxY+SV5eNgiXLP0mm0I4AkdlP/zBgIz
LjojuQZiNfWmBN7mRHUFsGI+nw+1U92xKy5cGG0+lmVBRlWFEBeZ37ZBfjhV+Mzs
HV+vXqw0945/pZzVhVP3Qb7gijvGjgRcYXXyV8m0bU9oLqQ8wBk8Y+c+R9/FrvIt
muGMtcGqkdc46yNhwpFrf6VB4wl8SD4+Ds8B/Nj98O8mpccC6O92C4EXBk///xZ8
n5sut/1zRKoYt4/E4CMp2b2BUrqPkWryzxHJ876/dDhPRxOpKaKiw7p4IwfgqW2v
Ai/eviFnkG4T56yHN6yBq8rcXTLBiwX9EJFDezb6ciFfTomezcXIKP0IFX3KsglZ
ynIAbV/u7iPzLUP/4GErbGO9i26xQ11/gKHDFMDTsFPNQ4HBY7bHFr1dCgZcqAQ6
JUSKNbKIgYYfyXOXpcnr5UkcR186+842/SnN23kKuQP3O29IpAX/p676G5lfuaQB
ers187Oo4tAW1qHafztThuyXVio/7rBWpsszNFxQiRHJf2oZRtjG3ZyoarejS/HL
Q+tzNy4GXBzxZqPj3FghoEYxflB1z5yFZfT4YlMv2OqYo6CKdGXqF0R/NkezCsqS
bfeZz94GHvzvYL5hJ4W46dtGqtNrSOvRkMh4L4BrH/mbl3kWe7E9Lo0c8X3QfH1v
u877e9Cj7wL1dUNA5hMMKuApeFjnaGGr7YG2LFQfwi9o7K4e9R84IGM0CCOt4I68
BbSli/oSxHz+JA5LcjlhgDvW3BGFkm2huPWglR0tp2NGOrVs3BVDJ4KFU9v8vS7Z
9TF1Q4Vv6n2AB1yUHHOqNnVXsyWSdFFgWO8ItxxohVDsCKrRu5xrk7VoG0GgbYyE
WSXRLthOCJejpZVHplm8PaFxaaUsB8nM/oHWi/GLbT8ik0pkip50hii95KTWA50B
PJT/aS85WNSW9LMZGSpLjUmK4ew9o8X0PwiV3Qx1IW37nQbbHfRl8Zau5Whyu6Tn
MDVaBxZU/MDFgevPpqKu3QQSKL1vl0k7IEfTapzjWJP8XhihM6Lylc4MP+3yhbJl
HoA+/GRJcUy7wNDr/SQk5k7+4KntI411fOfMzvX8X35P4mYCv0kEXdE3QvrNU01r
FPZJjAg/ms7EVyaItliOumbrNxzcaZyK3XYUUz3VOOtX4fSEBgu109Ys6APS4tQ6
ykExvqJc8Uc/A0Iz1m7UjhzPhF0gVcgJ7c6Unxu7dpJizvsixA0SkX3dSFKsqxcs
FGCm49aCO8gKseq3b6LRmyKw+nrp8BCID0+tmoMoWAXTBIQC9PWq2I46cyLi8X4l
ptX+BCjJ+hSaBM6z5bkdNuXg3OZXFnHv5yReXexo2n8WJtkUos5AB8x6uE7bw3lX
Gde5UWY6ZkWqCf4gKKlEij89npqrIBDSvO1i0NEtM+0h0MLZTKPu+wEa6o0DcLPa
vbRa5OylbyGWNgi5SqghXbodfOIvHJrRySQ2OC2UiHpmDcgjJNQ6AVpM5JCZZCLo
xQ1HNy95tgnawrAH8Nr/CsyjsEOh/Zv+pKMPBH2l9e7QgtMbrzwGE5fo9Knuqf/o
gARgPRBiHMSI40OHzM6WLmc/P9v7+HtE6DRnbF5Cktmjbd8pSmbsyyHGkCF14PtP
vXTsR+QKTT5lHTQ2V3AyL6GI1lPazOl1z090/9CK93V24Sr+F5DzjFW7qHGw8g3y
BJTD//fgjIFagiCzXbsY4HThAoxIqaulprrKids2h+vOaZeINN7oHPcgwucGAPpD
DNgRwRceRAH7UOfmr+ZdMipbq/4ISHtJR+JWnNrqquThgDPACUly+3MvzNfWLRd7
f6AIEOm2lIZ+7L4xL04pGCpSUwlbrX/ILe7pFxO4BmKgx+iKzpqZpJ9P37Hg7Tdw
OR6evRZvMOQxGSl3GXlS7HmANknoIbgNRPSDj6Hr2oWlZkeLjx0t94fQfxaIqN8s
6GJjFQltw5eexPiUwGInuwB40NBX4WZj0S+7jPKhVIvnmIEyr0dFHQiz6ZicK9Ga
GfWQkeyG33TXMU44/mO4DG4r7iF10iDUwN1gsEjuP0EjIWexghqTNJ2aqOn5oJO7
ChzH0nK65tzopyj/ZLrNc8LeuYPFJJbJWi3Jov4aPlQQv3zTKKbDaJ/k350B2fzI
C2NFqhBhbfjL7Ac40rZCCG5ReZn4fHWClMkMdlETAsvqeIlmwFtyqU4JA4THazhg
UXNqJLEyJwF7PfL+ze08vTeLK7mdhsm8jwuSKg9dvZqZK52z0Utv+c9RTuMWuP6g
Ih9nvEWUkNeE0T1gb7cYEI8zQQ/2L7Vm/1qNEhJcMC/drfnTaX7NKlTDEBkySbyn
ShaN7Y4mGBu0m7+BVyDAP6dY+1ldv5tdMtRf7vvHaPTM4g15DPMYx+sOMgIf9nOQ
ZW7xoTFfnC7Ygj//Ehi0S8vLDXCARXMSEmJHfKhkxdcfzbmSkQ0QuE2QTc2jfj+i
8EeIM6arlZv4TboXwXGlMYAavsWoOoRDhImlcRJywqp0NMbGPcVRtGjoM4qSqRDO
GSipXfrcsJ1jZgz+53I6huPgLv+N3Vv81MmjiWepl8ebIRqwjfSETusXMpiLmUGZ
qo4DSVSW3ZCpxwPkXT/8TeIaXyE/H91q8TLi3ntw5CUt0Oa+kw/aAGGX5XmLEy2p
l2WaxX76v2EvjR36HOdhB2TwUkxI8km1tzalJRCDLrgXMKAfcns34flmsSD2kuTq
ShUdDkJucl7MQpinqZhHMyG5g36zxTEfsmoYY6U3a9oiWIacssk+KBjF4kflC/ds
GjcqqYq+dBX1iFECQdyCr9vdzAKxd2b9fBHLfysvPZPHAs1U6AFugg9/Rdpx9WFF
r96nd0z51tp3pee+TZEyUObsnEAC8Yo2klcrJxSzv7BvfdLH1pPGlNOQW2yMbAH0
ZS0UwOVS1qzryIB45kVbRHqCduLukMaVbTkimp58+oyfaYk5CUKgGpm3UDibyFqY
DQROqohd+nz/pZXuotkbEd75GBeuqh3W5iAcma56vTBAkrbZPQL85MC8/m8j0XSy
1w9YI7vntYtg5OGoh9+bkW+EcVzxppylgVCM9PWlahUWE3mjtCnAjKfmgceZBmyv
z9WBE3Ych3IFmsDzCpbbtPCsxJTzbgXxfd4qncTMm+stNSxbATUMlTQ6dcTtNLaF
GGbBF8QvH3kLqK7uCt3wBgBbyh9qn0vicB1uN4xsDIWVxz4IYLwDcNyPJaAQ/vkw
b1gkhGXvNKdkHcN2X/OrDmFeG4OZjagNpGfWkZWATNfcdLAwRNwg+5rJdLrvQ+eR
KOGyckI57QvDh/yqPuvqgJ9OALT+forhOV3tip7/1HgeW9Vww8EHl2uupYxWIq92
tB/GLBPCc2NRxqMR6JUuZxIn7ONYs6JYc2Kf1rGJlj8pPr95Onc+HICTUtAyc+6h
oG8PCW6syBego6zRYAUHLFNgQQudTtk8VOJMJyTNwnYKT1h2/ni12+Ccww1H67sb
68YzISfWeuowh9AAm11EgIa0Suo8YY8KHiVFIEWDx0aWkx8YzS1pVqpuUGpRuRGM
U7bj9wkaaFJ0EozdyEoOb1IGyP4/s8s/BXiyvD2eHwigT1g1ObWIA7y3SJhqbZKi
Uzh9rpzGZb+Us+og3iaXConMy8eIxcQ5ZUg5aOvLI/dO/LjjMk3pAEx75Pizs32q
XZwO8S13hviwwgtXCto6y6cLimivDrDcnOBFW4bNn4kXW4wwy5I07Pgk3Cg7DHo6
y3MVgy1aSzTpuuGXs8cMOUpFMyr1RO3JiKci8WD/VygJwByynnfpk6OaeoLq/O+C
MgNgk69T3MaFx4if2J5KYNIcR6PxmpNUpI4R7Cta3Tc6aE9aZbZy2sEJXOEA9puh
UFGjk5ygAzoNUd+h7O3mUERPBbLj6hSdjW+zb9g1U16l0iOXBt8s1FMD9j7et185
iBPKnEjW8uzeIWptsQYkIEYVbWMk6dKNLkYFpPdGPiGGKQsxBtrZRkRpxV+oleqx
96XvtwyDNP1OwmMnKXOAt5XaRdRayDyOuHZs2UdCgj8e8YZ1U+e4yW4nlI+7/aVu
b6NHE5U7AgKnImxZxsO2HYLCb325W/t+O2jXDtNoO2Y/KlhIg7flN6TPkOsvAdv4
WlMdgb+CEarNvYrBP+W++r1RY7xVrmPuHeiOfCoXEiXztzyAu9Car1iKdNARL8tp
EhQtWKJ3kekdXiLog6UWA6Zh2wOJtIgnIepCTFPG8utdGEap4ToUnMmZrwAtHM6u
mnua98difsK0km/bGoN72TcKeTurTbASALU2snUYDZneDdal/vnFW8JSlCWutl9r
NZWl0qFSUSYdMUSLoQjqzwNAycFC9198cNTJIbIMkKBMoB7m2JyRi20VUDIf4Cma
siqCi91hJ5nh6pr8JrsB8IYtNMs8fSdCn5PylfYR3ULGEvn/UrzzupkO4+G16SHU
0IhUeE+asFy+UggJR/WmDEK071fEmUKkckjT4H5pfAXrIkubwpfdnveLx4tgD91G
DTwIv55C0G3FO0y89O7Ap2J+tCJg/UmZ0yMvM2aQqfMqfgypBFq4By1+VNFWkGz9
htLwO2tmbYdyBwsCIYDPW1adUbojOeiuZ1ZAHpq9agPYS/33SOuLKkghsjew0RoC
81E6l0QJ45MMeUjf8Av58kdOTbKsjiqUprZKIpV3R/bcFcfq99UedkvH9pP9A5yq
5GeccxZbb75E5XmVq6jxTLTodYQ0kra6ODjLTlkcXOen/S88HsPJNM3YaHSw/jb7
zMtRnk8YR5x7xQ3ay/hJia+7+iztuxdijPTYfU1QJfH2K0X9GXibMziENbK2hHz9
uhjD2YQyJa/CVU4a0fFsvEIZVOXDPcXoFLfF7szaBRni/j/If8g/JMrN6JZOC9Me
KtyCFG+gGKqncg3tSm1VeAxlGQx7vSAGhb7vQqJY1c+E6a9UHyGM59a2JK7VpGxq
Hq6MiLLjKZkgg16ay0Tt5TlHuKug24K3OWVFkUIpb+I6H85zZ6btxyV0WCmCo4tg
tRdsxb1YdwyIm3tyVtagLAf72gYZHpL+vT0oJQikznkeXns3BR/uy47tXBiN4jFo
26K4J8/kJpWNLiIz3V83wCzFUZU26df7AADsynex/LAjkiCjVxQhMqPuCAnQkd9A
RPMiTD817+WT541JynTRL1yV1cM08QR+l985sV+H2i1bvhYhL3AqZscOJyViAeUA
PFdYsCFgD5uY90wvvVisQaklnUNrhKTX9KPTnKJvQu/YB0rBrmq5pq4BA7T7PYz8
xHsVV886RScd8F3g5P3YINDI0PzAGIOqdOEDyVMTbOMpoC5dERTljOlUAHLuWVk8
3+QT7yIHmBfCRWvZDtDAX1FfOdTKvDV5tfqHSk/SNkjRrJCCiBKgnRspRcA35Je4
Jnl+f3afISA6WTpBqFY/KTsxFMzaQD8ogvRXCaIxH/GaBug05nPSJvBak5fjnp+C
vqJ5XYKABpnm/2lyBQRQePL2llx+lTh9G6Q1L4MM4NABWWeIhY+hSpsy+274Hh9K
IkMhChlE7ON7uAfoOcJ3vj8E4WIOqqKbN50M/kJQoBHa2Oyh9zusRbOB8uXKq8ne
3NvgD8Qk26g4V+NxYFT9dHoDQRCBxwtVFadGx+9Ev5Gzr90HlcHuEcKPgwvSWZPp
92aW1BbHWk7hu/kBCXbEBF7TlQOP/UIqfAnwTLBDKE2SZ31KRjGaAJm5ymsvMqqu
Fv5/pCCkIfkEUGHlMFDGH78ma0FmVeJKe13DNCGWhiXsLYCn1ZhEU+d1yE3F2vLV
M6zH+Kl7OvCQSsLZBREocDoWVwnfkUpvuh3Yw9nvFj23v6whOMi3pSi/paZ9NwOp
DED2nTqVdG9s1D6nomGBum6pI2V2PxNv5aHVd6d+wahtH81qXBW4BfWcst/34iCK
Iu4UofQcil08Fh6C1J8gDkjtOLH44wnWNeU/cHLqZy2b2GGDifeSu0XThSB+nFYE
x7tkyoKtG3kYUhzHDoVv/LPb9CMeU/hbFepkvmqOJRTdVdSktmLobYhsA621/YWL
FSnTEE3BSRJbM6ab2TRbezObAuPavi93J+C/4lr9Xav253RmoUS4sP38EHcYfKN/
Pxl2C1iKi+DV8sePb3IRlJHrIXoEyCi41lQVFBHfohcE4wUBHPDlItVFUVcCg9Y3
icoMHp0VUqqbqlEtV7qPtJcG3D4Tkr1NqBGybRRK1NoELXpQMqPPJKcIB3xQduo7
wyiEKWx+j1lPmVtmvhf2MCD+4aQyJtlhSbNTukecW9sUlHl8gW8p19D8OQnl59hH
GbUCGpjAR3qbwWSum1zUyvzdYSvvpZT7knli6XQclpq9ByiHfbb1WHKbt8FfCzbd
vP7cxdD7/Ir0lhB2x77GBEqbIQSZWvfwxA3xDx38pefWez8uEcDr7VBpdqQWyWwi
QCHD/Mwot6BEOjgwN/ii9dBtIbYLcJrXQnEqSyVmh2PrLy9pbfFi4a2/7QojsNTP
3wTLb3pYw97RwQGxYmf3AjKs5dT0duSg0RSXNkNABO69GOpM1+4lcxsGHa5kBTbp
4bvfc/MFkcGaDyeatnoIgfNYu/tdgsoDuRFPhQ+HcSIhuDR+tbFxCIv3C1X1hnpr
VSR1SEhl0ay1Lu2WPoq16r0btwBLw2Il/JErnD2Bmz16Un8eJoOIMcJ1ebBvm5nA
o26umdBmQfRGPk9nuCHsLWt0Jvv438CAsp0nAVmw/cHoxjAgbKE+UdGsVxPUmdjy
fhXGMjhlZZoAM1si1cPjZntRnMuOr5hIzvQpBIj63uhixcOBxeJ5mpUurZyxvSTT
5YFMXjcuswigRehDN2lgF9AcPfHzTD4wmtwCo7VHird5Co3CHmTLrk4/tNfjBljk
CDADeBsGZ+3htC+BZgsnl3Yakb4451fMNiaHae9/xIlPJuQ1dUBjOXbNRb05Hp87
eH8XLGPD0bDJQ1AGiD7ionxPoKU08f5dVMyiyNqBkWq0bRyNe9EEEacjNZ/8aCpi
DcgRSj8Dcv4dbXuYQTOQPbioY+MBHP1Z9CnyoS6W7rPcfZv7wV1nqc6Z2h4khGOm
DDOarz8Q21kHMP0WLt13H2BFBmIO8E2rT9C6I0xXziWou4kJdho8NzkdW4lEBMBZ
A01n6XitESKlQ3YybbUxlLtUXnPLdNcEpQKK+O3kmLzzX37LbnphffhDPe6ipime
b/a0zNHeomXwxddj0fM3QUgorPR5/QxrviLrR2BMxitwfradlwtGbf9GWxFrWmqY
Cizd9ykSP+WlW0Yl9IdR0Vn1ysqK8DmTuojgYzK6/UZuuuFNs70ogCou6W7z9V/H
0aE8sw+9fic/PTWI7MmpR9w3qOOyk1MnXU1ypeppcM4rrDqXi70SI9uX63+hpRJM
yGPdaYdX4ADMgfgvjJsQDNRNmrZaWcJYcZ0T0aOFfAC/IbyLLsmvFrmdNSONi5Ob
mtO60H60kupwLaVYUvZAOVWD++bDSsHouwMF4i4RmRAD1kzmzayvURJdR7lm/Ao0
qOGUWwf1xR6ZiNSLtnTNZshsjgO/n05BWJYg3TS65obnBl6DcIl6PA1BnUJvNCbb
vY56Z5hkcfl4NOs2SpE5c4q42eFWFyLaxrs3p02Yz7IJgBJhrw/9usGmFMurYWNg
j5yi/SOCsapsN0v4zVTRP+CWYI4tFhvHmhfTGp0vKyNv2lYd0z75srJvBSnceTqR
+vrhvomFOueJuH8cBA9Vw2dVR+xUuqSjy66TDlzuhA/vQbGDqjivFOrzYiTTrKg0
QdjXUUTil0pjMTkpZqAomQKUXzOkgHIV175akn1PkJEO9+9fCwLLm9rO1I88Vhor
OS2obg18wRVQN/YogghvWGjlMKTG03NIGc1YIFC0v6WQpo9ziY4/u6p/RbUOf73D
yZoOcfCrBOV/KXuvffxgJCYbSHjLyFPhzqRbot1C2GJJRAnTdiILTyeFNFDolnu8
tDjuZq70sgMIqMCg75wA90z2bW06o31GhLO2mpG88o0LLKrqM3uuhiHxjrP9mrh5
MNZa1RIts/JxoRLRibCh0d6GapB+L2cYmXbfznVrYPsV42LXwoCBsgBsI9FMMHAz
Tv9P1eOKdJBHUIj78WnNSeFma082yiQJXgmU4Inz49p+QHV875co0LKgOK3YLDm3
I76bpuNpsFDebDaBXj/Pya5XY0idtfRZCmRhU2tnikEyab0aw0g5Y0h2o+jCHzQJ
4K835PFgg9coJmubLJCI+tX+1W+6claT2yphm0+h6Lryiy133KQ4fdX3Sjf+yLX9
kD+D37P8qnUjwnyRW+b7nr2YJ4T6CrgoWe0LSMn+lrx1uVyQRClpE2Vw4eZENZaS
zdDz+0R0d7T9+Hruwv/b2jtdz5uDiSxNayB1hvt7Xmmp+MFXGRhdi9rHrxLchH/x
dCY2Qux2fAC+4L6XuBzmQjD3IVgQmjt0gVt1jkmVxwa3c5oiWlURBArJ0/Ppp2x7
JkMyl1zFSSbHlfSxH7GWMF5+E7BcxQsrHLWo6H7t91xUfXUxQHKO+RHf9XnoOVMz
Fx76LhcdQ+V5A/wfz6wAmqnyN8F9tg987bZe+RqYa0ql9k+Wis1qNQJsct2kegoW
OmSoDxOZzbHB0PvAA7LBpYbdWRmRjNqrLCAaLFjH5qmQWlSkGXb+Byvlcz+9BoS1
TFe7D2PVAuwsGKteJ69COS9XWs3aS/hnd8vgI5Tk4BZKaLJEcvgKwW1LnPXhU+wp
HXxttQSPwlaMO86rp+5/KuikR4BmNP40I6RQ3UgVBcft6DH3zXZSd86J7EhhFGk1
oQHwelIhi1iBhXmOcUPJcKRVA76wRU+X5bJ1YmM2/maD+NQ+zP65pkNnFKnqxJoK
cuNjSJxSx2ealiEwI1Ug7dTz6/DFVr+8ZIJiIYnecUcoExZrFRgLZUC+Ktm+Q3j+
yDSBBS2AIN2ICw0rMG9+9usSriRcdLKoi7jjhXrVuy/G+sftqwY/ozp6eCUCgV1a
5O+dp7Dy5Bo2SkrY0OVuOnSosMMsBMdQtW8/pD6E++DPXHKjHf8YUqR4MHAzZRQk
s0/Nv/jFhEaSe66VHtMiKxO1+SiJjO/Lu2JUkZey6Q4tJGiuETSqZcZw1LMP3W9R
ZtzAmGXdo1jRDrrhsRvrjBaQa7d8lW90VqcTj7DX67bibHxfli2vna9m0/g0UMk0
0IMZGxfEX6jOQcxu2x1Y8b8U719u2uuruET9yoy09QYh5/a0+EAKrQ+7uhn7e/Kh
vWf8/kdWby7ptb2KvXHeYQostl9QzaCLD/yHibo13xFReS7DMCT+9DHoz3n89Dvd
8CNxusQay9Hz6miUy9JGH/7aqvQ9twrBWUOLc0mw4dLHZUxoRgYIJJFFHRHp7J3k
jW/5A9Ez7qD9k0FuSjdHuC23pETimENzAWTWIkgL0uN0JvWvWViuxlA2OoAn634C
Ikwg/MhO1osiiUnmTCQvjDzooxXB5CnDsQO/nSuk1tiQXlPIBHvYT4jumNnn7Ymd
wyGmELY/Kkt1XEHygRzVxUfxeqbejZ9XOEbuYFs3Drf3FHzmkZHeE2Z9GsF/8n8V
mW/IQbmoJ0R6W9EgTkE/+zRkHH6GM2sqiRW+PB5jnPmqKEq5aIsfsSeDnLJxiW05
Qpcb66VC9xfOjIS1fMU9u2GgVgharzAYVCD4Lf0N0TlaJfeFkXNoAfChmVihA9Hj
gsSw8r+yqzp/6Ik/k5w4Zegodnqxs6QaOE6vQSLDT1O9XtlQkLrBYPECxtB3qoKK
sFvdfMcJVG0b8r49etThu8YnrMHLQTWCaaHp5M7H8EUiZs2JTsIdqb1+Kevon3qv
M6/fITbcErHD0PpHz46bRa/9Cq03xFVr6eRTNiKLLVYHr4TCR604ZO89XUBQDWxs
ecpvlWCjJeXdIxhRSMTkhDw03NnDSREGBiO7BzbTgFaMqzBlrg4DJWcO0gxzuGiq
PbwXcTQPxJ1rSZAZhBuG1M4SP5WPTXaIVEpnhSVTTI29amQKFmgKAQXDBmQpoQsk
mN4srAd3Vf9zCsPXgsjAAvxQGpEu21dAOwJPRpkMPGOEGgoxOlBrD/7dJS30Pg4C
eBeCjbmjxHW20gShAQiQFpPaxfG70K7zrqFrXQiMlkuZg7bAGirf78kfsAUGorND
aJ7GysDfFNiO3fEecVC/gIdWa0vUTuFesi7vn9Lz8ThaS5unZqRIVpMudvBXIYfr
OtcbCzhFw5hhRCHFCKHZauv1OeApAAQRhRWyBytpPH+VQ0Tfmhf+WuCgKLsw56qL
WbWHL32VIcIESBF4pSswE4TNBZlQS41Ckx32GnrEzaS+PzlVrOYcSTGXHWslu7Ee
wFJ7Lv6RQXSR3jpv3sHmAk3nYZgXMYrVz514SjvSzEqsbGv8Dtsq+ieMqIZ377ZJ
DNptHQGmdzWkNOty98IqAmJYNBK6f4NkPKBKw8LWzc6nqIe2rgViuCZtb0yIVSjf
tO3umAuk6cyz9XVFGQjkLMm2MmfYlQtjZAjRnX0e1GHvLzVARpJl/jAt84Q14FzG
Qh2hiBduUQVMNQtdHdpZUmym/maRweIISgQtlC0TpHcsurgYKWXvaoMoYb8YN465
uRBxlAw/SgQJ/pfTy0sIbtKquUqN4uli2ZiLXBAFE9k0nTne6H0VG9lkxJFFszUq
mjkwi2RVWPtRHKRUzR/n1LvP69eUsJlrHsUoVWXSmsvDQo7KQK5cke+MBkI1S70U
89fQ8nqFkUOIw62giX/qqM0CeLd9X4ZzK/HrVivQTaBuG6ev4FqxUGqGbxtTz2LN
G9P/zhcBciro0sRfNSL0RERbYtG1jjUWHRM9JFT+DltVaCwbjZBwdm6JKWhsKVZR
u+TEdNkLaUKWdw6rw14JXLp/qjj4LlwcQoe1J1xc85TNG2WP7764ex/1Rbrrcnr2
ePJfa9zsqS+K2BqpOMYfJn1rnPLi+HicFQujR46ZxM+R2qpkMDwrUkBJ39XPGusS
DPSZt+S4N/yh6tWGENqScFRIB8Y8B9UqtDZZWroZTSV+KeCjaWDgyYuZk+4cyjlm
fX2G+eMN0wOPP1C+ymSrWcUqjFr4irhEOT4i1tNOoF4ruLcaj3HN7fbs5dJl8M7d
AMr2a2U6KUDz7f+kO0JLGzXFeSGTfn/dt9CyIztqvGiboSskj8Hszb0H1eTwtaPJ
qrPhHZzvfUGoyTTw3JFU0Rcsr0f9p2/b4SVtVL4oFo6KH5WQvEjurXI/hPoMtvN1
kbcx8dJWEzjrS5nK/3ZF8lbDVXHa5QcxSyQmWz0XRVv4dFGYL4XWXltVETnHmR+D
GPmhGS09KLICsMu1PbDbCpCPL8OiZfcqpTipSI+Bi0fewYbsLuTEUH1XWgn+fh5+
yznW9zDhDZPdasUjU1hYK5p5pgeW+GROIUlI+UfIWLtbpKyi8jM+QwoccDx2Evnz
ZOQfpO7BqkWgogTO0gUMubdGl2wP0JoiGyhSvCw7iHYPl7phaHjeJEv9ANJSHQoM
eAc+awmkI7PAq9XO6CttU35dRnLasRdDLxmcNnWQeojl2CE7PbrK+i8e+l9ZId8L
4EWwAiPc9F4C8YlFGZGWkkxdx/yQUUJPG/DXUokYguKEmyhKW42uIjsZ3UQ9x4hu
WOKUfzrlVUDcthp47lB0uEheviCWhbmznar+n2wPp6ODBNGcpqlpjG7yAxKelYWJ
9oeuQz/lWwPNayIb7ZhXQwsnvtSqJaPjZTiipGYE3CvW5nFVSV7E82LvhssuAn97
FTDeSVJTaQJAcC2SoEV59Ezj1iQqmB6uYUmfFCSRrXgHJ+t21UtolO/Xt7T0osRV
+Zh5hjqlP8+esJFPzGxdzIl6YkxhcGHRjE+QpS+vP1ngjLNdnlouTTTyYBjPXKnO
42TDPefzlyT7bMb0ZNGZKNIaF10bj70UVavV3V62gSr28T5HZ2i6L/XeF2FgPmfn
uObfpJ6e3uLKWCgiEFogi2ym5kSVB9gxOBAt17DHRULUSzUxm3yB3qpFq52UJvWH
pvVnvXuWxJx9unfG41bXEDy82h51AXxhqm+jI0RbI4yl7FDQym7AyscmKlSsXEPy
pTxf/mHxZ4EFOHRcny1NMTAX59azWbckOxjdt5Je26ymziUuchqVPX1rKJou60rJ
qxm1spiKG73+sqpPHBcwAx+WTw8ltw2Gd6IIVwPQsA/2gQQ9ClVEMQNqZb+S05x/
Mg8RPiG+DREg1+RhB+JbAudtDacRv3X9RrE8dfgIqdZnx34CM5RywYa8jDDmv/QP
xepgdkdFO5gYPfQLxpGOB5FmqnriNFscKMahPflAYT35MLrtKSkLjW7W1CIAiFcc
r8vV4I5XOuoCS+SDMzU7hLWEFmvhxI8fBEm+3ereyNEgursXd3A/IK/vdhgNa/YO
pPf+6XX6JTndBhOECBm/FM2ly5OCrTERwUWbasiG+RHdFRb5WD13WpTGMBT+A5tt
I/pnYpQjTEK7112V3tZ55A+bYqTSwzeB7vo/g5t+cVzYfpVR5S8NOeT8Bmf2rmy6
idmLC8Uh4gDEo+6HCMHmkxswqTDllqU0sA1O4YZbGFuoBGxYj4k30AQu135Lt5JD
7+c8Jy84L9MiCEr6v4cdHIyKeb/+MltabdCmtMGMYhWwfQGopObF3tSp/im3J7w6
Ry9FlSdwUeBjLn5iYh7ewOA1jNYO4x66Gg3NJ7sRdITq8coi7mqK/Av6wVWz8NJg
q0zsuaxVRalsKImIekoYn7deB2PnGow3PAT1Rnip8D5LXcUA4pTEkT9zecwLuMx1
6yVYd9nvELVh22tkkyJU8YmzDMMoXS2jNGgAx807h89Eb7rv0KwxsExTa63hv0Ps
JlWkQBkuLgN64KSm8yfHNQr8x+gGW3NniwWExXaN63ZrQiaUAEVQ2Bye0+rdRy2P
Kdtg0J5XTauyJY6Wo59j1jFEPhG4f6dUnIGvQc761K4fqe5NAyUa6voPf2tu5Dpb
kBf+BWqN1xKI6jdkCuYVbZk9/5LqplRRHkNHAM1SagGuzcI2cgfE6qKZ39wIy7EX
rrQ36Nw0Ci9+gEuGWtJiGSaga7+x1DwFLZdf/kiwCfdmDiRmKX7I2Du+39VhOnSh
AFnBB3ulBQdVYGzUHqnp8czCCxn0bPuTtCvmVqwWFNapWayEnCV7wR6gChN6qK6L
csXiIts55kvq9rccBc6xQzmYomYXfffnDTt1hoTyvkRy6mRtcdlSbxFPIT91RkoH
fMc9trS4d89LX/y+xuOSqVfWoGkCuQpBZuILWBaKWInAZrKbaOiR0pou0Oq9+eU9
XFFBwp0vdoqOIkFNGKWmwppezk3T7Y5TqjPyor9Q+TZ2zrPiyXiAB9lPSuIxk5AG
Vx/+A7elbC5ERDLh1zlCR3+hLxEz8tKekjFjNeCsYmXdsSAhh3s9T4T4GC9ZsY1A
sfCKWGggs6fTxkOpZr3EFjh86Pucol1/LKMds0Npih2DaYDvkJsh0vtwseetIe5j
FMagHuGn1ceeMX0Bi1GYUjg0cBBfrygU12er17eEeWS3lCBg56CWIFzC/1/BXs2/
fEhGx3gU5tmNM1k+/cRi1saaBwfHQnfZ35qI3UOytBo8hyWQPIyZS7KztJbnuUEJ
p1BfKVuc22XvjJ7m+mbwSCDBAgOqTwToeItKzbQw4wSdtzNCTrcE0OXAgVLMWG6D
g+1z9uITrT4SgtfdLMgSeIty4cEO9yFL7b1OKtJtbIj8zAWlTMh/8okiJJX7aQmn
DyTt9jZY5MafvBCZsaPWhs/l/FDwnw5trVR8o79Q0N1hlglQStIBPVVGAJrT+aVJ
KorN/l+9xxFJoQD8r/FlzDeWqGE9UfoNbt0pgJOxvWf9qoMadMw8cnz3gpgKn6g5
e4Qc+bfk/VGaB+XbtRcluokwPjuPO4CoSUC0J9+Jsr/z/YqWoGfpVooAEYZNZGhK
K7upzO793cj4G7SKD7I61pMq7COlHmIv/gKntaL3vLpdKBXAXKad5lKYTY7C6UVj
17JXPEO0WJzSkY1gWhzw8HEH1eGdUvDYMxZDn+sEYwK+0s6zUC1xqUkHLrFTJxWD
HaBZWemcHzC+5l5/Efc1jRSZM1M5Fzk+Wo0ZoXy8ICcKwXGP95HfRWtpaON2oDjN
O5C2EJhumyKsMxbmY3YnesI4K2q8ItBp6FeE643aG3H80X117nbgJFrwt4VQORlH
k4uPxgFMovESvNEIiyeDvFBd6shhgdMoe9br+PR02SAjWBUoZ46klhF33nljc7rZ
EiiawPMvnZuQbKcB1qa9Iv80HVdPblAzTGs1oynFCG0/FLlihV4xIVrLe3bwyaPH
iHldukUK/mIE0it7mWOGc767xHeyJcVY8sFEC3x0SeQ7vDj7iARTH4nCoAYckVGC
MR/mGN7+shs3d+0nDctQt3UIdW0UcTr5ZYTEdx5QzRf5h7rPwUes5b4zDJq1wIXs
Vp66GdYIlxyLnryfBqzlApQjhgDYL9HAJq1t+1s0r/QoOOR103EvWlI0iiUDXkal
L9YZOQuGgtHWFck0n54/Db7zC8tc89nx8CrSavZnSZ76nZvxo3W9dFKI+bzEHRbX
DXOP86kj4gf6FmZjsWC9tbcEE3+4zi9uI+FMnToVkvbn67GNVSpj08TSRB/veLpB
uXo6kKptzRFuHHJNKVxdY+BKz6oArdJwUNSeGqIdsBwfZyBHqX7upyG1jekoxkq1
vlyZsxfho4hNge4dUep6UqnuQfKb2eAA010TPa1yJ8022wnkBq0qPPI4OWylaXbF
B/7VNhML8L5nD+9B1SMM0YI0wF1bDFrtE26cAcicbiYdwueitH2xSuQKa9U+sHX1
A1Dri/ZIy8q+/LF+cxEKFaJnkfhk+zvKUtXXzTPwkyMeHVK05ZwXrZG43gsyPv+r
jjCLD/rxLcSIkgLgxv5xiUTx7i2C5R+bE/dnV3e3U5eCue3TBG6zJUxnfJfFFKxB
D1ISU3GjDWji38GT8shrrnLxUPlUKmjYiFLLmMlmTFdhKlenQB3g6vewYTcIglqE
7l52NrS45uourI7mjObO+6DTVeK+eOLLujTp6L0hJkuCZgYRRsUD+Dggn4dZTfDw
xS0xIDYGwNvUIqBlPN2Q1TDhNQ8vp3cp6Dd/kyvvbY2ljbeu/ZZ9JVAPTcy3XpzW
2EmIkefV2oKIOrV0LuZOqea4/V+qpAKg9zajZqND44dyAC2qcLFld8KxbPYfsfW4
ywLcDamEz1wIIt1zbSGUYkdcmpQLQI1+9hAKT1DqxBfaFh9gseMOxMwF/pyf1yIE
xtwdVoeb3dqlcFG7qyO6Oq43lgkkSoSfr12tcuDlQOg+N1UTMp4hs9WWorV0OH9T
ndJU3iX57hq0joppIJnb6DqsHnTRlQ5ihFT3QP//k9tZ3u/cR5Is1xP7yvlggprb
R7yRbI4oeTMAkkGMefWgxPMSWnsfhzZGNltjYK8cXcCwAOyGYpxHwS263OA2PfTl
50dirHRFkgXNbPnPvPfXJXIWYmvOr0zz3X89g+Qbu6d7ti0h9VWmsFNJjH1YCISu
gb4ZmXqDSBHeZ4DvnvO+cliPOT1SnmAj1QYPpjx9z45CN2Dj3Hx3ADxMSLM1ifHo
TTjSKGfqIvLqSL3YjqVOGkpcT5TO6M093hUhiK4sp3zzq7oWtjQSe9mtMJdRWsSf
QOZs6xAqEKCY2Wii86GAHufbKN6R3/P7CP63tQBizgHHWnGubzPiR533J8Zd+g6u
EWz9E/HPNWlcEB6E9+uX8rUpfFIbQ9S2gwGmFRZl5NwEW2DVZGVzZYR8rNKB/WDp
YQYIvKauMGFILV6IeP+NMsMwfMMsz+fVF86Z2sT9RdSujiGi4anw/HblQ9r4tk5b
tLikwK3+nlyNXebT1bEDrb6P9Wl2D5EUg3f/vpyI19forUX0HCXZyZTGDyVaj9+H
Ws0lUV71VmOH/8dW9VoA+JDphbOcU3biWpFT3+FKP71IkHHleeMGnEoLLrOfJ8pk
+LtInS62GS/RLJxileRye1hWFM0F8ghdgOOoeJb1s95W0lipKlZifNejT/Z93YpE
zEgU00fXLnIawzMaO/1mzqe2ZqeT5L0f95R54dcI+LIvodKq+BDnGu/+RhpUudb9
GZVxDdMvhbamU9ITmLyYvgMCFCuTGc5XZhb8KO2eJNcPj4eD8uNEjcLatyf9OxO7
vYA4WbA6+0OQ0ZMdkgK78Ns13WrFFvFGWlRXrIrWnxZxjIl5lJ/JbqLawGFdfYfp
193PWz8xUJ71APBOp5vtHA0q6NFz9xQQGQFtSG1IflEGj8nrZA1XpcJESEP/o+f2
rx/tvdGonsMS+VvDBeeei5ELmr1O/+oEV2PyclAmwu+/JL3F8blADw0omnUbXU1+
txm4Y4sia114kRH4XJNus/vM/V19npFGj1Sr52Zw+UhXBXYgmgdEb3maC8qvGdRD
vkA2+KIAunU0B7MRdd2YxPOjHIiNA5WKplpm3Q/Lw2Wfhk/XHNh9SUHrQ0SL8LJ8
iC6JQWSkHo8xwiEoJOSQ9ueSTGGgGNBXNoaNGLcdHieoJ89wyVZBmjmf6uZGSjAQ
CbkNAcRRrThwCOXxt+q0zdNuP4aXiwFEPF+1W+N88zpD6YZmwwU8NMrUUIYQLDnJ
XHWISzgKSGVwAlPMDTpTmVXWjDav08B8cGhEt3RH4zPfZXDPQErv8+8GZzUletWM
VTDpxC/DJKq/7+uC3d3y2qqGAKyRSlpUY7RnPVzCz6ELHCJ2On7ebQrCFKW6sJrc
+JoEuGEZf5MbEGA+iOvHpIJ4lHRfeXLpbbLcix/GiCSLpvrH/eCKHmrO4sg2pI9j
MYamBqKWUIpRusriDK8lAPwo70/zI3hObgv9LWk6x7IIFFHBmEREzXYaPbMTvB8K
HrVOQVm+6iDJsArgzavsrSs0hju2FgvJuZzPuz6VX8vd7qtgQRlSSJOumGtdutSy
x4mJ0tXqrSIR3ayhC7KVjclRmJo7Lu8M7b29RVTSEzpedOvp1FefsWYh3nDj5rpQ
4qs9Cr/Xdiq5J9hlP8W1NMIuHleJV0LudStb4wMsPpmybFOzi+VpDAN3OV/ZYYJr
oaB1SmJSHLEkf6XNSSgWv1v+i/XtbWiBDoQozsrsL9W0DNpmmMwiTUJ/Stho2oT0
goTpmJncCwHVq/v/x3fiFGArdUwKIr0vG26C/NXaiAsE+gR+hzQceHotmZOwCkTH
7lDucShdi4WDCRTh7PM1NwMMCAXg24CZ2ku5oemFXaEE0qHNq7iDD8obkOg49+2d
Z1SGnpChgf3Jd/P2fjW0Epz+I92hW/nl+UbX5g1f9ZQE17wKs93m6Ukf2yfv1gzg
U+B6LXxCHiecb5J2A7pWoV+w1SrrHVz55fa0qhfscMSTVjbBMJPkcFCe9Kv5nhKe
iysfLwqiVmS/OApkBa74PmwrOyiUZBoi0zBUUTrIOYnch5qaUbndEvMPAPLVQmj7
NhW2O/Kjb3z30JgpOhMC273p4kCdDoPWV+h2MJkji3yQX65HFA+/D86Lctt0XBC/
jPHCbW2/AAOJ9l+UX1lGdUx7jDWsQhw61zjz1/0iJs5pux0MGm6d128+vCfLiWc6
K3zylBqXDEbg/57QdCrXymQ5aZlp/u+tfAIsCkeEA9KHPqVapjdosFGXbAxaCsHa
dMgV5JyuHhnUpL4GoDZSqVoGWGLL9KtzutuY9w26656olN8snlVnq2xpLSKQzXLC
q7d8MhjQtJbPORcBBgWb+spvrwMNPWJI7CdrSiQwcyN5f+QMoUj1ISoj35riIoJr
yX53DP03cDj11uEFeRo+aaGDib5raeEJ3n7GVh84zgCoTm4AWnDz1x3ru7iT78fA
qp3rEXNaW6hBJ2IRZU60wVvEDfkwkRwh4B5fP1/Kl3YKPag2EboqoFTUacLyChzs
8ljHZ/TBbo0+LIOdAqf+Jr34Wg7cW3rfwe00B9Df3WK6YUrjCxFNCgutvF5uuib4
ym7NMHMidJ/I/qmVqV5EuNvF4T5xyYwTzrOMKQPMfNMcTmMMXZY8VnjtqMl23utF
HVHTY/SnYYcRCQWBO1cA8PUwkg+U0zoiookimuqS2VQUlqqweybHZ4au4h+0s/rA
Ie5u3J6Ii8si1XkifYZfLAcCc+PTQ3PWVDUcln94ZpMvdnm1hZZJfnSO0QiEafgP
JwCupDKlw7aTeVrGu/f18JEpQbRYMNN22UNGZ7kN3kXDzy0D6TMDCfG9DZeYvNVO
n9r8XruU8xgbtfTHUK3sElNS8ALNvF6z1EyqQGVX4aPNxZ2fVoy+3+e+cz8Yqbez
tuhhVu0qzPo2zVMu8BiofEzJO56AXNe6RbHj7wmExaith7lPTpICvaP3kDxnurGI
k05ul+7OCBtq6q9U1Rdgp1nS9eXTJo6VPCoMPno4+ESmoAwvi3qFS2FP0s4cFSzK
wWCdLZmYkbC6dqfhnj8AN6IC2wrbivgKnYms0xqcBZ/iaDqt3x7afYsjkXUdtlOE
feZRZf+g+j8varFRhSE2P/cbBRDpBjNQ0PV3Jp1Tf+Nb1+1EXKTggCaoyaocBy2K
N8pt2IwvNVi0RLSSL6OYVAlh/zLDW0SKdHraKpSjs/W+CcKlUBosGknV9m8NHKmp
hZB/NhglNpg9IGWYsNjGO9APBya/QfCZSVb6YcKZ35/Oo+10I2xO3JMyXU7OjtOB
DRSM+3BTpT7q5y5dwL9pAFnVAQ7KaXt34syhEe263GVlSWAGUg37enoExHQReTAV
SQLm9i044zNo50oIeHmYZGw7BMihopBoBB9ejQDEDXNv9XjMxLElMYxTXvDE/5ah
KtKZSg4wgB/Yds97BRqfO2u4E5Bn5ExkmqOYLHWTn/Youopt7ryr0z3Z9ZIQTm+A
MZdWu3r1BI8XHrODMYeDqNpFlxYnwsPbbN7H/JqGkoEtiGTXocA3tYggrudhN88h
yzI+QoFsyKTcRgmFCME3Nug7KXeE2a6C27dYi9jqtN9diW0ki9Nlbl/J9Xpja8rO
rIlW051F6ssBpEe2SPmlKMCLEIrvjml1qFV69++2dCj+o3NDIfkni8aNy25hQrIK
bLHEy/7PGFAB6H6tYHST6ulajGko+RpZprzjUbVcUS7E8inmCZ9iEIkIlFN2UCyP
gbO2lfAlQgTawIaBX2ywwvm+BPQHsoADFLqC/s4j5a8azcgv6EAX5elamLWxFtV1
aI/+XvIzgTKNOKzpEGYilV8hlssdemgvuPQgiJhHCrpVmZTjGWXurWl5DE0FOcJn
CqVTtkrVURLkhq5lWoYijwmCweFOucMODHUE057Rz1xsWKQm9u41hy7j2ynvVguW
2R8x/k9l2ApdPKYkRfK3tZCywEB0I3akfP/qcDOGHCPBSKiDoLpjPHxAKZFyWjAk
Ufx22KlM1p071o25OnfoqRVmkDhpSvLSk7H3l6X/uKhdyH5hwvRrujTw3uHGcdHa
CZVU0BLowNPAQBrVkkB0P2VGpqa4plHggmzJjl3Zm4/jht1bh7GRnZQh3aSn7F/b
7mal8HRPYVdSmSs54ApaNo5vuV+/5C76aQoKVou4lZKCYIS0rfz5ROG3i0HMH6Gb
4JRfHuQslZsQFeGheeslyr8/cE11jkrXbjDAyDmuMmQqOXBMzSHM2n4ltYAc8SMO
vEfVxEOb0u6VwNDU9UU3fNRN0BFwAhDANDOq/U4H33yYIHcsRvCMRyvAfqXxJq5S
P+Tq2zdJSK2pIV3b7vfRU2OzBsNGcTzHWkQXdejey39DNs+5/uUfptFp1/fJOhno
8O2wLuRX9usWnKt44/wPsd3MJ94zHvuWEAEHlE9tjXPS9hgtTZ5G9K+NI3tdROHo
JTE1/+VfZVZH2bNA/U0xLiZOIwzVOe+RyQF6H6A9E6yhDhaxfT8PdlaG4EJThKi4
XuC53p5m8CENJyOvBs7xnw6A9b+KvDKYItdQMF6MnWPw46qoGDUW17xE3bhzg213
TPA2w50ib9Jep3dw5eKnQK6QLAipPUdxi2ede7BLn53WPHr+NcUtWrH+SeUpdeNh
hrVr4puFDAspvS2cr4GTdiKKZa4Nr1CxnYIvzVX609F+p9bkZojszbVSIxGrLiGD
0Jqz+vhc0OjAipAFzpk4ymCkz90CFQFDs15QNX8hwboCgOwm0X3CMppkDVZEKHVP
N2WgU1UgvDu2jew1paBcsGE+jqbhZkM7kBxhPEASZlBs8UxqUF5SDLF+bWLKgeOE
GRTMYUBeJLzYVWx/0owLwEmhOWJMYyg63J75xj1BHwXTgYC5JTycLLzRZhkW02GA
VXvYD5CuxramsvUyH+cz16WL4/8A/+4Xls7EmHaprr+f8QL2gnsH0l23PU3Qb7bN
I7WH1QU6iqhhN+8WJz6NILLhfU5iJtzch7LlN6+5WMklvWJh0ZgxBwrDn2mh9Zhs
+AAdScol4WstGvgTVQjylwHCt7saKGf5N1tgwjNVpR7bWJTMEzxU9BHqLeAog+/X
l+XyVJvwmDQp/YMIar/1lqUIqQpiv2IkOBeFmvr4c8k8Badc0rPMsKqMzHBYteD0
/6ABOpExF4W3oKMrbioG0E1pMtsQNiSjX/9cIkTL+Svtj3bUvn69iX3rRwQJpZ+7
bzmbBYVG3oLg3c90EiWGnDutOSTF/jCeSTMvuWNo+a1V+8DfBHJzSQRcOVspyKrP
fKgSP6dgwDacgq90YRCw2o3Ni1G04Plgsn24968Cov1tL37NDOuyfX09deeKSzn8
qY7g5VA6feqd3aiV23fFhwdwAOSSEWuXGFs1qWIkfZA/ofnJCeYD8susiPF5YLs1
/9epA4wDn+HXajAPBVH/xiRyajWrZn2aY/XFwf8NzxnP602ZcALX83Vgrqg9BvgS
+pyoyHGk2hwjV7rX9kq7LtpV7lM0OTHGjH19Nc1cYEqwM/YKuP1hMuuf4Syt98om
emJhUT+CuZrQHk9eUGTtHOwgm65eAjBDdqD2KJtvHu/1pg0jD2OczGNpsS4iYCn+
fBsPK6EoYTvhKmqwywQKH046QFQNgjQQMC/La5MRDeACecNApMCRO4n+RB7nAFRi
1ImnkO/lJlVDWeyy6+beQ2OGBxQ2yn4pfftxdXcgec1YVUDGiRXgn0H+le5J2wc5
rBUJLWXRGtYEfBff3Gnvy3f1Fo4bovcG2d1fdowUQFMioZIlyMg+yRvcFT79QRPx
rcjOv1AAfkDZHZcRT2gavBl8DzQCgtNOcuXm2yF9PevkCqR4oi9plVElG0fqK78H
HOdeiiV3UFtqswUFEDHA57BHU9fwa2DUkNME4iVvhErKfnAZWh3rjP1oNOP6dahq
uydtXMomC0kBdTMrgyQybFHnS6T00MH08wxEsk9krlfh7tY0KhOo6toQozujauzE
8w922XUDWp83n2KJdT2n5ktNmG12K3G+H7sUXPIdZR2bD2pNlnOamka5hhCzwn19
fcjQFat4tmibcgTeCZ6ab8ufTUOPsm51Y4Z0Q0mnrPv9sww/UAgFBGZs7q4/y9D0
x9uoBivJB4dEpnFpUtkIoqwoaMRS724GeOFU/iCujFrghsSryEzVVGOxON4X7Vtx
k89N6+RQ8VZr1W926IOqUjT8IImNHRdnf3Ig3xqgoqWUdXOcIui8sG6LKNtxE5lg
OqohtJVUJtoZKqgrZtPK/lgoxkBkAU3Q8zE0jRwvarZiPbrcKublfVgSqgz6K3VC
U738dRYLReowp6XampwETamZ+IZvfT/2g2OAZEsE3c27vmZi9JGZPjxQKyMGJ4F4
rvCSlVbCxP7kagzqUwMexJMo4OQ4csmp93fa+vNysr88h2EJhmZrSM/2wlqzsUZK
CdqBAHMZyU+GkRZVBzRha2qGCCP7oIQgujeRBg0eD8UpX5qIXMuZZ++Weacpel2m
IByWsB0H74lxFDiy5KhKBbH6JTGG7vA5HSOQwqBOIxdgCJ6V3xaVLaJ1d+YTJQJU
Vy7CMeXJlMWE2XmFMuFfGJXT3jXdbZ2udI+v90L+5po0djrbgEEm6NtYtCvCAdeo
yhdo5TBupecH9x+JRnHBGWeVaLnHoEG4TjCykPJ6/yoM2T3BvM7fGCK4Eqb7HpTs
/WYRwd3kFlyFyfkXt6YCTJy+k5/HXh1ZbPZY1renYcWOLu5zzZhhg+xHT5CkOtbk
0Rb9O+eNLrLuWI7pGUJyKgsIqYavCZVTjk2nrUuPdS7ddVdRxOV+en1VokeYuzmV
MUrd7kqHst/nXoQL0k5lfUnAIofuQ3nKod4r3Gq2t641pEyl4hipnWg6VObScd4P
mSrb3GfFGBhHxKBimtdHyVIiATh3utOtfBazC1Oo2kMoAG0hWgi4Vqd1pSYroml4
RdnVi6r7wuWLOVrN4x0PLwP14jXYLBMrAbC3JGuPMXs4chg0Rku1DLW1kfxIGAgp
p4EqOybR+kb3TeL0hb6IKr7BsYkCdLrFOTdJwPJ9oocdtVAHyqqSWl75ayjwol0s
T7w94LNzpT+qqTBy8Ue+sm5vnUPrNoZcWQsjd8apE7ycO8XEvfSE8aX5Zt3OMzFJ
EV+pQk8QraywJJoG5xbratQLks4HOe/fcyX72vjlg/471Ta43it9HaGV+H/eht2n
SutTAKZ/hJoJHnqAWH8WGDt1aC4rGoH2gN1r/bx5R5t7XxiT3IdWfge+qGN1XlHs
sRwU0NK5RtOYFHSdm6VbsulFAUgr1JCo3ySiv0k/baIzv3rGK8bPC4MyrfptUGK1
ychaESMyiTeiSKkYvVaeChKRJ4JrRgWvo45amUJed9mzZ4DQS2cFXm26vgqFB/tU
xoPILlbJPbf9DzvCAkCMwdMKcPZ+KDCjbl6fI43GVCB85ci1i+zSdMEoDel4+l7v
OL3rSeeHRpTPmZZ4j6+VTRkYFahnqpckIm2w7/vwDr6g61fZ8s5V0qh1fIserktg
827jLLh6IW7N5vX5joqvH995kW1D9lZ9065pViB3qykxcLhB42q1Ge66Axgyh4Oi
UFyVZAV2n289U89udIh/viVJolj1zoxDBSj7VcIsjEs2lpmFuaaoo9IDpiO1geTC
kYuh7Vzs1izsYH+ueG0D2QftB7upBsze4U2w178EFq8CZ8iS3AQdfSnprHfpxpsR
L+29a/PIQu4EFDTO+fDPG9Vcz9FM/hC5pCWD436gdLK15dxukob49sswx3zQ3sW+
OxCpuMBTPH2iWC4Vn/Xwo5AhuBa6n7nmGx47J9kZn9lFOIpicQ9ZZSfEI7d5S8ot
Rz7v75I8fbkPEYs2dpwaGhBzskXc3qZAVdRUty9BnBN6ZMbroSGCY3sU2/fDQYdb
EEkv8om4+ROtETl28S4GnT3tH1oQ+zEC+oU/RNAhCCtT9W21F0W8N0z4x3Px2btG
nkTI+7807ZBbwzPTk25YkL8eT0Z3O1l4uNnT2VughcSFA5HwIolc+iCoa4kmrH2o
qkRbzqTV4BgGisOEQ6ftQYvUSak7xeehCsygFwXRz6si7hLZQmREB46ax5QyIpm0
/M4aTEapHRQPve/NcTS41xp6N9BdRm6Gq2yaXdNht6fCsKqm3BkNsMP/gXx2XgHV
XTMhEPTlBC8MAzl5KVMsOiKK1BzVkIyXtmktucgGqKukLptsbN/df2fOy03aMDlC
xoOlOlnigyxaK2wri6H0d+kyhBhJD6h9tahhQttCk0SwrcpLufF3p2uoD5VlayF+
OJ52gI3st8RY6y5133VBhAAyH2zFGrXrxTRs6o06DO75p5BWabKg27ewtjBIlt5q
jOM2+Fe8D0DWjHgBNZ7FfXIAMdZF/bdZ81Noxn13aCrz38pIs+Est0zwrcZawBRH
PgpKwbPpR5CkcjGD0fryFt2fWe7Wloket4+RG5tNThRtFT1rlVVJtuzPG1R9IYun
RaAKthld+9nxK1ySiTeH73fyiwP9tPvmodLjfrG2kZiWNVfUulXSYv/H2uHKc0uS
BSbjgUEixB7ow8ohmguoWM99CTSFpYuQoXPZwA6+D6jpohXV+Vsyq6OAsRtDf8s1
krH3O6JbWM1cftYCJzRlNcXBNNd9tGLAwhvewxVXWO1LuQjy+1I+/5Enen6Eu3Yw
4Va1HQN9hWyzu0BUIy7XvPjI8Z8o4B0atthtwmNw+XZMK/Y/Obd9sYH8+X7b4awh
8u+2bv7HbFRDSYRjfNRz+eHGvc2QZjqZTK40hSut50/SMxe979TJRf3Z+2ybe0DA
IBuBGIWl8FXtX9lyA2a8DiwnEmEYGNpW5cysFUGwGpHWxeITxc4l+kNIK6ewtvcE
qPuep24W8mk0TetkFgyxlETSroAqiBSxqehQlG0rCjmssGT2Dw5UEpDFj8mMyERa
kNoqnbg2jnFTl/UpO+unAifFtepl8Knp2dP01yU+laygoaiWM6ZD11jeKL/Fis8B
VOOscZGcai0Y7ggWGNazVEY1aQy1HAfeEqAn8eosTAR71NmzJod7odUlPqIXLbzu
3202EGWSruw0n7TKp3KWf5N1frd+dQ7CA8j3KpEui+85C8AgZrJdEtWmDGxNb1Hv
/OsW352fUdcDcDWAcGKQIKy24LbadzcbHiky3mUNAVDMyYmYXFN7Yhg8LCdKLW5C
8tz63AfERTfLCf0djDV/k4pHp1FGEbLNLRWvtS780cQEOrU4C3y2uTvTf83gkDTE
jGZMBJ8r02l56DtPxYXZJRsXEteUUcgJCE3eBNguI1CSUqPiZZCZfBI+QqkIDTLp
qIGcSXjLpiKwzOXFRDvDiurqsIsxyqMwO5Pc/ZUSR+tN4K5dYKWymxshQLAJfKMC
wZf9kDFMmf+sgEH4xa86uuzf+9xQOatHy/KBe+oRWJM3gKU1OVcyNjf87TuHA1Cz
oz05/WvJgw1Bl5uiLUgvfX43va4Oz+FqrlHhlRAb/aCpP2Sk815KAUTnO+Pnh/vw
9L1IQ3TVG96UbLrmgxvd1KKnq+oQT7f8ULtfCckXv3CC09usBzJqQZmCNQX9m7Dx
Dqe0Y8ed8MG+Tidu1vSbm3+Cz83dNQvlvDT2F/xLY89kswGrFhaEyEX0lYYAHGb+
4ASQqvSnfLUkuPITUyoRWst3hE5jFOWikdnQwPaQVpNE4hjMYPFNbXSfsH8oUGRG
JfJkMMHzX6Kw4cjI0ZYpf9xBX7XxbYvVnlGt7PbjHhm0bHNwXc5YGws4nhzlDkGt
X4OaIZ+r2+TgaLf+y+5Ml4BiknIMqB9TwSZebxDu15bqBBTSuZbxd0bQlpSYxIoj
E4UbNOPq75l7TLEUdi4lNr2wMAJzTqTR5QMT/rf5Kn2sKshn+IsKLdmy+1IPIw9q
Jx1Yi3O+Zg4MnhWekn4ZvMHxFvQ3nue7tVQMr37PSDuOKDe3ZyxZj7Kgnl5bdgpP
F6KooLsX8z6xpBqKW2APW8WIE6UEZvasWKAzfup65AuiO/5H96qMsR9u9tQFW94o
fhsaaKw7m4KfLQqHCj20i9/ZSqpRuaLaI1hsOma+tnBiF5tPZFO1URhHUQQ4ySeC
/jK63DaGA5Mz0Oyx9GWiS/MB+4iAf0cJMzvbCJEQFMQWT4XY/avnsqPAXGrnOYi7
V//Uj2KRIVFmENNDKULpNJmQnG8RYKEzfCPelVuhl5R748A6lBTKBNrj6RxL8+YL
UJC+aG3Yd5b2a2vZSTXgO2/skI47KKfBBKsSFkCUHS0QIEV9f4e72xoG8raUjJMY
AHFjd9arLUK+p6OdfuOfsGY2b0e5uRfjNYQD9xZL8pCAvYmauSAiKXlHl1/RbwLz
Bb1y1IusP+ZKZYlifZteQGad+fk6ion01/t8PrypxPCDdM1cIgBuLtUhjoF+0FCq
RD2C/HqQnh/Mff6txMAOAOOtKFNw0AzSgwKOKvowoDkRYb1bE7zaZpjdWNjcvpCA
hfuNhIc6W2p4vkKer625h2x47orEFO+xy6NsNfDM1hjpwJa/7ujpuHewptM0xNPu
umcETzE+aa4tPwtKiahoLvJP7hDiF3kmnxGsC8mgFYWKffOO7zfNe3l5u86TlNZy
rVPsM8nWjvETTYQpIO7Gmv3oXudzR0mixkG9NemV5na3XZGGyXIImS95PawCkdsz
IMjTDo+7dxtOWITjyL/f12e8wvlIg/1ChYwQWR2N+fQHCP4x6Jyk+PUxRCoMoWMm
51PvBKoJzR7cr2P6KJcoE6itGhLtqxwmzYVB4yLtqtGIiZU1O1N0qq+JbQrhf464
zzo4mCOg3bBjoZ9WdziExPCgLpds8/Cw8oLW1T0zOZ1bIPnZbFBCxFrMQQFdBYmr
rY04GEybedVurqD0F4264dI2vLkQfbHAwXzAt6j4SMP37GvTxotuxlgXD+IbXZJ9
0nY6LWwsUC/IDtR6PWf30lyOoYltmYUPX+ZtcYzY7qmmJHzIE+hwytRV+t7YXLJr
H1iSQkC8QqCcqdmhfi+79qtoehqwva1FvGqdUXOmYaIypA9t2VE5IZrpWL1db8NX
ObW8ElLEciFqfaeEOb6SY5OGfGnIBnyUYYy4/zXl8WInrqk109TTL/F9VVIgwohv
OsTf6Da8Ki9seBlsoYD1hEi4RkbBB7s7YIFfZjfK8MfJFf/0mz9jYexVnYNtZsmw
lIPEfljcixmNN9xMzOdGmvO+RkLsfoYxuaaKkhEUh6D5Rww81sMtn3v4caWHjm9v
XsYht07JiyQ32p9B3LherMSxxmUNz+ve5WsWn2OHnpwNg1B6+b18KiRyuFh1CGou
fgOBzE3vmIi+ZnI68YeDPgNYOUmUpjY4vsfMwqhqDufSabLNJE0kaB3+m33HoVOE
79JMOjzGL76OBnvajFdiz26dFgBllyGwHaowE7708j6DHWZbA+ftAkMbGqseWiu1
lU2dHvm9F2nHU+za4NdD9IEiQC8XXemr8ITZf7H6toAwq8JwGFD7/c+ZGPiVoCKI
OSlY8NKP7YyblAjHQNRvTw7vR6JtEk8qegHvo0MovRB7NtYBm+3hsJmH/27OJo9z
gZjQ06XjNrZu2bvZVym4gW0asOgCK0x8H9Q/DwbbGN5QLeCSrvYdyWkiZHNeLYMZ
+oyo11wP29ZvqUZ1DFuVfxZX1pmnGz8bhq4d9rkNc1xAHZODaWmSarDBdBbsP6z0
lsQjJVBy+2LR+015+apPV5tcythLuNgEylmBqfkP1c3tLrSn5ZpB0rDXB4NV66Ip
XHihUYLPbSAGarg30BDZ5WHGdW1lPKJ/QnG9yhS4rZAkHx9dxwaKppeVeWKEnuUF
QC8XGGoX2wuW4Rkc3Bjq9pmKg3cIn5AVeY2Ch/MV2pKJezE3gCx7reqMpVeb341F
j8zIa0Zb5IdcoIT9y23oORtgtv50IZiQQ6qzmabm9tQ/ISzH7peX/p5Cp9bK/qLj
lyhtujjcNSRBgTozBG1oM9ANevWLXte9U3DdRxxa2tvG5pFj3FP7GYfJqUneE7ju
tos+FbLKFt5QFcUEuYzV94K6BvIdwX4HzuNUI0bT6Lat3pBwZsiJfKuJoJHqPRF9
MIYhrcSvUNHtVR83rwEPjz4CIJngehJn/O7dDO04JuV3nnHk2w40lQEPyIvM8RT7
E05vFRvXz9K7gkiELXiPkd5Oi0pccpT7X98RgQkg9LSH5GF8N9QNpuuMrVrdfJuc
P0QGBFQqplXUBofCvbmRfX9L3VYrCU7/KPsz72Z1vj1hVTnCZZpdYTOh4uTBzTom
wiV+idkt799/3draUL/jnObEhUCb+fzMo8xEg9G8rxzWWWSv2cPwLiAZATkP2aZ0
Y4LX4fGpUmB+gdtvITGjTp4b4AvD71NO/lAsT8eS1hjQqHQgn5rtHjaGLqjuAaDB
1O34J0Ew+IHdhlWmwDEGmglYiL6JTJiMZv3I+kubMg44sRCZVLa4EdCHlkqH448v
7pS95v0wo9x4SqqA4rEBY7GgvtAiaoeaxI6wKJL+683xfayufi3MZ3AXHJPKt9L4
ip02dbByUaG655wMnoXO6fh+n19cNdcNDwHSGLMOA4TY/hsxFej+0CT6ej6+ehzd
xrfb860UX2N35lgM+/QLz4B5Aa3Pl14E0NalZiaIDSEwOEnAY0TbMC02NBbZleDN
YGA60lKuT425figUCNiMOUlRz/CecYJiG4aHtsVT/i35q1coj0ZGoKoEPBEA5/6T
iXb+9JME1gqffCTKA5RgiertAAeCSCekLCvzzVW79Tzzp/lU1DC0GHMaLVceM09K
ZZyjlcA9AKOOO9SokkdeMScf1mr3jPaQKvsvFnBuIEft6kiWpTHhWPDr15vAMipi
d+T9/s9iNX5gq1adDxTkOxXOpc0MXLUdTEBX4ghPe6ysjMNWV1AaYoxG2dA033Wl
44UyOSjvO+cymzXeS6RCPsW07f6f2D8tMe9A/X4Q/l6yZmlww0aYotdCTF+uZ0HP
szBFEO4r0MS5+pUYPwINcnKBEbZMYd4AS+MNRXMu6E6r8EvAlvpPlhIZxypeU0Ia
052jmRuoLK25zimbQEKzfW9kkczi0abj8cbtCb//0KlelY/tLTHeHfmUv/QJ0d88
eaX2YwUTlp+io2FLgHuRWRZlwlt1UTZeV4H5FoacXKfPce101FDCwo9MJDCefM6Q
lI0f+BpGtKmdAACPfwc+E9EY7sOjB2fpVEqn4IxT6XKvXEmfrKbqWbQXw6GaXECC
xs7MhTEdvPEaJIgfq/mufkougvtYkXKaPbWU/BTkj36ZwvQXeziqORQhnaSyF3tE
18qsxja6FlkUX6erUhL8rQv9iWLhhYd6Cit8b1nt0kjdfo0GrAVIAxQPHZy6R2Qu
tsdNg97m0nK8iZNbW5Ip27d06nsqTuscHDALkXcXLhMuT+UycUr+GcP4Puh6q7to
WPsSI0wpMd/xfmN0aYUKOXE/WiHEA25TLejcZxEBFcWJ7U12NKhEk/Fm9wGeKBCK
fJwv8gguS/M2OJlKBdcjYRwVDhDllPby40ZJ80VIw9tAkXYR9d8oW5RS0Jwq8M4j
8nGpi7m6au7+J+0Qn914gYJrR3pINJnfrJMKYYy9RhPP7a9cTTtdRw2n/eVAX8HD
4txZYYQAFbd6XpBL/NPztey7LOVxeGcR4V6PTX4xwZpKucy9HdAU2hxh0AVBdono
h+h8+LDX6XoWjDMYzE0RfPsb1NwvYyVAlFIkPyv09j7CU2MSV30BuWwK1FHxol3b
jM4YXHW7+64csrBM0pPozAWaJJhBZsH/HENOmSe1AVErMvQoAdaStHekToAiWZFD
qDFQFUb3YPOv/s+sEKOLfMzWjzznBkhiqQWIKjqyp+q73GihixT2XeoSICggYWZW
TuCuRKfJoVwE7AO81wZBekXU5BYAHxUkB8NDTAUjzvJHhBiNEjBADl+01lJtkN9r
1olx9GoU6ycnArUuPbS/Wl8GxUCL6DKSg0NxUXVQcY6fcSWm7t3JyA74e/yupLP9
qzrH3OTd11Q0SBhlCWr1LTqImFje9mKoDpc5xaNBzB7bxLaWhlsxB9IE2N1WGytD
hAHhQA+gr5HYTiRo1ytxNEysmVcl7ppyY+t1WubcE0nkmC87/TSR4UkGhmsUosdy
s1JTB2M7wGC4F5X8HJWW6GDjfmtaFO8ZIK8zY5cqQrA7Q6z3Je1DAP4WjXsZbL54
xcoXNrYkOmtFOz9GpwhIjhhkCnT67JnTestpNpVU9U8b8P7WNbWZGMzmGjiYfJbE
FnXy9b1XcPl1z7tnQH8h7vmmVXCZsXxmIgIMUW7dGnHdGx0abZ5ElADdxRmM909/
389JLKE0jbLqkunfwDVsEPHXgIkWMVYs7QbBOuRNnzUOUzgxaGNVZiRJQJnhqA/N
RD4NX1i60JaB93XAWVA1xPi8C6dwt7h8nIAF4M/au4wiua/TnBAWTaVDXU0FpIoQ
mwXKMbxjiEiHe4OEHIdknzYNRBt+GA7/zzOeuI7h/PrsXjmwqDSjAOO6QB7wIJCz
CgFx5W4CFSsw01oHbhzSbDDaC3fkXxvOnrUIRIKF6vVZ5MhOpRRcRAZaNZEgupvn
gpHP6FFE3GDI3gF3sZZjkVYlq5x+QaSmHdWFb9AG4vD/Nj611NvNyZzqizUs45bX
Ujq55e0aHJQ3FEGPveVGXOnviBmPfj1yJuWmP9DeLUXCQvKReOfD1nc8S8UPM+xa
g2RaCPjKhvSEPQU4Av2VVxkhjoNNgiLVghaAGHluz70/5F7U94WD371LlHXuC9oN
Q26DfQ+AB1wuC9YZA8bOsPrerDtBz7lHQQq3DkFGyKGvW8q4fJR9xxXTfjPuxtuP
kK/3WV6/7TqroIRUA3GnBW3Rxlt7MwOaDpV0FO2tNdun7PEFkesaL7pOWHtKcRJD
5ngG1VVzDDqKSFFZbS5jCvBHryigowG4bIHoM2eljjVMjT5tph9l4fmuCIGG8Ipb
IHF1jBZ3bA5SqXKY8gWVMot6sxQ6AFXtVy6zf8DFqyiwtawPus/1DiAAZUQtHkRx
M1x80eajIg2fpoNBabGxdPg13EUGm5G/F0niFytFAVyxh8aLLYDyef2CneUuGOWn
Subum/CCAbPr+PHPfsebGLv3K2pzbCOTCqyfwFjPSHsTm64YjlVMFHf7+dPj+GH3
zSNOuQ5lzmKw8V+Q2RjiT841kMj1wyFvMfrWbtIWgKhf5DdTkYjrMU7imRkD4iNU
ThcczmdOoVclgv3RN44+FHTSlyTjOsVZb0PnD1dJ+TS/UUXfW2wE/hgWGWG4UQ0/
U9Y8hUgcMoBJ1OM1HpaL1EP4XSpioAVf/Qe2HUgOZKnSfTCtrHCZR5MvuFSM/hd9
Khq+qWes5ASSWVHa2ssiS0TbDwUOWAVowIO7kJBiYic3WsiZqK74yS6P5XFKtJBx
2eC9fnPem6yVxOfZ/kcfBYvx1LgjpEQfvSbDNKDhKTzCNMfoOKOEzGlptAfAmcWK
EccmHyGr4rn6eR67O9t0zYZE1zpAn3WcEYb//jzPiUA2J27j6koSJ3pPRjwvp4uT
hVydR+YChIwNy7rccpNMJgqLDUpduBoaz1oVHRqs/HQoU2ey9YV2xyqR/hbCwQ0d
1lEKhEe+y0KBJSaf+MnwQLGqkDr7BBKlolYvTD0qvZQJxfIP48vMaXgmu6suxuun
rN7P/Fe6VPYQWQQpbHFh23t4jPcWflr5OHc698BI/lJ0FY2gZMvOK+H9J8BF9Z6m
2AtQmtJMO56n9fe8tdIQS2EUCwyyNUglnOQ+Wdkd1AL+B44wH7T9wECVcBItRecy
33TnPVO5A3K8utAEAnBGZCtoKr1LqZ2eWMBKbfI+pggzmMoeaGS3NKABZtpFA9dP
MlVGA76WZ9xCs2bl/m5FmObXTonx6zx0F1nddtK7fRE5v/ppJtHahvKTxNAW2u6B
vgCLKuEOnJpPpJvhMz4n6mpSizpZ2dcTYJZWElmN3YuMW7TZtDfIfY7br6z6miGi
WwMFk1N9G6OEUO7Mf5ODGutC1CYxaG4NFjTNishV22N/IaYmIaGoEwYZ8DuwsYL4
SGsI4nPQ11W+fN5zSCUlTs3RiFVblCyO3cqeWPSG/gtq8+0aIeHNMxcW+JdtVv6O
VYbq1qDtPFVN2iK56bUwIMI81kYO/H9U5Ctc3wm3MgKPKFupex5Iqi35roe4PnnA
+3U9nEZfEpo7SOQJQ8JHDmoQRNBgkNWOYf3I6FqIC5w/I46LM4vonJBmkuG1H5CR
ameiQq2L2yDUU+68YLHC7PdinY11pnrw+3Z441T6WlPkUyGaC+x5cySj2j1v3MdW
doC9j1/WPNT5Vod5oZ/Q6+wVMbhOSLGHJMSw0Zsm6ugomvTb738D2fOkLCo+yPz4
nnRBPVrs1IJBYxUT3zoGPo2Q9aabHJTMzqkcPPRoZpKuEf+2p2JGyM3jW+qjLm3K
01afBGV6WuDfgjTBK+ujXkaKY0YPtuddBwkZWBe9gMfqRlnMsCNYZ/yahQoVX3xj
zpry8NKpIrmeEy2c8fWqhJHirZOqns57Vlr14SKb5f9sYqmz0J5jXT/Zq6Ghpa6u
uLLcF12fIwL/hLOLheLuEBcCJLXie8tU4ruMl1zdfcMsqxwnsXneJ/CqWrg0x4fx
vTKJWiSsxV4P+ki8wYzbMRUJx/hwCtXK2KTeiu9PES+mGXGVovnhMNHXpyzbqnuZ
zMWAqh029WdIf6BANoVu0YMOqRdsxnXUAU/4nqhFEmlqBhP0kmxoSt4BQbC2j6qW
inU/ddQAsa8VSRyrUrKGJuxGTlkxFCTh9o5u+XCGi8drZQbG+C2pmcFiuLE8jT9j
X3XR4OZI/TAyjA8FxOuA4H+3hdFHqYFcD7CWoFrOi8BKioYRwNU2JxCTtuYSNyoX
1JvlOelwuEBs9HSJtr2gEAN7053RsdN7nl4EGiyDTkUZ2B3pGptdggJEfhYBTVzX
dgg7C1AKrU9KKn2gtgBQB9HZmkfvpfUvbwpZFmMpwki0QFBIYlIc07R0rlLg1c85
IFh5MW1QH9qtZMpyUjJBpwzIibObT+hx9u/+tPdsAfUNgViYwrPFX+asKYupAJpp
5+opvmrwQIWEJUDcICAYfRZx3aileGqzoH0iKWoBPKmGdYwwOC7+Vq7EaDBxrLGb
I2pec7931uvDHe8lCmeWmqC4V/b+jSKwvwhbqu+JbTSG3dGQtc8G8gYquNJo98Wv
uysQaD7CpjhlSclDbqhnHyrEYZVzAGmlvONm/H99JR7S81SZtzCXEGIbsL6/YlGn
RIcs38bjxX48taPpLMw82ZVhdth8F2ef2/G4Hz/HL7TghzKmq9YwILTiXyyHOYZj
I2SC0ngE5LvTQNcs1FXyOlt9xiRp9j/P+t8uJwbSCUHIvl42SWSW2TYnHsgvV7M0
Z7PSZjHgAPwuziDPvsm21ALWZ/VNLW1BQ6eEXC+dKM9sUvmw201wGupnxe1JefpT
/7f8BtsAlu/z4rvRWPK7wF4VXNcjwM5fZNeEY+ujtnAJ6I0VOnV9ZOpVHQpMXMx6
8DjHjb11nPxuymqDC65WWxH0e5Th6e3iS40pbNg0T9EmFsuE3l2J2V4rcssN3yXH
97acUVi1DXeql23Y10lEw7ts4WVgM0xPk7CRppxBEwDgGkgCrmyhrm+7tUXCtc/F
OTCcj8x2VmVn5G3Bhj7QboKj6NsdIWmBbMAVOpA9NlJiqc69ldZ1VAEnT9R4Vy9X
PZrBtxDacyG4cHJK6YWRsSwaYsaBcJdCc6JZM6R9067WjZdrp204ttYGlhVSEdX8
52u5jcDHLEpBb9QD/zPSNijjSxyS8HF4HAsczOV5fcBFUxOsvCQw/ejj+fHroZbP
MRjkAesDQ2qZdJ2B/MXRfwYPmYpJiQbKLJcQ7HH9QxCRwaRuV53uo144KAuf0mhe
ggMWf6nsupEODbSEkB5AuSzmSiWqEcYemhlUJaaeELUu0liA21YqTYJVnl7oWToq
zDfUSNR11PNS8v77GwWrphkeBQnE7xs6l9s1fsOM3JkMU9nuacwzRuVlaC+beQUV
1WS1DNg8XFmmSHXGGIHidRWDIKVwmnmx7KxTfPyfnzyW/ydFsSfNUphppThTXmXs
iTjM7e5CQkd/DBNEmIXk3xzq2xVYMhSue3WGyJFhnigOK116NEh8gjo7TZsBT+nU
XTtCDHLxGy5IlfDK/PuuWiLeDN6IcDKWY8zBlKay+jX2SIZeoRaVsc02cpRyxUiT
kpJQ/R5XN8gG75g7Nfdoi4Up0MUQwtct0D+RGNcfdc0fbT7+7cfBmeqCgbdEFkbW
biv9SWu2xbKufSYCGuZpVKc9j2sHJ7lb8Yzsde3PQJRCN+YPw8Kk1c/z3NbWHKwY
o7CLelJ1HQeyl4Sw+iZ6Z2wyY0ZhNoqmt6PzBJdy55WLe6H7BKUmAgP0lWz3IJCj
CeGttiJM0XqZo76xbl3qXUlxbUeivUeoG+yNEaBCenaCGDpSco8CZm4io4yAiwSX
/Lo2E+HQ1hDDLYTEurYnonCIZOmeKH3I7tdyujpdMqRmVzfMOtDSxQlpgh2uIRMv
ZO5T3irT45avnHf/VntnsUQScflMAPJUu//gsWDmUU+TkVLDvFL4khak2njNkaST
OWpkegllStEblwrG1TUE+31wCWfHrBgspudLKsFnAsfyza2YVfKPIQaLoMsHJPnv
+Iee52cGtvV/UL9fKFcjIWH8F9OR14m43qEdOxBYTUkLzhAmQCRbGqYjtOBGDJP0
2rIHBZOuEfBytkMO8QMk/Si45WySnOemt+O4ZbtzoAb8mtyum6Ky7crfx5zWOJRb
wGtkSevyGDP2DfazhcKlMnxjM5Rx7ZDa/aoKPxfW7Ex1EzlzvSQKqvBObxuJGufW
FJePcNt4ap5hDrVvDTpc81o+28OVaPOj4IZQwt38FOf8IDTPaze80sjKoxdSCXb1
uKilhK25EFma1ISEv5x3y1S9cse/MGbzngCHOELaLJWXnR7xp1xvybo5c09xalAO
KMVw8atWwjjg/78txnyBf1eRh4sTksvcXnEDgTzmbnnggIDuTBB6aS+7pRLAavm6
jRb8RKKr4D/vleKZyaCVY8ZzSdk4rWZhGLPs4ZlztqCVDfkrG4YTTwXR9oYhnVC7
A+SG3tqtPiOhi3A1cFowq4HGJlOLL/m/MTLFan9Bas4hrLqF6EgWO9ahOyu6ksoa
lw+pO1St0JE8X06KLxnJoL0nquG5Zfecu+gxhNGbsR7bfsEpSOrhkfOJDAvHI/GX
Og4MwZXMnUnb5lKOX5eJyivHfnhcC5GaioT7ITyT0l8ag5AfyP+qsLVAUXRFwpz1
IpfIX6xg7UwDBZGYaSsK7StHtf6JMha2BP/vu+wDKwhNwAMGLNEhc1U6+Retyvul
Nfc8AbzPnv9ZMFyG+cxJFT4xNYS3qTXPocDGexS8aa8YFC9sVLcHVDAFUR5iZAj2
MxDOQgwMqwHcHP6yImwH1EgrLoZqci9h2iGwNZdWJnYUleXPwTmHscL1AHIYQHc9
wBXl0w1N2WSJwKIwLYs6jnqsZZzyXO6AWEsE9IyxHA6zGWJc8WsBMsgbLi/eO1L4
oe9hGvNvniGTivoIHNgt4xDrK5bdTlflTuc0N1WSeDWE2OwLbYXtaOGzbzmshmRs
SnBecEMl6QAo2S7/998qxZfSsO3jiXJlDSD6hvU/si8yhFQMO/FihLORlq7R59VE
KWfA3P+q3M2WkE444XTUd+cIrke8GkDngFJa9NcmEqDcvLDghpRg8A0UQl9VjWek
ij0y1uXTou3Dn/KRcgoH+5ItiL+L/YGkCb9CeVgyMtQ/1Sw6k+iTuVZVX9rBoSo2
DKICjMugSvpwDVa17j6FMT433Ap7sQmNEI1CswINxUQJaSmepqIOhrDAcaKxteGV
H50qOZHr6uL4gciO+NsWvS13+WLJh+Xjwf7tnVaAS9p4L/aQKzJCiLit1vpkeu/X
VNh5k8Z12TNLLiZ960nasZ/KUEwfeTo0kqUt0l1qDbRzy+we/h1BN5qmPQJ1vJPP
CT41y/Fi8ZqShdug3CeeyVR3OxM2gdotqCwDNP12x9QnucG0wHlTkBo8oDK+Uy/q
YkHwDptEz/+RQ+dJC5dEqhI8oD31dMt52Z16GcpFqnuOfiITPcii98D3UKJXl4w7
u/RxsMNQ7YBakg7+t0FwUkE6PT6/KU1jrEc/qVb3DZtvlb+kSbAbAY336Zc4rB5k
dV1kRq9nXQPtB/MZvHmRhu0oAVCwQxD9RIeHG+2NVzFFAyY78HGzeG9orG7Y3nPb
6PtPvmo2toUJXMEg+UssfU0QJkQysySmwV8elR9Id4QMh5RhV2mdvZ7maLYjRC+x
wBsfX839NJjx+6ij3JcPttFDkrFnSJYTSHA1rcNJysefiyFHzjzjF4lOh7v0r9UI
y9NpJ91B8f9EwLLch6hRYHwGbLFgIGh0bR/bCkXWpw4DhrXG3pEtuabCqpq1vI7p
xsm07aAU/l/+8emV1Oj+CX15q1giHNlycI9BXb1hnXJltz/CIqwmd6G9K4aciqnV
hQs/b2wJ9c+86UnMs/OsA0afEJv/56vhOeLBnAJqo58DZjjvDmtT9KFjZZArtn15
RnQcp4xi01NRykJGUU2LfQ5LNsemzKQHiFudH5YlmgIgMSgpEEx+PSxmVC8xB+Le
U+AoYIM1kTDiErrtHBgb5gbzfex1nXRw/z8g508zhhN5GAglgblf7T6jzrpx5HSX
5KwPyQBb2TervRD3KkZbx41Edncv03sHDVlT6/9pRrct9MGTkl5etEglOui5w50S
wFGmyIQhQxm8s5jHAuCSVZN0tQ9DcK0aIlVqdkALsUsJj58OaSuCwezjPFcMooh8
yRWNBkpoWlEJRwoYwuwWZGZ9iYQptTz0DepLSIlucFJChb5bc971jN7anFlWiWiQ
M3d+XOe/qLTLYGpY/3654zxaWdN40eOQONvSIJCns8obOem5kxn7PoTClZxmA8aI
HEHSrSsdvwhHEJrZrwrKTD1vICoSnpHgA/2n8m0QmV9COPD1qtjIu3CcSDCsEUhB
CjCq7wU3+bbkpdinCraGeZeQ7HRN9OjXohN7FtVVN9j2LxGC4OsWHyyAPQAUJARh
C62JNIBQ7npS0yQl10oW5E4BDX0NnqnLBPFQpOBoH3Bqgi1PJBZ4gf5QYbE19rkK
HP1wqqIVRlU5adXJOZ5Wre8BVE1cYMyFI36h0pSqcwtgnVGKkWAQUUEWcGHuF+cX
a4JesoGuFSJQjXZ9CYU3DPhc8WPau6+Ooe+NBTXoXDjaZAcfaBkjGZuWIxOC+FkE
klnJvTYBGNrWUscNnWQ6kURG+vFMXY2BAqTVUUdG25SwJBKBgXfiHfYUJ9lorKIl
sNfo5O3l4S5A184wvSl5yVlLRrgS2Q1KMcztoaFj41m9qbWPP4dOClSFo7KG4+9B
1x9cXPqKyXqAIGS7GqW4FeQ0/RpZWAwOmGljnk7YQtIuSURNIAkcCs3hkukLImhV
mYG45UHNOaiCFWJpwi5z45sEuugeh870ubV7T3Wdi9quPQv1ZtrDG4wAH0CSzlZv
jznwCYcuC5ZWmSKmneiK4wwiPlGCtG/QrM7EXlKymLcpVr0g+QNEKk15Z0xM7/j8
PCpLcJSYj5XCqzSx2feQs7hC8h32KZ0KJzDqFkQxU4CrXrjwnH4iY6o7tu58LVKR
aQUYTIQerjtoi8dKtZBnodnuXLt+waRAMmrWcAVJtARMOaEs5/M6hUgmz1iVnSJ+
cDQ18BFv8+FW0Iy+KcSlKi1I0YIP+gre3SnVmg/58yYKH0nUKhDJkoNsAtF606l1
rlP06aRyXAwlBv0EnNTr7LPARA2obqmLjQ798zLfg/+jvnw2u63kbuL2/DOCv+PB
3WaLTtwurE1YAQyEE+ePmdpIoZVizorEvUvvCwK0FzbYOSavmWjFG+x3A0L3Osls
EUdt7bi6/D0oFp/HemUnGqiQd58qLVFmmo0/4HjJvzoPV2laoO4doy+m9fClyq+Q
4j6o89btS8XRNWcMGjyqo1sOCCyEZz4fjOqR9Yx91c08HbCeyhG/QNLisTd02Uo6
q1zBDrAC9d8vCXx/v6kmBTCexfjonP9zWQ0O2VD+lEA3n9HW4TCXleprV34RnOCI
EKpDyvobjQ00Iuyc1glahFuO+M5qKbLtzERlXjuzzECKva3V3tIAtrt/W5BBk+uc
Zavapu9n48jvHO+TgB1GOXTsBAQ1ePkkaLlXKz9if0SkAIOwkfvoMUbSoyeUUSap
qOJcUUhIPpmMkkiF8VNmfm373Dx4qjq/9EfT2Df9peMQqOHbXBdF9FtDhYGO/Sa7
8clxgNYzShH37oYRttMc/Fek3R2mSLWavEbeLydyG52Lwp6WWA0vIppXIj2tmIz8
60t/L61BmC4UG2U6CRBm2YV4IgkAopF6nF+32qYnSULwl7Pg9vXNELOd8xmi/+6r
aebl+JdBbduXthW0FkyiutPM8/gZBZrCrv0T7Zop3BEtTcJEV7XiIqAolqWoveKw
fFn19SvpsadMQ4q3IuaMmyonl6jYd8oPqH+h9BYyWtOHIEgWE7x4BlKaF8PZmy1I
jAt1fncaWAD+679QWjePPDZH8zhqxn6x4mAm8SbCskkYpVxhF5vc7gpPCBZjishk
WMJKp0bwtWBsFSWs/b6I8+Y/pMyYocosB+2dBl+mUiNE1nFTaPZqsMtKxZdTB8Il
iRFs6ZM8R86e8oh9uLH2W/8hhws+MJlGhmOsWRYzu3tPH27eEIfAHhIa2+S5Mx0H
WK5dsK8pY7iHMBwPPSdcKzLD8FZOrc0vgZ3Lkw+fOnkXcn5ZxBdx9W0nr0G6WHNA
2+gMfgWP9W7Yv6Lr3pGIK443eWZO6XYoWMuv8fP3lqhNmGKhvCfWr6hrevu4V6qX
kTkngierqvDsa2fb+irW9A7QmoR8NMcVukorVm7f33b5l+N+IWIxO6WqWn4Gf+yq
cP52sL0/d6VIEgkkEXFt206DZW2Y+mu29hsHvRiLaJ/BFDr2NP1ZA8sLFaHid6ce
2qz1YLVXfRmWVYBMMSub27e/JSkCPu8yFptZTmD3tjFTFyI+juBcrZXrVbyEIYDV
Amomuatky/utVLqO5eSPbUi4FAhYolKCSsoutwlfPzmDgTQSU6w4iStcEgOssFpN
cg4HMauNBKv59Nz1VXCX+B4w6ezohKu0odiB6DAhqvbWCN23J8bg+zDAhzZ2v5Xi
dCoNECSFbrnzidn92yBUzUatLm0dDUZS74eDtIjT/BpcvM8Zju0jNwOakJxi0yWJ
9vqGYKH/NJUW4vpBPHomnCh9LzjUvMhMKAJ7DrGk3FkfIoRlx6ftI1Fc/RcD1j2O
UBm2uqzI3mhHQMu8DqaTrZTcKnYYucLrzaKgQqFbL4SgqnsAuKU2sM4FjDB7VS7Z
LWEyBotfwywBJRpD/vR6/GoDWAbG07S988HbvyTC9e+KXE7nH2rmuLQ8usOOzFMh
935AX1LBlW4LHrqxDxY0U1XDNYRfS3uh1+1WD4wpbI3ZCr1A0lhsTJFYHFygh0XQ
DgoAoUt0Bh0MJB4+1AnUbhyZRx0XzV4EwB5eCFxWnzsdFUjOqktVV5t5jtJMBQ/7
gNohVrLnALbVsiaJRjWpG32DTkWsyojBBrLX1cYjTG6ubQ66tbk4Lk3kMQBUjI1u
fJICpxzeszVlK/zmCnduuKMDquTyvObOlvViR0fAj6Pwh3r/hjj0NrqmVdsDFZsE
Io5ZpbEMCulaoBC7ot5783PbRCk/uhOPiMnHAcSs3622tcUYkACinTEspIvYKX+2
rNCzMylevGtfduZ7U68Lj7zcgIR03Himta6tMj/0ufp1t9rsJecSzM6uVaiG1tjI
+oVttkosHeOjV+OakgEvjLWHAxazeHijJDK/3DutlqR1zgsqvzxJSzpUVVUZs2ZX
TPqXaKJ77tvxQUraWPgFh1+rZ1ET+QVeKzTgNXLXobzIGq2DT6J61gU6E4PIpn7k
xMk/GMwXcnh3LL+JulKy46WwEaxz+NQ+6rWNKvr0zgigxZOtsqtG4BPouoEAHL4n
9lI377xjEF/fVsCTmBU6A0EX59CKgY+EjxGMmVMDJjwfGwR9xaanhRwBtmOvZlU2
tUqQVT9HtOVRTwc1NSM7sW31caYT/ftT1mXsz89+QQ82nSbJzAltWulo4N7I3o0r
9DgGeMHAWcq+DXyR1RNLIn71Nt99FpsJjTe4ZPd2oCwjQVz7rftuCJIX/XDW2mTi
VqMPnkJJhgHu/ozku0eLC2HzkQKMwtpJAtKrSIRU9Pr6o4445BEzlj8PwQaJHJJC
SmiKEts4THoDDdplp3n2TsmelCPl7PNNY4bLix++l6bny0ZswmhHrhI3MoMkMEaI
QVtqnIhoaTieTIJA/1TD04awYQ+2M4eXyq3IMey5zPAv/0BLRllhnhJRF0lI6eUV
FsHsB1dBMgqD5K/GND2jiNUTKn8N3gU+GK3uS8iNVxerQ4XtITcytWPhcQ7lIOlu
U/SVwL9CboBVm5fl7Ktd5vk3k1PdtW+a1XlyGl//5JCijm+mRahNb+vPffkMrY5B
r2xmIYM/6uj/k6rmd3N6xmuPghnjgj19rMT5CSoaz1IfYP+Pd+oPS3YiZS/dGNzE
hipN+mcSWxTPYVuxhrN9kSzLDT1APJY/NralvD+z3cnaXlM3riuvMRfj7eEYZ/6e
giAWc3Mrn6bbU0MAyId2Rc9MMhR0NPDyXyeaPyxP51gbreg7hkhngArfdXH+OnDe
mSTuOcbnlLn2BjYvNGw2k54rUE4nekPwlD266TLYIC3Fs9F2p6vq2yvuss0f0972
kUwzQZTMA/+vLjOD6wWA3IPV7wXPTm079+53kejkpnUDMduHaMrB25LgDc7+yftI
wOYC49R1bhmahdl428sMDStWiRNOtL61S827crRF64trwEz6Glu1OR8ERzNoGkm1
5EhMAvb1g/t0fEm2JlrsbW6fa7VYii3Z8v73uJRQL6VfxWCfjJawkBGK/oA4nnpR
x0+5wT+Ji6imnPwfxj3usmrZmhsMATmIFlCCNuXPQwAdW2c0rgMUhSZjvt3oIxBq
iTHl/ucyMojPH28UVTrxOyDi9hDQWi5ZV8HZij+d8BxTNnH8BguCV/teBQvJZccL
JheCJD+7LvAH1hNL1Cx4YQHAP+ZYUP+2ckPOcJ7enqB76lVAeMGDG3pRECIoUJ5q
bL4iqDs2dzI0IDUPv1CmBCz6rYGCMeebb+pmixNnJ+1eUmxUU9ig/wCBqCplqssn
KSvGg6WHacn/yA7SCb/DZ9V1F0iNbROE4FkPG1XvnlPBVJgC8oGD7qi9lFk1Wxwx
bSUFhfJQ3eDXVPxgpHKeu28Y3/pH0JRoci8OYT/5Y0nTfvEzi4JwJVySGSDzK/rF
rlZg7YS/eJBoj5mTU2jIDqR91eYkN9j5Gb9akcqk0eDP7u55BLh1pRaL/xDD0K/B
p5pLgqT8VYWllkHT+zKCNYaqR0B5LrcBSj383p20zm4pXV9cDssY6f5vSsEu1esF
GGpVHun79jeHGtzYhhq9EuCPPSQjYuhyaY5+h+O7q5RO0bTJjpRnpgdZM8oZXFv0
GKefBU41YsVMQ2z2taV34YnLEQ3KIvlp562wQX/xFWj83ZyT9h9dURGOteIfRhcU
XE6W8AiG7gEJGIm+AsfqMK9Hqld2d7XonD/K0qCc5iIRb0x/nqXSQUw/lfvPj4ps
r+IkVfrh7jwLRV+fpIbqIC7eTIPJRMxFkfx0kxWMs5SzeqAJTGhPHzleHx/mqeof
B4tOMZvcBz3em7ZjkSaqJcpqvoJDRUmo+l8xf7kyJoxL0hLLMbJvLbKs8BiL11zz
Dl9Zzvc8tj+btaRoZgbiSDGqbB673SP33ytq8KYzKmnNxFZ6HD2kirCDNiM1sf4b
X4+MGGq8ZhXpedk9uAmAsZs8JRQXlcQQ5Vm7yY0DFqODGt0q9WhOCkJVEaN8EEwA
I+igUsZ16LzcGJJdCy+G+c5bbzX5KQDG4NkYfeIYS3/AheUpcS0zaziluijtAnm9
ivWJNsPMj0ibvz1A1hJr5+XMLA+8JPj9HnlWzd9nfeY0XuuZZkyueeXIX267YKaZ
3U7KOipRUYTAX5jPY2IHydVyOAF9cSnZMKcrMLErDK9pFRhD0eRzv5rhYxvag+Zv
394D8yBE9L9RZ3R2tJ2Q9vfRqs1+0OMPR0f1SXhDc1Na1Z0h/LfpUNznUvOsbiSd
fvPRQwS0IgnUrTdQ5/L1Qipit9QY0h3JnmnAfImolDj2DSuTi5fFolZq7bOJXyvZ
Fjd8ewsMKGr9xyxOkO1sho3TovgxhFnK7yK5BlE6IF15gv7geprs7U1eW6KEw6iR
4aDWkZYR9adp1RNNiWCjsDhVani5bJrsDMcz5sFYrbvujnDmzFExGnEr6yrqkSdM
k3UcxLyNn8XqGia9qg7b4ZKm/K4yJDGiAOOdJ9NSdTrQVHi7Py3sbl2fszXxSCeD
fSEd8lo55pWjNr/5K+F7BEvrNAQAzyKWiG+ElDUinVXUCAVUi0ui+VjC2c8IKAYH
5/WP4jvMzWdY3dLfNeY/5y3nyDt9/pZpkvOKFp4dcLgEBZ4ONHo408iDFWZzCUKe
YfZTyEpuAQMbtUBY1UQ11MJ56iu7B4uTCC4+v4lXVpFjBAdpoQayXdIMHVLl1C1e
xehuWOjrqPfqbwtkyaAH/PVd7zxyt85qR2WNBBZxfcPmqcDjS7mQB1ZZD5IFHBu8
ik8ysVTs/Hk5znX0+DeC6b2rEPGHDDIfl2Fe8ji6LqwpGdftEDgj8/BwGQImSPjl
coD2S09ADS1nn8vGbja4Gv68YA5wSq55IE4DCQUJAdmQqsYdhAnCXuDur//dJaqB
+QQ1iaw2ZZQiHFKqFYnBMt2z4oKwFCbRxRfzZYGjIrAb0RPWB33WleJZGm2hS6V6
WtZEo3Eak7c5s4WF7Jxz9v1PrzquHPQfUcniUye8djlagf71s6hcgSyhnBnrBH+n
kARMO1f3+btcm4bFneduzvIM2CaCXNXtLviZZ3g9NBGkajY+NcnYRMEOXDPnvpSv
7HetrJnUWZsWht66vHIy+ODlSB3WD77tSSOwJLx0c74UkFzWtTTTfi4EdJJ+kpD0
NhSW45nhypnGT8JCunv77kLkdHbZ+OQac54pdn0Se003zKMO9b32zKbRK5leMJSP
6aCBouayvXO3WLMS0X0LPfpW9Zz2/C0kCt721f56h9d6uJFz0vD3y3DuGiUPEsVH
r0TMR6YV7owSBiqcnp0qkryz2b7owbBIr6PBvgq2H4bqOQhsjfGBXeMFgyxEJgpm
nKEAOosaGfj+6G2VEtmbFUya8GyWsfxODYtlVsYiXsfZcxdrxMlaUb2+VcLWuA4y
RSHy4WXFO8CtV+VjyH/EoyUkb8HVuIvN088Mgb3rhJABWleesR7Oy/Ww1IjF+w6A
u53FMaQ/0jGLvrvop6J0wimKBhUnoP0Rpe/3ILqlOns/TLap1SmSodVPbdmu9Ldx
Pz/WPlXutdWrCZ+IgaNt1sOptKCdyztD/opDJl45JhXsBPSc7N0uFTG8E5XCBVI0
XgRDqkHh4Sg3uFvKP40uvNxQKPNhwDIAu/2AzPbpgCQELTwW8nslVK0fAPGVzRIg
dlX2k0HFYdz/dnstMgAZTUGAJba0Y8x13RAu7xv4pQt4g1K+A0vvIfomyEWwymzY
hqV604d14gSXqMSI/QcyeCz4pCi+YibE/1vB3SZ6t3VCXo3+sfV+r4k9xWbIbWfz
yPeJ9JNXxxyzgCRSbNUaGDuNg4HjBlJwtrEFdYjxcjqcIp//qLCUJBuLOpMMtETe
Rb6LnY2+rAdIAd3Amvbjh5aQtYf2WgxHuAM1EQof1z73TauFSwsHsyFCvMiQjTHh
IX/OkYmmWm43Q4AvQaW9xPoTYXwuSWRJ18ZFWqqkY/3opKmd3yk/MM7q7MNrZMjz
RHv1M/DiswQHyzkXWVw9F4xmXl4A48THHVwgh7Oj83ychEXYHYOC+1TgjqmN0kQ5
SeL24ZkE8FoV/wI3JbBI1toebMoFJdVCkgsyKERcwcM5w3kIzaGxDg+EitBMhzl+
L+LZO2urhA+uiRgbsrOjoHzOXv9hlJV0Atjz4pcBz7JQnDsi/ZGZH1LkV+CjMmLJ
hIfGi4pjJ9eUbjR0hmjSlnAq+iRfR8e1bOeo8Tem+q7vlV5PWZ/kdVTgp6ES+E35
LWzRbEwFKR2BI+EOCoE9P/4YdHFbKKfbQU3kodqU4Swj0Ac7b43eMkE4ZN53wIDC
J9sX4TaL6/pnz9cAn2woTBDxIF4mukYWA9qA6Gdo6ofdCxEXqSy+gAAvfqNypHzo
6aq6lHBdwHxSEvjwHJLvKnl0XWArfy4D0BmPpXK6HnfqQ2cihuXlQww4evU1jrEz
dIvzETzPVbLm+/VIDV6LhEHRIQcNkGKiBNdC3OCjxuPl8lhI0MlsBXVOwl+1gnX/
7B9Ks/YbvFP4H28rOaZ3+7edq/WMkeC/dl6tIsZK8bSlZ+yqOq1h7fZOzO40BPfN
fAJU8N8Hvc/NqZDtVoDLIwqK+jc4FKOLmPRoNbRDlwx+R5e0mX4S8EpFyiFNXmOD
418SBLjHrjwDM6Cyj1JMiQ2i3ZkH6Pjbe1tI8kNH0vvMZIDIBoocs9DDmAhhypaG
O2uc076eaDAT2STy9QWjbuByAPtXhh3KSC3ZTDRpNcZZo3YRKjgB81zUFnK9/dyD
lYFdogzJeOD5RKjk8xJxFJXzlugJoesX+KlWMkr/D0N7MSQPNAfekMjyw+0W8ojv
K9ulPLswscMv8t6F6g09dhGa8/YsGOGQQ8KTGgdnfUgoTAp348JiQFbw2rGtxIwH
QLPkzuQRiOD/P5xw5wB2/CJ/XlYoJ2zSdBUi8arUbtleF+TglKh/vRGr+k60RN+C
pYMRpGws06KSlhy+eS4Jjo8zFvjolP3iUQxmS00ulZTqiKYIH51QFCxL7nQFr6a7
FTHLokJ9XTj+L09Gy+5J6zrUMQGb7QKZRBkvLUtihPGNRR7yHs7wCcn8/etFo7ky
Qa05a6JCWVU2Gi8fJ3WMWPBgwOepZDdYHlJvJ2IcbsFoKE9UHGmW8tvXfD7hbJjd
0RfaQ4FTEU5AV1fEDuhyrLks4k3BU0ImN5736d3ZDc7NfbdEyAeHkP54Bs1gNQXb
PEdJdZb9D3kjALyE8lATIfc/eoByByfBNRkV6SoInXBcUniHd/+yW15ZWItrj8cN
EP/MrEV4JsNsGOoIqNqa+OxCw8U5SMt5kMAuripvV+v1eEH+2BucmXeKbQyeqfyP
CBQouzgdT0IM2xrxGUgS7ojxXG8DB7Nzj6bWYV9RjlVswk4GLm13uqmocjNGNWhF
WUaRxcpnwGcNIX1Sp26yB2C/39vcCieYsVGjEWxHp7pSl1g9WLya0xu/jer6la6K
HCrF4ocbHonr9JyDyVK2r6kKTLEvaw8A1fek0tYnSzpdi+TGeHiL271NkyIfWL0D
QZEbkjQZpNyYXcUHt797BRaLvjgFBdBmPzfiPLGapCs0lHlvVqmZK2eC2LY7zbmx
azvOZhhmmki5lPt7xZzQ1f7mfTKDpROUtmh0T8CzK1ikH1ckZJ6sq5WbN9A7p9q9
yeoauytLBo3dBq3/85uO/DQ42ovwVx0FcgvVo24aNGxYzdeOkfmWPvNHUkpgUhG1
X2Vsy1dgWJOorSfP+no6uX7uxgBmnPLfsu9ieyhAzqh+SnRn08ltc3UL7+Qwp5Hb
ptRBGAcRVoD2lEbB6y9r0JUwISdNACk6+pqEOCC5N2NJaPs/AzkoSfvW5ywVS9HT
WePUjB7o7jyjpAnLYoKTaRLP2DIb739EmwmP/Zvcbp5SwZAJh4n14x45CD/Gg64j
rUQ5Cf1Uji3LL+oBr3C2Slr3hpWaxJ47UQ7PmOn8vcZUhV/TL1D0K+PJdrn7eCtn
MIK3Ak8hfnE/xY8ZQnxMIhPfM8UaKI60cDr7D2Fq/2SYz9I7AFIqoeHhvAyrn3XK
o7gynp4pZbk0OLdSLlzvGysiJUanvTnF7E+cg/zD67tozL7393Otzje/bgklBWqW
KsvaNlDBsUVD1x3kSrOz/1tE5EWd1kBmOJz5Obsbv/NyxrDmHtHc0ZNBVJjPcRvS
3+PfBXnrJdU1NXZ74gPaysXO8A9ZQb1OvBy79TiFG4phwGvjGayHVBfXS/g8OQl8
ChoJTxi2Qqnjt53bVL/2rxIgPsCjcS3mr4ON9Oi3/OGKsFuXnW6re1RVFaH58EJ4
N/u6i3vg+737hpFeuyOeZPW7cvMv84UctAaNN3Fb8QhgcjjA2EG3w5gtq+p1muUx
hRzExYfBNYqZeTleJLdzsfxmsQr5jdpaMAGyHMz5sTWm2vbaWAWgI9E1cHprJf7y
O91e+nCbqVPlAIWt9OQHCZoVcKVrnChtc5QMJBX8JSE+ElGlBIi4uK00lM7hzYX+
kJGW7cD3kLfl5LNp+bQCCpYN25E3xQKwvwPKOqD7V6ekIEsNEkYKYV7p77CAMxcL
cV9NeWdMzyi4oHzW9NRSaFuAyTuvyZVdJ3OZOmQCvoDAoJESl3BotkxAYnu3mFEI
++CrlHTDtem4+24dZQK3yQt2ObtEKFHt0W6SNwxaQ2rfo2FtSLfGj0zaO1gqpiQB
FhQjBMUa5D4JB45Q3wjSdt6zCOyfpKkPVjR/iq+eMpMyh2IDPfwvBZQ3vU0VZ8+l
lwnSZmCCAtdwfQjlscECoQ0i0Nc+u4gvag3v/0POi/7DPHmZsjpBOeTMOZpFEY3g
ib9AlDYnUW6k5uAOq+DhPtu/+kHbs/E6MTp/DQYvqLlTNIqhQ6cbYiBMNrhcZEHm
rrS6fMxeXcqvSLJ4nqOXshpeD3enEZLA4fQouQCfKqZbPwnEknDWBZE3HsyFYFX4
T2mUkp+7/QNKXVPzrEHGo18B+0nbZFf9wdqoQm9tLfxMe+cnKAO3JxjQ7jXtox4V
QLNaP13csjlequNEPv4Sfq7GrofFXV5nmPabEjRh2H5I1J49r6LjgEIJOBHVlbLk
lBTei4nccYHTO0ZmnRoJwbP8QSScxk8KqogxV/HaLCjTxwSmOtShGlwMvm6hNS8V
mf7dkgCQedVl+aYK8homi3EbRd0QB58mPdNe9u0FqxVLGliTnc1U03jbuBDiavvb
J+CONyTsP/1gtjPxEMPMC4vFfat9PLah6DDjrI48uJ3h5Hh6ZJhK751K7j0/XXd7
rT936nJXNnoAQZOXRPsjLsY8eYgA5aGNskvfHPTkLKiobAUnN/lm+3uPv59z6oe/
UsnZRxx77kr6nH7sgT5CtHMGpC7msSfyxVif2G6Dy8zAF3uoz0OlnNWn0uWI9lDf
h4YJlXzDDpjy3AEMEOrVSjwiyJZ/9Kgv4fjz2VdRagZ7T0YRNihFTUTQ04f+OeEy
XGb5Eto6L9BJsMzUdiec27PZRDa3gmijlPhKjzLrfA2A3v4rAUT2kjgVRGXOnUN4
dBW2Ljxy98jHBAcdWXOlDT23eg5cRB3TIlH9GIxa+4aQMmQeW+WyqRiKZlITacq1
SRcEOBp9Suc6UiLVBSKQnYSLYFFJrwC4B6kDSjKS1tfQQSayZVHo6gLlLRyXiC6u
XDymrL/jz6IDvs9jTODGO+plqtTBqyWATZSHaEcHazG94m/lBqV1QwhHIpLPBcHj
QWBTD3JUzUHib/Fj9jyww0WeFNi6UniTBhhk4E5a7n9AvfUeHg27BgyhCFx0+KRc
UbanoAAukj23YtSyheEnlCH9dCrUzSa5OEFrMdj26z6Ds3FTGywcx6cEWtAtVeFa
bv1tYFpVfL2x/9gbzIaiGsXeIjAscDKGD3rI/kmsOira/2kPJK4J/09ItTP++tXq
LK8E2HgL7mRFm5qC0eb1CDT7uAn20Z2ggdi9jEWn05H7o/AzpPD6xLQml37gnqax
uH1rnVyensCuNTGyhSh2QE7XfGkY+uavlteEo9KjwEIKaLkS00JBFYrPAnFhCanf
13U7vtnmcEz6CCu7KXGZvtgxt2sXM7SMyhcno+QsQDZ3v7piECPpap1cl8WVI+Vs
RsgKGYGcR4cUHI61cVDootOq8lCmblr0icD062qbmjJTciHAT/LkIg2WBAZurr8m
RVtTk+kXsFwNNGYXMbjyNhYzWzK9ZxfcgQ/eUqIYXgSwdIbv1+cn6CCsZ1C5f+NR
upiVYE2dRTmYYl3bT8Pw2LtWyb9yCA4OgBlUxPwlWFApm0QQe0Snc+dFMxIX0dfs
DqRvraEW9Uc24d7K2YyAcgJLO/sq9qaPvYKNMy7g5qBwKU1MuycflkvXj21Mj4Sa
YiDxk7Md5Hq1lPclIxQmPUwwCH+C+8HX6N1OBgh4f/X254NDm12m7o5WU2fdevw/
Rfc+E6Ym6MbGsUCCAsVRjnWrxVaMF3l3Y/gAZaLyzojdUVw/7pmqMEpINK45X/YG
+HM2PBYufslSwWPTy5/dLDEUJx6t0k3QZT1cHNZrh6QR//h2dlReA3J90yXCS7Ai
z4Kp2jfkiq2vMij7/PJjoRQWGvc6rdj8SjIKrSehgk8uNc/iN/QrDO8naDhlXOGb
Jk7LXO1tJYprVmeeU+vnWQSXMVl/7+yDEa0ie13cNEGQ8x6v7sGEv8bOLp+v6bgt
4NyrhQX8lapf2ljqp3vKq1NLqYy4DK3nWVNOgxp7Dut5ONs5noSH4u53j+4Um7GY
NT1h01Fdqf7ps9vphryuQKpraRPwq7cVFEkx/xMZCpfyM4u02oCJRspp7n0ZY/Yu
TZbkyLzXPUrGhTnqfu0YapyqLBpv7H1loFbYIwiH9FRqIsEWfWqAs0l6kK6N0u+g
4ASDUviSm1MXrYCCoQuPx66hjYF0G0LOT4fn5rZBwG3Ib0rvwQeNsnaWlqaZUEHJ
wiQU/la+8ulmqwCiF8OAVY0JD/MnUqUwLHXIZiwrs8j+ds+usT+QMtNc0k/0bt9c
BEZ2Pviqc2BIjSe1RSrw27yHPcFpSa8Ib2xM5kGuEYD6SR/Q9KJOTPMmIaCLmCD4
NGrC2mypRheuLcT7OhXPj2rR6Mr2AkAppvpXGp77K0FE4ZAkPYiX9w/E6LkZ5r1E
lexNTZyOZuwRxgsUSyrRmBYEQxi7wRDfnn9ENwv2xo+VaRnXGcaTKb5yjmgHfrBq
cdZy2rtFUE9VxTHCJKOROuOYc+tDTiFPLaUsQN+j6Xg3MRFCu1idVSV9aoiiROyu
Es2sTFd6oF2crID5AYFK0lPr2mLS80UiDyaemgjgmnJd2cut9dhdpjZBQhZWhl8+
gjvVyZ4FJZ6xBTlEO3r6SZYyQYG1ZvC4fJKKBFTnKxArQi/9qdKpLSyQaZ+r0QQF
ZthCOo6p6q06SNi4ENuUJRCVhUbY4DH3cYrWOSoL2iH+UZepS0Ul8wvcGKo6fttc
Kv+5fUZWkp1ZIEtpzR+MF2TceCMIEFMo/zmEJDNWR7XIL4+j+Y/sfjOD2FjW5Q18
vjNby8DumGEl1RHegQLbFR+2SR/pCvTYDQyeS7SpOu+d9Xc++0THTn+LX3crBezb
bW5IXkXqcLOPq2uZhoM+YO7DDJAymNuOEF7GcM05oUcQodYH4UMA6waHsMrlsZGM
EKra8HTk6QjpD87M92t/MkuceqUP1UTutALb31fKYPMLj62rpj1RQrxw8ODoUlsJ
vmy2qaBn45ri6DZNJU0uN2RvGyf7BniekjDOIsiE4JtCmtdKfDzmMoGaBwSxVtZX
cFKX16PBDrAhWoyqeNSIW411m/3mTw8a4QR06LXP6McVW4ixdPZ+CXwnGFmEvPKj
Qi91WHaIaxTWOVHPioX0qrSE1sXNWcJ5qzVYcGr1ph6gkPueM95rxwGw4pF+ex4i
BQWCPuD1by1hoepnUhPOKus+TjbRPvFKWRP7jqf59ll6gquk588J0bYVSAw6UUni
5SI85AQeQyT4ytPndLl6g3XUINmiu/t1CS76OjBDjF+7IxQ82JRJAtALzQ4l9RFo
zl6JaTIIg6SVZ5zSs26OlZeU+Cgwx2sUtfbC4yqhC+8152zFbxNrtj8H9WZ7TTrB
H7UJVXmwxBhjlQChpV76SS/OepxvVVej5zxzpzIFfPNyBgXQGXj099CWlxOQOnDo
sJ4YKOnkMwfPgFG4EAqbwuDKXjIN3b0B7KH6MhdECaErdJ6AHsuyFh63OR4fsTXJ
CoVc14iIRB8j09vK5fGTGmy8o2AibCutLafvw4SREMLSuQU/x+AoI6bBIl55d6NV
0nNamAugD9IruV2aRn9XrOcwx0HPRaFaw9z1ErJPzP5s4kxJb+bdlW3P637getmD
XGrt0CQ6vm0u5PzrykPCNU5dBgxQXQ5LRzYUDEvd6pz8O6Z5VY4zavbHew92eQrT
QLvMc45+wYqrYGQrlCZyz5b/UT/LlhX73qd+kjEVkmtZhrB6myWigdMkqBeVJ6+o
/0d5zANt7M4Yny6f0t7lx3ffbVlTTGm0Rb4513wsqTWgryjeMzriQ9AFGo/Fzlz1
UuYt/TJCjj6r33kmSkLgXFp9Ogd0EICIqnOIff9JKKVa/WeyOdDqC83d6cF+Oep6
K78Ybl5ogmtTON1YbH9mPaO+w8XJ9i7UK8CAk+Rpr9GcPRS17WKqotmCuMdFSofg
2Z/raVTJfWyd8ruvZNPzSXYU5I/unC+R2u4e6DQXQaYcdxcrYyP1TbRQ7cn34o/o
shC5QdDO93kletsDtQwa81ylJKapVGcTxjpK+XLiMIZPVxlBwf8Z2gzi9SOUI+Oe
71ppJ3KzZWi95BzY2F/NV+MFEWv9MvoJE/jEOTAFHUE15dsYFY8oK5bx470gdsgB
KsnH72mqEVgPftXwUS5jgNSLbkoEu4xAu0cF4KuBeAJbMj17qIoguaOXluu26UIt
2RHg8+iTRviWajoB3ZOtm8XifG4CkqJPGyuxuZ/R5QKAcymjtae4HVeXsjoHMWBn
daHlS6+pGZiH/ZXrk8osmlpd9gRgYvWYcGvZo6017BFTn+eK4Kk3FeCFLMw/XBS+
d4fv7b/hh/ayE72Dej/k5k7WgeG/kJ4G4vuczm66YmZkbTRehe6fHBI3nTQqB2YO
eeeJNzOyZjmeZGwLi88GtBQND7/6/AjrIcN0peZums4rLT/AjjU7WI3Ky2qomYaz
DRnjPQPwaFOVkfWEn6bYi1ZAHZ3sv4jdqjJ1Jr1RX7S0VlTiIJiHw+G0M3Vs9l82
i9zZR5HyM8tEhIernXN7tta+7hZOaAYx+Sy2t0SDR5UjONlqSfWV/1Cltelrsipp
+EMj8H7Zb3CS1sBLdWYzMidrrfrjPuHs/4nHf6cEtVheiZU0/1X74uX3dTvu5eCy
+aLfBv24e2yPQgB3tsGLchYd0JSqDoGR93j9VAgr09dKpRnbITZBqXT/US9eCkWs
rDUMAVGShHSPHPbg1XI744zZEYp+dPdcJdM8sbRkcy6W1qpUgKLFp2LHWeKIsPCs
FiJIJ3HDAx9/GZZDtZxNpbqouV3WIiqhpkNOKHKmB6flBWkXrzy3AYD+Lr/w3QSb
cSOj4wIex9n6fig3ytnC0/2DirLpb93IXFesqw9mcJkI1QQZo/YUZeO7GUjs3b5g
yLybjuo9cjCQWpWpEOaxIqaW80Yr8nBP2zXS+UopAx6ndUuZfYeB9pbg6ZdR1R/P
mN527NBGUAUpO+cP0XeqZSi0GU2lKpo0erxSo/VBYZMOo6LIcmqoxhIbdV4shpt8
yxuy5zyFRcMKqpuxslb+v8BQkN8hBaPRgQO0Hx6X6MohGvqYVqH/b9taCz0L5Jnj
aeycE7wxUg0VmFQv13KlabXq6bX3Fr+lKW5Jg5Xlj+89lQxkBogzgKiDfnq9r2hU
7WlbDqBsN6tIkP+8qEN3RdkIvr/F3h5mkDsXX68IY1GkQPKHaYi5Fx3fs9Z4MbMw
35l7hsXErOiRoldqVmYaW6yDo9afoxqCRSugS/cu0s+TwKfLXe4MRhktvnSeko6I
DnsNQS/o93AR2ZC6Y7hIXZmCIVYvPPuBk2OMvGkzOybyuBT5v3ahj5FobnfDK8Ld
8AfRDxRv2ghKRz0LxV/BwmrxQiCyfXJS90Y7phttV99MXqvSFtYr59t15pHDIUrp
Ry5Ewzy4z4OQyWLLzebgy0kQZa/hSvGzOXcyk4Ep1fkMpMktLW3m2ugTd+MP0npQ
VnoC7xpCAJxzJ/JdJ3+PF6d6B1550qrnMvS1kmaRKLO6jxunAZgWXj/6Y65g9AVg
3o6agvuWK8GuQH8BYqd72tfvQOI+uX8F++tHJIYdWFuCaBYHj4mqhYUArNFSfjJx
LtIJEs8E9ETM5UofpW/SoiWSdi5GCLWRfcqFWXW+j/EuuzDC9kisFOFnIMu5mgR8
BM+fODBCe5W58vISOm06rRnHI+gDV9MggxDWwnjno/WxkBGbrnw0khAJOWwnaF7+
tIqJ/Wfiy8IKZ1CnG5UX7U8tA9f+CCj2dgXBThkVpjo4CTb3FRvhtME8frHEDsrM
rS6PmrJMvif5CSV1fw2dwGnufpq9HoVVhPMUDxTgP9FzMhX8a5KunfEuqhEtB/UH
XcM2EK+NuJySXaOI93JHjqqEi00Gl96EGlscFPypI97VvneZ2eIBm8pEcMWmSO7O
5cEuTU79/fc/f5iQlPRLpmC9/7ax+QYOOTfr+rDV5z57UbXHYrVgyoIH31nBzFv8
3s29XVut6PlysODJGKTBEa6IfVkKv/2H6tZVn3pC1dm+yyfZZIQxcGFMBzhKa5mI
9RXw/2ZHieh7azPDZ2uA0kHaKqYm71/lw6mEu3CJE7flyUel5g/Gha1F5M9Zw/PV
jKvlrPMw5ruKDp0MJrvDkJK6t9eRv36yYpMkVOj7Icjyajk8rnqXMlWr21XXA/HX
Boid+/86yKTUaJVi1Y9n3dh4b2H30eDKNXBpUlJogKeJpeZ1Jp99vd1UviuUc318
pv1FmOGwj3BPU9iHOXyn4swAoFmaKOfIstER5ZV6kPRjWueKMFwSIviV8b6EOcVr
T1030oplvd8JNPCf4nnvThg4jcgub0C1vtv2Gz98oyQ7YRsTm2iCkV1s5GgDXYV2
JZVp43SdVagPIgReI9hgcLErVaXpSNH/QkqrCEobD2npS+tyWxacf52XXLJr/E2h
HaEFqmcd9im/GaRhOMq9u010qWhgm7ujHK3Y6QRmr+SbiSLXU8VZ7yVTkDyyEUk3
8T4rryEcboc4tijkx+99qCa5RZF9J9/xbSPu2jPxNID93drB4pzkvyez7cyfaN2+
zItnVvwxFU8Hf91NxJ6BeM4mVPvUveRCTf2vzTAH2ZPq6sftihrXGY09psSToKIt
QUmhaotaGHK7UOhdzB2vp7GZxH0Ya8/HpPE0wgOURsqxTyy/l7ev2t3MFMGtC8a1
e+Gddf+xi+XyPjP1yrx1lLhJMyXNevKRPkO0yeDjl2sxjDV/w+MLwgenwOwplALm
hCkQyfvSz9eUw2Y6Enrq5jYoCKXS4zBbKEU2prQcfG/E63tiG60iylxTMq/C6cDm
QSjRpkmJl4TP8og0du7vW25T6DGqom6UJLsgVvBMC3ak1fowAz5Odun3CjJ1qsZx
cbhUXA7K2k/7gpLeymz6nFhPxCtGag6j4yZd1kaRwkC5RPXd4BiYOFUce0gCrujF
R35N/jnsH1IT+GFxvYyIezcgR+hH21XV95re6E/lKWvhX/itVJ7NUgaDOMoSuspA
QeOD+nI2a7ETf+JBZpAWMM+UdkfZBSOrGcyu8G875oC7wdsvsYOYJxhxzrzGYVb9
flkQ2T/9fF/ujpkb3I9E6eKKJ7+BrQBe+Jh4kwQSbH83vyAlFxz+jTVR9XRGRO3X
1xxBQbce2fFHxN1teT56rCtbSfpCsbs5p/6rqvIlEJgGaXeexEw6FIhFexdobuFD
tx/CnMlcsqxocswUKHeBaKDXPBuuv5jCg4MSHWC6j42PEYkbsipHTduuVALt2jSM
fIy2C2mb40fNAGqfRYbALi0orAlxQrJWWxwNJ+oNggM+shRYRzBh/4uVPSeyeSxs
nQUlYccjwkQtb9bnOCAJZZrmeje6NLsmCS9X58slYfkc5SkqMnqKULaTw0c2+Vwk
BsKUIIITmx9X/Q0yNi7cHIsFh2zo667bSrOFCzxtyfknyIftMSDXy/Bsbtdxr5j0
A5qJMu7WiA1AyH1pn68JqUEo4XdlbNox4VpY3sk8v16U2KfOuqkG/pXaWHHPa3e8
qWYPkDcRBWjL0kvAZhM5zs38fIXlinVDIoJLLQLgVSDQ1QL4Nm5h8t/ftok7rTyV
VLGuWTbUHwk7BTPZCDNMnaYRprUbEgWBGU8ym9L714ZCdV9jgZ+iVMb/3NX3awHw
9jaeKQKfnSCTeD/fCJgfi+TYb3wWOJmoLJoD+GLM5/JFU+PHjj8pRZcQm0/VAee7
pnLH2TqiGpUKiXmCcbB12BFStioykfpk/bw9gualXikXbo10ClKEtHyM2HmU4DkL
AH27PkSKGV3H+v8lpSDazsO6zzo1vjt4dRJHcQQcaltpY9qlXVhyWeU2KNQ6y5OR
JJW09DaPuFLBYy9vtiTZvR1sqnEhLb/fv+2j3rTNOkSKCds7GuWpc2CyEzAQPN8X
CJiT7ePcjGjrxZbuYL0GQ2BEnF0lXT1IgxPtcRM0wIrHMF6AdB9KzJgd0hoo3F0G
/FQ7a7IDaRwhJ7OxRaRdo3lexJm1AS0eKXgo/ydZLuSmkWDFEuqlbz5K8GSfCZEB
QcpPcPbWQbF6Z+JHhKiHFz9GD0hFTIKmKEYjMB7SXaHYked1Ldl2BjXWm9SwT7hh
3Zjfha1llLdwjBqvnTjB5BBPvxEPdAH9fUldVyOVM3qetlYtK9dklzcbZ/rw3X+P
KaLyTnGGTMlD2pOT5W58at4dq/+P1+i5vub1uN0uujeWGBOfmUNkctM9wzrR4gcN
ClF0HMJBytfybSzxzo5luovdRrWpGfflE9/TFUVwp+YU5IOhspglNzBAUAP3DQ8t
/blYaq8CjNz03Vrf5kYRphInwyYzK4rd4LWedk5w3K9DGf0LSKgJl9SYjz8XY9C7
fu5+Ddzwyec3reqY99fi2p/z+ucbS2vyRlCSgByTgwjCMFn1LZYg+GsVE1omWTCf
odepfvC2KXQJWTYsIcYlMhoPuVdOz6lCBggsg04mNLG6kIZbCszEkszsLRMFl7NM
CsAoywFZmt7IaTjCnZU4bt0SAPpikiOe5DmRlOIkqSSG4lbEE8/1384ivp+wtbPn
FfGzH+vZhq4ztMdhP3lHCA6PZwWkjQbxGoxgMF7waa0ro91uPOmVRmBzNwW3zeDd
jlMxk3SUG7wzqhwzp/A6shy67JS5GV+R0G5q4glFfaCEfUsH85TKJsiMZ2NfIrJt
B7nEa+RO637OS0b+CibJ/j+1mMFqZcBUbdNEPecN1ZwuwN/tDdhBDiBpwzrzN0p3
ygkYZwONGgxxxZZGKVMoWKGhB60U8Uma4fZQ7T2WYNw7s7Jktrw/YeTyBQ6kJmMC
obPQZ6hC42yfY75NV7af92yOl1wlQGIRUbGeiAd/kpoLsWm2tSI5D6w3+Q7Xhp5h
v2uV49T3EkjO8Tj8P5q5WbT97305ox0a16lWH+Iao2NLdaXHZ9WoEK7CgCweHzOu
6kL1wi/khnG5k4KQnf/NlHROsmLIWi+CXAvoQswO3Z5XH0cEHgDt3FxIs7XcgwnQ
rGEDoYCPyXknSGkCb9cmI/fgrnG2JEWsYo6a7ZU+uuJvH5frnTbwn3zGWHVWviu0
5hqCqF/j6v4Zui9sQQYci2qzrh56SQ4LYvGCtzX0fW9JGzpcRCDxdODmDT6vDPhF
8AeBU4vhELHll78OWtNTyViErShbqkp81dZdcfjmxzcJ7MjNNBApORsUDFPMMbRA
xWRtQhOqzSyfihOPGhc4enVzdPteUE4wqURSJEf+AjCdwCB9jnfIB9UWLXMMDv7R
R5gQtUKjqnegwR/EkfxFq6IvBKQMrba32LrZr/XbZpJ6LeJve9WvklOYvQTTRP1P
a6dEFGOSXu2tz6w8IS3w7RBWHRfCkU2HhedavQVEXsFNTVOqmnj+2nGPSHQe4sKm
m9e/DVbQAu996UhwjkRM9wP+8zCeEhGCTuSzxLq8XheQFX1hbj8uJDv9iwj+7WCV
xo+F4WUXzw9muUSsixrBzcfJE3H2Zr+Y0cD+6NxCLtVmKYYH9DGMuHTlutyQfpsE
l0gunldMlVO4mZwKQODpdmzHvEKtNk/HzcKVe5fZt8SYjeKiqrJcE4CKte+TvcIi
H6BRjV9LsMnIAfQGC8f0p6dKyhw7zDcaJgMjn0jnFTEttdGV/zXOsxzPmBfyjUpS
OjMawj2FHsSII+Z6rIokc5SjBqV7/LWzgOn5LM2cgUpFP/YJoBUGKToZ/Sr9WFbP
iLMehgWSmvxjzgCF1JE20wE8xPVVe5RWR8uVNgdqwiyHb+i0JPqBkyhAvLF4qowU
zOUCT1EwCcb/Qa39mB05q0s6XFro276//lORUzSYXw8Z4bDmhvMIm/JWdHUufy5n
BwZLwQXhB/ZsWyyclcYtS82ZQwogBDC/Cq/3EVqiPgu74G1BSncgTb3PtKpAFKfq
rl3oWBOjMOrw/34cD6B9qR1j7ZCjsCCgjdbuYd4H3+YAylE5pi2ghy54NvDAduM1
v9UWy4jnV/vJMmoYVjx4/tR2VtSGYVLvEeq8VjVxc+puOREJLCsmSpFg5mzRkMn6
EVmGjDzhtQux87xt9GI9SdjSgVmsMGt9RkYXs9JtURfKy3lJAVaE3j3+uaFfOOPK
2VKqLtEYySa/O9nxKMssQig4vRqv1h/3H5EQhoAlAxqUWyGil5M9fjx3UjZtnt35
iximmpQvZ3J1lORpVIg0UTi1tFOUiuUUSa4D9p/ZG4SBvQUaYJcScifi0T6Ts8/l
pWlzJIWIqCEs3by/727zz3C12nzf79HADhxJboqQ8eIvy1+RY26jSHuXmuVacNQ3
isT7Ugab1kAxLy6uvCVHO+JrwxyXq3j3a/HgAezGSizwS+I3upQQ1+afjAcE4xgw
oGBreVPOZ5GrOswIit3yc1u7OZD/wgZ4Qf5RJdHjiH4efXrYJrROSR6NT7LXfE1K
AUWrDnQLBqYEV5DLZjt2q4FJP8qI77GQ6ZRlFRaTdOsFIPoBzY1e6UKrso6nZuf8
3MhG+lW3LaaQgv2FIX0xgexE9qb+GiMeFdNuK3Evtz/2B3W3TQrl77e3+t7v1YNN
YX/+MDyELDFwHFq8CY0YdFAZzgmHrQU6UDUuYCrA/jIh/iD0RQK91P6Le6hwSZ3Z
bCsNUGVAqoSiR7GZBKKwkJ6EaZlZidqbAF+GCM/WsqerI0VmLu0bC8LTUKXqqG6M
Uv7J+SmIYhgm7gt5PTe7BXLKd0SziM4AYqRL5ry4NXWfnt9jBt6uYOOsUqXtgVpT
K7SbXa7Ly3stBAzA+gXelYNRiQuWosPnkFEZ704Srrv5mHCGrEjU/EnH2CdoyPtF
8/lmREXAorgKdWG0ZHcMyrrA4074b9Z2Fns8ybVgqjmsYCaIHHOTlHhguAq78wND
D52ycazvamfxUJejmJj6zT+bOlcsjZfT0mct50Tp9dczueo5jfN6p64cf3lXjL0a
dj6ND6Qs61AIz/yZmzaMt5w8PL1K4ZfO6MWIVk4JX9aMFBiYpGlZ4Z0djbf/z3jg
P6/rctJKdUktFWHSAs/BezOhUFxW3v8T9dmGxqYJteEH/RBc3Jz803PeXkE6Tl32
Wlkcg8gna6pPBq3Hb2xWopCn5Owq16OPpZxMOWJvJKO2538S3T5PgooAEiUu/nSR
r0gVZi4f5Gg5u6GGKbbhVOYqAYpVzSmwjZHscCecEo5vEK3dsvniLvXbCdTgiQKQ
v5au9nEWVyF/kZ4IaHO8k2UHCpq9YxxRfH7MIHM5rBiGifEwqUaB7uNPLQRQHKtX
iC7xIjnbfEPNFhhtL4gdAaugB8EiKIJsqQqAIUx9As1t9E51YOOaJR8SL4nNXGHo
lpdKWamc57X4G2xS32uPJBSXR2iOT4TYAt29XlhldUXKs5i1BIOXVKlKuLMtY5s1
6t/ZY9ZPw3BM7VnWbFnNzvshtGBt1ToNJRxH6pSCUWinsMf3zicncMbnxKp+rrij
U8Vtkr7G4AKXQGSmTrShr7YZkJ8RdDC/is0fCV6UqzNtbmm8y79A1PobvUPTiQV6
PXe0cAuPxdwLRe2X3yVNTB/S1BYy5OhSnEZtsCyLn6m8H+OzHbrByCbrZ8AVYjbO
ZXNG2At24fUFabEU2wP3VZX13+KtIYF+X9uRl3bZnUOvRG1JZtLq/t2wDX+UY3SD
ixoC8f2kC2NOFiPlxYZLDRAZuAVj9UU2dWwutxcvVFed+BqU6dO8lgCg5klVhCVI
HtBSmwRD4x/bmOaPzvhnwlHHLOzBKkBjfpUNApUMWzxKXi0Y7JfV0qVZXxN0Tk4n
Rl6aswC6OBGCK31d6HxoKNj2Vc2o1mLoPKxwtuVYSRkAp2RqwgBFTZW6r8e7ldfM
kMHMSCIgTjiJNT4lah4HSDsC6g+/SXRjV0Mog0Zqoi+o7XjPgAkxw309wfdbkG2q
GF/+q1H0i5SRHsCOeCkwod51ustra+x/pof7aILjJAyPQGAfplBzmxDNBb6VT7CR
b3XBVahBCajkZkhnS9/CGinHOUSg3UBKJE6BLScItTgifFC7eKcrAC7xKqjRrj/F
J3TPXM6qqP7FQe9lS/Q41FNKnPf1zfEqZYV+Gwju1PDsLCOxyFO/HbUwKl+TnWj1
fEjg6pVzfY4QLMgKSI0ji8AM4AnYoBofrlo3uavEDy2aM8y1MtiybiT+gQQEbQS1
1tJn/shEQ1j2/AoEmLGQrb+6yp1b0bD+TJTkgw7xYYKkSaIeSz6NFCLzU3RtoWjH
oNt8DW3U+zxrARQF/Wwyt3KV+z7i/oYic8hapq5qm0GWx3ljNmodvpz0c23i2LwY
Wknpga72/ucmsf2Emuaun6c97ED/CLB2pePSiApeRUNNJMRAH2zhMTz1FEkVTWDT
gsHanDumlrPGjTdULEAQxJZ0TOfCbnd8uVp11GPfb22K3CIdFMoGQiDvHq4vE2LK
jpE0dum+qmL8rRViJj7uZW6tl3xveFjKQUKW4F/Ly8tniy3Aqee1WfCFZaiT+bIo
v/Czpr/to9uiDAqimVSwY6xFAUOlKoo96/BBHJYD0xwp0nMtkXJL8Y2qD+0wz67h
G1lkD2XzcrCrrGLu5tqx9Wgy0trw/7lU5y4loEQs12akxpX0PwAeEEG4cy6bTwXj
DFxSvp/EyCL2bJCmnvUeGqb019EqZKeTs8lOzs3cLyLyPGHMUS+CH1jTddAE08i6
aa/LNyV4MZaLhLGEVNbQuhqeZDMt8d9fOQo2qwAv5CpMfjsCkVVSENIh7MjgNTyO
cgw5iZpqI8Kz6Frdw4GfrnKcff3bbwxlJp7Fnaskv/U3R41SoUn9sSb4UZtcttN1
cYOxs7bD15hQt8NY1AAlV73BJg7tZeodwedHXFF1Y1TGdEh6fCDxHqkisIbRNzrZ
8ZgNoSy1WlZd7f/fM5RO2a7X+iZMWQH8YH50aw1/GlXqZwHZQw0X5DDffwWCaQ2M
nzG8N4h7y4JU8yml9GrYZ3X3Hdx2+BkQMBHTFBBiLRbW5NLL6sJDPCOzFf5CtvAa
fVJU4OptjQK6fppnp0E8fFyWJLT1ijRJp0qVyGwa1gNhtbXy4cbojpHS1o2hA/Z7
68puKiW6o7+PJt2h2DdkEFvT0s1ScKl49wMFIi/j5OUiuzU/6c/jJtJLHtmqjWpM
lRg4pRY8q4bsffjMnIvDk3LtSV8GVGIHdTu/iyoR2w+QN5j9GNdNxo/tR0M8uAwd
5awwntmcemHdA1bwGTQZfPPcC/kYHkou4tBILAENJlgghqBeO1ozdwh7zeuNMatr
jOs72IxzoKCpOPNam/cT3hHvDXbPeuxzwYvparSui6OBuy6ineVgbtN5bg1Vsbq4
UO0wOqtFCk8a9bT0avLsNF413hlQBKaNs6EIjObD6f5pVV9AwU82AYLuirw71DJ9
+nIN8Ky5nxoX2/vd1cIaBQ0GuPIlbb4AJ3eLKnVO9REW3vmTl5ZTzEjcPRM3lIO/
LGhAqMtjbfqCaU6JqO1SG6adWSIDwnQ04JqdZTpYaur446QIUr8xwhtcinir5PSL
hsy6U7frXfIa6g2JquBzYxQ42U+K7aUeWP833F57C4aUKCMk2hWyDfKbyWCwc92i
AY4H5LwYhoHXKkE6xNeVShdg6dAEmGUxusIi+4TLApHv5BsALPT0vsvjEZpgNLLd
33D/qZlandaYOwvjGWNA+n3wAKj0iePxXXOO2FkT2RmsvB5sN2gw2YgRghiElrB/
Sn7q6VuxcVgg2EyZI5/K+zbntrhpwEurjUUBTZyEHm92fnXoS9Dky/jDMqVFXJvJ
1F30W0VQbCrgBw9G2wp3GT+LfByXCNVWVpaBJlnfPGO0q7WhWxaMvbV+UmoZh0cb
WgSA/g22mbAGPpYXZz15etVX/V7Og/TGgI7p4wgwYlRbmLltaXCBFqN3sKjfvyEm
eY5PtQOFzWkHaZc+58jSOzSW6ZaDNoU0SLgNKnKSHfaURZBB6cDoAKqGOhUgEVmF
huW7QertnRyzIMllW+qzZRbJCxLP6lzWTUUxz5NlRytINXVE3KYpqbHNffgCZZSe
bozicnbxXINQlfZ4I8df4KymNCHojZdINGahTMjw204zlzYwNG8BXB47Ooke5Pyt
MShSEKHX6bbLunq0H/OE3LdWz7dpQMqDWVaypAgoPtSFStWKwosk4V65FIhxJuaC
zeKtRl8YeiI23vtgUl+lBfT2UA8N5HARk2GbzzCT6plJ5hqmbK5BUvv5ludzFOCw
qIuV0QdU7Y5YjJR8q4zi6mhGsQt+PscZKvgWuAD/evNYOZjXOPbU+I/wBUC5WH74
RTvvCCftTeKfx3sssp7PZuJAqdX45iXCbQTab/2KDVxNJ7GfVZMbiBUgHG1jK+Vb
btQS4gAAIlEr1mG/eTjbvBpmEKZp4gAgts37PWSySK+UWq3kobfkI839UDihyWxx
ONmeptZitrOIwaCX8eJn/76DB27LFmhm4L8uCPb9XjaQt9zuV13q5tfW4v82gUKp
5D3DX4iCWKbO20ogXfquft2s9qvSN0Yx8nBzJ4UsasSAIG2tuzri4acS7ghwt4eC
arr36DMchZAW37dnhv8sYI3KeM9mP8HJZYQdVJhlda8+4ibGCrnl7tYe0UpWgR0N
Dajb1IbHaiMTxrzZQByXkdt4fKQXXaY3XjTvQ4SOGBxZG1jmR7pu+f5zFqtznf8F
5Jl6FNkINf5Ussx7sN7YwQdsVQp7KnvAmtnrgyE3v77QX1oaF7Bcl92QOkVjKB3I
vjSX40557/q6S2PzrW+704LBcYo8oPMYV14MKy0TzL2Py3HKnfQJRd+Tk/QhmvTu
zWBX1Y1OiG4lPJ8M/LwYrAPX/N2K5LwCJ/NQ7QkT+U7DZtlN/XtCoYiTmPk79XSI
04ot6N3oIAt1trk3W85eMBSIV24wdSfgzpk2C5mE/5pICZooSgzumBK2h4gu+OOX
OGr91XW9u1anBSLHEcPdUzGQcsNAwW+V+oDF4uONMt7xf0KREdBNYoTh94vAF7vz
xkr8PUXlMLYZ3iAm3wTF0zDrrrlw5WRLmCoAQCVzV2O+rmcdyPAElLIFC4p/sXcU
YEHwCtCLXVR+9oiMAVsvRYz6Fg7Jq8aDmmxPfAe0Am02yt25Uyl56TbWexeUvOwO
sKVjBst+mggqEQP1OukKEYeAZAShSboJ6WtnnzgJow7qCZTfWL+kgktPa5fnRbMw
51m0B8xdr32NQeqHEE9PGGfgxNOS4cZV4qBVtoAvsr2sfZIYxDG/un26zSHenqre
TvuKtm0m/nljJzYwdTmVFvN7wXmItLUJYXHIwDy79aQ/NjXSWUuAkZMC45RaXrbp
izhBSXRXL4UUJJ+tpR2Ddj+4+Gmx3Sql9kHKYA8KYR7zBNRmRc4gQgrPy2oeI655
sSsM3j4g7mNXzHF0Ar8wqrP8uMTKCi0JBUBGFu95Jio/bRsrLX2F69HvyVsNpkwv
WAaGUCiemL+stqntYxkosKwTE8KxwSy1PYHJtx+0LzkgoVmcUzn9yQ2ZZDO3rW67
EsH79YXhzw3AjFjiXL+ITokHcmmfBRq0QhKUiFwecE9M7XywdxyEOSJswvTT+56f
oohzv0ZcBM5j7yETUbZE+Wg2kF8y7Be57h2qYxxUSsyla6UDAjl2x0aSIyol9b4c
OuSfiDacVRpSvixyC5QlkQoI5NfAKUjEDS4WJiyIESn/Z96u9IcIrW5wsW5DXK8l
YOmRe5mJLM+bPk8YEOi4yd2GBlcWKh9wqRZe8pAOnrw0xQR4CZ/VpTEgt8XXayYq
LScQiKLk9/glLH0ooAEBhHAKnnPG7Skl0EoXftqTeOfgPNldn9kd0OBsz4qOrrUP
KHGOzpVfIsKAQdE5SlAjEXHsQRnS7s6q23dSbl14x8B6z4f8hd5EdX3qWfLacSnj
u/rYYXv6xq+HQXnyOz09vP1RSyqZxOBVSSxpPI4MjnA4FqaHlC7uas1BTduYN0b5
Vbr1+i2pMpl83V5N/Akn1eqI01Gjl9PYBHsF6diaSEjS60RmhN9SUgfJVbF81EFi
/oIkWpAe4BJvGrl0v9JbqexUQBDvDnTgvjG/zb6uY0+5T1GCynfJ3K1D+8gdIzIj
1zl5egVPvuswtV2CMrjkBEKf/N3M18hZOEI35E2UsOZ+WPsNv9mhCj4mpRKsxLDB
5jrB3qaQY1gCBtTyqqYJMswhI4hXihl5mhxCvqrfMeox3X5XLu1g8wqbqdU2kBay
G/3HI9ye3FawZD08EQ/E38b1BI2Zbodvwa5tihWhvOmatK3o532uLneJ6lbr+2fU
AyqxZ4bsJOdGPkUFRaByDlNt4vhGCbPbUGFJR7cuu5LwcKSIr1jNT+DwLad10jnD
22kH97Ml6EepV1osKJNrIQTz7dLO1+VI+ikCHLytsGIgh4QQSFtWFpBx6vriziqt
jZmwJGBtZt3luU9Oh4VUAikZpLPT4e4ijwNPQvjCuMyxVSfAmw4RmzH/N2nf71on
0smDXJ8pZAERXXZ9kC8pwWmg4lfKbXApZmAWDB+U4Tfyk+eACwVPnSUWHYzWgEQM
vQeV3+XuzlqQUdB1L3ipWSuijYdMNcoN2l9wrZF9AgSt4AnQGOfz6aTxmhxOMfT8
Jt78BBgpSPmDsujpflUihzCLhy0I/+W7EQI3BhPMstRvNHT99D0oJZJf+gabeI8g
wIVkHbr/xt6u+QNH1Z6TCIx+7cIBaTAqAAkY5mw0PtcuIwYCVz9pI1Cp5L+Qo2AV
69WMWBOq6ltgMZm35zFJSR/xjjjb2PoBnRLoMvPADh5+jVHeku4gmeApsBFnPw4U
qK7EcOv6+m613mxMzsF1TTVh7zxTcbuQsnv/3+LRXEEXqGCKDEFEVgfU/1nCd5Y8
uUQn+iw0P5CfJk47H1/0odRvk5G4RxCYGCijGyJG3I1VMVM/eZBJh1dMnx1/PE4H
dQSaw8Fp2xvwDDyzknEqZAS3u8Kiu7E6a0CjNOqslolDgN6S/JBm+7hTMIYaD1Lk
/4bjls7SmW7mrVfT77ZZkUO1qUsgFHw9yiMgYg8CQJLUBJ9TPXE0/MLTnRSQ+bhe
vFEV5VBJfFu5FlfHrdBe4DrZ/DqPTyhzgZ7zRk6XuIfT90GmCUiK5+k+42T6lXHA
Yc9wQ1EyuoG3xDVJDDLbWEha6/4yNNTWbJbWbrByvtmZqZYCbEoRl3JO4x0kWoX2
oaIN1m8Kp5AT/ixdFLbfxBcncP0GRSK6OUcHN50/ysl0oUcouBIby0Txj+NkPb8I
TzI21wWwSdcwRgISlxFTowvvNJoGu6F9O71wcsO7IM3USdNrF1HtOmXmlnMx2LVU
dPUolNGBVxba44OxWB9oNGcpCB1coIOiRMM4gLQ+emR8DAxN1qZvDKjb1bDArBUw
AXWzTa+qgG4gMD4jliehByEAFLOUvTxzQvIXJM1glmEUVSg5n0DNCzxVAW53nr/+
6r6bAMdee8hIdyrX0buHuzkyZ2yhMq3Up+wWbHf/IVOYTQ8ZMK/ygIAXLek4/UJe
ZJaii045u3uLfutii58nM/Ns2munqbtHNV7Zi3VmfyqKAY3lA38BVBe6enU4oFAo
fDXt/9hrtmhlihU7X4PWTAz6Ml+iXBshsOVNXsEIhs4AYZCgJRHG/sY3talmAx74
MvEYwVHtaOr01svO60LupBMbzEH4TglXeZcntkj+4ESwCITP6JAKnDpRA2XjsXtA
0jhP2Xp9A/+LWrIc0qlRkL/v9taL++8JH8ZW3O6Nhb7isZcAKBPgWlqPyt3+n0G9
FhsW72/137NHSZ3cGXrULS4ZdXX7qTHEre/SmPgShadIy/1FLBJH6uXkFcXFtQdO
7vpm8XoTfPUJNnIMNW0MZUL7PwtxmUpZdS1NmPQZcmbhuNiyHHlHVqsy6x+x2Fsp
/jehFSR63wPQ5ZQv+kPIBgQ+kkncEq5Iua6gUlg9VSwDEoKRXf5tbZ1Vrh1XbmE7
bOupi329SLYraXQI2HrMVkRIJZxHWoBG3WaQGUJq3fCFB0B3L9Xq0dG8Wi66OQqL
zYgu/B2LIn/8OWbeZaBt6Vh0ceGGiKr5cRFQC4a84OiXxPLzcabkYJxmz2ODPIw4
0DprwLmyFjDln8cK9fc2h4jZHL+ro9dty+0zGjL9i/Cv/Id+OJQWAoGBqRj+aGvN
1yeou1bPHWsp0bdEjly8Od9sCN/CwK1Mt7Gv6X7O9GCSp8D0w466NaYDkPWA/u4H
6bptyYIZDgJqHGvn3zKEcJlpbZawgMOLzt/ViH9Zeivif+ZfS5pP+vz0a4P88kpB
8HxOCJICOa/zh9onDkteUf/F3dPAzQ+5zwKeSudPdkqPWGVNSndHMNwITJ+iLTOd
aVZ8y1ZgrCJn74CsBYVou0ug7QRtAMIGKxRoVXauGxerrDn1Wpw+l9ippX6u/bBQ
8BbAB+HBHkfwE1WOOwqbZ/8U6+jIRf4yyZd1Vt9PTCUb9jFvv8Ay33Sz8BryQgUB
r7UpTETJrtp4tcSROIhjuw3F35cJ5N8+LaBpGWEaHLKn4Q8zppGhM2SP2qP69Kp/
+7XHXRSqsJgRxnzXCXZ7PrskuIFVsKKFaY50dvexrV9LOQ4crnMvE93oJA+HjMku
JUNpLU/dgn/K3Wfkc6+GYgJ/RjURjxYIJ8AzVoAPZ026aA6FtVYxc599CHQE00C+
Lfv7vya8hxkrcTemd7nYflmpVDIEpK4MH1uQkYtq5ixC3CmBnyocHU0UEEVqdfUT
ZoIjD8GiiB02r/ddK1zcL1FVkRpvxx4EW9Y8I4TcoJe/nzBb30kPCi3wv/Ha2CpV
Ik18C9u5KuRowM/vl3+WEklG5tEyUniTJGTnxWV1AYUFCOXrN5QZb7zy58q49CBw
KKZp3QmXCfAjoT0EB5mqAbDDS2tYqQ4cg6uttT68+I4ysVzFiMNOl+/52hEPH4Ps
UzGxWnE4+TAI7GZmMngGx5YMJpIiiBkIIj2RN5EzWyE4WcXvMZwR+hX7Cr9cLqTq
XnaJKpbGfMAsKFJQHBWY5QH05dhZUMkQ5PcQRCIbS1tXne4IXGIiTb9h0jJ4uQ6l
L8CJhJZqKLj1rA0kyOF0bMI3+I+TUuvx89DSrvUPVG+1r92H9y4H9cmZnj3m7KKN
0dHK0Lqht1CVdjWPuWpBpBcRpSfajmPuPJjN4VDRtrI4ZeedmBxwwgM7wheozA5B
8HI97fEpBcWdpwULGqMrr8pedIHSffdu1c4i5QfAkbDLxgzHOgPUizUp0ng0oyC6
PHOTcRnH+1pXhorbfvML8kVmq5kBBE0S1o0UKlEYN80Us38z8UMDzCsTcnPaDdtT
HE99yOyw26tHsBHqjddGgg74diTQsT53N7tH0GkvstGTV4vlc4BxHTY9EBG2E4HD
jImibW30R+g1yjoQdawLzW3WVC7HyEOG4U+NcrMaJEumunslGL4DqVO3E8dr3n/l
kE4kthllWKKiaHpiV0HM4B3+VzCiCoBvlPAU4DVzVWDROfNRox8JUq0ZGDkRBSJW
B9EoyTNtDnr64AA+AKCESLtLuSYdEcs1rQHtIw3X3bIdIlC+/HrBEE6og3PU34Zf
4RZf4M3GsitbW4OM1zMgLp0BwTs5H12yQk8W3Pn/CFbs+hA8lLN0jhbR2K+xVM4n
SX9itOgWJoOrFkp0KCvJSqF7+oNd+IDKw3CbfAkrvBaz3AimGOHjhFRaeOG091gY
ZWcSHAy7uNkNkyItBuHPDv/NAP7sPyE8GnfVF0N2fsYLv2hKQyzvw32ONaEzgNI6
1GKY3qp6iPd/BwuU1uOtBuA/8ZcHCn+qz01wXZIUk0Gw9gfk9qOfGmpRN8L4Fhlg
LiNy8Tdc6uAOqfnKWfv1Vq1OPFZpEXwhjcGtKiNEIQ6+Cfz02YxtYV7VMECW7rqE
+VuGaiUCi9POYxlxeVazNmYMxYcYrpSNPqK1NsVwJlxN6i3DVP6q5SnWROobYXL4
4KLJZp3rIZiuIjuqo02Wks6zTUsAhf6ys/iFpQyRSVdZMuNbWh3ozCKYWBSieYWU
DYQMxmMWzX4nY/tSdtQ1xOQQ339IvnH3sEXKtVcvH9XF1x+yUCI8GJPeCOUbz9Lg
+cVgIgTkyS4rrzOmjGT/iG2WyZ4bSU5fIzm62SYpf5AlWSteQCtdxaMex99+pxES
SRjKe2DNE2brcdtTFFTvSWzREipjYmFm1gd+EkxYftnFkcQipCogVpyI4wtrLCVX
qEOmsVZdutDsOSGcJSNNewK+XZ8Uoo24KNuilnv2UoGvg8oO9zegkh2lDKQrUVk8
o3nL1wQ+IOHrIp5ozRz2t0VnEH5WkkWVzlEprzPqAGEkSGF+4XieO7GpdnlR/oVy
7zYyRWT2I8Y14bHs2Hiu8kCr6CG61QcFbwV9gj0fzmZ+5QFznK2GoUq8q/lUVPrv
LYXKOdTeSLT2vl7h/VqCqigAod76aVGFKjU1roZ9wXXloszqyzUInu+kxUt2vrAX
1j9FUM2Qb6Hekyx/EuezKXliNJqRDonzIYn7RMCQNhTtoruzI57zJa8xA1Uzhf4J
v8N4Xh3wkkIm/SDvpC3Lq1rt/lctr0vaS6ze7M4XkV0uzfcv+omAogQcwN+0kZde
Fx1+XrUGz862GzZGtTCPAJhdXlg7ok6CtZncV+BgXbZzPUz7HfoTH2cmJG1wYoiZ
Dveu1pv+mhJIcKN4VAclDk2Ntj+89OY7s4/Bga62PLMaTyKvpaKexp7hgKUgzIB9
7gruRhPvDqRqaTs3hdi5avEjFI5eMx24cLnBP23gvHHK00NSVECRaLe6Al04xbea
NxhAUXUE/JwWcKHErkrqb/4CD5HY7PtxCfQZLk98+6EMzUtXjXwxtiuVINwzn47K
FHy5fhNlUF8b+wPv4IaBuuv4vPqmcdPtgaQUlMXiDrTycUoqDzG7Sqc2RoSjIImD
EDHvTTifevrqgqBW8jOW+hWLCYV8xEdwd3inRzSLDPuaF1g4oeS/WkbxezbcEoGu
6oCbyVZWBLRe09nHbsCPpE2nesCCh1rr8pLJsdO83641eE6pAq4hyxjr1MDFUTG+
iA3yLvLMZUi2F7JyfDoq54jI93TRju7Zn3LsdZikfuvrfc/hrQui5QutrHlBuNCM
MmliL4V3dPsW3FZz2+ps1hq6F03oW3VtmevwlmEL222YBiyVyXSLJoWJ1OzK9bHh
eeGOxa4LUC8e4ZjDejaiRH0328Md8zCDJg+5spLubtNEZMPGuzLW4B3Op3W10b3f
v/QS5MYJ6oOxJ4U4QDbCxJsjUIeN7WfoR+RolKnDNXfEl6HT77OY7HuusDYU9U6a
TMhgbOVvKnEeMKGVfG+m+JG0cuLl4xAbUVdhVfw2aaE7XH+z2Alicy+ym6c9CIeO
k4igrq+1K6zD4uhiXSv0sK991p0O164Imr4rND7IDK0BeeBxvME72MN4ezcQkpLD
Mlqv0EfUmv7o7XnVYnhQdy0QyaNyoZZFygVWVT6elFrkHGUFlK3311CsnGwWuEOn
pp1xE4emspELlJe5WTRLJLWb+AqXEEoiWZyWoPniRiPE7WSkXCzQ+nfxw2/6ocNs
zy1duSUaAafOlpLxDmxL6v/ak/BXDZnpVophsSI6eUjD8ekT9sSwHxThgXCjCzhm
aL9gJqDV9mAgGAhm3XsTv/Z8UwXlq5i0bpqpEB2cBZNczo1ZYVy9yL4u/kKHHzZ1
e4AD2gIYE0TDGxDOSuhcHBwL/FDq9Wy0+45tPQXfEXE8WkxljXp3qJuV9jEHzMUH
DmHPf2caKBETQCu6OolXwq/DByET+ujpt9qptBoCe5kQ5SoFkh521u547IOAQQ9C
+4Pnnil8expXJQ37iwwaA/xrstyfRw4o/QWRVVbXGn57MCyosOJRy/nFeqRcAGKc
/2ujr/r+z2ScHNM0ipqbBLSPqGL3f3hjS28PX+YG14BlG477n8lLn3RgP3nEZXwy
h6DvG1qdmh+EGDf31P05a1oxt7Nr656vBmBsrRkIDpOQRa8T5uqTDi3qP7Vwhzuv
v+g4tn17CJbewUfSuRkIDixQiZ9AceLvmNYgJJAKe/NCl4TO+iv+JLSZaUyaNk+0
GJ5elfHp6aCmFFUggrwg5Dk1UDSsWAmeHV3y64qXQXLrU1R3tZUm0nyQDTUajMX0
LzZMeB5jz9DEW5+SK3s3lddcwm4EiO9LAZAjLepB+PFQ3vSRprxSg1TEPA3A0Ec1
yL3NRLla5FMVEDqCda2CnnAvNhP1Fx0pT+zG1sLt9mO+DH/k9GpGT3rCFOrVRyMZ
dvbT6Oz+Tm1kmeMBdWCgvB0YTecWXDEC9Zb2N7OAE14fnVRSC5CC3KxFqH7jsIBr
02VfQYQqqAU8//ykd96GToIcng3uLwIMfHgsWG5ic7zG8DY1dIAWPLeP2wyzxiUk
ALRGiS8XRco+kc7i29ZDCJ40DvvvnxqSTbhRe7N9Ne2xyoPhIR4nNpVEKd7kZAt0
0I9rZQDg2adBGUaJ42s0LQ+7wHZGneUt1IKQucmfFy5UTbmVpV01W7tKd0KUQ+mg
hq0qp16PRH/EndjYlCGo1mhHQfOb1HsKjo2YNQLda3PqYVZTVxIODH0qbZuSBAbV
N1ATfzkATlrbSmgQfxyzYE8TF6o3Iv9KilGhjQtBdnqQq4ppHW7ivIQTbFM0pjGg
iDa7x9cLRGgj2MtACNssbqEd+AMbH8xmy91Nc9O33lERoXRCQtA0GSR+o0zINwnO
3APvMReVVOfQQ0MtqdD9g7/92XUPwJd6Yyw1quvStEUGy1cZLcT9wxUG0n7/5uT2
RQrIPCVETlXbmsfbKU62CoZ3CJER3QJv9xR2Xrp5DYh3fchWdZb636ENGuWcuo2i
B1XZFP9ObWWxHjPgO8mBohK5t0nhdstcXWSePZmngIXwULsndbQvG9/QD+b4f1Xs
24LAfqXimDhNXtLghRVFQZjhgkQ4PVGObF2VRrjcAf/KFX4342wFHqfuQgj81sG0
gAZuHaB6WaJYjEAUgwQvOsIXzGldB8ypGv0ihlH8+JAmwu1o0JLa2YuajB72TgaD
66rb4kbop64rY+ayQrIPKmgiPeg36f58sSTI+I4ZkNQ7s0TrhUPbMe09p7Mv+3NO
zXitTmPXW+pV8kKb8RKTe7az0sIyRC73qmZ8Bmu7dLMSJ9O8FGz/OgPgG5x+yNp1
cX+ZS6nHx9vuboqfQU5QhalR8bWktUmIb+W8w2lZXMqRCXotn/wE3A0JPHcT4mBm
U7FQntnKd895ZiypFmmY1o5SZeKYWpiD8+BuEvnEQwp1WDt/kLG44PAaw4e7uExd
Wgee9Ox2AgqwqJNhcCEsRUSlxVkX3kjMqUAI4gD+DxldE3n3QDLiFs5T3W2bhbG+
gKfgGO7l4IWPk2kB5OEkBNRNfl7/l27Ec71wDSddpGMTU96sVebZmHrO6D4GhPVB
t1XUtmZNC7V2gmDV0wHP6ueIoUYT3A1hsYqNYe0DIRUFGNGT0+8Hs+9L8r5ZQcNS
a4nJv4BCQ1TT2AlxwR1FiEYAAHJucTwm682ZOkG6xicOIB/eUOmGouBWkM3HL933
3WhRQ2iCdoq+LlGnEld00pJm7JWo/OajlN5ZC71OA1dC/AJoxFxvosPevgOw+qBm
7pmpmXhblO75cQFV9hyuoiRBDL4M/F3YbD0vmb3S3nGMasqM1m4uI8NDR81H8yRd
gJBXljAV/UOLHQ39MjE+mJP3t9kxqXI4N30+zCzStGWlNvsH+MTCOSRC2mPjf74v
Txt7QL5E8UxOLVcFhzTP4J2C9cyYsdJy2jyZnVYs6Zre12IfOU3jaPnD4EPuOEiT
tMot+wXZyt9ZiFcnsoiNJCqk00o+Lt1BXORuR73L5peLaj1TXirdn3x0WAaWKxf4
WWqXAh0WlFH3Myg14EV+aHJYa4kVqc53GRA7z75nPurChOJFpwX/sm6pfuNYXWqs
JfP29Y1tGC1epmIQ5+3d7V3ovmja0n81NnlUjOARM48QOgZ4SJOeKxa1sJrk6Pus
TY38ZZhhY9tdd9RhVKF99KedE5R/GvcauA2qD4FAUU323Tfp4Y6lLWyy7C3fMWRE
Am2+bVlVrzzKn32iPUjecQOHOF+/0UN8NQmOwUcUJ/dz17IfPdjG+eI4tlTs1e+P
NBDlTFJSBLiENnw6UoIOdWfzrP6+OYhYfbfrHTq5a3qjxsfXC1Yc9OImDKyIUS2H
4s1R03kipe06PGxmR5DC7G94jhPOzLb1JkLp60sYJ36rtEiyrcCQt7E1zN14/hmd
gEjYISBxK4TsixOEePdMiOjwPavNVMMsmFStfysIM1ydZFshM/zdL02iD1HU5NxD
cyk+xSsyviVT5oKlRzYFezmLUAOlKFBxQyt8ArzUrIGZTlxN4pcgNOtVjCAWeXIh
1k9c12p8bS4x673AhWeLBhIwS+BkaPQYQDfk7qz8Y+cZ1keiep0BBMjS98BYcva1
O46CHkthiwK2/QVzUgsUJ7J5FbLV5LQTNntdwN2JumyMNdpyWSBpcADS/i5b8ufn
zvWhtWUlJrBoAzwICLrKJzlwLIBBEv++hHIao925BnyYt/ssRfJbseR7e884lhoz
k4OehZBba+R+UH19wNX0Z1i0SIltuPEIb5Acj79LyHJGBKiwW97DMc+KbTguwR79
cCuB1YH1eTFJP6NpZPx3XMHQkUPBHaYjcID/AenQjlxLEertdxrfiOuYr10CgUgd
fmSLrfG88XnVb3PEB+J4wNcQd0Ic5Ac++kVDVnRWfo1pAWb1H/CCMDbHpjYcyyz4
t5IPlrt6CWhSbhO+JTTJ6joF+CX0CTSKx1u4/WlOu82PiVaqTPvDuOJLcD1Zm3xE
K5VdsJe1DdRrnMKsxbZRUJbUxjZtZhtO9nQ7v1cBl7/LPdtvnagT2QCi0abn8U/M
CuNGmYmNc+LpyWboWz7prIxu6t1aZeNP8dMQSM+HYmLXUT5D0Id3Klt35Wpmzy8w
gJ93mcyhSrpsmjIlwCOLChSZIR5cALwIWSZ//MLSHDtGBu7M+O5Ow3gWqWT4Ybmx
2kBKHIZ4L+AINXEy8aMowOeJ7kdy+jOsUxOUP6UsJqpmW3NYOdVcwCMOdYspMBig
TkeZJV5Kl7uGp8w5WF4gr6Mlvzabw2SShHMM2R37o+OiiAG9bRxpVh0Ey7UX8wt+
y6Z9P1r5kq1V/pVZbjaVH+6eTmshgdmW2zrYmKDGx7aQu2oqIM/x2Srb3az88At9
qYusp2LvRLnD8ArhyWZihNvJZxTa3ZLun3ReVxgoygwKY6KuxkbIkJ/GBYcTbeae
gAePSsrXCwjPyLWeZW6j7mqJOCp1A/mSgKIo/uCgVMeFlKCS0OmD80K5iCa6ZYFH
ZIURW2hwUItAdoPu/zaLT1DoenYpr5iEBWgaarQIPcfrFlpU50Vah/8yLyDmGBaU
q/hZuKL+8Eexqnh8dzTRNyzci1K6qr4laeNEulFI6bd4N9UkIUvg8yFSN3sxQFkh
xZOXcF+8VXAFju7NApWpbgMr6Db8cy7tyOr/Z+1NsyOHnytVtrjeHVAkmBlbSLjy
spAZcnArTQKyxtyqO6oFdg33eqZMBKeXQ2wgE2HR3dDBuEQaA/0YwWzBVDdmZ8wH
Zo+R4vjO4G1QmPc3w7tNoGZXroUkU/XMNt3SlgvlGygCtwhQ09sTmy/WK3q+1Yrt
YeRmMctky+zZaIu+Sf55NM4giSYjGSteG1A63lnzbYQAiw8g2xsBor6VmKRYzFgQ
kKRAXhuK9NYFi84aU1O+qXoSaaco1zLEWOy0T2MsmwcQupqmKfmiRjG3EP4ias84
55HUC9VST6FRz0AVpq1HeEpVILZaMmEobEtmjHRbZMNF8pcdhfTkICzH3X4yde4x
ILhUXNnq4lEYJ1a1yASnsaO9Sr5w/5MptKL46VoHKEsJo78y5VXYWnn2Dh+1oT5W
5E45emo8Sk0tzMl6yqBUUo5D911SX3gTeuAwI4EMDnuCIdWl6aQdiWpPY15jUXEg
rh40rFblmk09j3bWZJ1JVaqiwtrVfnjuA7w9iszI0Rk/k5aHgCTjMYLeivimotwO
N3Hf8f3VrLGt0HjGmljRCOrd7YQXayN9s3+lrMOHdq5UfajOVA+L5NWRp4jL6+hj
Rv7YnNyTaA5Q2rYWkOPWCFohHWgELEt+UrPGZa1tfr5Np57ZVoGeqjNiQ14IEjiH
gYRS7XdjPiyu0m7FkVcugRNLFEUfk8/QePINytLHhO+yM+aN/dY1rtgU+rATZIos
nBbfXOLJYLNmvp1RJNj0sgLbTSLEeZq+Pmu0sIi35UoRL5Hujg3FvHBnv5dNQ6Fw
wh8KWjaYoQ2n7xboLdsjRp7DPQM1LspIgGKTM4lXuM3FAV2j2c4iGboVHxFtD1bw
eu+E0MfZ6VekMBR5EYeaeqRfdfppcpGZ3ej5s2G9XNeEEn5cePpYkxcPhTLXYrUY
B9k9wJGBddBgMA7RvqPnNNE+I+V0fU19CC8y9QsKVBGZ6nJKRV6udjNzSDBeOyAw
2ZCXtd2pSaxd+Z+ZN0saWwh0HZkZfhJCAaDW3hl8+boDVAS08zKvm2TYmlqpZydd
wt/nvlL1COXdFJ5lH8u9hjUGMpYHBtOMGRTu6d1hiNycxrTCh5RqNj8zJzXUeHTU
Plcc0A4X2+LTWCLSFALPf2NoeuWeTFELOK3U7N+o9pkMa0DYSVQ5B51Rflq4pvJg
OMHMTnoDkbt0t0hdFDYy8IpB6SQDjQNXbIXiKGta/JTpJAO6sq4okr35p4NWvDdg
6CHyhoS3U2vx/LsKt4FTE6ovAWYg/W15BfpR6ackwkoGsAfn0EJwe0KmYXrZGgbW
aiSPZlfEvV/CTczsmp3xXDud1KpgBasBI8I5dGNT5aRPqelS08O+ajjHrId3ou8l
2EmKLcCWQKsPlPjFAfcLxcj95LpYIycPbjaIa1WIDQN+5m2Bgyw2fDIIMRQwv+Cn
QJ8fisyn7h+bNIQZXKA4Q/BgeMbGlelovkkQxQFQ1ggJbvUNeiRY3rgJZXGxdVOU
hlo6SdsSw3Qz58zAbVRJdqM24Ytyovv9mS2aPATOMq/Cz+p1MeLRve4hxOQfTeNu
OPjUJAAK/aDVkMt25dcdNhQrLnQWSdvSkh8IWsLsmo2mjDECNbhcAyo2YFPyd4xg
xWJSYbmu2pQ7pOKyRFAAA83gPAytK/gxVRo0ASjLnax8vzAoC/Y+LlmXtAb10VF4
ZQK6uqbgfI0HsiUp34KC6beujQkcOX/v6Mb43ppfiDzALADa9X7vSjsacbbEuVbg
K63woEqUM6zEVmENisTocQ9BxxTfP1qdztCpx1dLY5f4BeH/uD9KlAxfK/vU6clI
EX6DqWwoMWlary4ifhJ0g3X8PeoRP32QDLUGZhsYRuFp+S8zlTCv6fblp/ImVTin
WlZV8jnerwg8SuLjh8IkBAGvpuV+bc0DjjwnJHaTfSRrQh4cWEGnS+m+hYkRYOnv
BD/WEDinqdhfvU/PW//52aH5S4xBzKAtjkkO25GicLXhukjvD7lF86WR7Nane0Y4
gTJIMPhDycJktItHiOnrpvQBtf7bCCVouJphgctGkuOs5RmG9mEqNOBlywObapbb
okmj/aHJriIyZTE927JkyKWadM8EpMV5OisjDSoT3pF+jxzNQ8h3ie4k6R1lbe7d
SD1H0VsFJga7tj0gTJoukusFdZBNYTc6zBI1zfxucffGrJgcQMvLV9rT9WJdrS/x
nVQ8HhiHRBoV3Iak6EPrTA0Rqx6HIlPI5wC6/UlP9XYRk4SyfINxwKRCbEAFxVCf
gZk2UQ8jhlJqCvFzQJHMPqHBn8ptxEHEwT5lphOtXOWLO7lxEuhL/zmmPWesJJ8h
Vvu9XIYHeeVhJ361tJ1jzIdSi43aZxVCvngw7MqHuvrPkNzDdm4HS0Iypiln8oZ6
P5Wn0uSw2JTsll1CEWR2eQIfGywsfub3QQXjfelRil5zT65QmLUJYOeacFQxyyes
9SBRJAqx4pPbElAZr+zht5yu0or+j4sB3kR5EUyPcSf7wdqv7tPDTaxq2FXdQr23
hajNwIxoB32hm6pN/Ht5r1zEHFfvRfE1PlE0Yujq0sf5YMr6zvB21roiOjYbOxpY
hZP4OlJ+PKkES0mo3ghpT43PqMmSdrAZhqClt/CYHf7IGKOej8aX44JatMbigAoh
daByPEXWDbVnGd44ruopIg3TD+zyJF7YGatrKfbMmSNXqmxP1kzqmnxlIgaT31GW
8rE4B+bmfzoJbHD7QOUe0WvEtsq6qrwusxYq1EAoGjDxeS7P3FADUcnOpeci1DT5
AYEJb+CSVeIWnaR3Gb5/3fESKsnOZIh16X1iTesr/DocwSe/65VMYSFYNQQ22dJn
fDPzM/EnppCADFd6rcygc125XGuyRH52nEaJB3cq6htbh0MKNgYBgFuqqH46XzUG
XmPy4lNPUmlxsN1lbtJENTDNoJOLIoM0JhmhrgtL/yUKtJyW1rzEFCAOyE7AsfTJ
smCt3WLFutQQOZdDV+Bn34/wEIrLwXdgknJosmONpCcIna7yGrGWppWOptjz/PAU
G0MrIm6MmzNJ9OpYkaPFFPhSPv3VbOrnkDc+p3JNeWbi44D8B/f6001Lj+CquoUV
1EDN7z14U07ev8LvevS5fGotfdkbDjhng3Fw0SHuxPOthG0WbhBstZpdC/9Pi5mi
tVHOAtQbn5KFUAIUVDCsKzeqtoPJmZDcX27N+mxsj7aE2LTHKRgCZDP0NyR4iyZw
Ndxwx2SLTuu85iP6DDGe+C6LYzOMKAdKJJy6bCZc2BqF9Y7BF4EiRfLbvgJOr5We
yrirjhsH3xgDOANzWUp+8oEDrjDRQ5H4p4cXUWx2TfQGUIOZ1JQly8mKb9/Nzz2s
9IMf8Nt64O3XFgmSJYy+e8Yk+yyvjgVx0WCWsuloevni7w0JbToKZX9BURNi9JuM
xYcvFCvc+C5KHhqb/A1PZBxtDs0KyFg8a4pUUyfiO1SJNoNzLW/SSh69ho5OkHIv
clS1UgCyUMMD9jv1brqGBlrmwmHFCvmVVAJzbaAQ2FsJ+pDfdURE46U/V0PnRWVS
4EudI6SGJ6bLlEHswEhZNEnEDZgHgECfaweTKJ6HkL30fdY6S6x14mmikEHLOBqq
h5BLCegGvrO8drh1L92BjxGTFvN90ErsW9qUpLrLm7dwM4x9g1veOMYLzxOIqOtr
tkiCaSlXUzD57B8D6KU21hlBX4iN+CTUI5MoygveORs/r0z1LT5+w05EfY+xOnGG
Y8HMnAQd0ns8UF7gs9UeqctTEuAkyVSURVM295C0HcCVIQdWCbYCEnx9KPsqLMDN
wa55mXYLS+gg7i99mb2iRxPTy/t3Y/Gkpb2BYd2vMlX7Z4v0Zjfb1yQnaJwTqJSy
OYT0TOANqR59GISimqM8osAQAATNmg+YaCaVR1cC6qCV9QSiRtrSbMj1xtRdj2h6
UTZlX39nETfa1TKcxxUqhNabkZ2Wbho00xDvWsukmkLfPtQMX9vWQNiQOBWNYgmj
Ug5t51Zcd65eMnKo39zo8b0bpeRRO9xiSy7ANoWVvTiLzeJcxPf4dxzbLk7ow1/z
H/2Jr5ISMG7sgW29yF7AD39u5D45XVihNhtlVAUjY64WIaH5hkTnOaM+ufG2EjEG
96qzyYcRKtznl+9CcTmQtJc/6Gljxtj8hlOSsXk96ZAvWUu1IosPA5CkoyQGoKqe
3FKHwf1ga0bue3DodoyuYq58fa7iDIuyfiYoNhwkVehAI5q/0yOCZi/GRKJ9pQIh
gUwQuRYz8VlN9E8XA465osH7lEUZUdIXR9d2OJGWjvRC8rVQjYUUSzFtMnmmWslo
v9KdhkKLtyTFHUDS+0/GDmQl/wB3cPLfTaYSVuhMBLS/siUZVO4geac3nFrEPXcB
YeF0NN4Vp9VoOYb2CIc2ivp0kxBqk3yCjpThPaaYRq0Vuy3pfGGe4PiZdVEZsK85
koC8RroSE+DB0Rd3qv4XUTs9W41+/f1xGsizkJNYrQw9ZG2Pvs4SpzmKvZdcEO6l
uGgES/kQ5VWCvfkWdt28V9RgbYEe/xspYOYDeGfa5FLULR8Uz4w8w99X9Ah70Who
uLsvTaA7KdoExUdXeWrR/55mqXa3DxSksqGgLWFyzixa6VaAMVn0iTP6gWsdz3g8
UzmFmLepQ7eazlPURuSH7CViUFFBTza8d70Y1kTrLNqFA3gGguNBgxHRY6duzeT9
DA29iohsdicqiFeq8GUss6fdwJIJCv2L77FxqDHzX/e8Q5Xc68nNudsa7YgeeSxJ
NpuqeCitxn8UY3o3qYLqo8Dj+TVY9GUhVqLIQc4ogYdUtLGaZuW3VSx7M0Urf6j8
bta+UPq+tbRILVtLDuPHInLr/mVPoEpMwisiGKdtb/H7ltLCOuFn3LTXP30pmNfR
DJsDYV0wdI8gEEahCItrUSZxdDIp7OQrRA0gMaXXVQUyd0mdDRibtY3RlpvRPNG5
/lXxj6GzzkK/U9tzRO8SXCsJgqbHTTR6YDriOOPpP1veRcRpSP/XQsgM98EOqV8k
uR0+ZFVsJUx8lznVN9LBBRH4vjAApg7qNvJCJ+qNQPxuujt5Dxn8mG2iJkD0MSzy
jQAEQ5hWg1i0tAT2QKEiMwxkkuTh6OioWS/8xYoYEhjTbdpA6hBGFW794oEB+Ry4
I1fTE9EGMvYUPaMpi8+fTZBnLXds3N1SMrSwKYF8/zjbon6XfxEgxf7mo5xSQjiU
4xBtujuZUsugAsOXeRAHZVO8evhF+K4xIyYzx4quz/PsuON/xsEM0Fkgv2fxVm17
SlaF66gFK+6Mi2VKL+FmldJivX/lC4/c2SzT/kVw1n5mFbCUuK+f0BT76pWAZEVT
/Q7dRD4D73yN6BI1+H8bk7B5hcKBVSFwygfDu6zYJKJVuODiLFjaN4oW6ca7QKfK
RNw06M/TvmAagx+EbtOFXQLBEJHfpWzxi4RNZS6fGjHBccu2Z3HyUp00MzZN0o3W
BUKBqTsfkeQgi0vQ0HV9EWnpULVeRYeP2yqsUZNJlKI9Ci9gAeVlKW8K56jyzGCl
xn1vhGKXj0NtyBnDEDptfxiSLT+R83OEeKobemYwWTupF7O+vAJzpnR8eIEPUnAN
GU5WLqW8ghuAcBELyXSDZ6igUXz85WBUzlpoCXEfIcfluv4mQctJNNB2eA7GbmeS
9J2/yCLitUVDxtimqCKU89vRAPKGJgurOkov51iiXoihEAOYL791TMXvtABQXfkJ
Ii6Hs/BwqpC7oE5v1KwDzSX4mZw3ZZzRVL5YDiWGavQI40SaYFu1NG5rclU4wPNj
TKIH6hLQENiGFylozRD8f0H61dROTq1vEtlB/O6Ydr2HFkyvPMKl35RmRu9KLZ3z
zUqOyZSyISjuDO4VVXKAlQk2zJHBKZx+4MInZD9fJ4zZ86IdQdGjrVo100weeFVu
HFF3V0pFNFBOuj0VFWmWU3N2xhNaVlJO7SSENEVgH5naclp+z737X3nbw5Bf7yBa
1cn/9qx0LxchjBWP5kSHL+qMq2qc8Cm56cIdF+uol8UT2yNdPgXz410ntaHT/gES
Euw8d6t4zahAVdR+dVigUSIICX7v28x/ZRyaCkxIWOnzybpZN6xII8Fjksz5ramR
V6Ah/gnwv5ZiL4y06KAKlXpfr7oufMYWJMpSfr52p2h3hi0YMC1U5VV6jiT8WtO2
bgkmLtmxmpKVhyvXd/lKOvdgav92STlTycjGnGpWnbOcwR5vCIB6hcJNO/41ddTB
dZQCk+ibB456boLmbc1sybhHW42cSBSPMasq9tzJssCJGkefSkDqRVTTrwUvQ5rZ
IMGtiAwOr3a9TcIiSg3vMIsH5BRn7fwwHVpSLI92pvTB3/ZwuQhHBr33ECnlKbCa
7pszjOUvrPR4pDINiTAjvu9Sf02UL5PZmzhe5CPq94K1XsbkmDMFEb/DiMjDIt2j
H+1d8xnJYlDVRhIddYysW5isOa9OS+eQFXQCcZtyPMUAtILTuhTzelxCnsHidpcW
ZBnCqz55p1Hwb9g066V4VSCHL3e2Vi0IhrQ5L3SusSGl/IdYlprBfbDor7c+qYkI
Z+Y5OsmfiuonQfkiwdVTVtaMkeZGaYKdK+HyT52Vrira6TMW1bj0cOvfs+GIomfD
RU3V7NBm3m74Tb1TQ5wdp3V2s0wVpptpmbMNGUnZu4hYH6nytGY+CUoVxsWRjjii
G+ECTsHKFNjX2zpy+JUA95VTPk/juZyrxAC2rYGEpvriaN6BiKEKFj80AuveC26e
ytIk4QTfOoaEN5SBTqvWfT4VkhJy0kkweFWeg2s7v+QnyZp0VEJfWmYzSFzfetwH
toqeskYWqavrQpAEIDMRF6HZbsO9O4nIDzjVzhRsEY0Vjc27d0M8iebN+F5M8P/t
Fg5ZjffjtnxrWQdrgVAd8H8QaYnBrzclkUmBjBCeUJFqUi/C3S9RYuFZqw+tOdtF
KSB2CTaWiuJFAdZdDIxkZ61AnGi5R5TC29VsWWWoAfFqVXctB68wRmUl8GOUEYbk
pTKGSHoFyd48MUmJ4yyGVbXQtcmiL+6ayWKbNLROEfV8dEk+nmvdwRLOORiKLWBa
SOPIks1vvY3Rq4ePPTxZWcQ9Ob8eyvWcfqqCdzAk9NCA2LDczIGWUYeNiEpURyun
dmUHDjGnj91TfeZpiitnpfy65suWDu9vvEBXY9pUn0mmq0KPN1vLabpEhV6h7o3N
rUhjg4hiXNbiYZPlZAs/XSLO7wM9xBwbloStuLaJ0hI44ieD3phnFXUQJaRT6RSJ
Ae2RUe17oSySJOA8ea3332TX178tJmhF5GzxORka8QvB30v0S9C5Puh8DYQxZRbV
B2GfkericqNRJWzNqcW5TsUf7XbsdaOh3P7jBliNJqachwnKOeGsOkc69HyfWl8b
QGRxjTNxfGT2WCJ30t+GsapWi+QlzHoA/xMjEIpWNSkeS+XGIWj91b/OQzbGybJk
560MPzUpmAZ0BqXWL+a0wpmjNw5oLV3cCKcqX6BUOvP2uxKO17yOZW9r7w06O5nb
E2KXAniLeChlwG2Hu1LmfELjUg5i/PLKHKC807ubGb8t/WTrqEOlyvU2ZCa71Db2
DMjqIjG08Smu2mGU+DI5WlXuRKFU2wp6GJE4yweixH7fTkbIWj1UzHjkismxeIpt
mORQ7ZW2Y8Jtd7sFKhsGfjKYPujFqpFruoqgpKaMIVol+5bqYFQr0IJPwxLBrEmT
eq28MYcKkQaCZR544Svbl4LzONhlUG62Lem4c9R8MDwdmhIC5FQaJ17WJFZoSLH/
JXHJOyhS1ySH3rzWiuKG0MyzGn1L5qDDBN0a8tmaX2GxEVCt4uAG7CVWKnuK3tfg
bKRiHaVcQm+ly0LId9FyVXdmcWZysasci2ho9CF0R1NVivN0p0uVJHQzm2UhrR8C
1fftNz2I7Wdae/E4r/cCFKIkvyN8NxLdFLEkEAAVsZEmR9DJkPSUydLWCJi/yn0J
6MYteXr3UwCHIlqqunO2cEr0xRv8I0j3yvsKRya31m2aj3Mecu3VuWssNVXYFcJH
U3TBcUrAfmT5D2JJug/q5fk+qh5H/qBcntKiS/5xv/tOeEMgT9Dh0YB/N2N0mgNU
OC2YS0a//Y2cBXBSbPHW0BoVLEgVGYfNIpGrzfo+OuT9bG1O8QcWPJOFsnI0Mayw
raiUgHBqJ4/G50r72ntBEuQXZJ+0Jzf0V4FJ2uhN25PyKkp1rNwJ8A7zspS9QEev
eukdfssG3W2eMQiHTu+wfb/YqUA37fkVZbYEv4tOR+86YvphxtyNgkzhcRCFZNwt
uSgejJ8ILQBLgKTaSW5hikxuTt2rnTuVcy+e4/M8x+T8uOe6oiNv28AaU3cg1CuV
ehk5uKMdNNrHtl/EXycFqNlpmwilvhCfIclWOq6iNsmY/+rtjW0o0Lg/6g27Jf7w
/tRc6zqbJLXTxRphTtlkquGm9zk0dzK6F0gychdRbAsv7juKh8Pj7xTckgCcU44D
rJqWC599RF8NIDI0HijCc/+wjoXq6+jzRLuluYiP1pEustbSyZvFHFdb9zchVHmd
KGwaB8VV9dsY46uFvlB/FjsQ8WDl9SjFB/C8bhZVyF4aMb3lLODH/1kXVcoKFkXH
ej2EkRXwu79+siVx5uYRSYSOZNAUlqe1GrXMNDvSqYTJsRtjff1DZoJfGwFZNjqh
+RuJpHNNmTSbpLrY/Y4nI/fo9JBkeKaw5vv9qq+x9Fpfv/9Us7run0QqpdKJ4njh
7QpALS/9a/KLFNg9mi8JjdRuvWboZU0/TlKO6Xe7fATHy3Bja5q1bjeaCbZjuOAF
/o3gEG5KLt/BRsf2EXIbQ51/D+0pTDflWWHzJ14mGXRDUSqFpiBxyjALfKEAV9YK
PP+qg8/azTejpaNNb4VhARAAxRxCm9PSFT30cajbNcV98XZpiWpxu3RzwqJHttRJ
0YGYveO37ew+IlurwfZcEVb2u2rdx1nTH/f+EmHuk0wL87kGpneOxlihlCMXj0jU
T9BHRn0xKd2Rzebc5iG2/CpXs28adJQ1TCyovDLoBFhC+jfbtCXk6uETEcMDe8vN
Tg/MkRnISiWj2pXLXwaz+xPPIRqdEnEJa+alh5BegfzKJ1xs00dO5Kb0FRuNHfyF
CnvGKcpe5uYRxBbISIkYX745QJ8f/VZekovM0my45OFSUL8xdffqo7yX5QsPfOot
5ne45RwxsZz/l+Jfgh6Ksgcf2DqL8wqKZCVe8GV1EqehYovdq+mettB6HgoTlUgD
7P1wUf5YvTBNY36ss7TV1kVdBBIe1zKGSjIDDwG+j9lNAkN50Z9h5fK3NLx7J/MO
RpBKhz3CXsfLCHmqm8N+q6A7yrYYysDutxvBT4MYJRyJu/sMxrvEzAxu2CjDGZ1m
kh18bJnlP741wXB+bq8vRnmkHZKqoHEWH5nFhZNYiwJCcmHw1Yh65muBp4OxF3BV
2KpHrkf5FLpoaGJbaL8d0h9lalSw21NaJU22/aRUeQzGj/YzYDbMVeKXR61oMBqP
6xei0ijc2rqHsS59ONoLCO5jihuXZ51a7rBqMnGEzn4KFdN8Lk1Cpw1dWqQ4T3zn
08oW16gM5L+Tq5Km808FirHVTaDF0fMvOzAfi/KV/RsRz2KI/ht0d/tiV59hI7Jh
9e4MoieEchhR4oazpg0iHm3Rs3rL1vIT4Ba0lkjy9N+Qptt1AIWlL+t/cJjrVpZy
3jXnXt5b4QjUHwh+Gfo+R6McyD+RYH0LnBxnr7bdyePHcG3G7ttZHCtJr8urJKDO
zgb1acsD9I50L7YdIZKJOcGBVjBrrwhGuCYB/0V7Nwfmv8LE26GtxI2Jv8xPL4xY
pjYjX61u2wwgxYXxjN61zsNIk9LCYRtkXnPuIPh2ag6jHOIVwPMIWg7gulAazrlQ
nsbrK6/LSEB0f4Npry0a/+0ZSnK3Iye3fAApXBVsqjSHVl9lcS3wrsOafEYgGy1O
1wDjA+dJOaK7rnwTBStYsJM6W9H0OO87fqfu5tjIyMr9mBHtwo7Q0SMvk7Qf8SXZ
PlpqE53yiHBuxn4PkQn8ar274wqTln8+98f75PLEIXVJOpzyiXM10FyshGS/1aU1
bko4ZtFzuJ65201dDgUCE5u6Z65TXyh2rnXw5kyPORb54aAbY7YxzkeSkRVEsq0f
/njyxmQOnjn5pgOUTfo0CTWD7t5j6Kcm3MygeCkCE5sbG7F20N9BG6uZQT5zZ/6Z
gFp0MDKlb4WKE33R3NV0TTsBbv7NZEMzTiDUMcpJCuZQLcuFlUVdXDiHFsTGPNhP
m/d2dXQcsRrR1P0iy35IBVHP1y4+uQjPHekbH21FmsCFIM29NuxYSg/DUMrbPNbL
XqcQXkOPyvkQuTog8if8NK74AlQguMryTD0GxF9M0BccFOO0i9H1neOGQgAgusLm
Rf/S5D6qEFayeaGXrh+TYbD9do4RyTBSEB9CVX0S1yxaBjqgbPN5diIwM7H2V1zD
TSzMLCHB5lPHKCl9O5ssxDiLSaT/3ee/VxpaHkaMiCgcXLD9oBE5BAEZ9YMxabB3
1P+Yn6bWjDIlsr7lMLEfpKODrko4NpH5xcsXz2fU6U3ONk8zkl2Mkmk1JFVb0HVd
6kVHMiJQc1GWjsGdnr51SooWkwGt/OZbG/L98d2CQP379LiQ0nDv6kUXk4etO1Nr
Mg/EDpkveqkTUexltDr0HQ2AzlFvJURQ1XrZ0EkPqALqu38UJyYOa3J821d2GupS
uHezdKADIWNLOHgDBXFZpsaVpEeasvZ7Zk+4/4/CgDvCjOLybf7HGyaxH0693mTE
cJfQ8+rJXxatL9A9vQiyuWqnyr2CK4yRRkAJQOyjLUABOaieHST034et7yb86UT2
mZEQT/MHvFlLHZQaPlDicjF03aLhMa/yfXjaVhpdLBat+xLVJOmPwglUtMXpeAQS
vczA53GFcMaHCGSR4zL9++ZMKy2DplCoWLzvodLml7cHkfvwbnz5xS8hQIsg62mz
mDUDrnQW51HJSDU9h03BZqQkmwdviIeQf5H/Dh9nUghrve9NRCszpoDbpsov3hQh
ixdAFwMfjRWHO4D8KeeYCRwczF2E/uE4jMgX3MrpOgrEGzoOFqblfR/8QnqFcxj5
ulsTgUt6UcoBfk9Tr0rFRlxSZnFpYnQ4KvaEvz8tLUNCXpSLCgmOgpP4DfYr5m6a
+d/1a+Jzo6pFMHTbZoOzsUwNpz+Ws53mcX9XZSxSWwKxFC+wMNNNHfvjM1a2ohmJ
Z0/taYt8+/JvUJWbRpfRoHJTfIC/3OrQyWGyIzMnLcflFiwZDQ+6QHy7bxigASP0
nYPsemn3UdQGxWW7qW3wNp/EzxI5//I7RcwkisDqK4Sr+tzHx5z5pQ1JIMext5np
pMIhP+hXJrvZT7P9eWgLF8lVJ1MDbQTAuM7CmMEFHNtY6MoDuPMKu1F5N0XBvuY9
Olhg37KJiKYPv2DC37j7oymhmssLS4Rxciu8oKY+zil2ovxMMzayixJ/mpCXCHB3
pM2orFz93nAg34WPZiN2zZwMHU38SmN/brC/4vPg4WxMZa+h9zZzm90OlEnn0lON
V8nHKVD3p8IJ9BxwfyWF3qgmLh7dn25WdxxUhSNIUiuKBmEpiT1sL8vuV/Nt85FL
HvM8TzxmRLQoKvjIpCpO0o6AUeV1j6fQQ1XrAt7IJshCrLB0h80zwmGCWXc2VxGB
gH2Y3tbczqA02oBfkrvZAbOE2GVxf5WJsXLibWBoWjSzW+HmwU/KLWpTHumvt19z
jCSPlAh2Ol6X33Z6ePCpOufVo6fahnwAk+hSWU372vTJrLgzfb+XEM9Ye1yHZj4O
tJ4XWKTRjfmDNkjfj0+UncUfFhBFeoAOuAKe6PzveCrXkXgPxF9iC+bouoMHlU/Z
1Ikg6FhR/e9Fq1fdsnkwAvq8Tcy0dsaqlFC2pLO8LcfxZmUv25bEef0JTECnzWqK
fuyVi1zoxHHV8yN5AkZt+fUwECTeI48xVH/zVZV3hRWltkdlPmPeDDsyczyV6+QP
SN3EGo1PgHohQCmAJ71/FT1q2URZfejpgZNb2jCKpxZpL2GD9/1Fe27pAMxx91E1
i0Glxoq/dHfxCMwvAM6cWfo79iQpVkBnguqY2SeJwK2Ju0+YCNp6N0Kaak1Zk4Ul
OqIsoVhS6Z94HtI+JDOHe5FFZ+UZWinAVeidiGdDRwMfi3NbW4TXQfizdFeLpKRz
4OQg2om9vieqYQyKMp6d5QIiwVz5XWByBYlVMPIOKXkNRBhQHEzAFB627g14nP7s
wk9RHXQ529b4coOeMd7kuP2jN+OlFZH9D+dOw9HcXsTfvvAXeK3jLzQGXHFOOsOK
6UBagUTQB5/rPmpQePuavKlDbY3K6lprFiZwJH3+kNFTJD8e8JIORWKw0iOwtTUe
meKAycuieRW0WG0Fa2WQxPuSS8SITPnexS3Ck+8y70GclCqztKeA+Msep/x0GS9r
lLaJkj1OoFHD/hDcCLKD795COXixdubLDfqPg53U4WwSkNni4UFVQfbMrmZ5NNYw
ogDBV8BPehMVdOB/X+HWg5i7pPYpDb5lX7DT9bEaP7W7UE6vo7/CwaZDrRVarPNE
/jEfWF094TiDF9CFFlrIijEDedK2wJ2cmGFH7Cs5UcqSeOAjzLYNhM2PuPhNiMqt
LCjGmkIDwmMoBdZGBZXCYhLU+eXsDtX55PkTo0Xts+ATEyCtaPgLOOCT4rKgDRTw
JjeUiKUlC+7V1zAJ712CYgf5zc1etB/gQKT0+mX2OXl5vo2HuD7x/KZKNpAfVwC8
2RukPXKs7jXKyKJC20PRRBD1FhAS0jQuGsE11ceGyxN4phHQnwo34DFhVLAQyYlC
Vg3ee5rNnt425X84xf78qSaYMamcCHmihj7tHfYCowuixwVdyqxuga7PfB8RIvjD
vJprMtrJDC4H4mLqm0agzTau+qO9m4vEifKMF3Q19obt2Dq8Uwzs1ieQEVAytqMd
Yw7d0mwK56coM062dBQ+F+F9Bw/KA2Fo++n3dRbKl24pXe3w3u25dvwf9OBS1G/F
pAq5lOq6P1rQuWi7eBmm3Vr75L8ehjiY3Nr6E2jZo1rDRrX2ZIJJVCqwrBIAO1Jo
ujZpZd6DqnvrpcTcS/ePCUY8XdhUuHNBRFKpSZ1221KPggOCnG5zCY98dcmET5ln
IXZxGoJVojoaGr9z17TbIEb9jWD9zqkt29TzQxxrwH1oPSW3PXdpQ2DCbzZ/F64i
ijeVbtxbzhDt7ICAqp/m9xS9ZbEaCKoOJozG7G8vdpZzFu9WvvO68EtyAvH4hJG3
04dc+XLTCwczjyUUKue5YD+RqhXBQQwEkXqKei6h67r+OGM5RZdah9+PYAo8nmFf
ZwpiQNQC/3uzAq7GvHwOSX3KvRmc8SIg8BPtdmzIJ13qGk4IFt1TkgIK3mXO79IO
ZoEzZ8wGu9/ZKaK97kfAkLezZDgwwBu6dLH02XmT4Th6duS9eHXOQuozOkDTOdqe
W9o+IZLptu5YmKimUE+gQrvJhHj2svCw6gONTsofBYwt060OF/A+Epgh8Vw9gwJg
xWLZ/9cUFKr7eQo1yS1PRUvXvAh0NEiOnj2kqfNefUHqgAig9o9rTVXQm/tYm4wk
a5NmqJ9pqhvA2dOorane/8TW4hbHQpz6WncOdAYJheSUc/EgkSN2i8DTubfJcJfJ
sqHbgbOUqrreL0q40xDAZkwt9A7Ai+TvSkzmjCJlByZwxwIKQVhmV0TLqnRu7AV/
ksvWYDVRO90NNNM4vb+8PhoYNoVXY33nJESRtWvcNLR9JLj88PmxoniYu8lA7enK
hp8yyKLxS37nGukf8bSY9W7POV9Rqwg5lRRS+hk81Q/YbmT2YauABxyy1pPQRB6A
rt8ANGo36TXIqvV/qeUdfwKbUqRHdNlZWGhHnChueBFT+YsUZS1QWxNQvYffrycZ
lO7fJl6IFe1/LTolgskhqhqr+bEH5lEYjyR7Mdkv2n3VVzbr38jqX+f/4j5Cet41
Agzl/VwtULSmsYtJzgF/fyc1DXGaPF0BR7TeGdiWktsMOWlzFeODUTpuAJgabS81
8jhv1RlgKoFixiHeBHnMz0YT3ggddvTxIw0LdIuHPrDq4ld2/tl3VfTHVFYYnJs8
NdjMu630eW9300wmjU6kyaPk/aec88HKSpIlc4TX9RbPiv+OO77QZLhujwI4q78x
zZemoysD22yoyIHN+wvnt2uEsDRNFplr4FFlNANDKbAvmgFUIIZZW/2KNYTT9z04
ikNyQAFC6JNsgez3watlA/aLFm+ZOZTLyCDBhsy75d83ZQ/lHccb0C/4FaynzIQ1
gRQCxqiRlcXE1kAMLew2XE5IalSIz0RWcxOk9xwW5FWBwTMtpNLE0LkeCu2KQ0g4
zefL+LMZob6in4iRNCApooVNckwK9zBid5Wsra5OZeU9JMd229NwZylcMrozWIwW
bGDGO/mYEzl6NySZqgxPo8F8g7hvztk/ScOEG4sfZNu5Hd9c4tEKpLR3GdUbuGbC
s341uclJ6aurR8xGQh6tvJTE48zfb7QLUM2GVNklUNLDuozW13jbgpoO6B5uMxbp
mZqjQJb9pOMSXIYd3UlR+Qh14MbELPLlMv/0EelmInGIGgL7ilXf67F6gyhuJK76
3Hwgj97fTAKFEVWu+t0rYkgQf4EyFAYdNWsfvBtXnG9ZXsOEibiAwh6J8PP2jLY2
RkxAxPtvByHLYS9oVkbNkZSMw88cX0wBVlCyMm4l5aErErRGF/aHuxCXH6SpulfX
GWzv15RiX2cK+lVL4YtFUN6QVHeumvwa/h6XXIu4KxXr7wdy7TZMLr9234vgbwAR
CEk9ryAAbRuFqbRlIvrGy2VqP/OFhQTCZLn3kuXJZaedCASFbn1NdPXOcqSqO6ib
BOEHQ2zqfeQFYOiADjz91uceVpRW4sVVEtJnDzR+nyTbwF74D/dXFVYkv2eO95V0
KEUoyZQVtWAKxuMqlvzblBRJbA3Od4qGUBjGiZvLjJ6nx8b85ErUClB5c66LV4o9
RsYGGvyqRuVPino/lVq9UW/vxZUwy8ujs3I6nN5CA8sgY6Qgk/ZDseVf9w5bqiwv
lO7TNBUBsGi+/+3KVNWgbDajeYRE7wmsTTKMQVsme62063mglTWmy6R8ZavtdFd8
uNBQJK/wM4e/60gGfpcBrPGnRzku2UPnX1rSEJDPgFaD8A4OxtB9olTbWMu1RJ2T
nxPbNs58yOnINTPRWNDhLceZRwtoWT7HrmYLkvx52PqclqzikZ5rlJ7I51uHm66E
BNYiW9C08vJ0ivSqXVZxavQK2jzvZPfaBBB3gQGsQB87feWzlgivzVZI73qRcJiF
huPJ+suhhalOSMAq6IQsLbhqT42x3NoZ2brYAHEqPwCqcf2+9dIatgOFU2cW/UTD
gM2OsRk3ntLyjlzW1EA5FYubDs5fmBIU8HIS+qH1EfYFYvK0Il1siJM0pdqT1xfr
Nc113kU+Wl7/kAnJjzQ7cpebiXM+otRFtS6/QL8uihiczwW9l2EyeIozRJpbBK+v
8ypOJKih4FzCPZjcFx93nrGj7VAEXH6eN1+a2hV35DgjGMqTxMijm0mwvLt+aTS0
WKX6g5MhIWg+RSihk9jrZnHXhyGtNf9sxgTgTzMGvDQI7SyXZMUuX00ND7J+gsYN
8profruiNSc+FSzJuxIKFwXjMI75mBhfsNd9+DCz65/WknZJn+cCyuSqS7ir/BR0
dPrGdAcLKPq5xfXj1RX9Ac4LkXl6NA0r6OMIMa4N8/IpveOdH42MRGXOwD1BW9Fm
R9WUkAa64y3gbO10ACBzE25jZDeIlxNsLDzfrh72u/buAcqngD8Fl9Wu6S9zJS9d
6sV07gQD4a/OkadGcpd3vYcI87ZS9Reiy4bVhdP51OLpGz80uLvVj564DjeU5lUY
e/901zKox1x1eeruJVhSbVi8P8/H8xB7ufNrkpgHbmrCUMYZGYp6pz6c797HtYNg
Ojb5n2iJmM6516JTljJt/TlUkG5d1QlEYGvV6W9wnAuUOq4g5OX+ZZYJPvyylc5y
vddNCuRH7aVPyjc9+mHZAwC4xi/GwDY1ggxuOLJKfmpBqaGf2+yDTmnss7wnSdwG
uB7v+sHkNItuQ42kGdl/L3zGdypNStl2jYWAwLkZH2aPZaxR5730mu/g6iZLnfz/
uZEadZ9623yc3+iscp6lclvLRnVfYkBRxZgsmb3XjIE9hOu6xsmhBE0KwES1bJFA
X8AVXPwRh/RwxYYU7ZuXv4CcJ2jEtJtpMARnZExaJne3Zg97dRrXp5pprqVnpWqX
j8/QL7hHkFxkM71h2prWKt1fuSkBi+EeB7dd0P8GFOTsdW5hrkrlm8ZjbuwjxXnP
G69nEg1AuoF10OdFngkDU+/zpF6gJl49AbvexPyuGLho08R8NUKPfa0Bdr+P7beL
Tbjng3ST5HNATg3+5m7Ue5RSU+WCYM/DkMZiQysg57q4h7ZBfnR6EivvXNyioq3r
3aBM8Lj8rq5/k7vN0iJes+/4lJp+LxvmEIgCIuoouizxvPXLWD90P7SN4IsXpcE4
I4AfaxcI/O/cLobWvV/m5/rL+R6MlSqKFBzmjmV+B8x6zNkMiHfb4vrq+jiwHWsC
Ca9/U+rmnWhIq9+QSKbMDPAjyxcRfT1c5tN/VA8PT5qRkLMsO8h5q7OmLIa0PpDR
ORgEF7ntYPs5nkSFXwCY/K11Ubp23g9pwvUuuXTZLCwTGNFNhUiD1Yq4hTvadam4
mztajVXVbHmuziwPdKndYpSHMsbiSEvM1hfeNGuhNRbFqkwh4aVR/xX0iP7P7L3I
akBiyAIbAWFZJtWFnJR+IV4bz+MGNZagqHO4MSL/bKKAXUejjx5Rj1KhNYdFujpT
I0UqGeOzrAHNen/F4AyD3qJyulfxEqu6pwtNH5nnEB1ipb6IvQNPrmnUFqq8cr9d
fXNnxkZd/b+0Z2jjNhfodc96LVGj7Blhubt53BEqaO98rRipffddOpnM9aRd3iWc
FqmOqHpbWniVJ9yntBxqiJkz36ae+Wh4OBtIm9J9bX+gj2MbAi0w7QHjhpM9WHUE
wu5uMv9iiv7S/iCTVokiIt2qXaEg5bsx886ofj4OixOpNb6UNf1cvKSMU87Ya4iu
2t0CvSK2iJBSz5FYtZGXWkoqUnfPGqU9CNHQ1TKEnT+Gz2/oX+sJBm5YulEob3l/
gdHJ/pq8Ouv9Tz0dEM7PnkyCCKEaq2+SVYJv0PJBBztp8Zmnf2N4TezSsBWo+EXd
Z0PTKPUAkSh4X+EIk34gETqMkYtpaN0LkewjJm1hunzI0p6RKvNnsL2++Mr+2uR/
S/+EzHes58UexWkx8gL9eWiInGCZEzYTt3C1zCxlJsEq+Ewc+QN3hBQQgD3eN/4O
41RSAzN8PdTEm51tcroFrpLmV7n2fdgciUzl9ZDPsy1+m10Wp5n7oCMQnM0H/5iI
y1LLICfKrgP5718LlJ5pZqptAaDOzi7aJ1GtU/zI9F9bjptVfodJ6qKUBqwGSCgq
WHgPHuqh49fCYcUU5yzMD5SQ513Rcf2b0M2udX1r0nVA2hGuMBiCMjxGwQfNYv2E
+D9QoOtHNuadvlp4nEfBwPGLTBptiAQu7avYWdJPEOJUhC28JlM7o6/SoA0iBCAS
t2O++fdX/H52Cl7EqScaZW9/U7wlk40wY0uKAaBhtJhpGvh0lhpAxrPkwLzXi7zO
fUgQHZbo6zB2VJvNxwdscmJNpqZb7y1QS1mLBun81oZaVJC2PfFEEh+NrUBotD/0
riyePOcFw5MCXnhU5BVzNRkSRm0yXUVHFpbso4MO6T4BnI8L3vLlBaFsx1MNGnh4
wmDxyxf2GYotomzzkUjo7QF3EERKHasIg7X/CO80hYSbcX7R7/9CVoA7jrP/cSF8
OWgjdvgZ+dYA4aFB6p2iNg3Ho6q/ViXvZnJ3JIx2Y+hMrugzpgVoPC8U7yZ1TxJ5
2Dg7af9UQGVRa7jHxRN6vE/fB5UEA+8d+ei1bUm0rE/CxQ4Xj+q0ZfSX9cFvLN33
fMeeeMwdj2/x0YO1KtB6do8TH07Xo9g/jLdcKblJKeuSxGrqhRMWrsjpCnPHly82
bvuQS3E1x0acIDVuMRbRwfnnlRl5bIPDbYp6/t+/3QYBaePt7rwAqj43CX50fcFh
oif1yXWgFvfs/VEElBsgXBhIGWDkgYFfXtbIp081PLsFYqb+8X7c6pow7wLmGoDR
Am4p7enZ3nFZ7RBOikev+g/tnSXZkZjXYgJP18S8zOZ6bZjaZHCaaRUWC9mUImy9
KM2OGT3G7cKssyzgBbFCe1kQ+sZK5R3/udmlSUf7ot+QvYfOPKGo5cyZ9e5uhvVs
Q9PIU41Yq3TLOacEikwOUWqZgz9+ookZ2wsul8iRZ9KpEi+45FuHRBHv/gSV/1Jd
2RE2Eq2yfmzBkuM/sWaUeXs7Gy/2EZUrygV9Ck5zlgdrhomRhmtXRLJtofZWOmCt
muiwAIJv0OLiRVbucdMoWYrmPfR4T5y2FImXZoImbtAECSuXN1ZC2JhLq51K6qdm
sIUyo/IRd7Oi+eUV3nhrTfv4ecehzAsrgTcu1299PKCfKPzJ6/sFHKzsN1Ip0W4p
nbUfCQmmwJugW4KPzNKXjYfq+VWwe7zEXl4m+JQwsF+kKz8njowAEYKOXcUi65oX
OXW/inn6g+XvUmIWElQmwPzHN8rLtRR/Um+Ik9aIaMzIJR9WdNjtFE/+Ew04g2+/
8ZMyggCFjnV/so6BTRYhAta2Zyk5Wvj49eHhN2L5EG8cvZQE7dE/VhgGTHIFo5uv
+kUP6MS5BAdr9FAnJHgCHKWVfO2Abddxpppn8+TNxRADF5o/SIpbLEnms/+yrP7R
NqSSvHgT9y91gmdOBHxiNQu3qemKLIqpn2EBTIp3puQblTUc8CAq0MHaXw1C5oEh
B3lCJIPB2H8bNHaoK0LTLQCK0s0KbJpw62gR1TqyN4JInCdKh/4Ll7No6dYxBPwd
fynHAl1ngfEXj5Xvitz7ZPziUDN7Ukx1kmx58a/ChMLHoErnngjX3qkytpZaBq9b
NxTPdXqJ6QlZl6KMsJAcZ/fMF6BV1xdEn/Iuj2qJdLiHkUJDGs2PGXInlGOoa8Gv
2YJ8FBj2lrJsi0XdXBMMrDyl7uVwpgGwo6XxW60VrmpIrNO2Yx1UILFcSr/7doRg
RwyN9OVEA2NY9jFKv827vl0YPhoWW8V/2KJEb8jY5RcMvMfYYIby55gwbPmkko9W
r5JrIR5Flt9oZ5IzosOEnXq+eFXkP5KRql5GHOgQUFc4R/8ILuDfoCU08Bou77wW
laWjpPQrn2TEodFlA/pzPbwtUxGwX/BEfDQPbD9Z0V6X4sFlD7J5Wja7OSeMR707
vEXHA/F0XUXo/V8Fkcgo8B9fUODNjyojxcvgHF9VWF/oUibyfHfPWxC4RxPsjrsT
U965gqy3RJ0MSUj08RSsJKNSEcefYF6NtBpqWuSQXtLHi7Mb0huYkQ+CZt3KCacp
BgzxfqugFC6jjdpHqmYjbHuT3H8cazRlfb9NP16lob94VQF9pvs8PdKuB2F7QQON
NAW8bwL1ASoRJEvzD04DJAObv1L3EZQh03fKlHJrnJvaOleDLxxZchDV5/wd0kqb
WuEazhcuRRTJtsrKcsQRqQeKG1k0MipLSptcgQgy3t0ULtuS2pmDSpQlxgcA1xgs
CoWEYcmOQ8eW+++5Zi1US+C8HeTPyjzSHHyq1G5OjK2Zr5Q0N3qjfLNGlxpYoR0t
iCLgSo97/qZFIN+ojdJgbaw6ydUXpmbBWHggEbAWWL+x28ILmOZgbtilxtaDaARD
VHqGJ8wcHnBuqZH9iTRTSJL614sM58tQhY3y7wy+Amof/eR+0czSeJ75MjlWc9Zb
9KYDKsBU2CMDIhFayxl/U18+ytk8ZSaa6VqqA8SJACBcjU8JtKnPg1wDc4YA9k/L
O4pnkmtBXIPYYyOFcw6sdNHT17C/H83k13/F/DAcaGXKx0wR3Lpyd6FkMAgMyeAq
ciLTxbKZKCcXKVEGGfa7PFFjmrFZMUsrMYfgXXxp36nSDZZwfWqUeDwwIp+x99ID
L8KkfiOVTQo4CuCC0qDDnE/0kxaKQmrzCfsO/ZC1DOBYq0PTlZknRdz9vsk4q5QM
HJ1bo3UQa1zMBPtNNGAUfkSkXxoA7I2G5SG/hG0wxg17e3oFeCBMhj3p8LicESTb
hC99BfwX9SZcxELBlTEg0ZvDhB3kROj6+8K8EJPBbqqVF+3rq1Gm8RJyHeIKPSbX
61/sajuVpmAvgdrDX0q2VLGjdZoFA2dgxQiA1ykY4wB58EWMsJIWyiqnR//NihqO
AYF/8mzEocgeruHp7EowLVCY/hEunxkHAlo7Ajrrhgo7XzlNv2L7uIX+GtoO+wH+
JklsFRudciqaro+6f4EtyvwtinoulNflnpdHjnqjaGRxL+ZxkSi0QObTFtPo4/5e
nCQr6HMokznNtxVbuZICWz6oeG/irtwoNnEBBrT9hBLPtjVDAb1CW7VwTWXDISPO
svpGbFtLA3qs8KcVVbC9zuQdCH4pTSLIVCL1aJ4sDlkr/Vt536L+mt/J4AZ7UeOL
7C9GvbIkj0EOfMwgYnVhH8h9kMvqdBjzunwCs4rNzgAEdopVN7vacCWV7ImaVdUT
obpRgzMhl3g9rpOM1C6KhFjkbGkZC7VCB94Zo0lGlUXvmdS/WmkhUBOscQrazygr
rlpWRARHxBTzdluC62hfv3pV3liojJ+5mdWPJ1kLC+ssxZhb/yzcgQjVRgjdNS4y
AsS087qcuIauWxdqqfuY98x/PVfXj5ZjtV0fegiPoU+iMozDDp/c82Odh3QtWZnc
qITMqY8rW2GigpyvCT9mMYNtzw+YJxoTohiIG76gxe2QNXXQX3IUjd6aWnRUFnup
kS6hFGz5leeBaZa0KhQdt4UvIhWR2CD/gy3kVcmzaEPNmLn7+Bou3lwuRwm7yN2n
+o3++8oC03RpfaRUcgkWTjWjnwChnlDMpkMYohqGxjCZxahH/dCAR/j9T5moZxiL
0rRt/FMZJ9fwXPNCisliH0qLVdpHU8YB3KNly03e0XvmvX0wImK41gJnwLPywGT5
7alCZUu0QGfJg6B8VKp7cbufDIvpiRFptf8xSlhL5fQQU3/imauR045ghHT/vrIg
d213jXyRPP1TUyOr9Ox5zsg6dbswROwVMs8l7uFOjx7yK0k5BBZAwlZq2S5eixGp
4pq1QEUJ7g3EBjvm0FhD0Fkuykz0gll+oFPCTGs3u/n0TNemw2V9uQclaY52AY6j
oDUPPjut0lhMCTT8p8qdgNubs/k++qToO7zDuRyuk69qct3RAlULDIoTPnT308wQ
zghYYgmkS+KbdJGBNQPNX+FSXWJaMBwdaekApLUU36OCshj7E5VVEMya7uL7+cGA
38MTGiRz7+wtuQPuNTwY+VHgsBjsv+rkJ784s3uVIfEcMNS5kiRDVAimGijaTVc0
2hSWfrymqt2p0dBCD0guis1tnrzliOpyYyohLfukTAH8lQb/d6o7DrN0CJ5ecb3X
CE6BLGMeonARIwz/+bixqcNwd1wU7eptdp6JA6SSskxcS9GoD5BKCjpEc8EQutg3
ft5S0YbzHsvJZwyf5hR8w/dofgEzE8OdJyFR45mi33GDpLPWecTZFxHNmKZfNHP6
uMrO30A9PS6ehSTLmDg2/xv9Kdl45jOdfg+4OsuuE8ZiGevFPxECsdim9qKURUEM
9ui6YUW1yBs1OYPqJbR5smQzhtCxyj8G78b2ecMQX1vvx4WFHfcGYKcRgpAcYY1G
3pZh4RtlIL96ytwLGzP8Nw4g2RPJi3fiYCsVElNWysuYrot90DAHK7C4silpD42J
+lz1o0ky2lmUjGYiJ34zmU9I4Vpq4nz5+41tIw5SW9ZKGfWgaJd4uftX32jaE4tK
mz6aDyScqSN5gzmMoTttz99ZocFOYwu7A0a2xEVnFiR1HztWq9A2LF+4xM3IbxYG
YlfonL1gme1UaK+m0WodjpiRIALpHo3c4ykcaTAXDD9WLOA1xkihWVJh63te86Lx
5f3s2G8CruZBYQQjhOKAYW74tLs0+39SujeGqVHeuzfzPkof1QuX74tsxa/XKY1r
65DvGSh08BQyco/3/KjK3GUZYABedFVIHoZRcrPpCzbiYstOVaH4FSc/RY3Cz71e
J5uqGM/+3zKA1PEG+wlsJW05LbKSLylxYB5iZ/DpIq+vGvZLsu4BDKcBcVjITyrM
akLmiNQQ9eL5l9GnQP3GVOfYB6rIs4E74A/pu+2R6OVX5R42BYBR0w4HuJk2ne5W
z3QEo+qEzGvXZfUX5VDO5M4kOChIAg7fhf8YO29cuifLJjOair2WqJlSwwMSy9jQ
XRKBNBDIwMX8v4SBiq9Glthnnfv7o+HWjZiL9m6IkYbzQt/hmQE/D6zbDxA7DvEj
BghJGPwG3GTsjj6SFWFs2rdo9xvBabyar8/5fC3JOIHTcrM3NoVXG9POGEjStBse
OwB7502EhPQXluw55POabmhomkpKc29vNmEPjN7GSYLz7FKNwatiDbz+FXdHDcOS
PExfOJ+lSbHlYourexvUV83/fQ9d7ui7l6Q3EDqhCPmLNpvxX8fvPfiI+T9ttxp4
NbDbLSJYDZZooaubPGzuBiLPu5+NBrs/zpjWEPxjK5j0Q6D8vPGftHUyU+KqxSrw
WVmkkgcaFe1teK7aQ7rzDnssEZx2CPTCcsoIS7SUO528zrDCrDXcG/d8OT8v0k01
x1yj1rCsRXTYKpuW1TjCyqF5ySmNisRomco+xxEGKmeJsPtmscHNpYe4rj2nsrUE
heKPav+Xiz5utr/Z6q5sr+eeVZC9qzcvQHuyObiPImQtvwV+k9N7SdyWG//GdUiS
zR/VYjRfjhiEkSFREN4A+3xQruFA6Tg8JEnhgWU9FxTnFIDqaP8ZtuFlTcbNkekm
9DnswV4ebOJqFm+Mevp3vuGPxy1mUcXo4R1TI7KY1AIFrMcsxk57m4/9xAAaLstK
zWhhjVm7Im5jwmKVqKta2b44ZvdjOHcoWSF8OoCW8vOo13tH4xa16NNPk1Ypjbzx
8CRLk/25jQQqi4FnFl2P7qktuxZzgq8tdrt+pb0b+N5uqgKD5Hmmy3hBiFUZZ6DY
erJqQ2wRPTAZbNTZMwTdb18dW2n4j2aHlaR5uD6Bzvq0oPjbQAkEH50RqN/ubNtX
Mc9YAOhRm11hsmrRqUfSHu/1pw/V4s5K9doqEZC4zJU9IcqkWYBk98qCzHGs+3rF
rIgVS+8ergxTDu1FXVrAhgF1i1gvNo6cL95wz7CYI/xmiVcxZCu1XYqkcIb9liHS
69FMQmVaicY1KouRoFwjDJoxaMUymNyOWkYFnjiiUFlZva1P6zKSt2ueiDARCzMU
7MurLsHKm2nINFvPGScvdrYaCIiX0VI8GA8bidufmE2sr3ZHJz0UFCWf3F/m1f8h
iZK2F7FRbU82jCx5CFirdYynKkHplqu0aVWM2EvmlYWg02/TD7jPD8FOksJ6bB8q
qwHJW0mSv/txBr6vw4HEZsdtFFWsJbLR4o2NYfvdDYJH4aCDjde/sDVxDigX9Bho
Z/UZMqIiu1lMVapeiGmPMJOEGw327OWzWnmSLV9uc8oErX3Zxi2HnrYkEZnswiON
1Xr/TgXx1IQhUX1XSdeoQ7hMMrzoSJ6+LMfPH5iu8u+y6II3xu6TN9UGq9EH8GKf
nHBsBSMP/U/OIsl8X4wC+IKtbaxerMCfCalyMthw0uzKGvB2PhnOCYivrFzfQiiT
hUgC3a8Z5jH+48ZvbHt3mjQjYbZEo2X7otJY1MnprRvCAAtym/+FU/acgDVA5VfY
S5fN4qd4j/oFaj3jSNKlmrWEnVYbGfbSaYy2n1yUvtviGltNndUQeqpe4eX49vOa
TThS5OEdlTFWVUMHFEHag0pGKA931sXaIbrYqKHKOOTYULTZsPl4zAJJiuYXn+ES
31r61k4JWaMKtyLPFNOgTJdgcKMO6ES5SvPRGlBT2TzFWZbZjMlN94K7bzZxAMc6
3Km8ofVbThbHxns4CicChcN+DtmeGDRjvL/rc92Mw9VsmeJYHJol+Ewb37ke85G5
sm460cgZZWBtZgISdG17IiBygXSELkdTM5s+rT2/LqfskK29PEuF3LcsAceC196b
F1Hm8TbqfnV6x5Ps4WkV2w4wng/t3LkRPjQRXyUI19UqstVRNoRpb19FO+/cat1J
ANtrYPKRyudxDPNoOoApBDA3UvzyhW4cEfcQSGyhHWkD5xURm1hH5wIsNO5oFb8u
ejotKRFiOUvX+HjdZMlg2Obzei0HeIxjrmI+9Mjk09O2nd0Q6PbPi/WNcs2R/dWD
uS4OmnuBpqGxgLxFhzSinltkT4I5Hj6pcjTRnbd/wPMZVH0N6iTA/JfGd2N1ik62
YiimH5hmZ6vJvL7W2Z95/3LR8SsRJmBQaiN35JZmq9rBAJAiDQMb4bIEVjIlAs04
rNyk3b93ldrV9yLK+fVSEC2X6YLX9bDCCe8GW09phQ5fjJCPJlMrqxk1JFp+FH7v
AH8Ml4f7z1wrQObPBkAKFLKz+LXdwRLpUG4kaHuYux4rBOezdp0sIOwkxgmX9Y6a
XMkPoLX6b50PadzOAWI2yZWfP8C2P04ENqQWvuk9P617Xz2eJshQfJKR2IuTE9Cp
2SnxkZ9T8rJQUH0MlbwJXOb+6/J9XgMnQZhKBg9cGiPHbQ3fFArN49YCjmoiV8kC
Y4gZn8Izd6+sfjBp0y8ksHDxPNJePtKR+vEFgnBe0MR7ymqTwLTph6jrlNUuO4rf
6wzO4gedJLd6WYu3fhsoHUNjUST/oO7I+j13NbCYIOFXBzsBAF+4xcaik2XPpP/c
KDS0ftv/r51BGfKF2d01KU41b1VdwOMH9UJBjEZgbs6rZN4v+qn47zkQ/WgOrFht
YZmX0eNkZWdBnpdPjfLidTLF1YRwM4XXjVQC93Noe44lV5SLC7FmTtMvhM4fODvo
ifjnbtEaqWEDOyW4vh9FJysYEZseLOdljeoemXUDqWzdflkReb+pvXAt0a3ONPbc
kcHNDvS+BPKaEVntcETh7vfJ8/2ikULqYHPErIxXQfcf80omytEPQVsgZNpEnkb9
f48a0FsWUZUMOwGutWbc1djo5pe8T0plY6i9AnNIxZRqeOF60gaVM+bJNxEMVrDE
2LhKIr3oKt9+/IdWvTbTJFyS7bciD+EO+eIzVpM5Kw6EerrD5yZBQHiuvIxYmoXk
9b13akBRzi/d1eop9/nDqv17uAIyaZPKobo4Uk2XqXl0QdY8Lp3yVL54conoueiY
S1TjB/dM43kY5/JFKA/0uer+vX8RvkRxIVRiZ6v6ccXn+Crs1YcnmU6jPgp7NvC5
BSumAsh8kvDunuXz5rwkvScq4e7TPEMhAl6tNgWjOtbV3c7wSafwxZCNx+piIm65
MCAhyAacaixB6o6tXsSUnc/oKrnXPu9oh5GwDWfhzgx8U9IuX2YL81nD4+RwPskk
u/3n48sazcic7FsQuQN0lkMihO8+qJLQJ6xJzmkF2dE0HCfIhIneVcnpdp/+sv7K
uV6tUbGmhBYV9eEk8Rzj+Mr0Ts41DMlWNL1bH+TOBDSuPVr8Klq53OOAfLKD8KB/
/truZsVdBixkWcib4wSe+fTwZT9YU/eCnVCuvAcDFKY1cQuS8U3tnZwGGbxN5LrA
JiTNk4yp7lwFsQGCkBrhCniVAyDYYRo2wNwZ7DYtf+ATW1hE/RB++8WAlan/MzZV
t4teDcefs8YDOpmYnih9YX0zG2cF4i2O3UmXmvs/6mEbkoHypxHejBaSmwDw218+
rr6g360Bhifrd4FhjLHJmCd6fCBg2Snz59rsUdg0JHD/j0tteCbf5QvmFp00qzlN
5jGmUI/4rjXDgzzw8GiAunAdn5W1HamzMwAkrV5zLJzrMngP0Bby/fYv7n0grM+5
lccx9P2o45tAgfkmCQw+CiS0+6k3jaDjCWTV/Koja1OqkvJ2CzUFazOnCvliGNw1
IgRAivDYnY62swNsQxGO5a/6WpYCG55Df7EU3eHDSGZPL7zqxahLaSiFeVzb4T97
QDX2AhiY4gEy6SST+yYWXConu+Fk9L1BuhMWZ2HIab2HLjheIQ5qqM7dehjHVERz
xIVyCpLyB2EeLGfzPYkMMp3cAlV9zNgS4OJsAc571cyDXKrDWX5pZWufX4ndmVbj
Qw3i7X9TqopuiJ5eHpzOi43r9/p2OK3MixIZWhLL7YDaM6vOkTki6nTusqkMz8b6
PjmD/izKUBwgDTwSQAWZ0wGBiaiZ8LB+xN88Vymc5OmcXZHsNZWDdwP+Z/r3bWUq
4Xg17L00HnfuCCOpX1Vuhh00F4RvmWM7pdoV+Y6el7YQb5b03X3H3BCDB5qSTfHB
kZkthpZboBwit5fRUC7H4qQRSzk9TVPuR/iWZWhI8Tvka3fdfe2fLcxk+QPWy2Ct
nthX11s2+pSv62o9tqcyvwiuYXCE5qDE4jqWKiSHB1bdB892k3/oDP+5HGVxNR3Q
HURvWpGcoL8zZBVIqw++IDR8kSU3gge/eXvIvr5w84fyEankooBoE8S8/b/UtTBM
Nw6wRRusRbZkSH+WhJQpMfqQUYAFr7B6Mjsyj7p+VK/lIQoW0ml/eMaC9BFYODce
tghvmixbiCcKs+gl2NX5urTKK16sMcMqNOra2vEaLxdLqrOxT9Zpu9Xa+CC/D2QV
M5tABe5dYkiKeVqmk6VyD0MWTFdDJVvleS2KAJDkOEYZlhuw8fNfUGBZhNBoUkUu
zt4HGJLyQuhRPpT43PN3MITZmbTg/Pdf9L4CQgcdNKLjZPsS99EFn4Atdz6PXQrY
mWDsQzxr/rWWjl1ujUkpxw7HQuG7b9zSGnq+3fWYE7xzYmJKRr6KvUSlXgxhMrwQ
lSBaO9cwGENW6mqzAb6prhmAc6Fv4TM8W858p4se0NOOkHvTs8UsCZmsQr6ny0A5
mlMu/PJ4CELOT01zBEhEymaDclusFszhm4XuG1AoVwO32ecxHYDzCr4HnxqwGTZA
kett7DlTby8ynDB0kvzxHwXBLLZqfN4zMhPMREot3dsKLhe0645KLPYpKIZBgzop
cSMGsJjBfGMOH1ctS9m+lDochkV2MkfxULN0N2CmdpTvKal16SoR2PO8VYTbqg48
8GUte0o0lcX3vrKxzCbeFninn6IwFZ5JMKNaMKjH9sN2x+ytjXq9HYR/69NaS4+S
Vo+U59YJuIiDxNuvN+KGVCKHYo+/GFMAiuuRgZ29hh1KMPb8Af/6J1MTUqebFDXL
HZHKP17xwfOjRva6YuJvdJ7YH7ACoe5pJLhlNVHldl5Ls5FblDPe8t1/1T05W7sD
LECIairvi6lDYhTBXeaS1AQdQIQXzMZoxOgL0Dp9HoelegdmLmT0hNbugMZY5FQ4
Z8TioHLSvlDRUUJR7VIAMp+yiVKg/lQW9ZI4MPra8PKD7xK/D8YOHGMw/P7PkeC3
vBYWqgwbGljOlI0ncKzHG+VQ8RxiF249qI3XWaw9b0tReLMPAA9saZUAQUKx884M
IYxwloY2yeuEF0en2wBtMB51MjDXNtHe1IHt5KRuAt1kOQ7b/U6kXnzqrzlB6zj5
PalJD1wEHg02NTsPzfrR5Awp/3MW+9W0w5b0IK8Lg/kfU88OVFO1XpLKMPpKQ/GH
GBfTpe8kjSkTosY8m+4Ll3yscHEQNRh2woWoR76OiL3uFyrm9ZQPqBbMoRN2FOOg
tIpGP0yp4dt/vTpQ8A+16Qpd2zFfBQ9EUEewDcZ8Toohc/lCzqGvy67QWHTipaQB
byRqwm4yfo/B3g9m5PqNZ0EfGv9yR+kt0tQUi78J4uxWW2PAZFwDy1clrLsZDnIy
HtiPqMlugTg31cHhjpnomlqk8/rOCHwVYiACaixTgdj1YEnMDFLnG2148lmgO4HU
GeXrFyeLF2A2lObgkX/qBeSD2WIwnO+lZ6xAsLwavNyszqzp2ng4LX5FnWgbRKYt
sK7r3txpKzZjI5debcTH/sUHQsj38DBhg7OVULjvOKPk3lL8oqs2cZ3emNgaFMx/
xlyhIisYyZr/O5XeJjSIz7bCzs2PFnyVS58F4GihwmvB5ZZn95ScxyRt7AoF8j99
KBHxtqIjJD78NYRNpMT3NTsltSH3Oo2VmW68SDzq01yrkZwCSdICfDoDNIm8Om4m
MDxEU70ItwJuT2QK0xD5AlZsuCrUCMOlDn4eE4eLLqbEKIKfxboeXbmSXuV60hUW
kjV+Zp91/C91DMjVIk8UhRQikItVcpMPxHbPDRM5qZQtosXttlOtkMjOrWw86tfb
SL2P5wSNCNeFyMeBIFOy9DUzKKstIEsmRmTTC9BFuC5AO8xBKO20bwgVBOksefJq
lZTbDvBzbOnhowSSrg+WcpO/eskKYaID4IFmWzaVnriFf54ZeosaT8iSs+Xjurqj
6d9kXajTjvQgPUqqtFF6tAQXDpEDGVyM1VmDXSrtQc90x/KoSkdvhoTzNrFEEG9b
rFTO8vYhzCVIQhO/IlPBzDuaR10LDJN2rlPjuXR+3wZu24Pb5X18iGK/x3scU0Xu
H2SJFzrBpvhX9CtxcUJoap82MHwjWggSi1FtRiBZ8W1u5sF6m6kYhUbXcZOzaXMJ
QimreDPk+wsm/HLqEjgOtOyWQCHtBzH15rLBGM0aesXLqH2eF3WtHMBIGuGyBrmV
HsS47kaQsbEBiaLyoDwuXuYmX/DH91EwrGeUVNjTN6VdUBWHLCS2s0+ifMUbDo3a
HfjQuJMyJEkSFHTRDVmWFLOyqzLlW34CQ6lqafFxj0hrxCFoRB24ZA73iZ/JJpbq
aVhpN93fBCcPCiiz83LuX1CWGzg4LwqNxuKJSE2P4awEvx2/qm9AZaRmyd3yaa8n
hY/PFeNwifaisqXv8NQ3LvYLrwn1hc/7TQGsgB888NaSnzrAMwqbzXfZ8w0FIQvL
DJa38KYLTZmgHu6qJzUGgPxOOpNufkdPS+8EjqsifIU93VEzs4iZUt9V48f/Scwm
GudygrjbTulIDcfQXUfF/WHJF9XHj+igFHhvpk1I1GlWXf8fMsYTP7hHjATGqYmw
Kv48Yrvpl7FBOotJNGhIS94vl3jm+HjTQPFKPj07RZj3eh3ahoBbRv4sCjF6YwJl
hEkZLPfRvr2HgB4YAKofkeqKqZ1f8KGu7o+zvGBs4ScVx4QP4MghQV9ScKaItCrd
ALP/4i8sCLk1izC4m4DLwnu8pqagWr6+GZL4SagOebnjqm2mb6m1fjmmTNBIyBka
M/wkK+kE85BoTVfmkH4QW1fYrrR9IZlI7L7UgBUZoXW3vpMPEbAGmDNoqiobpodI
A036msIlniW7Vs3wLEbB6MhKH8rooJ6K6vxSuLTBV0ycskYkS2bevHn8oyvn1l0o
sTVPuAtfBMiNS/cRLULXkCGl5Y+c3OV0GJKRSAEZK00KWeNsFumFuKjFVLZGZNDd
86TFv8XZXFlX0Kgg3LGcnZ65V6ti9NxJs2w0dEJSg/a8dYp/KTBD5VTVli99mznk
tAUSP4WGLfebP+eog6pENvxp/l6Y3vfmaT/iJO12ults2eCPnE8U2twiAc+huqrR
pvdN/UFoOlYMDU32fNZJL4z6hJrw9SUNAS5NFASXHqEXxA99+olwySO7BKFu0xb0
x8REl9O39j27oUWDuj7dCzubMvWKcchVg75fVzGjPIyCrZBTHg/W6AZEFYmq42nm
vIo+/0tr9MkPmmbnBqEa8CvcY/PuWYCpjNsw0xLPPM9VxpYbHmWL/+E49UoeEUw8
3LUk240jstken56qFdJ0kXIXXnkLTd3vBRYV0r4V8nRypazq3w1cwy2zMjtQobg3
EUlKmuhJyABIZBruTkHkP6u+zOay1S45HA56A8+STKvJN7cttx2E7buANqzmEAhw
ZDLY6nMNAAON13J9KxnC7e8KTsE9YooJj7YCqdEr4x6tZ0FtXi8pwPdWo10VL874
/BIrBMBybbvZFX77G37+Bwt4gW3nGvl42HShCK57cxcdJAHGlsYo00BV2MsCQWmq
PmWxfuPc9FGaS6AdZnKGhyCLm6TIq+LTUdCY4iZerzKeDaiMRntq0YsX2aqHZ7Uv
nc4P0r5JreAIL1SF7guBdF2/3y+zHq2Wg3WonZp1Dnf4/zR2m+i003O+m8YJtUxB
JlLVn9pnkrye2+sbTKiTM3XHRy7gYVaWAhXaA5AHCqs3u4W5b/gbp0O8BfIPm4iQ
7jNuL2gFwjmr+rgx2UNmLA1+1aDzsm3xjKqmPJoNifJFeaFc3yyYQPYzkC25PEMD
dMLC2Uv03x5U20jsSNjN3VJxqMzkMYNvgNzZk1lW31mBpuAJljCD3l+OPV48wyrM
PjoDcSKuyGBIdKv1ndI526HPnRTR5ob57EMf8Ugdv5KUDyeAZ9KOHQIgfIXGK3IF
OgBRTAd273KtrF/xhJIvnql6p1EW+JVkTdkbQUcrzoQm6eXPp1obzxDjvC+LfAjO
/HlYisB51yZlWfr2mH/95vzCW13OmmSbKazYRrsgh8Ope9w/YdwjOfMzYWFTXqTr
4JSAdX13d3I+vJqwv1w8uWhmw+PBWqF5ZN3aWUde5k/9cCWMjJAJ+tqgMhHteFBm
qHO7H0bcK1j3GSHVXXJvfP06lAJ8B7m8LVOShvClGxSmjk6NzTzohyM2hEpWIitT
HqOVtWQbxLyRTGDKPWCyhWVeRZRf4MuamT5sROnmqNxuzB5LF+iETFGDKxLOfLAh
tra6xpJpCCzgcVHQ8i6HXW+JP1psRbr5IdGN8mIOpG5nepouXNK//lxZXnZjF5td
4ksRGk/YYUfgWU9VpI7sEMNyVFGhDtPWsP5U5CG/r9omK9dDJPQyGX4g2n8JWSAx
FUsfkeyvSg0YfUa987+wu7dzwESJ8qQ7Mz/uMVXa1cgnA36xnH3/ib7GB6IaMElj
9rE+xuTCihKzSUKeTQrXU9HcOp8Ua33owtEGUFWK9U+cR1dgSFIWKuqwb51SRLub
V34eITKJ1+3VAqD291YUsMw3rW1/Hjzd1GtwVz0cn9SSWYWM1c8pl9bdEzF1Cwcu
X6l3U1eZmlvRgaMbwwnVkiOLsgQSuxfor1D6xyjc5z2+g6vKaVcPD+nMhVw+3e8R
MbZXjV2n2r9+Ht/m6/6nO6BvXRbJWXfpiwAT5b3MlgF3KEaQE1Uj3c95o9o189Go
zpLy2cx+nhDF8k3DmGmNLquWP8ipa6s2MhwZGfWnfhdRArshat4nnxbmdPrrX4m/
zbit6kzp1cf+k/APuVU0AodDGS7+M2Qzcq/6BhsFd75hxgIXWiLiN/1pAECGQXhY
xThRfP16+5ThUCp3reQ4htcRsW+Cog/5MiU3MHfTPldvZvoNjAjBMC6ELtqxZXn+
QT7mYdCUfsZ3KXnM4WkXMpAsp0gLb/4USgeJEb9SXTB6S5LXqtQvY+Bi2Uq3G/Hq
35m0jie5FxbZHABVX1sL0wjj4exHe1OrewCvXKFud8siQRCmbNY4KodujoCDDPs+
yZRv9wSGJCNLOm9ShGbCGC3Getvc90enV2wh5lAFRajVx6Wxz57y6t2QusAmwwim
PUSvHrW4Z3U6I8A+qrcDTKlEnCa4bkmGn4OCXqtOQKaKY0kCLVqcF/kKsmJTXqhN
gWlL0XYNwXOmUXhM+kTjDq2qh9IolZQv5YLQ4nuSl+wsZROH9iIZ0XVchUaoddqy
WH1pjYnmofsIYuONgnQGHHcu5JL7dVXcZ55BCUFcgGHkMQPJAc0Rci9VCjfaXwKX
gK10buzu9lFe8MeKW1g/toQAz/jACr/wiB2wpRkNrDfJjmS0T1cpI90hsWTw+Ohq
41kSdJ5e36Zd/XCdikFMYi2v4+18L1vsVV7Xars0obFwm2MYMNXqhSjlghN+UrxJ
2e5rv18M4JXkmh/Zylufva+40rGp/Us/K7vMtUXAk9sLh0bgJgssAer7zKb8xQf8
lcsNVxBUuO2VXKj/KG/J8Mk45WNPpysXgiJ0aY1Hb86Yotwlc3piLzE4wybVs9+M
G/kmx+CseIT+cnfRwqfR+QhzrkjSw7QzZBAbGDXW0qPTEsx1tiGYoP1xOfL0ZtlA
MNeOuADm1kdef8y4LF15YlXkcSm0J9kr+LueU+7tdsYXFd6/i3fb7crY6Bgg7Mci
+EOI88F7+PaZEcerABj7RtrvWZl8pF3nrl1zSs4PNB22jl+VbD96NYn8vyp/UXSf
ZFdHaClVjWTNRELv20o8GyW580R2oLP3jWEf1wmjXN3it60MZWlnXAJhI1p2puY5
J3ZNiMwl4miILANbv7HtdL+uwYsQHqCytjVe2MhP5GiGP5DN/T3Gq9ehsnb28L7G
Vm0gNwAh/nXuXAV/tCZSJSZD3h+72kLGqEj5ocb2aeIAqKF+ZqjAvy5uV1gMXPUr
cg+q+yzF4U4iEj3iOsXMX6g3ZGrxG2w/717oKhZV08BJFzZrpzmg4xpYhdb8seZn
CmWmvD6l+x2QgudeR01YYcee9fIajXC7XYjvix8whEBdZ3aZouI2pd1wLnnfsbiY
PDsZMCE6Qs4Ay6b3Ns5kwJiuX5yMwYgyHiPTp3L2cd4RKqX1WPqUSGvkNvspXz0E
oKPpd1/piVVV2EPl9gAX1WgAZ6btvR1DqwSAZ5t+SK66MP0FmGSitKQ9BRzorwK1
NOw3GewPZdHL0ojVGbtAchvSkoNegULiu6bqCXcfNyEmB/1qq42XjSyW0PUbrVhX
zvJYlyz5w3pF39g3cUawcaSPFNQHRfe8kO/8R5xwh6R96m/VWOeeD/qs6NJHAC0/
262tpak1qJb2AF+WNa6AdxiWe6SXN0i5DyN0PAwVjOrafW8GkGCAjNch1IQ2vFbS
cYWfU7RUt54w2ketMIFCOcYRBrKu/WOLDIe0UThTzFeZKNcJRii1VkV6ZUe+0/R4
OglKUR8dXIPYfzsnJQxE/XOwfrBILGm4EfS7p0TcZJWfY4+A5yeDbpu0fIpwebd1
fuSt6FnYLTm5d8Rwy8mEF9uEeFzA6MJFRjU/touJN1Rus+2YWm0TrTyRgRXp1qAV
eolgDmvS9TJPJsxN/wNofIr1x505xPvJawiSXmehy7XjDFNnFqcb1JcAfncLDDmk
OFjaibSmiWM0NDYkr2XSQIRIcwbrEzk7AKLZFelxlm01NWH3JfMBPWqvdvKd6qCt
pr5+2VrnUZ1v9oiW3sadaxiCcnAp6I7SpW/0pvesu8fqi32u+M+AbUtdaNldSMbt
HPHGfbIG8f00w1SIMeqIcQGOn94h9NFvzpX3quf3XUDukmSykDAXU3IeS+qKTCgh
mJxpN8DDiSuD8g5dkd/RpKTzWG/79CcKLE4gLYsE5j49Nfvwa8tGiwG4Xuttre8u
m8YQ8dqAlE34xecihEFE5b7mrK+QYuHCs+B36BlFRBCS4vPZva648q/V+oJ0tvLJ
FLHIpMLbBgxVubyEZIKYlMeu8yuf/9wMg3msJiYEL2Wm7HmYritjd8cYvgdWswhA
12jcLhiSO1UnEf3ZhWKHnHkqlAfUYzyTAMCNMu3kCvAnr0GYqqaJ+wFm0nEbT0td
5b4H1IV0p+QyB40ByeJE15jfHW6xwMsw/wLNLFuOjWQ5M0+L9iIunG8ldgRpJMMn
jVOAius8BSZi+HYvjdjV7qj4tFlQQSZI1Rb8EUGhOnjfoUPgFwDhgJWczsCRcFE3
zNqIaMmFxnPWDbeuT7cNus5LezmrCrE1xqjzitr/PvbvKYjw6ctwCbi4tcoop1K/
qhppeg1In3BicyaOedzw7pxnlWUMegNnZ/5j5A05MJ9hhl/NzECt4t1WOjX2T8+f
4IshZb3vQ0LAgN52y3d1JLGptP8dSqTnCDwF4VlnhWGOBEf2o3IGMkCX6UgmmRI8
WbKAQPW1le/s14HAsXihbY9laUhhENA+gTDGB61gm57Q4XU/+sXxTCkDG4nxemCw
ChmF0AWoQajZirIx0i5uc3EhAV/XQp4eR4FKIvJLielzeIbB1HVF2TETsHy+QGQ7
xJfWVQZTkVnozVbbWyrwFCOu30NdClL+XhQY1XwooiAI97V6z/M3cQ7TeYQKX/s6
eWUAS6kJ77Ya7kC8TgBZ+/MN39gKfztI6hzcuAOMvBS+hOIwe7OGUGeU882jFI1F
DipbNJ2qF8P9EkmkKCbwPuMsw2UheBll0bjXimQGe8ACve2lHHBLDp71rlQRLSxD
ApPnv/IY60K8ohgTHQbQThclcouuGqfUCRYkirWM58PqR4Ht70Ow+Iw0aPUOdY7i
+GQ6plVgfG3ezCQPhmdHgpQk8gwjsJB/zbxvzZhAtxG4O/JVCw7ZJbS8etejfw8H
rOOXIVkFqqXesk0WV900fYReMqboomplS+ClElnBiKWYXycpp5LXZLjIVFhdelTm
23Pa3LnsY90HOBwgDoY9WkM3ATdu21Iv1TkPtUTzaoxR75G/bBn5p3iZvPaWQIUh
tiUYo67uiU+CHW8G25/XUok9uPvz0iOCY7hnPF/ZmCx3hnd3c+cAjwYbT9WXGA1B
9OGa5aOrQj5FHdwR/MzwgcWv9gnQul7q5kZ9gEVEqnzmLtwKHzBrZObCjH5EwA0I
orxCkc5zZQCy/zByVQSPAACcrqdO5bxXdy/9E6QL7hInvd3jPMcY+h/Sh2K1jNQL
Veeu0FkZrTf64ZdoR8kXWl1qUbApySzPZdFcYZM6dbSf0O9qAkfWU9cAim733dV2
bmIgkVx3VAlz2Yh3OrZsi8YuIiXmCIxhIepQyX8cU1wmza9Kyr0w0G2Uhh877xvX
8TndYperkC2sKziCHFBb3LZ+bPQZjzIIAfmTnBO9arx/PJpfjPiVvsU7wiEXPlPY
tvFYwGQkxuemkWATdzz0S3elVfn/WL81CfoFNIBNwE0yeWYEkNQw6i/aX387JxBI
T7XHMCIste/E0ojLU9Ty07DTOnjuUPY7UP3Bg5DUfIT/ERbut1j1M+aEpKZYGzfn
C5lICa2tuqZHuTnWUSM6DmtXiDuqQOMoCtPL0fowOET0wzFZ94yh33bitK0f/wlD
aralhs8c99P/WjegYmBjq3vKFR2Fp0jn+ya9uYQAiZcn7KygA123VexeCD0qS/L0
/cMo6aNDutkk0KknLHooTeCGZA/Hd4YPmrjX4l0Q+TH/yR3NsDFvAJ37rrDWSKTi
1m8KbAASC16e9/WP2xE9e3DsodX8GkkoIMrFq3gWOVt+wr/qKP4llaW+9djhCZRx
RgodP+rINPZnIi/I0RSuA8WQlQ53V3nz6x/3PjBjx43FDUPDwFlHveNYkhFc1MS/
XYlvs0lg1ACO7OKCrPE+tIb5EjlvmGXwARst3e3rvGIxc9FfKa6E3a0Y6T/VM/DD
HHpUINZ7ClBuz3fbYE1KQ61a3FX9nhpm21newTRCcaaaBuZeJkoVrk+HaXVo8F92
oHJ/k2JEUCSuOH8tOgOfs6mqyBnfCaJ5gL6hSfJkgNTriaTOea7H0Ldyis0swsnD
axkULMCfzIYqO6HpynQIY21qxq8odZeWWrZrmE0SBzoTmdJYMPUBGBXr8KBS9vNK
tIdwnkDSB1+8P+Yoa1iJx75B/tf3oP/0rHiJd5F7jmrrmXOzAmJ+OmGFs1fe1AVK
Rn3mafXlW5WnjADZY4IjZ64/3vGoFVmh0jSZQfd2di0iXQaV3qZKPexQocD7pDS5
Fh5YBaZNwCYR3LwjeP87b/SbLK0Zei7SarBwhSso4KS5yjbLVW6zghNhdLnRq5l1
wcA6zTTTuo+5zL42qyZKMEeuZ5LhI++LzK8bDEzVz2gl0gedwl5PAxB7QHBkOuWz
mgz4o12raddE6nX08g6IlKfd10sCizqNr/Qg3uSLEgwPceAIkGm1WDQROK1BB19z
Q1O0oRyf+oJSbEAKogvVQWyLe9Ov7cNGhkktnJEqe8tCNAKxmg+6rU1bjv8ycWji
Tm+m9Dqc3gkEPu/28i9VXotb67p5mX31O7Aoc1a3JfmR3Bev1854qnRxYyMTFQhY
kfLOJtmZR4fayuYmWehGemHSi6rgzYTk7Bf5zhnK/0sjuW37T3jtishHet6EqCnO
NJPADgjRYd9Y13dx+aOEhFQXzRC08M/FIg8hh5FDCGnWzV7PqVJ46SMC3Cq5/vTf
b/PTvu4M0YvsP6IO1BcxXR1Sk0QBp3n9IhVbHVARReN8YdfRs7bEgLJ79UQGsn2M
tQA+6WCt2phMg83eutHxGrLThINxO9TEGOYYFoqikqfVHrS5G/ccUz3lB+A7wlWb
ngoFtAlpjfVZJkFEEceymfXUEt5RsrhC/IBEBXfp/h5FHb9brlfqUnJCf/Pz6PqY
gguTxRbjXjVpQRMBs591AQzax61tyoVJ13cvPcw6JWyEiv7BD0gMlMpc05DRsMzl
tRofdF8ckaOCpRMahEIWtnWFHMadTG8BV1hGJ5P8jJ3FytE8afTCkvO3RM4dc1Vs
zrwg2pAW2pVXUVYBtO3MKmx3bK5v9Pzr/s/K69IBsQBLlog2yw6Kcz8T6NDrQzRA
Vnt/0WRzm41D7GbaP5HZY8rYKnZsNd0CgAUTWYWvzD2XDABx8oxH4wz65bjsN441
ixTUfnZw8+JUe910KnkiHRpsoSOMYE4OR5p6zkkUp/HJDk5x4uxhyCZJwKd/KSp5
wsvwSwyqHKe7aW+Z7XLFOfwjSUCHTeV4qaZbjXXsyOCgpjrzfrYmBaOaVVaNLN8U
csCxnVmis1zqzWIjF+KkYe+G6rb2wM4THxeMzMAlZlkllctJGM5lKw+NXaeR/apV
DypZ7gop36zB4rb7RxRB8h4BzVKVPMiobJMgdzxvZfBapsA9LlP37aYAlpFxMpUF
8TV6E8c3znx5iNJfgK+A6jp1GBeowVTPyM3oj5fUeHDcIxHobn/mUOvr6z+SVS/2
EWGLCHG0qU79KxoOUkjoj/yfHivvviICjif/65jwptADlHWuYoM5xigltmxjLVa4
/L9FzPzlBsAozfMVuFpK6rH4t3cOVcx36WspBIroPH7bV+vCsRuImSWGXE9BoDdV
JdKVXXG32iX0fG1CcOJi0VUD0iOBbBhUFGj0h2F14nyct7j+qjvI5xhyAEaXShz2
LGfFdai8AX0+WWGuuEV5QWU6naxAxXODPNaBSFTPtQEGMAL3wc5SuS4BooBl51s9
+pfn6ogHxFx51fVuDMq0DjsKdCRoZY8L9MHGRIQMUCoLPcYOjhwGmOakeImCeM72
W+q73TVJokP8pGoyQdTS/+V8nIUD/Vwe+mZb4pk4hY/KpQSWhL18j+oSKZyF68lv
DsTzuw123uKhnRxAI3MU1FivfU6sclR4ojsAi139NzaD4nRRlql2vGH3g8E4m8GF
oCCARop33arrJf9w7bm+noRdybh/sahVV/pR5OwZ38zJSXriYNaIT2CZ1iJPoAro
8VT2ATlBfJts+iA7lmzm2ETWYZzbB83mID9iRBeqU01Deg95UNdHC0BiU6ZwYPGg
hkhnmkUyL4Qejc7vkzDs3q2qfTgzkbw7C5PejWg9Je+AZ4W/vszV8x+bCurRR8Ne
NIeRTugWOmqmPIEJGVYRp0KfY0i+lJwnL9HeWfV0GuPL5K5fy03ydr+3tQ8Si3Am
pmceVtqGppuqndJHdK06oG5tJzsyFcqgcySC4O+fx90fBOnWzW1y1ejkI1cZhb7D
kBrcoZWfMzhJ2/920MKbngWC7ezJU/F7TsH9VKz6pnGVtsLkuurt5a5hn0j6zoOO
oRNc8704Vgwwrr2lfvLFa3zgX61Y2r3kRSB95IDp6FO5QIxmneoM9/+NMAitFkD4
gc6kG65fRssNM65JQjgl2qtoMkGt3PheaRHU/z9Rzdi3Dfvl0+cbReiSGukTlyTi
baI4e0w8ZQR3te9r2kdKO4czoEMEN+vOev21vB3O6hFTIvRFmP7AvduwH1pzbYP5
kMT3doRbAXNzUvU6d2gzv5Ld8eoeue8KjFbU8dzaZoQIezEmbSCpvM/nUdWbxM9c
NoBiU+m7INL1KUJ/jTonujfBgLurJzL5H6kAU50GV1fk4fxnH5jFOqg5kUMD38OH
WYlGG4KQgJZ7vX9NVPczXgzBueXDkLSiDlLpXeE9lu4d2NUO+FItBHIuUXtdw0yA
091eInsoKXb3gLzSGLkNSf1nYNdefg2AveuzqaTnqWTcqP5jR6SffZLa5b5QTmPx
LPkEpSB3+WbW6gt/YVIrj4oItqtgot0BxMYEDYkRiU5ZPJZiFEJJEYdVit7lw6Lv
keXb0AGRIxOq1ZlVdpHZf+UOR9eKTolZj9HFYvDpce6Qga3cfpbHAIUxaHxJmv9u
rm0H91BJRoI4isGwJ9+r/6mucvOo48OqwUFVLgX6uxaPQa3A3XZcHpYD345cNB0N
pQonJPi2l1O4Hv4Imc4trYbGQJiHKsLWL4SC0V3gYvYhNKvCScJJPgY1F/7nf398
OnXAKjTnY4RJPoFtrhj50TyE9HdKQliPZ9bJEVX6fLP2R6UdTHd0k0f4R3oRBwFC
csIXRGfDK7wSQ8ofIVJoYxrGnTSlGOuvViS2czW/lv9IV3DMxTgm8uuOk9FkyA/M
ttSoSw2F3g4PQ6Irv+cE0fZN9zSr8eJ1Kt8i2bCYBmYZW29+Migmltko9ibogXRB
+A/qO3LJdIWuHfR5EHv5Dj0S4bOAjuCEOjcB7Vp+jQmfQ9gzLiPKxCNhr9qcwX2+
OfRr9AVSRqxvJ8NBPD7tKpunPHG2cyXziwERHrwaGhvmK/5/WlAYlSnJK0wiqsbF
GnB1gIdRF1A6gBqfJOS98O/OFYIt7ITmvfLxpZAxF0gLRei8hLLnVgvRaF9syFIT
jH2BOVP/XPaXFt2a7JQPB9Z5kjQWD3Abtnea4hNPeMGx8DVdL4O9nm9kvErFr3ou
J7wPPYKgRPtbQvgJnUUAh81yyhRqq3p2S3oIJNnmZ7QL7C2dL2JM1LVuiNVrqYtS
pQnICNU7KIh84KtZcAIkA+mFpjG2rNq6DFpb0LzoADY7kA57+F8Xk+LULNy3eWEC
QqAQ9GLuYWF73gt4NsLTxN7R1LXxN968m+Rx2UC2WwvyrcjcREKyVRIoiSucgKcs
xGr2LgFo+KUu741rC/OgV6DrqABIzOZTdbc4lWR4Sz0ySX5xIBGLnI1nygS+U/TU
mNsFqUGrxDEP5g5Zj4bmmNu2eSj5Wy901fE5R/iMZoCx9t6fPoI7j0N9/YmeLixR
NSkQ+6ef9bWK53/ehuIs47RMWtjaQ3PaalQB3DFFA9Dw7Wm/FcunEjnOmY6mw2tQ
TisXARa0ds+5R0KsjW0KmV9udmdOxao8/fvNFe/9BmrxuuWiBsaixyri/jdwDedM
+cB7TffpoCci2xcdW8nOrOZRrCasty8gC1/e9Q5i0jvxm2umIRYpnfaDW/7xnMHD
+u3OdZBPMQt18hxBI8JnSY+bn9o0rdEFf/WGZjzB2ieoMvET8JqMUx24BWv19+u8
nSp5wFxbImivYRlg6XMGVl9pCZD60HAQU7r3xIBF2SzzrmGJ8EaBGEPXIoglHVJ9
+MscZQ84XxDPgq6f3QHBGmirocEAuAzjUvGoOVNlLTt+8uotZZQKtPKLuq1h3T0s
NJA1k8j5kG9vbPLwBMzGraClgkVFF/bphHjMuytq5F3g9XnF6xEzSbTI2aPqJjz3
7atKVfbgmwENlqH8IbsC38P2fRbsbQYbF0pVQ9zS7r5BPrH2/c8yRFim/Pr/5gnm
9bd4gFTqTdHsLhbMnnfyOaOyHpYqHEFCvYQZRQ08zsZPktsC7ydPtHchTlAokb4k
VkVtfBWoaohL5WQkiuiVhHEHrUei8warLSKcj35UXGsu/fG0x/LvuFoIg9Hd9xYy
iH/len+IRxk6zakQnh2ia8mzB0+567GhuqOvB5jnw+9nAnnVym1M4OknHW19tKsU
qfu6VV4RFBlXVCgEHOUE83/65zj1kONWyaSSJhmqFlWG5OMAipi2r1aVGyILuLhO
iDuSJLCJNXLzhLqvkwQb2z5BbvgjN4O2X7JVHUxLqB8K9xhPvLGMdjTdiWIjYBXB
POgEwVlhzjPQHJIdrfjOzWVaQCtKL1ys2D/K37yOo3/VHw1nomEbHNFQKVhA4lHk
TS0lwEnAAvf5oxUtwCi8lhkMX1kDAujGUpsM7BHN7J06h9wlZg6CubkbjFZkDiSZ
4vEqyy5EYaVTUYHI/Pxs+QU6BkfsQNZnhb1qyFjyyL+PfB05zKCo/3/wvmRWPumT
2WVCyO6fJuPY5R+LcANRZUOs793oXmDn5bDFX6i9fVXcC8lhTAIrBiDgZz3ldxdQ
7EdTP1Rco2tBi7DdjQKBAPpIgppIdePxke94imQ3NAOkhFyOG17buxc159BKnC7E
9Wq51b/SLSQ83x8lbu2tT4X/AWRPUs2dl9BIAdw8Vjx0KCiB6CVGYspbbb9bKz0n
/mrYDIbEWoQh6rlDpbHY3PE8yeIb1lpN67La5GLuBTX+mpvHD728tdRamh08GXH4
KltEyRlW1QCdccBkUe+nB45Gkvlkw7wYMSj10xevPq0l5hGBcCPBUyZDQuzpxYsr
3qwIUs1ERnJK7wyhIlzC5sYA5YfB5aMUBL6dwvMSzB1LlJiMCXCpjKZ8swihlgG9
bawAKRZ3mcQlapR1aLveJUynS5O9uynkc4xd1y1jh2W89fDSW5uLKwYCT/lej9GT
tZdP6LysCDmE+Ai1gYS+Xx0zCHvjUFvFerRqzSLjbUkxP/9LeLsUHUNUPKc5qaAr
v7D+p7QSP20LJwzp+/xuIsrECLGv+PQRO0zB1+Fm1KqXKZkrXdm8DD14ubWaDJ/X
lhlCNTd5Zl8nYHn7YydFSBU7JvhflPQKwKxgKo1qa9nxckMdI9LePy60+9qZrGK+
3qsPw+WPZErfsY6W0+d2YNiH2BCwxHNCpYQBi62xLrbWMlGq82KzAh72bSMiNUiN
Fo/gw5MUerra7hPwbBPYMx/yg/+eFXC7ryEfP0xOt2Yux17QXhKSOg8cw05gnteP
PIzh/ZI7CalBVVvemKtPoycqmI/hmT3gfcG3XQO7NJrLqL/x8eOCtMWXev64i/sN
y9U+8bS2jS4hFUfQHc2jUIIrvPnCjjZ4v6xyD/fdMN/OGtyda7kpnXIrotCBBEok
RTIMi7svP5/va82IcpTflUI0sZ75v3kR18rkFSvqgPc0XaXlrU9OI9MVo1C5xFh0
keQ73ts9cOP8XeaX9mOP+p42HePSfmawItEGAq5DeuA9gy4y25AAvfp+y3nzcfvS
PKbP2Jlp/CpWn+/u0UnUJPsDg/h9qCXvVTyTgr1y+tZae0vYkINe4upePYj3rpNM
A3FiPtQsKrMSODaOKO2p27mLsijC2rC4yhmFy3VJy64oDhRDRrYknoHmwEriP+Es
oUzM6b1r7A/Xk+UDlLz++Spn+tqRGQ0NZ2AaPdoXEFMIFRKWq5g2q/p7mTqFtOPs
3QGaB7MgpIlRJRseJGzRcFb8KMsIoH8qR2NKM7A0ecL0vp11ZqgKolw0rHw6VHsY
rKMcnXL7GSFi3Y3JKZyacNTb+XjpYqkC4aycAmUppyxAdfi7LLwoP/ImJYL8MepP
pNomdpc++UBlEj2nF+bztHTQ3rWZ+a9j9HU69xkbhNMgs9j09iFyOJ5O782NoYKy
JpH3cs+3NSCBgVjUPmx3gYl5alvvKHHSjp16zF3uQNmMpmukFji278xBl67zP79b
NtXoGe6CagA88Fh2biOTi+6R5dQgG7wGw1E/dzmHb9YgGKJg+2WTQCs/+bxDznb+
EbstEvARsrqHI9fBKELZdDXhzesw5NuJvuKMsdIcn1wDjcZ+VZVVgiGTlWarxkvn
OmTJ15TRqIAllzcmyrpoJwWTcMuhnaFn2QPE9ym+MXPBVtJ1zqifiSb6bgvHn58O
QhiagPvy6Vc+upy3xYdIaWIHzfBWlkybQq05z3aVf6Qftbaz3Vrd2xBLh1yECmus
zeActQ4w9xKX/X+7jaYNPS2MkP10nvtKt/P523FUBaEBpQrcN4CjNv53aqrro/gL
nhYPVftD7VVlSUjMjB3MR6Lw1LLFzF+nGobh0Q1W7a4Wq9kxkpTtRfGTJPb+gxth
CdJcLVBZLTKwiGB5CmfroOOFEaWmXLQM3a/qYNQC0yEO5eH5lnKin0pUpYjX4IHH
cpo3Ff2WqvwNPLrYDN6yRyD+uJU9bPxMSexXv272gYl28rosz9a6yPWDf/8ZkqBl
OIUfjZqU/L2PnTK1yGheXxvjoJ09UhZ4MP6kJpAo2WKwqU3PXbkQRiF6tQqgBH3d
sLsmameEATz80+Zu0NRkKHBrXlBy1u4dOoUdzzGSiVSz2ePkC8rdAbdUIpY5eHse
/mhhkaY8Nr8cepSiFwx5PkOOF7SH+5nnl4KqXm5gLX1aHJmLe1CyVJhwpXdoSFog
ybfuugBLMVTTRAcAedgSkGwqNDcF4vDOHFj2/FzPF0hk5zqvmwUtt0BThzUNuemw
mTCtIroWI4Cs5z8z6nkWixi3zSAhKAKTyhCjdEIxR7A5wCNYBd5JM1wgy9kAVpKt
E7/rTxZmpdRxDlLhVpY6WSO2Gznz9qMcdhpF732stNuKBVWInWbpNMMAlky8BUMm
Y9bRPCC601pvaNT/HPwfoi4xPt1TNVts2f9ZjivK5aQcaoPnwUQ0TtrAJ9qkahlh
YsclyooqrD3p8k73G1tiFDjYdTVQ8RKvzv1KivA2gVrN9kAlQV3AINxX9SisnG9a
xtNiy90F/3I9qjZ/R28Y+y6JfPq6pGMxOum3VeOhQcUBjja+PeC84r6l1j0r0Hlq
DFKaN9j4xI9zLAFKVsA3sNpvuidxnio+bMjpe0UqmLziiuxOEy6+XRAJiGbI+P2x
pjUFG2555P1bQkHUGGzRRZOpJ+QRApbSaQKYjXJHIrS0rg4nHSHrFb+qwdaLQzGG
Ln1A01NMFd2A9xghvOc65aTcDLaI5sdCh4JrQYlvW/S1tBOAea0sbTeoJu/At3Ym
dPXi1WIafJc092x1yzDE00gyY3XMlYeqF7BfxbAjXYINEpeVRapGAv7xrAXHXSbC
msletydH4b3XUDPP9hnc1rDbFePT7tbp33hD8m+kieP4qJlk80BI2XRcT+zsJ3Rf
HZEPXrZ4aIzw1YQOz6k1T3vpNPZnJsGpYC6kIa3jPP08+3k1I+yp+TTeaBHco5kC
YcLPz3t0CzlHF6nKYWtddO3H1v5UMuH3RawQ9qGKuC6/MGjpFR961XeAoD8NpTXR
6qwQ455fLTshoPztFbHJrJiHdFCYVFLs2fJ72dnOJF7Y84XRLU2lfNWcyAft9EWW
eXlRLxv5TMw3lLK/nttp/fYfNzEwBOvuCf47ztgEo3m044gj8x50SoAVWRGXj8Nn
idJknjxLXkDmydopHAWiOkKhkSMPGjD3OCYoJyOqCRPKDZmiOKuftzgH3oq4+nX+
qYm3ARBf5aloc9CD3jU+BC4DgjWv3I9qifguKbVKSaa2NCswHMfHxwq6F4GJ7AZU
y/As83ktdddNUc8DU0XLLIqhGpv7njaJilxK/PfNEGMCD45nLkchN9mfvoTRkY8t
iUgazeGL07ZG8tU+stxxL8zTcZym2lpdwaD6ek4x2JSPlYQYowTQTVNman5DrcDT
QR77A3lUi85N+nHZH0lfDwDQ9d2uQGl8pwDq9xJm++xymvEMaRKalwlVe5YxvyHv
FeUKHpBxG415Ros4DQLqGIndY3o5Uo2YY6gDq19Qh3EUGnXS0M/wS9o4Fx3fBEix
oYq2CZOO9faJTwOuajCb7WTAF0m7zoZ8aj1OuT93XER6rhvhsd/VY7+mKhgEwJls
jbzwC3+sOiha0WxNZKPgWgWFXVt8StURs72lu0t8AeZEofMNMFBj1jGN6tumNmSJ
R8DF17cdERdihc7tiligGYNmHGVPiRDJr1Pc2YeOrxnu7hdngAkMG20pKTFRhKcv
FJgIc1ReUP1ruQl7bNptqV2mYir3WN2UfU0gR1cgc9nNsYwhe7Hhl/aXGC5Gc+yE
d3xObWm+CSSzypxxoDQw67COBVP+0/bTjGsDwCo9aoX1ZawLfP86BTavpJ99w/PW
XRztELaUsGUnCSRpcGju4EjMe+feroBtI3jcBpnD1gwFcHQuvTA4XGI1x6NtRo3A
E77PwgURrnfsJea+X03FtbB21z2+krUsYqpeCuURtb9XowZp8Gs4f+WTY47Xa5Ak
Cj6hAHkvqPUBBoHRIgUqB4SmlVM0YCm+Jr+a/gdtoyJhEHgFWmsEgNJQFcUAbR56
CwS3JTVOuRXgNe3L159C0t2ubdf5PkBzBZAScfNev2eFKIXb4ey1ZqjgpKVajnr1
2mNFtc2wUU/SY33AOfW6ysw+5gB+dxOkwwY6dmgZfYSHk8JMMxAoBesC5u+Nvx3Z
a0wyPq8XmQIzCKT8OEEz/lUJhiaB9Q9Dl+f0KQsjgQk3rNdT1Ozn6HkrdJWX189n
aHIpzvLBS95PiDgP3TV/AMUfd3rdPDvQRKOb9MN6b03T6PWVwGuKXJ5RhtWc46f4
7cA49HEP4mHHQyhQiaOTcFj7AThfnRvYNoFVN76PEanqLFzrbG/WPHSmT/vQod70
6HylNgUoXgMP/FdiALVb0/3H2xr7hQlnhDfu6KpxP7+jIaGdpGWuyJoLi4o8cAei
q9RZaeEbK2QcXVCkM8bbm7MEM1UJMdYRG6+Z0jbciy3QoD2bNXZB7f1dvBTZb0ST
49OxLaqUjf+Qh9eaaoo7kGGiipkTDkiUhkRToGYheirbU0SZljXybKfWbK9g3wKR
ODMgmqgtJbHKXu9XEGFRk2qd4KJ7m2GCKLRv56Vjwpyam8H7+CjUDiYgEid/xP4j
v9GIvRNTeuSJzp3b/XTYByigQ+3wKZdqQgfEaF1MTNIICVR2ASqm1ykMqBLu0ksm
AoRE/NUknyhMwpIk6KOoCe9irM0+j47d9hWe/tLgyeq3CDr+PSQxYti0uod0zI56
LO7rZXuSLoE2+CX3UL+JGD5LEe58c8d0xqfI2bHIpsV/9HLIFZLyD2yamiG/jXxY
1/Pj1aaVpouN5f2mQk4LSRn9ZHmNHUxE4sFZoJI8htspr20hXdBUGZ3xFzdlvcnf
d10RWFhf2rR1krs6pI9C/5G4ERQbxcqPhDwIZU10sPApUCUYoqF2/hIaoBbkrNlm
ZN/d53Ag/KyD4afXNhtBXoZWgp5B+CP4cdr9HEhnq2X3LBfW7m568/UbuiqhWEEk
p7GtCnaj8eIegx/N8ScT+rSrWCx2J/ysaRK2BOP/erpv95jdWKqHR2x3dDnTCB2F
VF0RVoCNS+0jMixC49sTGnL3lS+2rTe6uDd3H5+BnsnqAlpAwk/7tMHAvmi9TaDA
OmHeeHaWNL9JTst0A3FbAf+rVYd28C10XqbD0BTCPFBh3UNnlcNldAzuIYk6++a+
nozzv5LstggbUVlZkufNYlPnWQc5omkVPGx8MI9QiobEDIS4Y4jonBzS0Z4ax6I+
y4T0fYRk37YvVdWcjSjw3iiT/wXp22QnM/OFQ1FtO6uQjsnVI6R9DV1hZqWVPif2
zXH5s0UKyGasj2T52IS5Lgfq5vZKyfJv3RO/yxufKu+yA4pg9SRzVYrtaXbO4w93
Ew+2r3soDzb2bMu4mOPFeHmMF0g9RUEJ/1TqhalvG2vAJCRKijQ9W2C+5/HRPgy5
Uy8dodApelBh/izmpYlmyu9SQn5ApDHZGdFNH/yOEhr6UmkL99w/Hm1n9TnmPx3E
YgU20RyHs2mOVv74oq73ruo90YZ7qk5A+6jvi1BiobAeUB3sEsep51e2CeOY+HMt
I4hk3km4LX37gWWnIwkiXb2hhG2R6p+sziEPTJscEwODlwvsEQ2DhthH9ijXfsHj
iCBAMYNf6b0xkt4gY/NWVAYe4zEzESeZuRBsCZBvtmDRM35WhFUsF0yt6iCoUdPv
KnycrXqOa6YAQexgCzIP1V0TvlPbQDc3zEHc39gsxsBH1XOodKi7Mx2UQ01JxMQ6
Dfog0GzLKejn4KT41XPKhWCSmp8NunAoPlxDw+l4iJnT6xb5KPe0UGBiXtbeczkQ
Kuuru1BgQ1LJ+RJpIo5X8VGwGsjnPe5bIKYW8UM60aEbSTJ8yhoSh87eeq24O5+N
qdV+/Wpcaa7dSJYYBNbsZ5/IrrNzUVi3HHQeSXwtXZe9fpYehERfe3MMnf2BqRfo
+WIRuRuWat6NIUAOmARbdp+LbUXo2stBpIPXyNjHxlPt86RGUqmxP/jNva7lTRa7
lMUUHpVnvS55ENBM+OmyR/OUNR6ga4FfMqHg4KoltL8p05+cTqIsueB2QiZGp05a
paRCqIhHju94+GbBLuRjFABZzff7Pewm3wV9WRMpAoGYwtOY/MUjxflApZLh3f4C
8P74tYNJrtCdsPNLlAkNtl99oLVap88eoDFkkvTuO8g6kmLTLHOyoKQ6N4NQTCQA
uCzLIA6wfp10HXppeQRELGU58jVJ3ndifKkuXwPeAcK3Oe6OFKEphytbKCg0sijo
ZoZnMfqtHDhynrM0Doe1v3KlIi2i4LCLi1BB8lfDJkAPwtTQgxZpeFTPcbDK9kny
+0yR+DG6sH008rBi6i5r3a/FLaJXDJV9Dbcj3EMfRYxzrdMWY1jhRtV1Xp2rnsBh
s26Dm2uiC4FbCgAZo1PdmXuBgOwgIvduoK4w5QOSfqrf7yvOTq4MBJKiW1D1aYod
xNa3MXRCZPY0VFq05i3XLc0fsxgr18P0dVE/tx+F/0/D0J9kLZi1hRoV4oOkVp+T
PWgbDkWn/upDuXx4qsNOfez+HDvMOpZolkYjWe69qefQAyfPdWtSdw3boS6yZaOL
aYTX/OJAKoAXAAE4ppKhKkwPEr3t4BClTXbJieHslfJo4p1QvWRvcwXbVNt7kZml
7kgdMLhkGPhSeXAnIWmr0WODi3uB/XXfhFistpTdldH4qFQwUUqA01bFKJxnv2CG
M2Z9gvA2989lJm6yDb6PCwgI1/FU3mi/IE1sT5Y15FdnhzL4hxlJ3pamS6yhbdEV
3p9Q/R7Qg7v68C6ZA4j/EkaFPM64AAAuQoN7HontSgRKHZxEOE/oRI6hCzv/BVns
0ZPdB+zkB6+Z6/WvN6tWSf6Sidv7ByUQ2AedCIM0IicoimDadWfXeITdotZUZzQD
ArUUr4TVvwDwkNvQj5AklturNXJKPMFeX1+rLyxDXN0+W6PXTDpbGeXtfR/ILFnl
MODe0S58MHlRe7T23EgZxeGpYWeQJay3Qc404Co9BwT8ynK5stbugXFe6PEpbeH9
JSxaVdZogHxuDNVlKOYnQWCpn2hszsZZxgXEObF5KC0hSsTfkJ2qjWBhW2x+FcuZ
zqwCV4Cg9zMjjjAXmKvDr3M+ABtMxmFXmwXGPRE4CEU+m2SoJDdZdeNuPsg9NXUI
NaAGEDRSoup2RBkBlvhky904maL0U7a/VObsQrHtB6Br5TMYYRgma9LfkrmpuSZ2
i6QmVNpW3NtIPVKCo5lbOyd6xY5HO3EhhyiWpmBAFs1VkQdi5WXcIRUgCIADOssG
lWXy1MAbxTTpFmxzRtNhSNY3nOLGN64/gtCugwFBtiL740woetRIbWqeF7poIdvU
zGWR9AVCBktyOCEXHcedjXRZhteG1Qfu0E8HXgNvCY8ezZhoCnZA8YX6J4y6uI0a
PAxkw7Isv7tcLGFoM0vXrdwXm5iHG9aRG1WVXn650J3Ouz+u/ywK55m9NjQ8cUUS
La+fqXA5/36p5aCqe+A5nAKd44aMPuHsSWnsXSTA1obkutYTfTXtEwpRe7JBprSO
Q9EC7QyN+lFBIPaPMQPQ9IxkqjShk/JhOmybCu6SmTa3tNTnmfbi+PuwnxNzVtda
GD9dOVj/3I1x0bVP/LK+Pdyy4T8oAhxStsZtgBCUotqNdFMLH+KBdsEwx2EZ4sGF
bJYbQBMrp1qCmiphKBfX0s2rgrVnDEjsnERUFVoPqgeMBhGA/Si8wH74sx3cQao+
xrNOc3E4BZTh0LuVkgUpfB3lnRMMrJ3f6VetVoovxYL4EnRTYM00kBkaG5VRY9vg
aIK+U3SsrTExwoUo9je/Ul53K0enGDC23havAw1yxgL5+GvR6fK7/3eHuDN1UMJZ
EmKdiPm92J9mrOgrER3KGak3UjlJ9FvvCFk1bdrhIN1VQQKIeRPeu5vA1WHr9RiZ
UyCiQ1ufHRlA28F2xuwVaSyy55FpghdZ1scPhp+CcH69PH1/5hf0B5mVVjsnKIvG
VMvP5YwEVsxIjAEsP+I/h1GETEKE5UHk4gc+4wKm/Mv3hPVv+fHEbZ9+IoCD2PhD
VLBWdvcsdfqbwMKMIffFSeIXoOj8FgVWDHqxbJU3lKf3XZY4yIeGs7cskrhhRgbj
5reOJ3T3UZaIC54SwwLgdahqA6Qj5v1b+kUj8qXB8p/uKrhzvJEFIG4aHB4f+tUh
4MhtmAq2KWYjyseJfvHC7kTXy8kMhjE50kBrnbZwznw2RvISMIkY9vCfWUHPvKJE
yD1vLfKxl/SYQyqxbiCtShM+U+QQMQ7+0Kb4HjU2OWh6dQNBqm2HJ3VhMV8fk97O
nnBOAyNqX1N2fmQdnWAPmGFvQ+jrm7d+txYr6UVZbS2PgdoNVZV+zlIwh4YdjdN4
41Wxq09xATOJJbDSw49xO0/PEnqoE7bQBHJnCktm9UO8c+ls5O0wJcIl2b3B+ekO
uU+sPS963LQnM7GJwKHqTcugaTGETwGeBRdTZ/XYomzwi49qTij4waEKWZEA0Wmb
eJEWrnq/4TEqiH3iRGpndDXRWh7GfPnCL/6+hSvxnGcE1WOk5lrVl91SuATP9BB7
yyjgPaCroYXNspIb83/JupiJPCKNrs5N8LrHhJIPD8AWpx93QEGZGSM33a3lrgh4
es3hCgI0yKmQ8I9iQ7i5TpX6uQRh7En3GioKff+sK+EZqIwpwPq8tj4cau1OD5VK
0oPPnxteGE6gsqqAFM+BGWbShTZd33Q1QyHzuAakuxp4WsjEMz7llmTuhfPrEKDr
q8fYnw938FLuGlnUciWF0EDm4Z1prISpZ1qrcd4lysy9NlB4UeFeEu+7joV2yh0L
zuUwV+8F+fXWtNsgPQ0ZA7p8J2kqjfjxveR4eFAMh3CBIeF49YO5WLpg4tHWCKep
dbPX5jQDngCa9roAhnZCbjOkaUjswca3m1hFz28DI6W0lLGAu5qb9lYI+Ok66N6J
8yDZgMnaFUJzeGHDDDQ9aG1XIgU36aX0owiiPprVdQwMr6cHdaWJ8MXGlzJFVVKf
RZ/R1L6ixw7vBzJAW5WrAL5mpxWGF5HswfhV769jrgLQfAgaWd2ZpsGqhS8up6FW
dzaLzfqRrSqKdsTDrcSk059zot37fyYv6DFErdc5CUJgHv3WFEefVseX4HP8MVbU
KjgaMJXKaUJYk8KIU/1c0uKQ7HVOr1FNtGCKBkTDBDaitE/hIEDS8F8tiNOef4bH
qzC5dJN+el4vVN6kqdRuDMUtQ0ZwuY+H7DlLI1ONMDMZZF5a1thaEl/aIBlFLn7K
n2yoRmwWW5/nNO0DGR5rK9S1qMHm0QcujYrdOuHS1hdVwGJSif/ZjCeqj0vaRifV
G/Ws4NNT9lT9zy1ISJAReuoliFEZv8TytoDvdUKX4LbT8+Gh5Y3jvpZjVRJTuHXe
LE2vdNGOYDtTlNBB1u2uQfBO/YWCowDIUktZYvGntmK6j1yrlGeDZ3bZ7i2P8hRf
5HG7fF3gMKHJm4qPA8l2Lv7Kkqs3WQWS+a8IJw6mmA0jJacB5GlnDBmFgdFqkY1M
q8vZSQb73iiXKYrpyPzPiT6EyvEsdmF2DT16cDDOzE9wCr8eN5unvwhQNcItdcss
lEgNvynwAgAjzkQsldbrCxY/VcswlA/oNetVycCMzYiA36usajvc2o4iAp27aulV
4erYH4fSRZyNq2whBK2oG7NOxqTwOaPH6Lii1xm7+We7Ws4FGVeexMoBwfUGpTEd
LigG4i+gal3ly8Q68NkwNTbZtqjOSz4/o2gjeoWGTXcP05zVat84D8FrxNIVm4ZM
B0JWHJnFB8JJ0JnL+jUlF/OdosYky3R3TtCtVH+b7Qg7vBo1qge1/jiUYlDrJ1J2
zgK4S/YzrxiGrKL3y7xkoHHtJ4hamG9RsBMZrOtL0E3Ytpr/RFWImsruD5HzdNqx
jHuaf5Ng5ZJxUS1gd9snxGppypYJkj5wAS84ewmGIWFCQj1kdSfTXJtDea2j9Nr7
N/rq6oM/h4g8J/Kjo29fPZKlQJDL7fEsgeZeccucaM6IUuWqwtS7ecpm7CcwvbNg
F1u1mbQmf9vbCNqfQMPJhi7/e89KP1LUfDCGxk077f0O285qoBn0ByPFOtbKzJ68
kbN5x+mtmfb7bsedZmrIbNC/g25/9HPcHnvZvmWvnSCSYjgDaqNUbGwo0VpB8xZs
Fa96UHOH/+rolsoZuVl5AE6j/fzhiO2xfjenky7o4SJsU3zVodMfRUOzINj3tBB8
YqTP4B/+0WAVbXQOAt6QYzF1F7fdGnIpklV5xsh9CzkOe0amQZjHvz1FyGAlW5rY
jY65Bp1v7XLwRZYHl0HAR/H2HiIjWH2h4KHKIPG1iFrRWwPBQ9/aJLhf5ATSfIvF
aV9nq7Bed5NjpeWyo4uBhmd1RClb3GY7qbHAQ4NuSByFsTbSY0rPpLgoSEZDp0t7
ZCH3XNYZbUu/+ijq4fdb7hytdnVvwpjSHGPgUCO/i0LrlZz8qsirisqf6b7AfLzo
/3UDxcrjUG7N5U5gAvZoODCppjuDWJzUPcMcXTcMDpG6QyyZo5+9JtKweNIcRFwP
Af7LywEYOxig1Xf4TgBVywuUiolGs0UV58D4oXqKWbzQbVZ3nr/fSKdzdTsBkE6u
3V2Kk0jZ2BefsXaIJ43EhoTi5DehG95wVkIT3fNfPt+Jgh1kcUSlY8VkWgM0mvb0
YoZWjTYgzCM/UxpSpJ3y3duBS1hvE89x7p2djzxNkL8JN0TAW6zITCUrigeCv40R
T691hkwxODJKvXYQvZHrQF14+JroO3+ZpgtMWeJrEjmNBsZqh/hc4SzjcUxRY2Iy
Zvi5XRobV0dLbWsyq08WzfX874m7DKjRYq49RSHVL5/u/bli34Oh/pccXHuqBWdl
F1vIOusMQQVjVDTXoKEEnzx1oYk7vQg2UYKGXcjRRkZTp9i9rEaCT0F6WBQTp9ml
p66AW9sbCrZUr6mkzIG1MnR8TzxcWOtpibdSs92Zl1L8xNmRjKggEUMBgQ9rsV5H
J7CEwvShhvajMuMZuEsVCW2PRBxLf8SbeEAU4qIGC0qdmQ16Zo/b2mdgUrItGQAw
vCHtLuYOFb/++jjwcAHP2RSUpdX6f+zInIHFm8HrH3upYNQm1yTuAFVK5E2EYk+L
MxzNeiEgX4k0bcwcpTfLGt1BPhJXdQnOG7b044IZmxc4yb8UOdTt0fWS+lxgPz5O
KQd3NF5cU3efIZkR1eoGkJPqVG9Ia/CXT6/lLVLoti4PVtOQn62ScT3QvUSctcgQ
waV6We1PFo3G0lNeCXLiXXXS9pDT1sW+KWiFd15DFc/YHKlFtYz2L8xSn0k1Xp7F
94secagUiaRgJkF0kZXA7mYCr6smgFiGBcCOqDAWaH9qNZUA89mKOcnQLYT6+jZF
wzoFroojAwAir1e52pXVoQwIyUMBBR6JQ/IYkrgomLfs7EXHybHmG+lBCOg+MPuU
kxPO6MZhKqZFNcb9FSVBQJyirSWjYfaIvunXk+uQ0UdZZLBO2HpGldU5Q5piwMuk
OPXfoLE8gRRgBvPp1buYLpB8qsQs1KqdJcy2EnUQIkUgKfrd6t0i62NqvGsiAY9D
fApzDzWtzdGPrx+rXsPI8xRa54ER00Xs+11EhNoDMrsrW6FFn4roGQ7eUq3AmdNZ
QJxGbJA4G4s9V+5KJJl7pBE0CuUHswzysqmlxAdeQijeHY8+euAhdCyUSDS9RY5C
AZ4akxqN6SSwwA0K00GExoseXJoZOf5fJ0WkOFBs2E+He/gkUNkNRWn6BYWZFFgh
6f7+zwDRoox+ajwyIute8a4NaV1YLq7ohBbg3f9GlGviSkvGErzXu8u7d25LzVkF
kthz1R0FfZWasjEgNNBZ9eZcaGQ2GDFvDC88EuK1d4Tqsp+uWchUjtNMNmzqQ3Qt
Hzd5dmzONRWcRae3uvpmGBMC9tTVfQPqFCtw4bbOBpnMKAzQ9ylZKZmuUPchd3Q0
NwSJ0fFvTPfiQVP9bLDvHL/54rVjLKmnOBaWfggQngR/Mwwa51z4aDZFssHJCdTH
b9u4CyNxfp40bxisokS97l0O4d/7icXJv7McqJLBTXrkCkoVizNgEqeVYOzXArw0
7VgMjHK7eQILa5FVc046Tj3z+yKStypzaYRhwCKhy/d1OD0+RvlCvPoHKzOYPSmT
i4Iu1Tlg0YA69LcqdiG/xDOhshceJTx3IKoFEBqArpv3j9pSiQVm2iNeew2fFAMo
Va0vRFVyFX6FHb6UPTcGcSgTJDn9zvNKVG/qx5eXEjeMklfItYfijx4dwe8yzMU6
DXXXfjbNDvL1mI4JB011NR1YKinIBtD56hENIbJcgBKikTX+DRmfdb7yoL754OxR
HTp/wgjH+Cik5G6Cza1llxlYCw/00fvNhX62Zo5a0X+4GWmT4bM6CX0LoEn318Up
xXvq+Ij5pLU2xguYWs2C1DQhCbUbZKXaRfoCyK7z3/+c5eSn/18UWcfrtSgUKcN+
iXOVyM4aljQNFbFdX2WqnhvtLXJlcj7EUgbZN/g7PDTX0SIq/pD1OFEvkMSgDO3q
fZW40VCC9tqnaqsWN7r5RypGJeXh78Wx/SQZwnox3+WLgmTwOnBJGwYQNhQ2cUPP
NNYRwMtyxpih3O1idhHhr4xlWfcmVDNv9/rE2qaqO2Ewi3TFjklYorOHyJN1j2ec
fmIrPDNZwIXdfGFkCQ4NIyUOPjO6Q7pOLulKGIXTRIPrC1CyKCV5hc4WdJZ9HXkT
6cn94SjGV+7khxG8QsCLIvJ3RKcb/Ci4M62qKwqhOgmTmvfWm++RCi3qq4rTRyDA
rDfxsY+FR8zJ0CusoMbUc2RxjnzMlMNGWho32WGxm0gv/bBalOBuX8ez3GXCmOiF
RZfxjmjQSKnES7Mx/vNdj+4sPB5Cxm0Fnmk/KuI+fCQxHLlVoRY/VAVIYWz8e7/h
FKupQSWaXiK6uxLDCNxz5b4I0YBlgssnpCViF3B7ccyTxr1rVvDcPaSG0O+WgTi5
6dg3cyJPksOTL+s+ZjvibMmy17BDbGJhHo/m+fcxvAJ3Wkju73lQNlsewT2Wlzy7
ANuLguqcNDOXVKDwYFeVF0AgAHgYb9+PwlaG+UGZOWLv82sMWwUCeo8Fs9Ocoona
ga2rYkpNK3Yn3uEC2ODrjYITRt+goBeR/xD3gYxrW3lhjUsebhIeMIbc7qnp/I+A
W3gTnR48ivUtZZS/YJQjuWH6Hvyit/QSVC+ziVA83r6xWtLe7jbyi/ljiN4+F/7e
ktQPFV7qB85OQ4KzpMwS6ctn3J8T9NsgA9wPeFQe80O8oG3vAilpARJzK64WFjn8
vJVYxTWIm5JozWX1Lt0U+cNWf8t3X8EtdyDf3JACRemkjguCKKoysmP39fRqIciI
vUgL0YHtt8W0mGMsgPifxcIYsYYaFqdPyOcOoyGyAUHm95Z9xMie9QhL7UnBytt+
z9Ak1OnyRWzMu4VB09cStnreHXkeHn1branvieH6GBTquvMf58ZcLeW/S7qdL4hV
4yxdjqJ1In/9YeOL8nzgr7KfJwLdqkMq877LKsGP7+VWg96eCCYFJS54vCBe1n9j
QFR3SpCeBKM72LVC5ZaIODQ4Ftd3Eo1MakRfzoVIRLKakf1mXcfJYAigUdkoe06m
tpbMuaKJeHN2l8BoYro+OHvyJUkhXxGxaXdbrDCIvLW/118qFU1af8hD4q0wFX7C
KZrMRi/S6zs3r0+DXUOkfB7OTA9foHVD+GjKRkM/R7F0rdQKp8H9kU0YgOfzfgN+
Qy9xQWSq/8KQVr/ird11xtV0vx2oMqdx1q4fyahHc3znYwH+q0jRaxDY9sDWnZEB
8nldUMpOZGf1aU63/b131k1ILF4gucSvLvNDAZL2MNTE6hVfDgI+MesM+hwaMoFA
ZUY8vVcVP1uMTFA7beM/hf7EI6/FKrh7I/gCnrlfX6lTu6g1On0W91en+jz/yho3
CIoRcBiME5JG0QJjpia71pjfTKwSoHQvewSi52h+99y40zRjZnoeOe/fqmMfSU2J
1McsOl/Xs1BMlhGBY3UhQiy1jw6G338JN+I0plMf7UwpX06X4pBjgcMkWI8BAdRW
zcBr1VV0sfp4DddczVRBX2lIWrY1g370eT5pfHxhGMwPI4y+5zQyqqKuaKsGBAnS
jijtlPkI9TfB5Oobn/wZPYqrkkffX6GHEqYB4AFBuWKVN0GvksEH67H32GWDAGmO
DBMxvDFOXEUCYTEg3F6jwEDVbeCPHqdCfpmqDn2u9SIymWDYUpHZB2ZXWnRpo9c0
xVI6jWyVyRe7cGG1PjscagD6MFpyftUsH8gT4y7/0KmsMZbqlxBQlsUnPStiaZ6R
KxtrLC87SATG6tKg6yCgBJmbuj0EZ7cttHEUoLBjcTWUir6yP1VcL8PQhaDBUUg9
xUQ8w201Wh+r2yoexA6F8hUJo2R1BTXxKaJ2qbcEA3TRS5iMSdKT1toS4maDTgva
Jl+jHlmtcqP1ET9QdkMViX4d+TbyVtApBX2OrXi2C2aXKhEP7WlIgw5CLjAySo13
8dnhaVef7u1XdxlEuz+FBNXPaH9P533ILBuFXY8oaeIW09nx7bfNty9szA3NRaK3
hyT2mVN8EU5KVqTUN52qYgm94ncXJ16+LoMETDsFVYqcgs4vCmhuxBgt5eiGchns
z9rCckQ86g9ToYGc2qBmKKhvLRJwfnO6koAlrYrVJfpu5l2S3FvnRD9kWDz0N69m
F6720cv0/OqlGZc8RAkQS+jwYTp+3LQ7EinMLdnGLTg8NcDGwRWaeef4igGXpmfR
SPmJHDV/IagidXig0yI9hgcbXNyKxszVi91f5lJu+WQXtwfFm52xRX+DUzexGoqM
zzdAR1WUwV2q59PzHaPzuN2MatqLeqN8D8jgwAczLcBeYxtYMxqNYUi1pPWHbEar
IQkAxsWOjAvfgUuGRW9BGoqof4hFHe8S5W+/CL5qbiKvEqvAzTy434XEzATDWHgr
ywocrjfgidrwrp0iP8jxqCweBJr3t3uA4yHojZctDUMCMw06pT1xZ6oK2awn/k5f
XmnK0WphtTcD8mTpkdG/ENTxSlCnZC8+KI66ESZLvKjYrEwIizUD2vw7KYwacxdV
QynN+22G39b7i5ngW9ASdd7RY8sQraKwFhZg7zN6Q4kpDZEX+97qtVW9gDllWGul
O4BXSK6rW38g+67Z4LEA8wdBLXCmWq+kj1Tt5JwSoslsRV6df0T6mtaWbXVQBZao
h47ED2x19I78ZbPnLM9N/XnaygAIgjegxwlpDsnkr5J2LDvje0wd+rq2MV1VPD4w
yU5oEXdcpV54LoRzRSrXQiAXW/bbA+PjwwHomTYtgCA2+tvC7+fWWbGJpFsjmSFJ
+rXwA8pSR+SBlDN9RHZAjoBCI865olPLd1OnfXIZwedaXeiUIh9IZ44qneSPsir/
Lr6lKV+liRBPYJNu46ozCfsjnK5T3mF3ugnRW0KZXah9891f6tdHqaED7yPH1ONA
DjoIGeuEib+O+c2WP98DZoacrZZrg3+Pe0UQ/me+OHEuf+gjwHy0mm08bWFe7fz8
rxMWx+/TBXmB+0a3vnnynT04XcgXg/XZLA5cx6NrxvqsiZD5QxXtnSBwIxzae080
ERgoEcAxEN7Bjeo1mBWU+6Iw2JG60O6cfIFlN0+elJFdJ/mipo2Sr8uvUr3JZqme
s47yEGaIwnNCOhUalOyl7eIK8eTL0ismn8bU6inR3T6jgritgGjRPWazo0Ej4lpA
01dCF6gN0hM/iKg9q6ZB8qiBCrSXazoqI2BvAAtUYBBpAjUqHqHKtEZVKow1PC6f
oAEFraXzTv29Lp4S8vELVzYfvtjk41xL2cVM7yabalYO07AU3JOedqOfHBYw0eJe
QhCW1cwvGZtQyL1SlGnvmy/E4arhgIIji4BIrG/pBLpuQAT4tZ19wHCHsn+7WYAg
Vbns4ln2t1MqKJPKVkqMCNaeEqL9SeCG44EXylYTXNk2lLTMBaCc0BbfRtNsF/5U
2CzjgaHukDPP5gbci8GLCkD4CDLD7ZPpFKOD4rLVjYCZqFLdaeUri6YDexgzo5G3
CObw5Xa0zkYLUHMzavGwSr5rVJbabHMNnJ3AtiWOO8taI2xEALcstOjMghFLvpkW
CligOfNRVlHfm/xKv/2sNYOP40xsDKkzCDmos76Y0ETwrFDZNiitJNR0b51NCEup
jzM0h2v6/5QVLFApLHeMJNPsAnVENmVCcBFrTYDO3UtoLHsC3d/J+++7DX6PsGTv
40saBvaQZ7mELISHpq0Bc3naK8BEm/yWo6F3jEHyBCTsykN6W9jKd3tnB5X44e3g
Is6xJdEeOQPFbIHoceoIZBDj/4eTCKBWp1NwPWN9DOfJuhCsJrSjrNjJ01gUeJC9
YimXUWBeOr4hXzjDQe5XM14OasqYYKkqQFOrDgkxT1K6ZJkPY4TXO8X0drI3rGBb
R/yCrFWpraEQ55QDovPxjzSmVCFd1LqEuo5C+8iNEZseDBfHRSa0Y7mGmyBd9cCH
wmjudNrJ40cIv/jWvQo34MHF8JbMyTqqwXQCkDCbYSz2sbvw30XCIEcSxuIfg0S9
YKMN5sNAhGAi3rZW64ysQzaIBuD2WBkjaLPiLzp2yeZw+gYXw2BGYHqBXLXvPg6N
ZTqNczz6dmBMuzq4Z6E+Sk5R2DXIIQKOQ8a1cR4wEgcEcyr+X7ky79r3Ac6CTrr0
HgJhjGvO0iVhpMDyDJU38zDXBo+nT/PR64vXhvEfLMTZrFuodAoCCYvCrwPvwlYx
N1vao/JGy9Kv4sd4ikBqqmXnhFKvpRN4GEW93PbBwfoF1K1po4H6HMbGkYHcCY+B
2PF6lGksgzmoIbhbtasLaGI9JYdS4tom92bR2abKzLbL0Dm7Uq9jjsZRoM5UbHYS
yjTh3ZmCFPkDZcM1DyoYrWHNCqdY+oOP3sfVPyHre+ExIp0itTr0vLU0k0MrUnXi
16eVhmXATlLUPExlfiJJSnOLaB2SJuk+61E538yz8PLKvxipqCL2d2DPgHDdke0t
eGEBnO1GFLPAQJGMeTjQxhdw9rqDDvAgOgoW5oAncsYKz1Ti/xouWixKlpnxo1gB
9WVI43fIwZXvWaVgOvpScih0ypkQsilVjLp9XE7U280c2XF8G3DethCC8ZoURBEY
NrsSHNJCnrL5LgL9+QSkevlaL9y42KPsbeM7zgk53NW+eD6oy170l1EL2qwEm3cI
qm4BVdax96bfKCcOaaDFqxtfnwAlVFZkmq7oVd86JnplqAAP2IcczYYrXy8ArHxQ
1h+1rCtJHXhgbvwMSBkJkpdMd9NL7Y5TgjLu24X2HLqRtYbAT8L4+bOrtSSgKMzr
msDFga3rwKR/nkxdlyf7tLD7g5c0h6YMtqdiwMUJlye1j3x/AF8xzosX386pdSiZ
Y9F0vkIwk9MmF9Qe4tGTqQ67DFpaEg3HF7Q/JQdahHSjr4PRT97QwAJQZtskGSDZ
+L7ZntIQPHTubiAg7Oax2dxYhYJ4lXgXGUQ0FU/bWJjT19H08hN277vpXirFflIU
yoCi3EVx+J99O7BONaiT098IkPnZ8Jq56vHho9+Ev1ATa9rtJOBfTMK/hwu62TsY
A3DZr2dnuYCPPZrvXHxOiFkFy26HYz2V/jeecrUPKWXiB3DtDbac37aIJOqZSR7P
w6E9gXqmPwT2ryacpjLedThIs4/H/+YxnAKN2aF5BNPTbVsBF1IAZ5iXpNAWz5X0
YHKvhSzkwq0p3+exHwE+6rybqdtj3vV4fNh/etvzQ2ZT3W3hIL0Pw6d0+2BGEeJw
9SrJe1lgdvGf+g+i2EbR5O6V9EDXrqv8PbO26uwWHC+0s9TLXcA2HpdBh8/5mUB4
wGDVsYJ1SJwh50pw9rDkUR43AXXsMvoe+V1OZvI3Gd1dIJnhXh5NctOK8fWQS//Y
tIlOTGdKhsxgUaVWCCvDzwNBbSCUJxapCybnDZl8zmjzYulxQyRuknBGwT5C85nr
FqlyftziAx1fMFfKWGgp/5IOiYEQ0rfWJDOH1Ch1lv7KwXz23X/mkTrkk7ylBXdN
oS8muamT+jRXrucfVmgs7k2oKRyfksXADSPxORFJxikec5lAaRPz5hwxhn6j8sV8
i3leBZWJmY4sQRQLOCfCEwUOT1eTKr+O2pc48bEy08VvHEjEyPoEhqBnF/YMqwP7
UOwWsbMObw2yzfi0FV127e5TFWWxsG9pLkxJchToLwsewx5JuBuFERmrjzzLJ3Ol
0BGF9e71Hyf3+bs7TWA8DXrV56avTCGYOJOWQNx0tkTVtArAWtBOyM2AZHH8mgNy
PM0K6zqZLn9bU4p9hmVMjFQv/bm1T6oWRxGSZ89geYb+QXGHAmFPjZbLIx3uYwXQ
+X+/ZRwqGuQWXIeXy2WQDXiTbrhysQxFHOkXH8DLOsqOP9P6/KkngiKbwR2Su6Ow
dZkbyFaHxMehnVctR1mgQc6ZAqHe2XNdlbDq/TeaT8W/lGVa0QQSVvdaurq7M1yB
HuuxwRoRGg3YrrbPAOYWKJnTsiLcrnBhJq8z8cULnc6bMb9snkY9ZSDfHkeENIjg
zRoyRJ2ZQ/2Let4ZFhovF1Tngg7q4lniQc2P8yo+353U5KCoIMy+hoZed/zks2+5
KFuUkjN6K0LTeRW2LQS5x+MOOU8iIEqRZfidQWVgO3KTiDVy0OejcEr5ZHbIcQ/W
yP+qqG2jyQpt78AoRKqOESiQ5zapR9iacoqocLIrjlTv9AN5cWtx0evCbFh/L8fS
LrNFBGWzTafYvzkULo4vey14L1VkfPplP8dQJMTz+3V55w3buBqpkLKQFoSzT3g8
iqHMluVXA0yl9MyDX0Bb7TqFzlHEY3yCKa63qzzmaXZYAXnS/NDDdH5sc8yyTu1P
kAOG30dXk1RNkcF5UNK3FHe0Cn+w4cK4nSUfRr4b03A57GBgVSs1WW7hoC+cZsBg
D22GNhqLcnVjMgVb8WyRxI1tYZnACz7awP3YccIvFufIPImkuDT0fXwbCyKW7WEp
K7qB/WVwTMq5Y85ta3aJ4dORq4mUnZ1qrfA390sSGJ15oBXCD+Oqk4Yx9e3Xe7Nl
w3XoCJORLyznicpIaNvtrwHN/BGildNzgh6sp+Sf14EnbZy7uI2iQxCbGQRd9d3Y
90wBKvUfk+E+Rwkix8vlUaDTUfJKGvtJT30iLUd+6XDBlQPElz6r+8ANqVepnuJv
V5GLYEzT4LeklMtTcXWUZiURpsbjJqz5yVNljidqhU3MspNKA608FGzbI1g6ACQK
/3mlUGLXCORaGGONkfjBfX/E2CUChbM5uP2a5oNvVEsQMtwv5f8jQAPQYlaT1eX/
JLhYwvwYUxWHpAaH31V0GC7TJhW0DyE42MPXNdHSXh+vwCYgZ5cJEg+Zcv02fgCV
fzS5dFuXeyyYoVLbeNcGBk41B4GGiL82tQfauIRIyyzwnszdW01G1sfyLs/c2F9x
HItjjoTXXJJaDaFKsR5GzsezGijr2bqH9q1U4oUdFgro4hUoIDcSl2z9wiBM41RI
Z2ooZwlXvijZPb+3XCInbON48owDCsk4n8lDTa2zJHPtSupcFMwplLWzvwOfsbm3
5cv7qVQKnGo91QMtgZupNiIPxBVZ8JEgkWd6FtNaOkLxPOGz+d0XH2qwWWx1+PfJ
ECzb9x8NuxkxIZh5cvC29/Iv0YEOM/dA65j/A30YEqCidLcmKocSeC5L2b1l9cpf
Vy2h2lgAOM4oUQVre+xwVDf0t+l6dzCa5yI6tdW7IR0uRMSyI3JRSEx3BfdZUn/W
yhcxhWhWDtely//i98MJJdN0tCJE9ItNYTmq7aYP04iSYYZmuVl6KFbae37WdtHA
dqAVz2V1WGK9lGEXrDuXP8tQVwYRZoqwAAhSyJLCh7wqyfMhzMXLNRWxKhMV7QZB
2S/LmC8rkPxbyXTo1/ooibhWedBGssEVJWWMl6uLT5fKj0BGx+wjI4WaRBZPKLYf
4MfaTtCylcqdQyjepNVMwnoC+mb0V4zpbM6Ur8jZSoIo/U9crcAegUnPkuJXBwtA
qtJzoIPGjvatGkJb8b3k78QcXaW0IqslSH9yYbvuvNonuUmQ5iLEDQlyBXHMl5fE
uXaglRIma1pyx2S6eblKpNCiPXBRD91pSIgr/pCYsrHEmfyPk57mDrX+ZOAt0PrC
XhkcgVn4yHt9M5FTFxx0Q4oeC1mwE7NLKJxhj79IK6gu+KV9snFVWmypvCtNGDCP
hjMCUG9mdrQAuvKIHyGJOd6gDFtEWBvLu8aE/HCSvlzK8Oe977cyiwgxxOa2aZ9C
T2FmuuQmqySSxxkB4lvx6Km6nXxbyQnZm0Xmk/PWdDB1R9NCFHDglrK+eWPSxEQ9
Cyi9oD1swTION46h/dJIr6SysqAtYMSRSEkbtV126qzcx0cjE5xfCdAxkXXYfUpy
nWfDGIP9UgG2c43ztyJUvtYbs/DTePFXxqBHXhoLEXWmPGDooMnufEpaGYVx5OyD
CDRa6gHH24izE+JhBb+jG+L8vqo73EKiVzFox7yqnEsSbeeJ+ZDmRuXgxonK1SPb
A7yZek/pWgG7HxQWX9JP1dgzPCBAVK1LT0IeFPzSX9X76II0ga66tQ+ah9CzRc2N
poisjEILnSPqspxE47nFTp7S8jVN/kzIV236tBZbAYAhPvZDqvFE5RLm0XeJn8PQ
touCbZEwo1B47l92LKYDEFqxZ8LcWB1kTC7CTwa54gfS7ivW0GRl47SV7OPfhF+B
YX5D+DjY0UbBySvEgbSWpFk/68h3Lmjz58YJC1rRt65lTJGZkZ2XzL5h5bofUZeT
ha22Ow+xABCdr1NkD5UgnF7tYiPQjid45BOB/KXykwtPUIKQ55Fn9H2Nlqzfz1ys
sFfSzS2kmX7C+u7eMg/M2ONLhwAjRuFJce80j4upOZAY+0S5nFWj7Yc3cPe4XHEi
wkTyZJxTM5VenC+nv8XS9ipqHXfm+vj6NhWSoVEItxpXPvA9lTE90LaeJfnsz+hR
kt84rst4+2orNF0roLgi9tuTUbCr8dVglLNDGfLtyVORKndIBrVX5yZ6675HfKEV
eWzm89wo5P55edOgAhWJNOEuyUqHr6p7QYMgpmzIrJZIrPDzv1OOjBn4yx/jcpy5
JDYBR2OPS5y31f7x9+CcCm1JWkhCZWD7jxq5m1GPsUILvj5aCRadd8ibOKsWw7fI
b6HVlYfIoF0zQOv9JRZIms9wCT1n82A/LkqHPfB98cgmMFqo3OKJ/HxCojwfBXzs
mddQ3FbhS18R82eM0lyCyF99FBNAy+l12biYhIs6HFw6yzsuyOufIWXg9+5nv7RW
+xTnhbIENOIVLTtNGLD5Ox04QrMFT8ctLDOVzJp2FhLGFpfY0gdFGTMvWNCUc49r
tzc5X4Bgl3p4GZBv9cbyFQLFeaoNXYXm3E49Bk/aaKhdcqplV/WKqeTXASuaaJVi
bR3ZYmm8Q1tTcHgCtDQzumZ0mznxLko5l0LYy1KJDyxmnvgH3rDpIpZEBEFC/f04
wPBgb/q0s3WqeCwy4LoXXCTvNWJv+Z9ryY+Q0JaawrqscJO6I0f19difzw5M7Sdn
TPwf4RZFU4g6TNQ1zrRlTKyYNK1PcuXjcs4ReFITiNEXPTYns1yAiJxCdBJzNKck
2r2rU5OsVDeJmku8ZrWXVuUpWNFmZqG02R9+mwOFZQBpm5xRII2h6uU4KmwA5GRy
LgJI+vpTScrcAF9NwqwI4tctbOiqDLcy8JuI73N4MC/ijQlK2KvgziRqP5odDQh+
DTONbZQCt40viGDLYPCLMpfnMMnIjNf+dboRbIHfBr+LE7F+MsJER2IkhcgqY5uw
XTrtcbq9rbk7JlaS5r0DUSXNqR5F3R5hPXqPHW3xhRevOLHnLai7TDQrGMzyBOjS
cE2qA4LYlN3Jj2kBfBQg22quOffKO2yf2g10n8am4OuUaTcylX0TPswJmU5VbmW0
+BTL4/pm5WPWzYNQIpHnMYUNp0jUy8HQZcBez3ilaHkXTH+UVdbVewbZJvJKyWgz
kFYcWWxFpuhJVWvVpbZ47u+vheiFKWqq4GjWx9YQOIRrYyLssQYvcmGyazDU6K0r
221TVvWZxy7QA2BS5la95uYCHc145btFuHjVAH0MP34Pw+DLHhY9ilBrogpuc80K
XLTnfNvCdYCcsQfzAKRZrKR4Yft1oYyshmhBySI1roi7UOT4GA4dz6faUr4XJDd5
AxPNbYSCovpOcAvWJ0swMd7qj2hp2HrAv955PMHD2yCF/DGERsupf8zz4cADnrsN
foiVwCTpZgcMvHA7c3iTA/F6fD+OdQ/b7e6n2aziThiX21p2jBdjVHCj/wWVcoqo
4PW8d1SBAgm6opc+OfrBWwwJpabXolKiPg7Go8czAcrQ9DZ3Xzqkqb90Ga6wunRJ
iEUo+zYSY36MvfAyJr9b7HVPjacfHCIuTMAC4wx8DrZYh+6ggV0Hw9QaPkWgmRM8
S3UJZT4dmmHT32BaiHZkfF2gaMGd1Q1gp90cLR9xVbA3DVxu3ReNQjG3JBlUvBVL
/IQq51qdZ0O7aS3PiQonM5sBUFkOMV5dOeRYJpUEdMsF21/XkMN/mFV6lxTYZQnc
Jhq64S9DY1UovtXMgQsFVzAVMQJKtc7FSVuDwGQp/TU/d9KmlfJbyNR70ouF0ZbT
GDpzES93ozWIa8TNYon+ejNQkmT+MpcTTvQY+ZwJhQrtVFsrBhcDIuWabakoSjII
uH2G/M6/3IOVGzuJoiIt0PtvkhfaaxytSpVIwQk9xw/Xc9hQ6erYZJtb5MlWP3HU
hjBph6f4jV9dHn2I0Z8B2HN0lZFdMAffF/lDQ0UeU5BNI/iquwJ7FA9U14pQzcbZ
EW20h1eecAj2BMRdOVgUHrWT5BmfLbytPeaqkeKX1ZHQZC0oDvG4gL1fzfHQOM2y
jeU4t93xvnBKJU53UGQPHGmVe9k7bQZvnKmig0AfJ3RY8hEkIsxXs7/Buq1UaQah
TxCPG24UJnxa4y8O+OPYv3mBtojHQFHtRvhq4xR9x9WNLtMHHvj9SnCeEu8xiDsA
f7y51e9gEWN5GilEgPH8wfXHNz+0/G7vM2l1LD2p3pVXRge0MNvP1Uuld6Dm5Ihf
0cR3J5dnzZwhJZ4qA0gyl5EpWPB6LPzLp4UNdFa3rKoe6iMJkPHkHFK9xfar6EpN
lc/myxn8/NYIvJDnnCSnAgB2FOV2fv2Fy9qi2lISsLZAPZ0yW87vHXOkRzwlD1KX
1LAfNAIq2I7vIp3CTfrmSPS+9s6CeFuxBEoZvV6l0NvMH/7TVyvvnZZksDTGckDf
hExEd650Ro0JYXzhEgUej8fCaimo2y3opCFdn0J2ta6GYr4bRhkQ/POHRXzi/xIm
v41EGRYoXYVz+TLQJWWeCYdh/EMHVb2CrFU28AgDxEnAzfdsIKmhUsVdpTh0MYqP
JMSx4bvRagHJH5KSqfeFz6/wfEHAk6myH69YPvFnHXkACJTPrXECBZTIfoKV9mKU
qoLde2WHnPdMguraQYheW2pzVRT/GC/4yuGU6yxGk9q7MNX61GjVlpygHFpYtZM5
xJi7RLjWgmMNITlHOurfFhBc471yMcoT0abBCViduthYl+HXDD3DRHfiZaGxpZct
RJ5IS1HEWY4at+KmKJqktU3IK9bkwyOLhLn9dTDQ3n0Ok/DGUM2QobC0DT4YE0ao
XOZQZsy+Qc42SSAOHYq8nO6/1sBWNDJr4Tyq0GrN/CejhtSPIIrOKijJ+jS+Dtt9
52Dqfy15D6wOlvGhiA7nC44otkdthJziC7NwRGQ9oHyv9oAoZPBjkFRsswR2Ylq5
bYpiTkEfcLtnQENfkxL0DtE9n8XWamjId/sIagXVHm5EqfmUicX1In3PeNK6o5Eo
mvqnxvqnfGmbSr73K8erhVGrrTkgfKwsDgoEokOhZwPwsK6ZzPCg0g9fdBdkPr6m
NBU24dg7Uf5JJ63LV/8T3KKUB5FvJ544IjqhWe8KrI1pbR/A+1NcsmYEOZX/N4il
Cq2GOrm6jLbB+JEaEGYY9ZrPN63Z+C8PJXIi87dj0eZwcZ+sITgwsKVrxUJr5wf4
PFKhDLZuOcRDl6+b7AozCsE6StcWrNrCxYE1NaE2DHUKx1UwEI5M+Qc9G7hWwUY6
ajFmY25xyr1H3WWr/SiRIB58XeiIcQ1+mu7qlTm/KZlDYw5pXd96+bwY9QkJEXYt
TXwiqSFlKFXTgKAAfDWPuSStL7K8cBVFsHr/JqbfMZXEx70OdVCVxBiIJ2C7BVN6
c03/XOhMFfgmY4RJL22XH7LMBqPF6M7+NjglFrlTIh2HoORU7kHHuZNuryZmkJly
fes4YCU0SfJlJ+fXiW8LQAZSaK5l2+PUKEHU9D3ey4Ifrj0Z5oKbOo/hUzEdGPPp
bH7UQcBPOYmMga654ed+I+KLyGc3Bk6tQRtAm02g1iHdvsuLO2XfdwfMRoEKHQrA
sqG/PfK0D0fG6bIm/6EdqvPhh5PB3c99NRJTeQd7zeZaGQFDPA2H8Qamg2xUA7o8
o7M7mrqAohGLKLW+Jm1EbqzrUncg8PRJBMFaiF4qgobo03NJ1mVZPLxA7/8eTMvT
WitOMW6NFDUPjmcp+mLWP2RtV6r4kte2ARnZ6TFewaj9pIS4Y3MFkYkb4J07t+E8
5qwi07jHUd2ciO3yM2WHCihPyDqMgo499qOT1F11jqV6OA95OAbu3miDbqGTcTHk
Lwggwu6cJtrPzMVrDDq6znCFjn069nHgR/6HrRokBKTdxiEpaD++76EJgSDQ+22o
cbmKl120RA02wEK8ri56PD3nGFT8HBgOpQEG//lUa0rLTaSrrZ+7cnhQ0VL9/4YP
J4p5V8oMAU9N40GcrytvhBBdSagZ5asH/X3wQYDvkceR+a9Mnl1BZxFfMbALooLh
Ow9SuyJgqKlX/a1dzvazSocvD+adVlMegFKMUU57xrVkXJs0H7Y9TXB9q9fwjMx+
ag6tf6EAHYMqLxU5dshpFl2J1uWhda/11Ey5Lvq2Pom3A/iCmCQdhhVM4ILR8EWr
PyfICb7UQTOnvuseORH0ZDIXYhtEJppIm3tIVR6Oo0IXo5ZqaK3d8ifSQANhw0+E
jkY9XCFzxU91wNUu2sxv3o+EmqGGPdBs/Zp0NH5N4ir/b4G4f7Y0Vf49CCK6dhge
G6ESXpwcAVrjWHo0Mz+mmGo6Idz7m6Zpd+qk1QtkBb6D+125l/YUFmuUgmQGDbqV
JBUprCy1Hc1Ts4HGApAaW5UtVOrCnrEy+FGgeRjyCTDF1LpCsUr2RUtkE6OB9vUI
wCJH8PHgsiykin+wcinK98O8N6uXjcIgt5CCfUoERPfFvLA2VKyRprGC8eH1ROes
flwdC9QfsPqxf3fqWxGa2v66NV6RkU5AoeNji1MCSWeXqAGOHhGU2FGiJSISQjDl
4QZ0gcTEGMtXAKMks3S2X1J/WazSGCVwpb8ywE6mtmQY8WVFLTGQuF9xvZ/stSPd
CQ8wR/6eIkfevxoxH7O76VUOHKooLuuMwAp3Mt/Cm5CBaHxlia8hNu3zWIaHHH9d
zyO9vsyImJGqSumNKlYDXICKIvrvkFAQ/ezAyIJfDlIEM+VoNXEut761hF28DF6V
qa9vDGUXE1UDsaa5t0bfl1gcXDupg1PGAjYUDocPX77AQJZz9oO44lW8E9IVgEWR
A8miUO5X5Ng9/ghpMk/sFbZiIXUfOxY58FnBGN6m+dMAl4CEZiB3P70MuTCA4VxB
1CSsEnXFmNhxxo8jxbRydYW9tTWyJLCLvyxOam14ccASdTqfkOZX8pcUl/wJw5OH
G/jugnhUa1Qm+iQlJUniVKWtyA6jtS9zsjjpdGYa65zWMU0jw+Xj2lXGOfOX7Zmt
Dg1LX3nd4TdF5W7Cepn1B1NAdKVpiwEL1BANOcffsZkFzJiAqFi8hLd01IJrGCk3
29dfLaqwag0c0otgeAL397GE0Q+PFmkk/E+NVCUOf8cwYuj981eRY/DXoxEwgRmg
7wQQDoVWpAoN/SOr5e24zogFp6S0BbcBAE0PfjN0XK+oH/qAGPN4hLZ3L+r40Oyt
TyRQBMN8DMzERncZALj0PjpMqRqc6Uf16nYw+6G2LQpOWweSf/w92YAzoGii5buo
L0FDx+tPXoXDPPUPKNLZJGDnZkg4bn5csYZZGpKoJzGIbILY6PYkb2ZRIV15CMpO
F1HFwNadFY24aqmSlGwr9gA4nvUChARYpB2QgUlPIUigyuH8C84913I7PKb0MG6J
H7/oCycavGKSYuZk0+Gao61AwvRnLeEi1HH3u5eOJTogtfYys9OZ02xuUKrG3FC9
tMQV0B4yMSGmUsm3g4s4DGUfUMSGTloet4dhmRzYldwNzFNOFpYQjo8geP40UOjB
4e72mehvPGoi+9JKiPb/T0MOkk3amJfvKsnvOSpd1hl+cieLnxUYvnzOg7rclIE2
GK2tulPJaTAWw6HqfBlKUcjFs/1yfMYD6tn7usICqCuFFVGhiBWmyOYYqr6f/hIy
AVtN3cRk2eJbVKoZT3hJY67yvHOTvjtwtkq3UKH/M4+JxkfOV0C0YGeSlmmTI4gr
v+2jVTCWE4nthCLJiJqxze1t8p21jovQ581OKl+fwqDSmGQmyo39TcbZDaSqpY7k
fbIW018XDBl8Pnw5YahP/jfnKz5URlFDTbWk9lmofTXuwWtqQ13U0db1mmDvf2ZM
3KNEOlR7/hIia2oq659nhFg5uo2BAVuXE1tr97ZrDdjRcjGyBg/AD+zuzmR97TqW
syJKmquYmwmfyIZvvYOpCA4Nf2lZVMJhkVzibax212YOhEfp4Ptl8GkQBa1ufRxp
XTToYidT+cMcKiQlIkqEpO3OoqloMtiBf2zIWOcn/7ijYsAisoXFe81S8M8uyESv
QrepqS6AFBPj08XSTWoMutwS31r1t30i17btCxFOVTuO8o1dyvbG+Ng8011KSrJD
UQtEomOTXInUM50gAWE1D17xbPeGYU0EpSpc7GXUTugBaeX8RUgfzprGwJl31Cu5
VlVHk9+DEAXzIl5MTKFYtVq1GY13BHGppn1wSGDk7ML+5F04NyELB9tdfk389WCB
cfzIGwgf2FVIklPBaqLDkChiFCQkqsxK5C9APz62mPUErtPz5aU90BWR422J4bzt
4gsAp8By2ns4wV2daQ3jULr2Kyrljx4sHxkzAL91bftLSYQY7K0QVVTzROx0PBqg
fZ6Cym8DEMxdvFllXM8wRILwAKK3WYn7ACehAvOxiBV57A3R+wATOsfvGcxefXaO
1npbNo8ZTMtzMBPH6lOsF+hNSdscoAp1cAQMF96pV2ivD7om2H1eLXwCgQKwMsGd
D2eS/sOYqwrdPPsBZD2hHYEI/4frxRlGydpErqcARvptXeXFL6FhoVLI4IQxQnzc
jYZYDosXwLAZ0gh5C0H1X7UbpppmSOYPV8hd20T11UmT8V3LnUUoUAYVsh/2C6aK
lfRUVEl6Iljw9+Z4kJkLdmnzbDfMrUBxQcS/g46/Zi36TQ43JMsdj4JizUpMnfj8
RGR370YJ/GoWGF7K0o+ZA8Nxqyb4EhgTY4XoWLyf4gbAt9t5i4SXCZKzffAZSka1
AAcW6VunqnucWyBC0DOLzoQAkF4NU0tJCqNZEHm0WrneNA1EKerzpSFo9MeV3Pya
5V7QgzdydEFccLie3A/Rf+ckYSH9Q7itVOgmK39VL/fny8QHS8Y/vVdxgw2WFdPQ
CPxEzKS4KU9NIIp/mmImoUs1kbX62UAtk5djFNwdDUphriG7ayixO+YOZKLp3txH
Cf2MQCQTiaQ55uamKGDmBxWFjlH1Bgk7kl3Df2c2/beG0BlwLypdPdstu8mMETOt
HC3PL8Bg/5TYNvmwh1Mhzbs0POkLTTNSrMAxVQFV2S+LKQ1cRZD1Sh8rK4XmzT3w
wE0jpd4NtK/bKOmqnqujzFz03dvi8r35QPvXGR8uo1JgWVF1g+Vh0SuDeHKYp9o2
50cnLe6TOGQ4yCqVvXc0aUu8VAcuVJruoj+KD0Dx6CxZtHHppGk5/yoG2pp9YzNW
gS7ahfpQNoerIixDprxsEDUYYMOJ6hNjt/M+vs6nwXerJv1fdJLoARtNLP/yt/ht
xGr6EQCt33zhBell3zyxOWL5ce3vZfNgJninMtH1su4U1/B3GhmwAnC2Yv1JjbyL
XPHT/swP9QhqfNVhtAd2YMVRSVR+HBuCQnVVCgb6nmXgZFBgx9ep3EyJx+sGHdkH
fCGOLhH3TxUtQsXJTc8v8oqnsK5f8aIs+/ANzDI0vnKaN2df+uVAKVbcLqT3s7oW
q/Pfz35E1x6r1NnkCE67W/EpkPKFgYbTJziupTk4ia7hPw+XA4yygPNZ0ZCRtc5X
DXT5RP4eXzqYr2F7NpHNY5pDRrX6JS5yvGIA9uLz8hdvwRq8cdC2Z5PsSE+ibXCf
NCk78h35fX4kqN2df3LxtjUmZIIiMnTZHM6D0qeV2pul2tTU9ogTGuPkJnuPCUqQ
ThRmymbRDBLTSmMQEz3aZEAFSKrTacUBNRWSQslnAd4Z92t84XV6FVWzZRik0hSI
jVZr666JUju3xn7Yi+GzmvZpWXC9mLgvH4CX27RUAmc5L921v7KgLGlKspI+77Ni
MbZZeDwdTMUqx330a9ZU5VgrekPzFd3T+tmKbcCTa6p+SmOlQJfgk5U0Ol0bR4GG
c3t2WvTyvWecHEQToJBwLOxiwg7H0fSk2yRUfsGUrLc6ZSXyAr+VcNqbsPIuriJp
DjH/t13CfNfJXXgeEn72HdHNqdHTCW/4V47vUy2m9zyDlXgIhPGhAWZklKeVJYoZ
MZFg/+yieM1zQSgeF//Tds5mz9/JDeMXezrbXb+xFmxZyF8hGXy1tK8+A33xqTsp
BXxlqRdO6vZilHYMmN3alw7qVizBtUYFai4XBrax0X7NAnnGEho7+JR0pHBCOH+A
gnbt3FUxba83cBhRpnJ2dpa0n1JCe6mNj36NL+5PJM7o7eIffbA/0VuEgMO1JrRA
co1Rn7owAfM5bgjU2g2mLM+w0fXQWufF7l9ODHKc2fCATfAFPpfFWdB4Vr5Szs9I
3j8DV7n8NC/IR9QSB5YJ+HmWNsNS1Kz/KjqlGfv+tApLgPlK/IoaiB31dgcq1E5i
/Nqr0Iz8y58F6jfRnW8M4SMuALoM60psnpbhqat2mG70Ujo+D/WeE7mr6LbkMUFi
EliBezNLcTkhQ+pFhyJ2hc25X6QBeEvdWwwFcEJajNNalRr3L9pZ9kjroje7htiB
qG/55rSkszpy5hLB4Crqznx2hc1Nt/ORhuurUmKXhFUEjoqRfZG5WjgR9BCvIHp/
tCVO/dWFDRi/hv4lE3nW/ToTeSrCgdppcthBHB/Mi4iA8PseD9Fs2hwIZ8YUeVAC
DwUJs4ssdV/vRZRL9pKcf90PSxn2uWtuAd80qqhRg3DtulCJTlNkeL7z6w8Ie9zt
/yiYqapbnbixJu2hBbKx5OkSpI3J4OJd9On+0zdvzZd6nKFPZFsn3EUxs2pYUt5J
o1GhFi+AYuS2+S+MmV6CSqUFqbHgQYzLp4Z1oj2vhciFTbY/PlEgx/KaXqTG96Uq
P09ahFtrONqlQuaSJ1y/4RHtbKGe5kYSRH/STe7tgUqdtqQtOA24tnwB0bcNobZH
aAWN9k8lwvtpmI5TxBd2qbs34oJoQJ875NcNj4Hx5KNuUICGItrup8ceT4kN2rf6
luXIAsoHQJ77MIVcjFT+vAJIYozr45vqxEnysnxP1phatLNX3k7d9K0O2BVFG69C
ei1sB0chYT1G5YbXq+puoppOP3H9wPvh7BtnGMftZVOSci3byTOn6/rkOwbAanLw
OI99B/7YiqHuqBTCWd9PbJbZ/yQ304YqApJstcT/0huJBndrJ0mzQ9OPo2AsyJCM
fczclp6vdxGy9vQdAsTqohaMDj2DUV8nAiH9YUf/88qJigKDLcYj4jQk2g7iRHko
T4P0xGWlM1kR+k9tmsIl+y9AapYdm0OYS/XfFyiEnI4vwQUub/fao7WZ0tjnPIuh
HJQa58nd2yi5jxeDFe5/pvAadocH6so44u1iXcrxcMq0UaBW1nAmufW/FOFkeNDx
+72fygOHJI6i2LDGYujVNKs/YQ27QfK28PCEjbhAHWm+xkpZUoHYRhvwnqKlG7DM
nVMdHrqmBkhmHJrK98QoLfH/2h3zb0cJQay5j0ulaMxZYMQuV3tOigEWRgwl0AEz
UkSXw9ela8GENM5e2cjTKa2Jt8MiqgkUZ0oB7alGnMY72Xj25AkE8dMsK2QjJWi4
LELTonD5sOMoIzb2M5Ky3n6uIOJYkhNSkOTMcjikx7DmpaE74oKA3IEPWVk/hd9e
amLmwfv+ktAimZl3XaW7656gmKdegqWEcN27uPAVk/5y12tKsh/XB5euAIry2Mwd
OJEDbDke4xKhKzr84/nPdJMpz71tBUv8cAl3Ch0VspcahHcwbqo35BlS7kVUSpdU
OxFAuchcN0/go6id4tdmPwCg3h6PwVeIL+KbIvxhxpFqZicnkX8jxtXGyYk9/EKp
f8j3mDe94B700ui0D6p0iQOVuZxQLMUW7xfpSIKUhRcqTch7LBShPssXw9fgQpWR
LpHjPgYc5twbF9wBYdYioAY/WSEY2KKP5a9IIbU7HWJ9JAPoOGg+iyCWuYYlDEMo
BijDMaiIqiC4AjSbIF1yWkCqYnnA6drrQ9xr0vLJf9yeMbxIW8VEbMKAbTph5LcQ
wFv70JB+wAhOF1FBcFXCVXyBvE7FyNMMbXHWD58GCgFtC4QTqR0fKgys6y70GcEB
OQGpLiwUJAtsYyaoxAvKWeDdpdkUZO/CINCLoKWZVDkfZQ9Em3yZ1RvLyosItLbY
aEns9A9NfGJFtwmDvRE8APs0VzcIShy6q/gwNng2BTcFp0Cglh2NQMU0p3ifI42T
cP9iuoocNQ3dMo3HLDSCXY7W5B45zYSUu/bpXvWojK9qbjCZ1fO3GKjEqWHCcF71
yE300ySyUkjiA7B2mrd530eTu7Cc6R9BOjRi5tirgIieJbvPiPfe9vuHhZYCg+fQ
C7eb4QbbvstApHrD7J8V0Y3DYbXY1/SI3Ymp/I/rO6R5zDaRM+f2dqNmcIoq/bjP
0EQcQ7fUEghyeE4oNPUf7l53CKsLNKPCbqgM55x1tf5Ucd/vWne4GZAIM90d1ufx
joWviUn6bcn9ccxoTQdHL+gac2BiBiHs42fuVCx/B/bI2DLAMWaPZGF5TOATYywU
rm05cGcwWg6gBDBmzqv4CGEEP9DbiA6pTYQ8Z80GTxOO+w3yQqevX0FDUaolqXXD
JlD4SjZW3qPYkBm//j2WpyFpRzqHLuK/OpDeb3xuu5vOgm7RjWLfQQwz1XSgMrId
qnNOFGkW1r0CR7IukOyplY4eFPx6Rjurxn/qWS/75xpiz6XlifmLStrsbYT14KTy
y2MwKA2oeXlPpr9Jdj+zeuSbGz9ZDTpAc2kLsorQNYDScsx10vGr4dxaDIqFt5vk
eT4crrtfOHCirFY5jBUFcUoCL3KkWlLdAr8mKBhpM3FL/u9jcyIUO8MT5HAGLtxD
UGmigKTnuO6Z2XFGaBcULuBZpESKGgENHWMf76yl6S/yxu2CLh8cuRYm6lQWyQtB
W8dcusWiqktpwyLjoVjCu68/xVvMEjb0G91WYjKJ2CYMtE4FV5UJFY+b4fOmRXcD
Y5DgbbBzZ8zE578FMzPKrhKuoSXgYCgqHKal1T1K7RwDjm6HgTTdDBoCkKkd1VW5
LHT+F8LG3P3A1ReP/dPW6x0fkoAFpJk3rcrtw+m1JiTolkk7iGEIk4PuapyaAJUR
aiNtr2mXkK7v/twSwTFFfTs+XtpW2vCNF/3Z4ZwuEgLqKctloJKWOmy1/rR6HteA
G/4VVx+LjMxN96HP+gci9OkLthUT6z67MgfQwFHtqdAd4SWnq4TDmgHjOIPh3zQe
/dFTQZpLLBX7MUwcRHzT98RmXVBmdJcbE7/Wj9db+AW5PHQJeLEywukSm9O1+ufe
SxT1bgUIoPO24HvNz4bgFh8HereL7cxRIsFr1Majvr5PC1NtChxICVxIiOCtO/xW
sct7RPcfRNAavJ9wzw/nEppa4pxMEDcxiX6YoCUc6xkzXrW0bvKqHWhmvqhyIF6/
M7vleSSbQQg+W8EHa9uGd4Al/Ap/2i5baslwjI9QFDvnpzjmkTo1kgZCBtX6vj1z
VFSrgMoRc3BzxOSurdw6mVE2a/noEdpjDJ6hQefwsZDTXe2zTsAZJJywV0ZDNHKw
a1SO54G87G6MIlnZgIrY7rlC1KrmvJ2LNGdoD4qV023jam2+20U48hQGnN9TOATb
UJf6+3XFPUxr073kyEbfLCpKiucOjKLEIaRAOnSP+7seXk66vYToj5rixoRPCeMB
FZuf7nWBl8WkSNxQLBHUC6cVtlHIZYlt90Z5XIfph8/UOHwENs4XI4uy8UMbZtVs
U2xLTLekY9Yw+AXnDR78ZCxpG6UKiSyAsQIxbCtLLe3yTAf1KGOzF+aVPgM3NJDm
LDbQ8ieS4YqRh6AC3ChD85dSHHoPPBO7D978ULqA2H88r0VlAh7yVR7SC/fIvsz8
8muF+xfsj+ZPLfrmaEFfMiotQ/fZXtemCfzM03ABJ6upD98eN4yDiIZxlOZoNlvQ
lUuydW76ui03vjT+LljWjrSsVNOql2alAqlkVQENVSJdQ3MU8lhSL2pYu6kvWvi/
XfTUx+2I5vwI9jer9kDJdBZDccx1zztgp4fFh6uNhTh/FwRcDM6o0wNDc8+VgTz5
RuECXFyvhnBYw/6hi+6QS8vkzCIiZHc+IQxaWCsqGJcBZjHh/h/Q8hvkX3Kh6HdR
4se6AXFKnKmAuCBSUblg8YNeiSXA2E6hBcXLwzXyQ4HynyDgcJrJwzoQEm4W7bgS
TqQDXdtfZaC2um1ycDVo3YscK+h6e4ET6GVZzAPMFXWKpR8yPl7144GIgSADhZgV
n+PLi4ni5dStat/5faQkvewwNe4srjObMNUuPVtpNChgYklQFkjuNsqiti+sRxHO
Ak/wQe2z0UE7vgafYtrhGU0V8DkDs/xnfVzQQ2lplMfeGwXyDKeHbtzPOemrK5Ot
lDw8ZvF84dThaCWVq50UJpzEO6+WCidW8DIvFxwkrmZUB5YEf7iimx2lRDtK/RqC
5egtzGOV8uZ+/8tIK7SS0kGMGCWmEgrGhTcLFcUwizPxglSpgiQGzEKVxrNB3UUm
zP6JEOlIgHkuthloVUAVKmGHQpydATM6we1ia0LVeWSnFP1LOXc7vwLN5/zXk+gb
NqFRL4sQqWCmMLNswKLluR4YjeTRfba7F++/AByjuwbolr6s3+PHsjUz0JPc6zWb
y+eXzggrZpfRW/atQoKq7ddtEa6hLR7V+3dQDWFYByvwNIdXUkCUXkS9hhjEIWwJ
NQbCkozlzxWd+BW5ur4EJ8aTzNVEAWOtl2/Jk4TkWpv27xelyZv8Kz42VM2detTI
hQH6+ZICaVxDkJU9j5QpN28zRg99btCIYfMHXq4Cd0WnfRTteG3uKlCraDw+w4am
awOmStLDwHYbMC99MgH60xM7c35gkRVMWfkEJj6+a5VTasSdh1kPTh2HV5ZbMche
DwA+LYgXbgowYs0ppoIk10nPMyf5JupBxiUapxNH3I/593eudwc7xZ9k0MYAwW6w
bFbSDt7HVU3X6hl+AHlK1PAWf9vp2oodwmXMAjla9m9oAE6Bst7cNEM1SLWyGH8l
Y0B6+B8IyT86/gI21TNMSmYoxBxFsI0kSQX3EQww+wmaXn8MBuoT35XfK31kEE/H
QHwoOa8+bwbgGsYaisw3F01inqxS/gp+N+LfTzyLItdNhuiXtfO2N6rXtatr1CSk
NXM77MLBRDpsgJfUDAphACciM+b6dCXdfAZAQV5lrE5H1e1XP43S1b9UFziHleJn
cji2zKlzlP5pkUIXmoLaTT9fmI7CKXbW/GIThgeQ1bsGdZc70BWfRmhOH2xYK8Zm
/gjgtzeq4vJL1A4DYf9JjI2ySXc56zuccpu7TNkHejdLir0VSbhSP6WAleQN/c12
hkqsJ/0tTjZX9GSnpHPiuo6xPi6yn2lHe5/RSC//djW6ywEwgBQt1bX4iqICkHfV
ez8oT9JqIZLxn3lUYikh9PS9jvH7i5jWTpvnR4GsXiUs6C78Y/8Ewh15YFBcy+g9
HCxAY1BmDeswDX6+47f6vcHQx8ge9T8FqUkSyzgryFyi9Gj5x0GB2tJZkohYNHCa
dgXrTSHyThSHFmgVrH82Hv9h84YHb+s95UFf6GPW0iBR/wrfew2crhMj+y9fMJVc
2uRz7Xfboa3+W+rAUeSDguv8ilRGryWA4vnhBU3Ij+cEf9sjA0m6VmZkNqjsrZ41
24IhvYASaxmADq3U0B8rmq5P3vBhOVGYKRX7DIj8CHkxyMVhhGhH4rD8BYwpc7pU
zndeKWqquiOaF62NdncQnp+sLKR56o1i3+mTwsA9Zbb36OrP5J6HN+xs1Nyay+pK
Tp7ZdrSrucFyNgTUYVuQG9B4MjtEm1gJUN03d3BjacMfcJ05XrOMBu6XFa3wFBoQ
3DrHSg38BKibmoUHj1pjwADf1Jv+TIC7o7HEfidevPUMRJWJ1QTuEv4Lnc4G7b5K
uXK0e73lfr1mfh2ufqYTTGa8lVaZYsbvE/HII5MmF7R9sLSP+Y6orxb3U8lcrHKk
B0prSyD7JnI9Xdi51F/6GfRQdFvBx9RCWG3yw5HdBKfiZvOiJ9o5L2hZojWTcQ2N
2nAo3XwRlO5luGS1YwJx0R56vDMadvYXvMJAHvSczpZcATPAOdloVGOFBMCjiFDx
Mb+xCfrLx7e3WG9Yk3LHuQGas0zCNsyNYJA13W4azdkYv7ADNuPnHP8REb91X6w2
UVOvQwyLp7I5CxAQi+XaZGxzivcV9zntWtUesUBFGIVDFkVtpv9jFVkV7KJ+dijc
C7/xHXo7plLOxBh1QlYPeuLIKMd8Xo6pxdg8CKqq2UAPmZhQ+c4wAonqftEv/Loi
ksovq3YRFa9iKXFOQrJWxvx1CYuC4zNVEXahwvU80FClu61MihR4Zq1YICIaf4cI
f2xyrl7Qr9uBHxX/MB9EGaRW99Dhtw5Koqnupg6AUPhjFqwlfF+cAJKiXEt2BORV
E1A87EGOzZAxqdlul4e0HPa3dAqeWvHq7cSA4YEEo3G1vapX03FdUvUd40d34YWN
wcqKo7c8s4xVpwpmj5XjkxUqsNHqFaZXa6dhw1kKmud6rVR3RHbwN9zaTixyQJio
7yVLN7DBYfr2S4MjL12BtpPDDMdOikwk9pNKyuwq6vukBZXVmUAVKkJKx/FbID0g
5PlGjMtavdkWWQE/3euj2Ki2U5MUjiYY9aVbuxtqCR27aysQCTGMw/Gqa2NoK9z3
fBLJHct/tI53LPwgsxjsjGj7Ck9b9sX7U9OLcI0PvvVGruB+dmrCzFB2qA033Lvo
LLnsDfRhw2YZ/cTuG/ThgBzkosQ5SC6klCL5vNtGnQwdZcEu+B0DXI+lUsx+o5ni
Rz5ck5QQaXTYQEZnnuAtL8UbQUs6gAI4Opoe6mqJ6ANkHqDYoAwi0KvN4Bht5NY0
NHiCMIks/++fJk6K/KPtD3JWX13P4LgjnsRrA263tjm9VuXukFIEdr4qX+kN58Nr
gplzFAwNPeKRkrk4l6lUBQ4YvNqeP7UPMyVDAZEKLm76TeFe6/cujulWlI92pX5V
zXJRETwCUTjebHjyyqvx2JkJ9L/0O7yaKegUpecCc9okVaQOgqjM944oMjVYtaG4
DHh1KaYg6o5FtG7f6AiVZ5+jsKdFUpa5U6kUAEE1lEtrgIrcxfncCy+mgeY0mv1I
dJVGlELCvDkZd15NUFD35Uck3ZJq5BVVDZ6xHDkzuQbCWqXChPOWlQuvmqfdH/cm
Ap3QY3oEtc9UR2q6g7rU5phQK2ukxSL4eLT/fmalZIGaT1Mu8byauTC/D+Su1sch
JJ0IxQkSfZeXh2fsM7R4HYccMQsShIHHHmpOkilVWFoyTe/z4m92rE1HdXWoljT0
7WuzUY4fAcoxv/6wO1I11Q4+F96EXPrY3Fbn3bfcD47nqZDfpxA4IM6RhOipBOeM
Rv58T6CaolEDVxDMubScGwyJAPWK/JGsYTrDFIr8XLnkbAo1juZ0sOrZTvjLkJOi
DSSi26ZUpo2RFlnjbYyXqF4TqSNt/4s8nZElJPAAkiE582Zq6i6aB713OKOmkKVF
seNbdkWWObVQwgVQsQ12trHqe6pirPfXpTZvPH1SMfBLH9971dol3eKHUuWIZ5kt
1zPSwHckuhfQiabaQjzjdqOlPsRCQL808F0eOHHYtPxx81y0ZSWET9VnlQ5kiRvZ
rqF8rJSZbgPYydgQmdOyEsTPzY4ylFHuCG59zkN1h0EVZh/4+TDAE0BHLqmCMu2O
87mZ+fgV3yqPTPGLYU6It8I+xf1dUEmlLp7NwN2QK2dXkQhB5KyJFGIofwPsvexz
u68y+9yO5wximZPDPF3clM7q1LlzKfWlFpXzyUPavedN4sqnKREspcQNAA/JF2NZ
0g8nWIyXDy7icp+aDCZig/utNEja0f9n2mrNYc7/e6xv0Zag9tDa1EgcV7tbuFV3
U6yEbObKf/mmftVpupXcnL79Zkhn88h4BPpM35lvhXSWsFT2zOOsD9pSEcqznpU/
llbdmxT2LaZCsHf1yOTVw8VK52FjTOCZnIX6ZdJZ+2trqJnZhd1LhgvuL/lXLje+
6f97D3ddD0g/SMIp08fu4PqclSA1rTGRfUby5ScgXxwpXWg4yHRVWOIXxqunVogB
dDLf3ZRvRRIqx7Bk+dTEf/AoLDt6wwg4bLhS/mtUxUKfN8imHPr7xXPmTj+6uJx4
GVP3ECqshZQShvm6GKuwL4cb6P5uRMLt6wRI2MELbK8zG83/Ld9yZo6+9HqB89x6
Uk7GnW6J2G0HxJ+9Vjc/EvuAPyT9UQ6814oVnVHbXUL2Iy32VvrSEP4FsSd9GxTr
jDmIKG4TGGYsX74LMhuhd27OfoOL68vLcvr/q7vYrBtZLOzgYzRyoAltqVeLHIEh
3X6YOLTE3KBhLGaz5eMibqiFEa/iP0Be/uVAUG8GSNYmEC2X36+HWg/cHn1AO3Uq
3xsAXqm0ODNJtYsLgaOyuMs9ZR87X3gS/hW8ICw3XeK8R3GgePSGIWwQkpoIpqJN
H2oLJH3Ob50HIf3VwSpj3k1IElexLGd13v4SSeJ/wcGOg6Z6Vrm2EKKKEUTgyFED
+rX1vDbrQ9Hkfg6FTr7Qbg9G4B3PGYN5Hvx+/tIOOS0yB/8Rn5+LKxbgL9GJ2lwQ
ygZN2k4BQTjocsTUDvcy7DZauuBGYyjFHaGZltfVn/ir72BSxdAfxi3C17oaXW7a
G6p7NheLn79argO06jZxMjo7jDx7S+dOQc0zr6ahHGBfjrdQrq4YOI4uJZjkVBmK
a2oxB1jeRewwkXm7th23b//NXE6y5mTU1aGtdwAnJxGIdAkMKd9b+nDbXmewx5Tr
MSAG12G9NewWXFe10yuxxicjU0iJMVWbe9PuN9Z32FC/v1BktQzTOTC8wUUbnbnJ
eKYAV8qfi16ecuuHOvkRo/kRGAQ33ASEpHITpndSZS7HAAniOzHlsU76WGnpUiCn
zzZ57pHlNIkcsgOAZQnPYL1OxBcpPlm2ERFtNlJHXajTLndRuVzPaCQuoAqAuqtY
tS4RtdF40B57EHO9E6HVAjVOhDpKOpu46WHPqcxtKT5Rg1bp1qg9JxAdL63Q/ML3
YXp1rM34tThv1aNtlUYbxvvVh1WP7qkOnEZBHvHCHvwdJCeA1z1V3iHFklIcD4RH
dj7AlEUsxL6gCcYFFG4I30BTzFkknMYYXn8OMgE0KN9psdBoQhWS2ipnUYXnbipM
OQzSt4NWapSIjRLFU4vXSZJKbBGSvtBHxu+6RTk9ndZmc8iC1nQ0FmkF9/vPxYCL
o68dRWQgtWE+dx9M2WhCsKR43D0Zms36BnpJ8j4T+eHy9m4V/JphyHceJrv5g6H9
ja50NuPhNhMVOifmrdJPZQm+DQxXd5wDPqfdPqC/eF+8w2ozfjNzgdlA7nzJgkLN
f03AENgp+ozt9LDetPaH2X481pi/LPtkb+Q6c5ZsE6MJIkKmHJKa+1JhX0ebGOB1
3N1KMBMQnJR0xRFMN6TSVOwfpOcqQFlZ2fO4YxJhjcdI1O/NNkrmgTn/gb79IzVo
OLP9ObX66oFFsTE35jXJQLZl6f5Ff6akn1qVZa7GgExe2WXgf4JWWnSbXi45Y+aR
wD2khvsJGvcjrQHAxa/tjnP6GgICyV/S0CscRN/8Uep5I2xU8GXMbpO5FUvo5Xhz
ucxcDL43zzSxjVozX0qWkOLkB+Cu8Ew8zuA+TLTl5pBgsW8Y1cbEpNbaM/mxl8Zs
fIVfxmuK3EsOvb8/GRybt0hLLBsT0aX0O4BaLFOTSZrrJm8tlWHpx5eyhJx1YJwe
OVv1dibfqjmOtusLDtdOL5GhrLB/d0rqtN5fMJtj6ZmDrrSHlcWtl4dYe15ZRmI+
acTyXwivlsHCMexczDuQL5UWgzHIhk3LQAYAIYAokRrG9mZjZDfJW9qZ0PEXK2kF
8OFxGZ/KX8RGsyoh0PjyMemM3inpn+rm+3K5aAYbkVTYg9JPz6VhVdLvsJ9a1Kui
dV0O1reGGzvUQ2NoSv/RAqmFlIlk0bGHjIsvuAS7gyTeWZk/Pq3B/DKtCxMlcY1X
lbGeD7WDp/neP1OXswiz9JwTLPSn2abE7TFXMpYBwvQ0D9IqFLuMFTZN2q2492rN
Epmhp+m9HO5mtPKUccNq+2uFEx/C8oMaLRB2uH7iG3P2VxOwGQYcuOweMx075zrM
gI4pgRZr+NcFY4gBU6r6XSQYFsmhu/c0KYIQj1qRMvAAsBPw+p1xSM3hTltV7bai
5arhpUlLrhzSq793HJEqz7W5SNJzGCH0XYxXruKkLCV7Zwt7kVH9geZTCpSUzCxi
ire/5VAuEsMaa6YMzwu+nuRYhBRjUC6JUls+bJudyO+ottyKRrkaNiaJQCFOBS8l
J4+pMsIZMP/PL3kAss1DyaMpwWA5Jl59NjAU+5PyPZaT500xhcZuDi59K+veat4y
3u5Lb6pAOZnS1uIxWipJuKi66baqNPH14Hk5wRgotjOeMjdeVAR8Q7YmwilRqLdl
ou0QJaGaE+/c01GhQvT7r1s26n8hrUcppDowR8ts7khWJmjKEXxLHyRvRoDlf9gd
AeJ4Tr2CDnL0lb/YCAtDHt5cLhVHt/ZoVMqaleccjis7NDvL8lcOq5lxmL46lJnG
2AfxGWLzON/V6z8zFHO6YVtxFsdFGfVp1UHM1PauNovhmleKprmRKf8PPpq/q2qO
4EJQKDruSZHXymD59BsnVr8+Ti0GPRJ7RyFEyXpv9sPB+Ff82gayHDpt1vPL35Zq
xbb6RYvWsZOp12TGmcXQ9BMlEVBSKtOhCLQD7FMKcAw2baLvKKofe0zw3ECjJ5ah
QI8X2I/VCrKPvGxflQUtYgsO5zh/WqeN3/3IZpKcsI4bbtJBbMxWgmeu+5YToxYS
mncJ0qcneMFsVcNbRPsjx8Zn8iyBtZbGQQVr2e//7v1C1/8l13azRRVLQc5t7MrU
pQYbj7n41o6YYvzZPr1kvM3kR1b2sVveojnmhspygMTThtvCEOkmsIKK+6DcZ2kq
s2AMvoZsmlxNVGCeBmTposr+gWABTnxHRg9AF+MvhVvtMPW1oJeVmiAnqEna3IW3
Hs46bZmVJR1JZjV6d0Ey036gwvgKmLzddct3tqOHejaH/I9dwOx3WjsnjS2w7oaI
UJ48LC9TlCW3avO+klR/O7lGlqY/NqRIKuQVsL0pYTn4ZXHP6aVDPHf3Lf5q3ltZ
J46IQbKjs0uxcIXW8f7BlOSiJgQL5FDsrxpaOgCvSTrFaQDEXleA58bxen5l8TWI
fQwAtXgpdcpk2cpFa0du+Vx4uizGn7wPz9sjBuPoM5JGGC9BbMkOtKly/aS3SOM7
f7yua+Yvo0H+79DgCyw6YVI3e9mYky9cZE0isu2nVPWQPooj7vx792oA3W7iOxG5
R8fFdqoeKPLVIKclmuriQQaj+QRs9e3fDqxiymDvhxrKnhCYwLvfW9VrVZXjFxZt
4gk2WpeRXfAjp/QN+lcmVt98Ot1CLGEHrgRexDfUm0xbdWCSrVQ6OfHI5nAWJYY8
fIzR6w0OL4mvCgGk637fweQ7VHKCtwNfbLX3LSaySkP1KL9HJdHJaNMQp8i9w6i2
2CvNo/hdXQZ9c8h3pvOSf8v2RSMPxCM/fXcCRw2bGUVYGz7hCqdI/JqO0ldV0SDd
OCicXDb9e+spd4wEkGq42U1Us7IuZylAeU/gZ4SmfIF/ld7vfi/kl1/EoVmuz0CN
Jd3/5DPIUXtpTYCnuKgbdCruKj6QiJF5atbMonjIQdJJPnZviNBu7ToxPZyHxiNq
kOWFX3qVGSnqxjCnhHO+jXiA9wq50APubDStCvr0hpVNiEzSn2mMGqFne0s1jeCT
tQVqO5FXN8iYcpLpN29CScCi8e4BnMqtirzgVjjvZ3f1fqnZBS03XPu8u4jIrsJe
Ks01odyJVuffpFpmkbkKdTtnf7Tv4yhiEut6RPyKFb4VYg7Ru0ETamwY0/WcrIbs
9Ftz6C9DPWTOZ58dx6l94XX2//yK1GaBbKYM1BPjb38IAvEsKtgtsXpSpQ5kKANo
4Ijc7W1TJjnJ1HRDy5zAaDasogtHVSLeHSvOtgBMuJmdyaUqHwCzwdVgWopyMjl6
ZnJGpwIMLyXPBMT3Aiv/bYBTXWOQtZEYfdogptGfscTmSrtj77pKKDj2QpvZa0oM
sR8qymLTIT3kBFUD5aqmU/ncyKQ9+rHtsDPXSoY4RrT93rjaKQeqqEF4gmuWv/zd
WT61Z+QsuSgP/Z9jjKyIGAL0lQXvmWOMVtnQ9Cd4rtmSaH/9VzsrQWjtrxgHCB+G
bBYe9/MfvodH8hDiOPNpirZ3SpiZuM3QOrt17wmfsJj1762x+dfTsa/AZSu6gos0
QiBBd72w+xDs355lk/Uw6PdEhGORCE1R8JPJkDcTLAG6sadgJ1x5jz6UAKm0mulq
yS5qeJNcF7VUoj/IajSkCQnJGnjB9IY/2plEONADmChUlckoE/xhsqBcqrzFvMsY
pmRDF6+jY2k+CNdabc2qdltbTdh2hdFuTJrHhxFRQakYgtQ9RWHjUhUKRB35ocLA
aaRig5AfvUiSjezTOxEaaByV34qPznh5afI9nllDYFGQuHn3gXnUCPMavUl1Uhvt
1EfcfUbBoZjRLO1XzqfG2L8tTRNZVHcspZv0PvLfKWYUo1GhwJxl112cAD54nX0C
b1D9N9E2jXoARFVyIccCp5Hg/PoBaw8HNmEbMP98+r6yxAtVjkmt8qj47OsXhR1b
ppe6Lmg1j1vkIygGnt/uEKdovdf6dZPT2GD2E5ymtxXCP6flynvw1qxB5skVCXjq
7qxf2ih08jIUINIVOFx2ujyFoIPUl1uw+Rvjh/pw8bn8/aGLkkGO2ben9viwfuha
ebd6auEpZF7bO81y8Iv1qMNyklgXii0bgFyQcdy+A21hpctzu90/wIIIDidrYfUR
Ng+gsY13Z0NnGfnK9KU/bjcpzQvQBvtTnDeqtlQFoz40M/dT+UwIJOZjpSwOYWxo
qP015vWkc8cnmX60bqkLaorpV+kAKKK9EQtwSKhD+d+dDS9LEbog+YGlgVqoiIrF
b6J3KNW8r1YM9QkMMDnqq2IfeVy0vn7SKosOKyINQMr63Le88FakawOkBFRpDMoA
78rNkuCiYgnxspDmE2cfPogKrKSJGdLL1+q4JP73Y+vL97O9f2Z6I+nckXI8cK05
cqJt4EfK0+OdbsNItFkTiKWAo9n4g5IhLuxzNqh/vMe2cvny5pD7lfRvkShwdHO0
8qCEtKOH/UcTTstRQPtTL4bD5heRMiN9lYG6hXbBBAELwXUb6bLTbGAtumcrtMXD
TZVKlHjeI9CWTZvCdNpChStJnhMN9F+mK7D2aeOmHa50Mvn5xxA3dSaXQKhNjiwg
SBb0xVW5ALFYHrkzV8mwdKIkcno2/eUpFeM75x8NwjUQrhVBCznxcQSwhSA7A2TG
PX+pUz79E/iElEC8zNxlJ1TSmaK5AzA8aIiK1qFmwkKsq6amx/mgbNfxbCmitUbK
NnGpp+wQv4yyKtTiDiES5Vg8sJ6m41PPMHhxs/7fxkifEbDPNsVDlhOF/N4eeNKW
Bv51Y0KE2JgBvSJBaSl08cZqXj29buabG6vOZQDTKAcnOamVIudF4nAEdqmlVQgy
pdHMUOAsqIZqXUaGf+cWRMq8E6klT74hv2nHTCmYzEtELvhWjYTZRdnnDMy3u3We
Crvgd1aLfFwe6iJZnOc6NweQHN8olK9tq/1s41AjZmX/wZLhfbXY6rVUl7XUK4Nh
BKMn8z/yAsU4mWVnFhalY0HrsXYm5GBhN/Qvjw67Y+bEzZVqHhkzddjciW0uLN3x
C1obg9Eta9hyiKg2Zz3cXSCtRIJ2+AlfJwvyuRuSC7fKxsjm3YKaGi66eAudfhAL
aXyxUaiHd324jwKxnwDp671H9sOxcBig0OdtTnpd/QkpW5Arl4iWPnjmp6cDxyDG
3Ipqmr8FIt0++pKODJltZTEhxC5C9VNAo2wnRhNZ9NkuCJzNb1thizgEXkTPc6LK
xM5RaMxmhrn+JE+ID677KK1D7cYGD1homS8M/sua2U9AgcWjzA5HoPVzbYKb4CIW
IkZL5xhSIGCJ+6SOoGe7mNgDSrrH7ziE9SGgFHb8EiEcoHM+yHDI5rGoMkHrFB/J
qMsvUGiZP8q8xpUMb0iJ5F/uQVmEb9Tcyt/GoTlaVccUwYuXkLDVZYIQBP4mjBB3
+xLnJ6aRzVVk81Aarh3UTuJvRB37/5XoLF9WXpacFvgpRTnee1zG/jkBld+JBcgk
97ungwdqP3xxgT90RBcyBJ7Z2ELPSNkvPxnvvJivfQSMU7gOueK4MFRV1VYTb8Ay
TdSUZvYur5Ofw8QLUdm9X25ckoUAsdO9OKM2xDJyxjkSOCJLmHdLiAvhFolHaV+4
fS527TylPPbJ5VUgSpbaRvgK7XgnQQaNBMi+rzjqJzlFnBHqXYvhuSa0vf2RwSFo
NJstzxF0koom6ynHx/jteTRtshcN1NdoghzT+g3HpWJ+C2CKPCO59EgF8lI9LcNh
pZ4qZTz8pqEVs8PZjJIOytQ16LF8FbwWUdR1AufwVRTa/nqPQw+cG8btNQFmyOoT
e04y0qs3wfZl8oBIux+L4E8ypODQ4Z5+V+IpNqJ6pZNF7Iv/UIdesJSHcBeA9tVh
JzN/3afFJx2+rAwEJV9gK/+qkd15EPc+d8jsrZhpzCT6bUgdPlYH8OzBcCmA50NS
FV7WD+F6hWiG5NFJhYQoeeytrAW2jQkAXYchILRfNvJT5CpKq0vuQzuf9qncPffS
0yCEBHhBlqrq4lCva6Dp+r6ufiYHhJgo/KBOexzr+4nZTYSuD5hopgh/g6NO/gbR
FY/xWkhTBl8ykvkasuuPjzZBc/UDAnq8uSl+jKTlsDSN1RCypQPF1z2DAQZbhvBS
BEoK0+XvXzKGL5Rv21lMr5vLC1vQ28lfVR1bthcmQz8PA73Im72PMsUQwLFG7Q5x
xI1zH04Ur60NPoiB738/cJO4cQuWeUsoLNqtjwsd54rklXJzCnEOYKNY4H6hlkY0
zTbg5WMeEX7WQViPGuF6lr/+XeiHBKE7QuiRbc1oqEUviyY+V9qqeel5yi/QxSAB
Q0jM9sPD4h5QQoCAqyDzWlEQYDPwBMAXt5MRE97x7xJTIG8akwXQHfu+kXGEsyRq
0Pm0nEFbKAnvnuvxGMp35G9XoXJgcYP8NJxkOjnjSxVnEvfH7wjtvq/h0qvV/nep
DP2pQ8atAzH/RkBXOiUs9LKF6FPTbAB6WOoML9GeBr9Mrka7APSyy0U04hsXQVR1
J91cWKMfvR0PD8EMugMQU1aNsaU6eqCTG8OWW2tsOqtGbtL8t3cGN8zA0GJ9sjYX
kO5VdyVP1srtnoDsOCbTUns7xvoLSLQcH4zllX3777osFrfuCpAFG+R4aWhirpdA
pGBxZdiw1eYmNpWDS31RWe96AXVjd5DjA8gUY29PHgFdGbG12y80qI5bEtxo0tD6
ljMvJDOeGiqVqK/VyBmIHRaF/65mdfizi9ZoecNdY/lsNZIRUdHo1tPg9XciFoQ7
dqECkuwaevzVZIXltjad560vQyAeTHGgzCX6tXFil0g3+4hvrCjAd5Xm3wYg2eQx
CuDUlpzBqBwSjFkARAz4szjQWxP6hV+wZU4OlnzwiosfmmdruEJjIVHz3ZlRubPt
naec7nzuuHOtjBbQs6HkPo3kBJJnKNRjLjCl2SgkeeF6i869Dc3prJRlsttZnzcy
53rb1jv2MA7RLUqgMk2kN4EpZKx2BnGeomDM/VZTURODI9rQRH0aE3PbF122vo8W
mmMG6dQyL2NUYG5ii4Pl7GOBlRndPSNQFqHnR8OZZxNNMjpNNtT27m2J+bPitQWD
OXHkPC1vzW1SvrRexiTOgzg/ExPb2iKIYTphFl+LRJ3ucezjTS4aMfLFOkoK1uDX
q5jkeEB4HRlFq2C3dR1dl1Br6TH+2DNyb6MqtLbtTLgb+8jDMftMekSnbsR/kD+Y
lt5RbQH4xCpHkyBlrCb4bKb76vFx0C9Dtr9fwnh3lzf4VskAzHjOOqkh2CZ0ToKu
kMkOQDKiDJ/qDWYl0+1n2z0Y+lwJXQsnn55GrQFuP3doMfCXIxk0F6ojiTOK5fo5
KSqI9WvuSRyOSujY859J15BKC44cwGUGPw8YaYQSGKBpBhuMjjF3xG2PkdtVlTis
K/8Nm7Ems5zTKUY+OkjHMgeXHoLVdb/hm4doSudlgpAFVH+OsTk1ciM10fj8E96O
s0giVV3t6Z7BSA4tRSrYTVVwcYRCRxUSuuFt6R4GxT1ZM5tNzi1AF7xtpLiYJrjZ
tvuEfs0wNeSKD9RNZRCpq8JaMyW8bwxZGvcy0fDBo+uOs433nOSG7vNh0miiQ1WD
y0SCtTbj3QKHQQntXhJJfLJZm6FFBw4/3FpNMcKqotXRVwCIJ3Yt2Lnxci7eOiF9
I2cBkjsom+5IMMm5oPziQPCo4f3P1gDdDsyUk5ijA6z8Tbhi04Fvzpjc/ZFAq0QP
WhcF/aLRquAC/JhuFZeBN0GaZHpOQIw1pQAgSbRUey4LcszaJNXBHPCdTYkuQSwh
nIpPhrdEPgzfWDQSC1mZthmE/IbhD3X2xT3PoHBKCn46Dizr5fXfPtWIjm+mw0UM
1EOxrEZc1R82lC4DcEgubYTwLhYcVMJdmUoiRxuUhcr6p4totOOLxU/jpn4FwDRv
yE3XxaRchouHshPpW83BCOSJX60As/GOwOLy7r6Fxf5y2x1D0gv0i+lO3MV7jxjl
wNdUibLPXUpJ0S7L1V2W+x2zDoTcLynYtUrHJlnrQ/MNLIPjn+M4Tn069XqWrjDQ
RsvhhiZz8nWE/eAXAGJyCaqo/LzVyka97Sfj7QezVG2OG/vMUkhKLSqrVCIWWbQ4
2yD/B7lCvPd9fbq/s0iW8lcvjSY0szZmZ02DiIMrMcmbVms7pgrJdapwYOKZMNpI
ll7XT39SeX9visNFEaC8iiT0lf3J4S2y8A1i69hA/CK6uCkM2mn19Uto52sx6mlP
MBuK9Urk4oVnW/Ik1Ps0DM03zW15xgteCScy7vZH/MNUKYHpUvz8qJg1Z6Qp4Aq9
dvf8aHcnRcFDexuogmqE7xnI9ZBFDZg65jm7Sxro1JMqY/noCL3nHxaHG0i5TEzS
+WF/QYiCfIVJVUvRYt7mQuq/mF+uG98j8iZagjSl+qUnWQKoMwTImCWyd/O5Buru
BOPfP9oADco4IsOpErssGshHOi1wheLTbCSm70s/r03R++LUcygznaBoiTtYzmR1
3jQzJ20RQV6uJqVhqGv2KQ0H07ZR575PP6sD98htkbsMW9CHsZG9HV8jLTZd6hy5
JT9tVAOxOgoGFCaGn1ZPlssVKiKqgMX6z+5sSoh3/2p4BhMltcRa1UHMZqJ73YJb
6bxdRjD9K9pgQ40+xCFGtGlacgcf34PdUUKxNlLlWS2vABkRaXbuQHwrsWiVm8DX
d+hm8pPhTGiZkx3/+3DwmkvZ8Gx+JlUay/MqrpKOzBWhP7ib4qOHAsucggi1ScqT
VzUDdA2HKtH9h87nkH4EIXiK3p3ob1kc6pj25R8q/OujykGQS7h0JoxQeUnyMo76
zvYXjDyyMZz/+zeQX8v/j0UraDo2WtxkQT6aaMmp1sulzsD3It7EQYEexAGCcHEA
myYc6lTBZxOWxoqrUqHmbrM+2dh6PSm0n3m+9Qc3f3o9hZsqBaJ1ScnkTKdWgLq5
tZ+uNKSSEsKOhJINFySD5D0QT9ee+aixx5uNwCL76JmzsXuw1n41KmPOFgZumNCv
vg9JZzKSXd3a3YSNd6sO9oee9QWnU3kpx31CiOIG5EdS9q/bUlJPTQrsdhxgS/uz
+HWFMm7Q2icmtooqcD62ifOdYvuJrvvvwtP7Pf0awfrtmJAIeobyo4HAy/iJ7UgY
Jv+G1NXO/Ddc8ShRLBqU+4JujeSkwtsHYIagPlBMXOQfy3x1fvMllh//5Ejsak+i
vnbHB1/e7r/CQNhn/aZ7QaEFMBdmrgst6VrDU60jjqbxmEwM9lQtFGz3i5bdyjZ8
q9D7biWP9EaZu+M6os6/9D12z5o46E4CEJY+DYnND9PhAXtFTGSurZLiR1qNcmOc
sVxksFWCHpWzfP0fagkCHLhq42seZ4aAfg2P6QUjYxztYqETrj2HfY8i1qEeRoh9
0biG+sRAnOEoQZbfjBD+h+md+kaUbcy2IEdixg78gQ9hBQkrZk8LBVntWC8FmHvU
nbC37EXN5VCsGmF9P+hE/s6kJG+MeMhdsbnEEXmf2zWO44/MbudZXzmHJJCX4M40
EBADjh0kGs+JZS2yX3Roc5lDfGDgWqoqwya9pq5VCTGadg0zhyD6LwtS6gv9veRR
5z3c/GSp4Bf8RWKaRsvEExt1fID+ooD68MEOHzF3PiDLMCeafF1BlP0/spuaK+L9
xz6dUnXNyOzVgd0+ciQkTf8EBCuHpyprpdxji3ZCVwlEqoTR93/5ZtYDl08iBOuh
8Jy3k3+opCymCPa35W5/GCeZgU1swpMciCf8BnUWbF8JrZ/PxXe+DvmmSIlwCltl
k2paW4cN+lwW/daW2tYVXJQmQYF/lwHWpBVQUFRKmYgje8F/WvrZKogFNuPPBlQO
lxuTNvbKMKV7EXFXqcSPtiLoOiLPNsC/QCU0nSjVHb5Iv0itRURwfYMco2+DoEqG
oHz8vJ5acCvulfEpnqeEe3E8RxSM7jTb3dcDx7YY48jaqbtPto3lHV0i+1CJcWqP
yjEGNZ1ta8dlMBFytl8d5Grs4pwl3EfIFe92dy/hgaBtoE/nIMGqBKS43wdV+wKb
x9ItUWsyS84G5b2/fkJ8TuQzCX+pPtysRGRqEJ8Q5HtSM4r8IG/3SOudoEBaQ/uN
XHz0o0coFVszsi478S2rFf3QnigWUkxjHN8RpgbbXMh01OKKX2jHRFxbVVJBR84L
SicdkSnFm/tzQq9XXGPGz10VGXkn54cO50Vk98+6jjHW9zVIp8Bfm9aBeq+DNg29
doumSXXgti04kwGYFmDmW/MT3qLvPhYjx5sT4TDLaVuvIbqZkmRNgXzxlkugYs3k
mT7Ne04B5Rzd3/n5dDgC6Q7rbO43NlJ1Z3UbtL5JwrQKKf1Ouy5j0aNZ+msBMWQR
RG7oegL25ksl5YAmjaS6WUDaxROBHuA7zPH232KU7lopnVEo8cz321o/Tucv06KF
q5JfEj+tqODN4uKm8pX2FlsZBPGo4pf68vtmGyfZ0wQrY8TD27hBLKYovqleBZse
6yVoHR3jxLjry5AnGQjJi1RDSorOpHyCgC/IbCC/r/lcs5jUT8zNtxaFTRC5nqVz
H9AGx/4Sykzx+d5ql+V3TJUvOjqui2wYlW2aE1+Wo1HNxGNYeyBwriRP3332XXyK
3DQKYmfLjOHrJxpqToW5UGTxRAj1HH7rK/D6xT+rLGL1z8jJHTKrs4wj9UsUTJ8W
Y3xAnpMf7oAKLxDY661u5YNCSsg2pKI2P9AV18AdHw2q/TxuReFGoo2PpyGiTv6r
ReLAoy+pwm+cknWP68qsM8D2fA4XatfefxBeZrKAMyIRAXlmABkf6jsOh2N9fahL
84405+FwXHgXdsAkjn8BMMBEqjPyKutQP7dOWyeQgiWbFcyf870TMS79IZ0cCbzx
SSoNSoBQ4OgotbMWxPvtHhQqJO8FUlYbLgTcVpgE8c3pi52/Ud1EUIBoN7d696+7
t602vsBjqNqnJ6n4lZhcazAqTynon0jbBEhsH+qpHlMENbELvNYfhyMvDZwIWgzx
HCs9fwAKXRDfZ8CVjRBwVotUOZe5VapNhZdZpxBgPyyO0z2JzfCrl8M7SMI6JkfF
Bwq9hWgFE50MojiBUNazR/60FEVXlOiAUJ/QaoOMKQr8w3i4j9mowj4MaAFGDxB3
OaX/7YYVu+kSqsW95yrrPhQHlh3YRILYj4I47/T/2iRXbJQ8U12Rc4oOg/V+M463
xGfHcjiKHFIFyvuh6H7ueFg3exd4YoDOPTUnqHpbkRj047ZdMI9dqQaYAq4DkAJa
PHFW4Pg90HlHkfE5412wXTRcZm5Po7IAHlgY8hT/8SYy2ekuoSIC6VPps+SbAjlh
XaK61DpbpEWnSAfo5GF+kXvfEDKw/x+VOUxxC3PZBi++aYRWP/JEpcwHwnIM1gn9
WS2bWWCfm2E17dUQsPcLxAua7ye/LNTA5R4lUkwGacIDucZ1mUnqiSruLGmgkVb1
jQEtOHBddDlSr5IWwk388nPtQNBsiAlDS3j1kclMhBZ37Sea0VirX6HAOJsu2sT8
BHTpuISXsqUgYM3Noku0p7E+gj7YmX+evdoVcpfDf67DpnPbX6MyKegYBFbv4jyR
v7Y770D5NtTI6K0yWohjugMow7p0Jy+LssxNRyjfZjpbG9vkEbTPrYbPtAyD7P4d
PWn4rQNqZOIgMQDrcNmEyda5P1NnWVLLwBA3kw01jmYOlyLpDpS682EzjG4nhbjy
DEtZka6DKvmEetMI40lxnrFWryToatCXE/NJq3c+rwTJ1EeOTelJ7RHMP2UGKTmW
1FFUjRi2XLwfuzebWjejX7YQZLQ7uNdgE9E2CXCtmot+bJCRNPPtt3pwvMGp6MHa
IUaD0J1xUUI9wJOI4F1dYQRqsvPHb/s7YD5iawJWHRP6az/qfxvw6s/EjTnT+cwr
DnWoA++zGY99DEFKHln2AVeiiRSCVfJZH7ZhUsaV0r/Ogoa/qA5h1zp9WWmpUEqZ
juymKTcCrXYg9QGBr2g6Y6yEqJmsAMs66HoqCW67bJwnVP4y7da/k3TAM+eyB2fn
6CFswWohddY3zzdZk8jsDMS7GJxHV9CtnImxwGGNc7vcfxTH0vJI5JY+yo9WxYyc
9AjDDGW55IVI4oPcCGp5Q8AX439ueiA2FjFF+h2xgaCuuyVQnVCmrTI48xVwPSsG
O65ECYP/Jatj/mL8e+O8e3fUvDi5GmukIHhQfc3YOWMnhTj3FsUNSzq73mGxXclf
m/km0TiSDC3QkxdN2QQwGi0mWX9FYdbJRLCtn8eLcEM0GPk4JfPk3mDg3691iqKT
pWSLNy+JPRIKTYFuVbQRGD0iZjdhN6LAOz9T2z+aCKNURNJiMy+D7N5Ht9gGVpvB
rijewIu0cFBo2aK5WIwH06W0OM67/W+QLwyXcSplP3wR+5k9+/6WB0d6pXQab+fQ
rGsH/HvWn6jW9HKzz2KenOBl7Yi7vs+51dWsOAENjVl9jm47NzUOKmYP0SNn1MaG
P2yN1XbursXCo9XhLi4OEfIJfO2YzI5Bycmq0lolW29rNSN4C2vHuNyRjmdSlly7
wlhAhGPGYAJBDUZ211fCKEgQTZcC+JoPi7+qYBe3ErM11504WNIp9uzr5awBIBZ5
WcJB26jofBJgPpIAXFq3nh63Mvd1YOn1BAWjb3ZDBeJbD1QPPDTa+ARAYxW/2HD/
gNTQdAzEh7xCnMDtCo1DhoTMxYE67c//mrvrV2u84EETQWzd4ZsukPQowe5iwX6n
+xEy1mJNWa2ooHLfKaUC4L31igr2LAInr09UXZ7ZIUm8ga64MqGGMISbdCV6iYUW
wP1nP9su7s5vyDfErW2n1L+ZQ5diGxiDjgLI6c8MB8EU/rPtoKlK5E+vJAQB7NaG
Vweyi/5M+awyLtUjT558I8/14yvLP0hqBZ6dpj/MWbQWsixDDQa5MgjUluKAuVRX
iSyDh0mvsMSwrMIXJ2EH6d8aGK7Md3ycEi9C7bMzUzCdK+K/6JaGQxDavB4lnztA
hKrFnVKwgoPGHauDNPkIZ7NwVJF6iiATi84/5Ya4d0NVtm92T877Aw7JB0yFAFpd
r1P9e41qXKs+ZmT+WCqNQpO6+ZvBID6IrrYvm+0C9QDblmrNO34PrsxqSIqejRyk
PYYNk1aUtSulpas8mSgsmcC43vqCI6RkR02iDLP/hwJQ6Mgh00iwlmQNQE6wwwoi
c4XGDkRKmKJaKLjPwLkMs3DjFQFk05EGeKbHJ82KTo8OBO3sgi9JA42zlfmvC7J3
gYry3BAmSSBiW/dpBhDCGblAqodMByJmwyrBZSfHf2rVwHrQhLIyNDao1tk9pX3r
2K9EYPYgSUk6Dq53CDYY2K5FFZFYXzvOcaUs36w6X2Y12OF1CoF0/DBJ5Oh6lc8z
5B/nVoOpsPsdEqeeBocG5KRZljlyffUVB55GB8QfaigdjP1lijcqdMsZKM4Evk6v
cYopiEzLIvKH5SXQASmHoAh2AomIQMqaPOCOYRxrcgq2OQVmmaV667EfS1QfEbpU
z5bORBfAJgsj9VW436prUzE6yVQXlwQ3t2cR4s9yTCNmpKhokzPcC8xpH21ogY7o
vRmp/6yvsKXAdIBAKlacEaDLpeRqgwPR4vNmee9zqeMPZtDNQOoIieCvI73aK2ml
3NtYozDwPUjx+A551oSCMFbjBBi3FW0w5u/YF8Wn9wwYfslEyA84TUBHJncpEX5x
UWl/Ch8TaBCO8GxDcOJszrAglJds9nuP2+VwUV1boCjJ4jpxOCiPifzhV0wyG0CS
BswON3HhqCAh69bBVZ+E1kU4Jq/G4ZeGCeuARuWzaZYof2OFt7Ry92HEQZ1b4vqp
ZukFriLYo520C5VR66GFCELV2lWL9nN/OdohZPA6PeDAr5mL97nxTZogYPeK4kCZ
qBFVOEtSLrlFHq8F37I9z0vamhK7AXXUtxsIkmkiOwOuP/HzmDNV82COpKGLKvYV
cr8YPLC3vQZAWzzt0uLtGj23rPvETS2elCWOatz54JY5Pa/wvmch9wTLBozjtRNd
kj9Xj5AbKMfSoMPy2qey/l04Ny/Ba4aRbB/rhrCvLJB8zdiBxE4KJydlB11yuG6w
gX36gWJLLj1YvgVyA/c75q57TvEH1VYu9KBnpNkQcyW+CZIme55x+swSVIFKZq3e
zGfN9AvdPfG/xJeodRZN6y8wnzcJZ8NShlSA3sB+mvdCJQDdCbry081bwxrI4fjI
83AbY5u3QEpYhVa287IYJXyzTjzCj9JsPdZZNSVGKeUDI4jl6UG+gPYVTdQynVoK
Xlf0uqRC5hg9hXaPGAkBLDZo1B/X1R1zy6zlyYskkyf27Qrry3Q0NCo7qXXrlBeW
L3SNAY/ioV67nRNWERp8I5L1WJpMxGL0n1qDsFxKpYuUapaugtGo77FvU4nMm9rD
NWheEeyjTc5AniY82La2gYOO82NaQyFIQU4TsYWtDy0YUqm9IyjWbWyN88y7WMC7
IMbeH/9mpxf7cIbx3w0/aR+JIviTm09z4DnOaG6d/s9WX/bRSJhijrNp8d/v95mP
/MVs/bPb0DiNmsOJZ09Ljh4E3mgvf92M0QLJaha3jfWRq/b4Nd1RnQ4Y3jcbI6uU
4rSf8vQ+XBIqSojM9BYa0bHeLt0fEbZTi0yKPce6dSSHn5uXI/Mi6kiVZ79ZNAWj
2BB7xmas3k20p6qMhDVpRweJvNHnd49E3sMLM63jQymtoWinMXLRyvEz8MD+siMG
JOo8HdpKChRVyE3r0tJfzR3Pv0jSIeEoUq4nr3+jcwQMmoMxgD7LvJ6Cyd9J6RgZ
itf1ytZH2U/4TZ9kBg7BC9cEj2bDBTMbv9o3BLMyk9p2xuRt3/TyHdLoO5BJ7hCw
UlEFuTIfGZlCpqhONepkTH8nIG8JjGiCzL3XVrI5TXoAfix14U6MUX5vl6YiRQLX
yrh6nSKqDLNh6AeliFwJY2I8drhl/swk0ZoBIBBrgjQK1ctL1N4x1BK7ReNOL2RI
5EqEc7ognfjwTDbLc37m5IeNps/f19humMvuEYa6WfJrpjCexCGg5iTcXoTVamZ/
lvnOJjeojYrJAVslbFZQ+EL7qQPYZNCWJHsN5XBWEH4VI9IBOmUJOUF0SsK6eN50
+kU6zwblQG/vf3x8xzr1ZuUIW3qkPLGq9zDl3mw6zaGzovr8RtB2oFsZuzQhVWd2
GlUjGJDlhYSEJKxqxKKbwNuUMGC3c6rAIoGXZVi/RkC1n/D1cpqHLawDw8Jr+pHe
E5ktbclWSyxENVDnSXzFzJiihiH4rEeeHehEQpwTGZgCjBT4gYdayTKHR9FcaPn9
wgb5EhBwtpjkDF7gONXQLiZ5agpUn7Xj2QzLmzc+PRzVy8sYPozmeHOW3Rl/2POe
NHnBlrV2yJi+1+ubVBO3o4ESnYvHKhZjuGSk9rQCkDBoCQNjX6+tfA25ldqaG4hF
oE8MBAQqJb5SZc8krCvWlL0CGBRXmhVB288KM1wWATXVVkIp69cDvGN9tqaDehkc
bL1jRjZzOf8ODo5+0SHO9+Fklfq3GeXjSyrhv6xGwLjpd8bJJswSAPtKdht6wzqz
4msLxArEaK0sZPQ7FxlFEKUQpuCIpWCKkXodEhIzNCVmtB4i6hQ1B4AbuMEGH5Af
iIP3Femlcow7SfRnFuLiBtQjwPUAvki7fwD/g9aAZVT0ezyJDIC1cUIW+qFfqu1F
nlu3g+ZZsq6Z1bjYT39NDEs6IGByZSySOvjXu7aogfHIZyW/HnZKPqd4dssHrkwU
lIx0WepkM5z0gMB3JAXpQF9f+DZ3HO6oLNYJmVXdducaVZUM+h+BEqBoVlxPuijV
KzFbSPeBOOEdab9sqS+RnIzehWmDSLwE5b8Hmxmh2krlDCfnl8tYJW1ptrTrZ6zy
sEgXeGJ6ZUbQZcNlT1sOT9uNKPjq0PUAhqc0tURFxU18RNTEc6xrZstPzA0f5iml
/a3jwxNksEBFmY4kC3PI0n4P1wnvxofiu3xzMeX2Pk5Hk+rpwqO7jTHweJkH+Kiz
9gc0ekqDaKsr5ePSz4AHOpdBqvFdR40GnpXnlJwv0SENf6bR8EFUzw1Q3oMgLjby
Cz7Wuq/8UUBK7ICVkZJxrfu3dP5cMwcyd1w2hgneMYNbAMBuU7LR4WmqMCQFRMSg
06wxzLvqjmlWo3D02E9sJUaf0KOFXp0U2/2UJGjaWA5gBDVCCCTiaC5MKvX5Ay3A
XrHJtca36GAQ8GykBIxpfYJs5/Bj+Js9YPREQlF/qQ3B95AWDAiol1boAHBauRf6
03sNLqJJKE4DzHzBxM794EYAfRUSyW++4sPlIet2y3sBpAOrCMpsZau8MZCmyzLr
VOw5jmyXxz60AbpMc3wOUVKj2Rsl+5uC75Jp38ZmjBbEuhqpoCrtmyBFdq8Cu8HW
DMzX/4PjNQ/nSvjk/EeBZOASK6V2IUefzZsZWlchUOJ7mCyKEYg1vpcSPnFSbNWY
C0HBzP7l2LMc0FjGYe7vRq6xIyCFMs5Vcb7dswqmj41e5M99xKLc5+RHzbHLRxvN
F+TZjQ2Eqhh5xjvkmPR3B2tAtts6sS+LhNm8V3DP+ojO+YUFToyIIyN/x0VPFqEM
U8LisqZ9exlXYALuHbjj0xJ+bNXduPvR0Ziqj8ACgKK/0DqUSfkPLiZWpF1ayBLF
pyPk08OBTJicFui6xivBBwYmhcNIsGSHxsWiRyAe4p5ux4F1uymTjZtTFrmC1Hrc
pZQ2akma75JUzP9F9bnQSGGB6dl9BYq5HaZpt66EEX4vCEGm6uV8sdQUaFBfpYRS
bWLQmLbNXRW6ofPRCogR/locZ8i5DTlfNTjvzziHY/poIhB08xVOLByf1YwMudIy
GMikD45t0wliP70BNLVuFtM0B0/004FpPcon7VQgzmkxyMMnFHyEcqiw6UPPzkiM
1yZG3LjeZLiQ9fa0tBrSAkifWHmxqUXSccH780HMf11mZcdBvjlL5g7squKYGeDV
tYSJ1mVrVyQAuOLs2p5f5SoHuhvqGz6udxGl0vPEMd2aGXdt2UjxkcNFTIAN4Jix
vpGyKTlbb3VdJNwIOkRpMQqo4+TPSTfiaEnL5xC+CJgLz/SYYG3z+NBY6yvlHhZy
Zk8kvECG3lVkN3QKg4GjoyicglZwiseDfD4ZqcQoucH6bRYfbs2QwuPXDzioqdPD
8JbvyCNYCb9kPOYolCRr9ubtggfZMZA6y7uRDIh3Y9/Cid5jw0XsJsG7CPz1yS1y
pbDBguMQLjOboZVpV0SPLrVfbLaFm/nfgoDGBCDaT1ChZ7RB4Mccj8Wm/FEBAXxd
H4tszNH2aiJFE5BhqRr14iXBV5rw/7yBRKbsNGENi87FTTL8ndzUzBIwln7eUZNk
vDC2IWS19XV9tzhr4iwjH3VEk60Phb9PHICMphNraAd5GQ+kBtxqI0LuFucysD5P
fjmkIny3VXUGqBl9xfVawsYa7j/9ohMZYouUr/QWoKBHFeuY1EeH6x8XrYAw16Dk
0lNjpBxcAO1mKN3ZRV9+kwyN4XR4zx4bd8moOS1D/rF71ddkc+024jbvkcnIMiDr
Kvo7uDXBnp16uR+CmsPOez5Zbe5QxDUpSCNpRkeIJAcR7O7FQ125fBVvARJM6756
uFqUJMmU3Cm/goW1Xv+f2SjUNm9AWbI9CH3+ioF3fd8JIbyhBbOWGl8sMmmsEf7Y
mf/JZksmysBzh7qiY/s6F5+xNjW+B3A57NJc86ogjFoE8Rizgc5qQojiJAbtSwbA
Qnv2FmS5eXxNZUu9c+6cTXk7g8TkgWHrsPOmbfDWXLHvLQUrPiYA+9qOzfyWO8f+
8Pp1zgMLHesCBRDnEpPWtvMsDWPhJ+nE1628eFeoRVfn1dz4f9KpxTjH3+bplAlO
Mm+6nSfKZDS8XiMzhPwKlY4O2N8n31D+0KdfCCVFOWhJEmPcgg4C7UomIQ69outx
TDvzGOBN7Ly0aU7Ms1/YATW+/BIHtRNskHDjzsTqkPfU2NXt+ZL61RSuEic6EoBU
6hmEVtGK2nTTGWMaAtpxeGVaz2HpU6VCZOZQwcImexFRwXldPwtKuaLiHtP1LXF0
gdxUJSgfRZTBb7j8KZxGe6i1ubctbz0ppjIsPepVBWhgYamPGyrBHRPp4cmXdIUL
OGfvjHE3TEYIWtEUfGaff2CLg6g8QfARvhvZFYoSsnHdq9+oi71aKO7yw1tZvwRf
ARojJG6xg+C4IECnYVXvjpFeFFrWmUqTqtDSKYeabi328NmipqWwNBTrMTay1l93
N7ccGqvNn8s+yeHwN4db9Fw2g2wc3ZB44l8CLs1fuOBXK3WSTg0csxPZ4r0cxjGN
vc/g/cS9IjRcoPFbVmSbL4hAORUxGza2xPj7hpAjgQYvqg8LqpcpR2DzVUfl4O9Z
2r0brydRkX0ZflAcateHrU6zJUhdOIs33GuNVtVCVSFXFebGW+yO9IIuNr4XV/7J
QLHwVfm31TZoqwkrlMBNiYcJQXjV256iOLncb/ViI099UNmj0VgRh8JWlbT/eoGU
PM3VCLWFLK3tu38HJD4B7k4XgWIKxq3CPbcxXyPpr33PzVy6F7wpi3dQ79Q171IB
j3TCVWsAu9I5jLRmrZt1BYzSGA+/N73T3sn0xZIEFGb7VvD4Ft18m9nJmmQ7BPv5
TCoB8inx+KqEKlFNPWRBZ9Unrf3RgQ8hQ+DB5kTHy/AxZiYQMEQZNc2a0dJYEEnz
bpTR7IZtBPHiSCNPwK+TAOkfOyrm8/6TRwOh1/ThMCUIEgBxUqRyXVmUjwzWjJJo
lDDKKUWAeZywr0JnMdaM5aay09hKSwWkDELHVJp66UH6ssFWYq9UCg65q/bY16Xw
LEUoYnHHIs/sT2IDVjMhn8cZeJsKtnRYzQUEwZeh4YG428b8Wjd6ur9znfURuvKk
NTpxb51EtUvZMd+YQdw/T0wBi3+muq+N8lSwLLvfe0KbmV2HHHk5bZu0ePIcxbRI
VwoFhkhVdrXMYgOvOTEkGzHYoZURtR+W7SCk2JeUwfasdsgfIL8rPMCLhDdT8yLq
IhHepYbWr9MJXE/nwxXFR/r6Nbcq73X3o2abRFTPTuWTXX1Ooay3Nh7EmSUzsBMh
Esvlu4l88wkw3quHJdQnrOzKUua2XDtwXH8z+5bEo/+iYwgsMmU+uqeSpNsPXXon
Kz9W9TOGSjUrCY4ewwMXq2UfD6td9/e1MeW6l1hxKttFvIG9uzAkiX6p7ONR7GMN
YgLWkMhBmr66SvCycBNyFicmA9u1v0cFoU8a9STVJSiGcWZEVXfqDxJ5G5AhDzQw
D0EhfKatbMspudOs4F3VwRGpkTU8kqsFTRFVa+deV0FGkbFwC3Iwpy/mKm99cdkF
W5+OHaDXeSKROGK+jTibTQaKSlaTlLev68ui1/EfVnQ/Ugo1Dcg/K1KTMK4Z5vkP
VxQOMBkGVh3EmqtpvmbqXersJO+jrLQ+LKPHXCOwjpb1c89c3DsUi23K4QPalhTP
W+SMlWKT6wR/HwrQPd5EEt6z0E/0aJl9qXUHaEbp/y+ewK1jeGRT+nLCNZN4sGF5
072voUZ2EBgRz8hbagVR46/S0ZJfEbAMxxxDreUCKPJ8nYg05FsMJh1iaKbOg9ap
HumsuvXQBZ3XalOgEMgniMnla9QSelqs/nCIHdL1vdMM/DVklGeYOa8Kbc4dLLfG
89aW6LenvlTNXqLrnHj5nhQNpiRU5108zrlw9eiTCaDFN2u9KXp9p30vkzyZUOQu
NmWt5JXwrizCt/V4cso0KOMhzeVQtEYTciABBP17+kM8x26HT4za30lwGPKt7VYh
1ptwQcOtk0nMPEqfYnmGGM4fnuHZeXGkpzpYL9VJQjoj+DYJ5YsM3sly/k2CdEms
TWSyYFjHIQ21hF0QupODoUEMcB9e3BWICmJPNAz/YPj6088uTqycVo1efPYrnNdc
2Cd9kCZVKSgAhtA9XMbDQ4mwXZRNVNPwEUNLkwCMyNnl47MKz1wThGEgSv2PMJj0
qefzqsh2rZvU5fo6Hf4CRHm5uZc6VSCHO55C3s+m9LiGJzaMcm465NyIGikgpseu
PHy/kI0gjS0mBQJhGS8X85gkIHzMAQg+gTcQXOppmpO0Z7qP5I9TrqJBoJ3WInUY
ondhBj87euN6kROOxgfirGSZR6ygePJIodtCUssBPmBrYc92B9WQ/xigc8hAIiH8
ib8bG9Vs2gN1TljxIaIE9F1yo5tpduiMhvCC1Uuriq5DfZwfJz4oKekJRkpLoXlr
mckzff5ZNZHkJKZc1jpZrcoDzw5hz7hxU6T5AFJtnerDXcxUa4N9WnHq+nl3HqaC
jDjkb0oVaHk1nKmEM5MoTXpOcyQnrXk1tnqECf4FgtGi2mfAIOa0zZE5+VPdN+9p
Rln4qqs0i/eNfu3nbFwM8CNl/Cnnv8jSi9Daz//rbyaUaxLvmyH32dnlc0Ayuckg
NWtkky/4sdHEuQrxzz8uz84e69itPxK1PGSwfhHAmHypfK2b+pONTZoa27NgACLZ
a4z3vUvIcpoWKiI6PlYOJaRXk4YczpcffkynuxCrqG4HJI3PsO0nwB1ggE+QnRZm
8TgynXW/Aynh0GEmaWOATv3UTDApHfWx3KLmVAK/IsLChWBnZwiX4uhVlo/F33qX
HnDSR5yAhqNk9fyc87MUwN85kRyaf+e4KfaZmBsy3HJjO/6uDfm2BkecY7VHDlmU
j8H+UiffSDLF6YSfSteJoKeZxXc6b78mvgeffXHqowwEirj5VtXyBfh8myFl8ShO
YngigeqgUkvDGCAXZHEB1x6GGZ1DzZVvVrz0oTBOvOC1h43va6WeSpx+g3CbA84T
DSfYDci61Jz6NFmHqfMXiZjlHE8/MNOdQFCTtUCjlXHt8a6XSg34G5oBMQ/CHBwe
2itsjmA0NHVcDf8fJVxBusDXSaoG0j24LUgBq+QKvB/PYnhOzcVmlZYq4QbbQXbL
x6QUQDIIUVumq8Iepw6lbHFYvCeioGQJvpr5xwy7h2p3XMLWKuj5sPxZhgw3gEyx
c9U3rfVeL92uUlgVFcNKRd/WX62YLxRpwU5KUg1WYAViNtc/zmqA+S+yGdP8RDwi
l6aBCq3XvztAOIQqopSS9cQL6KuO8OLkSU6SMnyOSOsQjHopqIfYgNAhK02Ochp5
4MIL0/xS/FkP9BJkaHW/Lf26NqXkuzgXqffC6yKEr8DeyXJhDbaQH5Jshnd6agfC
q2lXAb5muRRzGAUY+GqrkYvEb14NaLsN5Jl+h29K4Nw01ILwM5dHMKVmkeJnyOyN
1C7HcfmgWjWsFs81ldyRHoG+qeeuyz0bPXOZhHfYuCmtXHRtQKywJLUf0SnT37Vl
rGt3lPFcvU7hUph1gX2xAbrVllQz84ufBDz5FvCQtoPw1C837RJfOQoBgHBcRwOy
GVr2gMz0QN27MvucWOuJgDmwArlMm8MfYlL0QNNDKLcBBBEJIwkbmQHoMAjw/NSF
AgP+RNRQNiMBsEGf5lZKH9Gp9824pv+RZgiQbQYZFQiAF97z5nZ4tpS76dzFh0Hu
0VdL4npDWOYy3Z7Ara4GYzWKC3tbAzoR01AUrkrfuHzKjcbXyux0dfpYNDjrB5z5
TBnFcBUhxK9xsqiXZ0pu8zxI5JE4Zr8z9G52Q1avmYIy28BDl3zu7HOUHkmGCF65
G8v4XKegSn0X/OeancKF5DdUci9HReGuD07OVGQp2RRgW9xJRVtImQ6XDrAWNgzB
lYo9gEVFZ6sT4RUpBWG99eEI8I8ROBr22WhECtGB5F8rDwk4Opwg1dQb2MU5wYAu
JGgcf93kwHgf0bKaHG1TOzsyYkGEVJci8//LIUGL+4y6SDJICPOhZmL7cQMuvhFT
MPLagcFk+9NutgUwHDoJc/0Elj0PYFmFhx0GT5p8gzLVIli6g3FKrkRGYFuBmYso
gjWs2elF2mkqavHP/vZ9+adswAWmKjw2bfDVdKy/p3R5aDa/LBkA83vsZktpDo1R
6FqPwddp2/kl7U2FENnXAzvTgMI0yxZJOGK/ZejXyE+P0w5pQnMV9aRGYgO5NNbq
LC71hSMl60IcoAd3rZ3kOuYXhh/v8neNFcfk7TZBM2sjozy9Fp0RRH8pi13me8sO
0ipopA/oWHzF0fPPj8GM9LkKgoryksDD6E6lQX4ao4GYyioBE//HLM56CRHJeCgt
jlVXZX3fB5GFvq/p29loMnjnu4W+MgInlJQv1AoEtFvXWIzWJN8Ak/F7SaabHVbF
ayeOgQymQ2PpKWRx6YCYTYBPQUR3si5pP9B+HdakJ4nq7pH9o6XiVE3kqka7att/
3vIUmb3VSJhqncsGdF2d4BmeTy1myodNSgo+b0kDTUuQLB2mXT2InfO7d+qpSc1U
U1yJRZzDnfXOEyAupMAelyr/CrvRjbOGOaU7q36OmgW/s54Yn19TkkHf0tJUyR7t
JyDQ1Bqajl1OdwMiOTA5NTgJZNkwNMsJZ8KvWEpgRwEcppwaGL6xi3aYdzjdNs8m
QuF2fCRUkWqjShvjJT5VOQ9JSKK4NPL3vt8YX+tJnBfXRkn2JUEo/Z9lJXeZzBlR
3QlIL0I1AwtDL5+tT3xvU8aDWRIkM8xd1EtueSvTXDWR9OZFSU+ctztHucR2KYjB
mPnRM37iRv/DTFcX+MP6fj9tLIXG6iKihklXTJOCP9gR3Ll2r4JqlL68hVxddl0h
L516Oul2P9BnyxPBWE8FPg95c12x9g0c5KbQjJs0h8TWfRtImHNPgmmZ+7qVOyuH
JyJJfHPndSfk30UFJrbK62Ejo1xi6jDTVJVkdetCC1VaHrQH2Gn6SDpYpBarIQjp
med/RbWw6UXWi9DNaD3lvf1IHX+1PIfgHSxDFhENUTCCa53EL7PNf5s3c6d/X/My
2gE/T67xoNm6BDQaDNJ33NXOuN0sdKHe/rNSZPozj1G9MCAKTvtCsrP8fOkbdMxJ
5qhvb1rx8jVGjVNzj+rrme6YD/OhIUKmwpBLkFzvMlgPijRRAE/kPpeYPhGG46Te
85/Ctc4/R0yLV5ZV2VN8hn7Sko8NYsh7RpFioHRUQibD1Uer+CfAnkIEJrFtVJGG
yQFj096gRg/eJI7wP1yXDlXNE+xBUXJI2lD5y16GAd1HZsbt0cY0MCA4c5bI3xPf
j1/UdS25VMIAzGxbzU+KF3jSxlxX7WpQCBOd/GtpsSSSNWP6tlzsp2W/ZJ3TMxME
gKC5hsEA/o1gApPXldJ9E1kwQ1pX8mHHlSgbvl0bGNpO+2XQBwbfav76WT+BmVWR
iVsvrKda6jQxbZCEUUtTTZRuyIUA/lvtVQ4SEmmK+4d0D/WazDs2jdtcSlY3tLgw
FP+ycoOv3maWklkx6uObT4lJknBAYaO+G5NlFakNYciEDB5+sRUdgzLgzuVpDIq0
S4QdemRmWPFc4w6t1QB6FHA0tyed8LAEnOOCeYyoNOd0uzLu0u4GUjaOQuHhhmXB
hTK9Cd8GHoYSJ9r5G3y7sXTqS0TZRMyekA4Ta3vKQlztNY3eGdvOSs0l+3IjbL7d
gmU2WMoIdXJPfYw5tyuukWfIbV/FHCRi+u7vexF6CwWrFC7AnyY44lt4sFO9kJCz
sexslJ0FKgbMOVmcEgYI1epEQb6ziCilPHqY7x189c63876gKqut6wNSPdHrXk98
wfgcmUsNJ2YwtreZT2bchGsgt+nsqFAlULv3g3aZDIEkLpcZgqoGAoZkOWfXVU6H
RViChXFV/VN6fTZXjAPqDHfwa3yMDdfKS1sifXVuowRbUG0DxuD8iJrpRlvu9SGJ
h/Fk0GIboLxUulf6mR84pzLTYSfPjmeLvtw1sBtDZ5Y7q+0Hx65k8nszmw4zicp7
ucqjMvXc+j/xmUTMP+jCLFD0epUW5yJUWsCujrFwTFqjQKvoENJbQ+m5vTMhLtb3
9/yQbXhq8BtaQ5l8VuME6aBoFjTjenXr9AqsJzLvrMhGJAP8YWP6Yn488N/wTsaY
HxGm6OBx+tnm4gJDsb8k5MtsxSLPdDTgIB6CJVbZ4AA27E+tqBhEsMIGk4p62yeA
X1dINB+abSWuX+JkIEs26pKJCSaoIdmkWtoho4tnSh98xa5iFsq+8MaYh+uQXmMG
PHM1aKs4C7rKE1YIxCSKvehv+x8AKU5Ea0FbpVLM0ORlv1PckP6WJhdzRx41YXeq
LWGynl3a/ltvEwzA6hTCVpkccPJdX7WZujQTMzy1rHyslKlXI+WeusH80z4tH0od
rtuc/0ZEvIVS54e0KUMIrKP2kkVlQq3LBAPMvjkyZdJZ1j4fZs5s7icO3nl/FtqA
Hq5gz7M7sve3Qv4gpXo2lHUxsU/QcDtYnB/XAfHwb+Uxcdocxj+ujEKpvZYk1P5U
TprAQ2pEakwMg4WKUIq/TJyFBcn2qf+K/bBpEjMK5nvoUH4UF/xHRu6+4nOMVNL4
XIhBhPkEge/QzVMVqf81Q2LA1Oar1fsn1VJEsC7IvciKSsZzEeIMNg9JESxR8M3h
X3tKiSKq2f/yNADzXrlck2B0zjcSGqiIvpW6/PuzuQK6x+nMYsyVa7kfjlSZw+dg
0mxntWAr4JaAAchu5xxNuBthmBROLH1BiLD2jVN3NMtv98VsjN3xGbkYTDZNnUny
f0f1WmWaH3sp8GVM2fNc9huILFjpLXtDsX1CEe3gOrEwL+7LDffSgKp8I+DkTj1q
oZ4oSI0lQJHTUFH4P2jAxz69ybQTegH3DnN9wywnyk+Iok2f9MQk4niPJnM0O8Yt
nuNPjDs62x0FKVHNogyQHK0LBcxtaCaVNG88MSxZqdbx+IhTiIaPLfX/Bi+7N3bf
ddWgz4OYlHzdFioSYxW1jgQgJdwuDsdSdojKoyUGZZu6v0ddxcjxWPKBlUAfQuDl
1qLat/d1rjahENv4hMoT1EwSV+EirqplYjo8W7CYEcsDVthfakBFqVP0JjW+CPP9
QhzjpBFpESdEv54X4mHeS0lSfhKTgofjuFbryYwWzV++pfZfKHsjurBKmcitJkP4
ezXDen9/q2F4XZHrDhN9F81wx8AOoowGi+eXIXj82RpihInZWuToIacEjp3cMhqP
m57Cn82/+n1oJqM+7ZrcfNg8QRAB2WYsUKtoPxry43aMILL+yr/bnlAGt+DODONy
z/pJOARhRY4Kp74I+0b0PTGJ0quJTsJ2bWPVgCtGQFwrrEZYkIo0udvaA/4da/qQ
K+as7S7NZ/X82vd2hp4Ibc7iGS+Sb2MPSKQENr2FX+Jtx4dhtlBmgf7l5zWuSQUv
NYTn0oU2bWqe4DjoJyFJQfgFWRYNKTWwqRXVebozxs8azQ08DsEajjMNwkia0vGK
V/mqRTyWfuwMkMhKPdG/crEXbu//4Do7RbVJnVqNyXhh1fz+0QjQ2mMIBzdVgy1X
h0+rhpZpmTQw+zj/04jj4icZwWDH4c5eCCu5GiB37T9HOOJnTDewUhLCjd8hLXeO
cGGa6H4biXUQ0ZsFz0RtJVubZiTDRmoiwIlbcIp0Er76w8hSCYjT9Aa8TrQrH6+8
284xeOw/vChGs9lBeRw2XIylab0/BjUbUbWp3WMKtxuV1dT2ChK+6t0Rg6P0tOyg
5BHdr55UmYTRz5dNR2GC3I2iwZ2f4vEfbhqLOoblqPcOKJ0jpKZ+Mtf4ysjPIU+e
D4+gOCkRXgdIxirHUYQCaQ5CI5Re0jUrnAZLnhoPPddYtcOF8yW5D9PdrO7153zq
ctcjc5LTeriqnm/NyA8Frlcn/VcYeUatAEc7wWqT1rHnB5HsJzrMTJdMhubTfXkH
zgDvitihtAiVjxhX/5SZmFOKAfeAPzirRcI2APKm0TZH1RnQwa+YiA5NXc6VnzoL
ydm/F9LdJJAT34j82nfIfkhGkIwX6PceshWnPTpqePovOBcTtILELmWA7VjqQXsB
pe9SfR4MLlDY3u7hCxR93l/tqI7P0BUJ2GlN42zmdtogLWmTlGb5MzgzDvM47nuI
EQMQPyj0kdbX94un8Lf8nLXwtdxB4Gtw8jgTLo2dlYvqjqvXAvXetfXH0T+Ecnbc
NZFHO74RjzbP9Z1payhV08loL9GXcS0J3CkkgF9XGrY3w9+7gxj0p0D8Zjy2pGYO
yUzQgT6N1zB3DkPNzajPyJxTM182ro35eHrUbEM3gd4lH+K4LtKuYQsn7naCBSqg
Fb74js5iBsdCgL2k91Aj4w/khZWlbC7Pjj26faDDb5+HVz99I6FpnBjgtnPYgQxa
cX9VYuSG4KD21F0os4R5Vxt0TXA26qy8m7/IrSiHHJtkYMr72nEG0O8OvTHn2JDx
7cECPLX9XC+JD5ePLvBJXWBGk2q9dmw0NqcDRz/ays6O69I3HWD/6ck13A0XbEYs
0rPRPa96gm5uA2eAGbaQTQba1mbVtkVjlQfy0l7HAiYcHdjegn1m3yXRNfyDiqW1
768CCvN9FUtv8u5MrH6oyVKaygAjsLh02YJ2AEiBgGoI4u7vMvt5Y7Y88TX+PeBe
ZhznYBCY2ZY9kZ2gRml5IZPzZ8vnuQ+I9CoFGKhSoDS+/PXJoOw6DhZ9wfxB0tpA
yFrnHlh8+zymiG8XejfGxe+buDBTqfx3bfEa/6DmQdgHGet04rf6Up2lsdl97A8o
RYHqAItTzSe2f5RmtclqNreoFmY9LqP8EcCo9wriUD6FCYX13MSYkCutfB+ympe1
e2E9NF0xcIVf4qrBjOq16kVRWWcLuMJqAEa0zfK/yWexcUz2hgAVjHB2sM1Ms0Dg
Vv1utPNLskR0DPPf3mpRrNZ11s7XO2IsyNgXRijHSjtJMX6knSGJucC4Ttgxp+VE
WLSZWRXk4EK8w4rsBMGDiwqagSlplXdgC5kDyjZYWviKLTg0SQXW9M6ztRFt7UYN
wP+yUH+Byw8G+OLS8TKNkLNB9iSpaEx1gfx876DzD8Kq9je3zM0Oabsl0OGsftQL
F/orkMH8OhxcIFXjOIEBlMShipnFNHKvmlZ8ywWPn62o9nd/xaZuML9OjqZLw9Vw
1FqULO3+9OPa8jcL0dntat0BUkLdvFe7opyVsxPxFOPucAQi2H/w2NbZxxYQ2JA3
MFWRCjOLu5D0Y8ayEyAed25wwhwk57ByeSeNM5oglFKZoz6Mn7UamIzP9OiiVwmM
VYPdi3bpVloEsHtRv68X9SWyXRm8Zf00Iasu7JFzG+UORLtmq/RTUpQCOWy3SsMW
VfQDF51uN9a8b56QFQZxldeQOxCAoUGbLVhPNbfPW1MwsfUhtudtaWbHaaPg0VsS
yi2VmoMvxijkSTyDSYyQutgG5h0fclJYMYESLd70WDRsjrk7yrqxJFO0Oj+sLbVQ
ox6twLkHHWCCEOr/wBfcoJyxwmJB5Z3M8k1iZ1qb0pRUWTXOd6FmxRNFq4i9dEae
E4o7Od1cbsbVcpC2d9LqaAkSH5KK3IZrPUliO2wExA790dkMOXbPhSpC9fdmpSM0
lPDpSZUcbLBOVGey5pBUyjyeflrABeKBPIMnu7cDJFALNNHkkfMkBUCiNzOeuXm1
GGQ4EVoEMwJS4TpMB8VrIfGa4MuDG36TputvxeVKAf/d8PzlLELNWmZ8S8IkQSuA
sbqYpVYIPvvsgah8vsa3IKrA3+qtXwlxuYz4YrOhOOtMT50mQ2Yh+wSIJQbOr9VH
QbWQ7hArkKj+UEIfsRhZpOdlJoSTEdbk2TVpFwRdGyyvidqys/X0eauUMd1Eoi6O
RpaY4jyLuZshOR05zNbH+98VbZRhxGpSYHq4PVIp62OL3fnaOt5kALgDdEh6spEN
LUTFYPj4TsyJ9Mcoz1ePvNIah7W1xao3iIgav3JtGvAnPjOkD2j4xc/JWy6HEcfx
qEajYOIdao6GjUL1GZC+d914DMkbc1w5DT/5v6kJh38upNUXsEHQfCWsrGyNLPjd
jQsrT8MhxHHT8DPz/WxVLv+DUbNP3vEQrhhYlFW/7TDLkYAGtJUe1OTfvL70HUsg
urExiY4G4UbpNBPnkjyspj/8CXL40ZfnNRLErpiiX83DC8g6IdRHHPhMViMKaz4c
7vNJcMrUflqhrVf3iY4LiTiKxA68HjxkT0eqevjV6EB9pKD2kJlt0w2/k+vk1ylY
FqRtWjDxvh1PTeJgwHgj+ka5hHEXKDn3v7LBmPPQoJPdHfEBypQdz7avDn5idEzX
C5Q6P/Qjr0XoPtIhTnA14gZqfpozbsih0RjjWia+Yk5pgZGoR+3hSjyCP0+vny7x
in7KQQOq7z2O2qrunZh5Xgwulub5fm2fuJkRVu0eLwejVt7XIqXD8VKf6UdoPTV5
vquhKhlyFR+LnrKjkOnYLuN0yYjZF86Pbnutawgh1yap5eII7ZcFP7oUw2qXB46T
mdZZAXCyX8Wls6UT3QV8eRG1nAwYfuPLWqtpCsNPEDc4jTWuY/qErgx0ieyBvrDy
CWQ/yjJZRhAnYToVrDtcy+NGyz7nWylMOU5uMzAlhkunzcWb1zvoFI4arHf6LRIL
Lx15R4sLntP+H+VobWqiDSx6LaDSpvZ+yivnjQx6wdf0mYJwfJxpcGEM9SC4bN+o
7Wwv/Ky8jIG9yOMG68cnDpRVtWtmiukMniGQXjnEy145qVaekOvG6AMBR+JZDMTR
SH2Eu6cT/TI24PNHp/SxrR0Uv4QU0nuXr3LVehIMHmJTBwCcccfQmPPBFNcYEhUE
3gLBOU8Wmna8GUzq93U2zXAtubjUzzV+RVZViD1IM1WY3YDs8iDO76LTYH+1kPv+
nK1L61BqoGMsPFZoH5EcNTnPw9MvpQebGRmOIUCKgssZYACyQloL3Mup21mR9Er5
/cCUOKLvftw51vuJlapMjAjbnh1kwjcF6x5nqLL42Cf9LsYi4BeZOgJq7i0j9gPN
D+oIaJH2C+hRGTdx4OfTnnax2gikUqkhtjX4urOEngUctXwADJkgAUyBXTqI8a4+
ZfVF2IAKy2TcUClaoECj5mbTbHUn6/NMPo1bobDrVzK79L8H7ZGC7i9LOEvGYQmT
Km+DzJvhiudUp1tqWEd7dAa9F+Mk8broqsBinoFTiTF3M5+XB2EDhkKJRYfbWtSg
0h0jtBgHv2kRl1GJNwX1HTdhkFZMbVJAGx94VgbalDJhMeLivcsgez9eRnqrhRrQ
7bNkWBD9Iu4qctbjxg0fszBBqp0yxGmz16KaDr76XfX9+v7wQu7GMQ3C4LJRtCUv
qJ91m+RpAD2jyMVdKSx64HirayfOSPb4NHAz6zmDT/fR9Ru1WoRbU6Lacw0jWgfA
xTRhSvqMcw8pJCpUmYQZQXeBqjDtsoeS59f/CXFbqQIoMt1VNMPDp7I+b5bHqisJ
9v1bmpulYiytn1h/2KEqb+ZXxK2z+Fm8EUPVDHVkRcuvXczFASpHl/RClX+4dACG
TJ/NYAuQXXrg0gALINkdxpQA0jaf97RZSAhTcibm6MBZe8c34zFWoqiboTAF0xTB
xd1kI+uNFZ+AHmJQx7Rwb6JpL2KvNFyzdJQ1t/Z+3m4TUAMT9wMSODGdYU5/TZiB
xoDUi/yca8vOMJeebgc04Aeg0i5hxNNPZ++GPmBm/HYaeXAA2hm9uCYafBK5ARnl
LPDSeW8ivl3sd1wpZLMjiHGRjaxHNVU69129qtcppQFvjI+pNC+dy7z31i4Vt01P
FrG+TTxpddHuwBNK8HLqyYtkV2B3Nbq42xwUw+EoPX7fKHXa8cJtCsKcZaLksjEf
cbiXvnBPzHWprTAWDiToMhhNOg6CtodpzcyObm2hvJK9fnkgFAL9ZkHz8gfBmRqX
hIJzf30s4ZrseiVgAMzjZnJvRtR+0DcR+kDljAi30EeGHvt3F0r/cickIoBxiLlA
5V1p+L4alvd+61hXGJLEtygvVBvQ+12fCrNwd1Xr1cf8V1/uvYUN28Kl/Fmy+Tyc
FwCfLDD00OLHZPb6PQbAGtyVrHS0jcYtV/9CsGMeL0mlRYxz5UnN+eMKd8pSuVCg
Af0GBDzkXInGrCQeIsTZGZYOA1ITD3jUythsJ0Gc/axJJy3R5Gqmr5wVvDa2DSDe
RrK28Q1u2+ytpyi65ny4HwWMaQG+gTT83BK/RRWuQ6ikgUYtQ2/CXp1FRBHOfk7B
x+X26KFNxsEP5+cNyGHkHJTnHhQ/+b0PUWok0kop72u2ajvhhqK7fu0JmIC6+zTy
hSJ/JJTNoXr5qp1Do7f2qYQG8q2utOXFPzp7zWxMnrxlpyj9s/ptMIZ2Y8aR7H34
PcaJq9B21KJd2r+/HXoPX87tzKIZ+Fm5TScByJ8bUfvyprVqLasTYNZr5CxKk9Jj
wFQ4pj+aoOPhq7pn4GiJs7Ch1s2SO9xCkxenhwbukotRCC+jHJzhZOik91wRCZ8p
ZSjFFUo+SgbTHABANznXX1gsV1DwpKQaAi23/DdkWU26687Kd7rmFubngw4feLA6
Sz8C7ySPEn4gsaofo3YwD3JeDFIaNjRenWOd00VHhkjZkpjoxLJ5jfMSFp/C3RWZ
XtVPlvn6d/o6n7OMD7wY/AIaAm4jAdqBu1hvs7GwAqRTon/DMUYTGfUev4VuY7Wq
pTW5/AvoxXBYM9v/gn1v8TcNQszIESD028kejqpoQDOyQ+wpJAWim96cBuYhm+bS
7iX0DbxFlJUnsNvHQO2KyczHv/nNLnzCHHyaO43/iNi1fkruhN3Vmwf7cKOzYtpa
nWb7aZaYnttoNMAEmqA9cAnSzhIlUSq2mjKsOEVpqzN/mYOcgJoXysmK87UxTYrk
bQQjDVhkbgAqH4lYGk+j2hwdIUly2/kc2uUsBnAotVf2pej8VJSB7yu5wp1yZHAC
gp36CwNcpg3LQRXDkJ9nbiLhNz4nA1M2lrUAqc1TP958f4Kii6QVB8z2KsqbbRx6
n6pii+Opc/GcbwiRJEcvUJuim5UsL4Jf524gT4JBtFsxwnxb90fGcJdnLOit7Mv8
esYp8K3stUASMcL6nT7ibzYyoGyHLQVnUhrumSKvUeiooQAyX7zA0rLFvaao2ALD
iCUqGSxhX6X6Y7id4OTroZBrtEGH4EftrPqGLBIJZZOVQ5wLN2BrLv+4hlSAIs9u
w3k2FomMVqGZzW6fQAH5NXJ8zqtPrT7Xx8f6ohxlNH0iiMuF9mHBJhJ/MauOJHow
+TQBhV2Kc/EhAsD25H9pUEzdGwsrHB9gXQ8JA6p20itoAVHIBKn8+bvS1AeY9Nvg
CB7PwoLbaMdODjG0qxxz85rwBaGU+Zjnh81KZAv+Tyn+FXJwpvrcLAlfZTFXOlFJ
QC4DkfA4suhVt9k/PVVLVzpCcIVfsrJIB8oWgocbkKjnPkfuhOWNU4RI7F6OrA1o
rXcfruf5rwgbREzNwuiNbs0TgwSn+omdnA10Y2JLmWuwDcSvDE8jf7JYkqJaMNOl
4nBbwAH+7JlrayJ1lr0g4OimkCwE24al9B0RUuddj5pYgVOJj/lbeC8Up3vLu+Xi
djG0K4zTBLXyDOEEHwj+diRcNICnPeOtyA8Wf/Aa5BxvJBqO3dXxsAQxVcPoKs3w
ZodUwp3eEiY+iFdkzVG3HmwxxZQ4DkOnf4zM8efKf5s/XozaqvNHjHo+4fx2S543
9jtY3s03eTzOO0OsEDH6aWduWspQjl0660AVKNnBO7FOo4gbVprpvLOQnC7UXsQP
Q9NnMu47GOFIMcj8Tt1OKzaf1mpVNff6KBQvCDvwBpkd3d90kxmwiB4DDJsvcU2/
IsTweE71NVMCwNGNTgBZBe8MFXPKadZoT9P5i9Rg90lCfIyBjd38Mq3Ud98G1hUE
ZZ2XTkiAOjbUSd+sUwCmJ98MFDXkBG+UJ/QE0K5KBwLQJHsqYgvN6Mc2eoSVvJzs
O/iUasXjjZrsq3wlmEKxre8xPCcXwN5CN2sIBy0zWqlx//CdmYrDvXVsrzzIYrjf
I9WDIdaZMu6RuJRSYtSUy2ryCRHpWZQ5s5RxPFFFZKsG02qqWWX0d6y8n7Z9Zflq
GjHRVw1cERT+7dgE5sBQa/fTHMIj4GGNcgAs35x+FTc91o68BkeZAt6H2uqavb2R
bZWkWp/9+fUI6dsA1tAqY06xojdtjaCKn6WHrgKuuBKEzn2lL+Ihc+o0HA2WTi6C
bLmhsuhQDpA6HHa1ymyj13GGKn/MLkBZyzgQPxnUxWa2CSO8VpdQG64Q+TGtTZET
cWE1++fA/ao2EtYSd0qfWCOVggsogkj87PmRLdeAx5vDvPzlRU2W9N9gtLIv4Bq7
SqCcofx/yvNnZeGAYYLMaKkajHbyEfBJpFOxU1c6Pa1AUuwovSFj8wH3EyNtsac2
EbwxqanruUWoZ0S5d/0hOby9P/zAznZ9IrO4TYniOlX2QPSyszR0G/1+Jw3bEUVE
ps7Hu/3YzkNuXryINwVWkYODiSK3WuuOzQqMtinB+a9Ru04BLyXaZ98QJoPfLXAL
WTj4M9ZHaNpSQSZON018MGtGjk8jxaJzrqzMhjFlwgwOgPkSOvIzXxauGI+wizCb
/h7l//hlo1gbBtrNuSkzS59pJVZXq4aKRQFcKEUsrpVc/LP+KqqUUncw/+jevaFb
KBtb4+JzeAQ9E3Pi03vvam20WV1bQL3rA3ns2MEkuLr424BAcsiVO0nRaXxS4BWe
+M+/9G25ujmz2cbZck0DqxLxtKB48F6K98shxJs95n3Z1JzSoiEhSIJafkcX8XdB
vsLf0YoJHLjpKqxCDKN/LQC1JzZzicCgOMWSRzz3ntE2AZTFEtpKP5Z6aSwHPnk+
jH4r8LCj1D4QGFHX3kY3snTIj3klTyzWv2/B0oQ4u2adeGEYOv5v2G3/hxgBvDLp
TLJXxwMH02KZ9LPu77RBf9VsSzWwmwHH4wDL8lDv4Mr4SUG2BiJCdHTkrb7E4/EK
PCcC2yENWlbRs/HXbWvTYwvwQ9je/Xy/ZIVPmPw+XlGpIwfS3q4YJNymOC9mhPFb
AnSi1QiLOFnd3zVfvHGHn2srFK4L2yAGtGSXZVv5TmzkzFAzvzdt7DwI4vT5qMgg
vkBT7xjyOIf+Hs2+okWXLa7nTzyqs8x0exJjUmHRtG5h0/6iSE38Sa258uI7GmYi
onNIdvw2b3TXMfKAXh2RA8a2m8WuriyIx5TvqzmWRQJ1YjgpPxLe2K050cqDFF+2
AUCaL+fBlj+GCfaT1AtSUhTptie3EeP5N4SMzvUNBdbyNgireSCFPdxWAcfOdsCW
gl6ZmbiFvBbmE3ioX9BT7cPLd9SoYmRPz35QQS49wE5jp09Cz/67PVO7MgD9EfVR
IYIgliP0t9G0NQaQKpdXyjs1cyo6ScesvVRdxDugOgQBAKVte+Tiow8Mmg0QY9nZ
sVcLm4jOJhZXSD10Jk+oqjmcqd9uZOWwEQXnVV1j82QE4Xx+hyKFUQ7pb5n0ohFo
Q4Sq5cK381OVGtTneLcf4b5wMEXtWQVzf+4ADI1keNls93G9Skq0nWtXcLX1w3y2
P5UIZ7IN2NjxlPLuaPujXEW+G0YosEELCwYpGlLQXAEbp8+TXzAEVmaMpj0G2b5l
oH3aTm9fm88VngRL3UoM+WiMomcOuVA7a3um5eL6kKRx549tNwEBw4JGnpIooSXI
4BAtQOSq4Gq/AYzbZe2w7AtkcDhVYAlJj6vFKstA2bonQ/MqzlB8gCRbTs44B9p4
Z9UgU4ksrT9+3Jo/Fo/lj6WlnrhIfCUSBk5GFlXXK8fuJs6kLkn49p9UI53AoXxt
6taomyFACENDL47QHmUnjk4c+ce+8D7CzCtgqAX0dw1BkC8l+Tbxg8zjwq35rMm7
wZqOB7JAfhRK9g3fdU6Vz+ol8c7R/AWnzlGcXagw4ZKTWad/nPcbqg5wBYRtOQ3r
cYC7PJP6LSSJEeIcLSPbfq2sRpLxkxM2+Jut4I/nixhxQzVo9U5nAyBqLYItqRo9
8jsbUmYl0Hp0thCCXBLXxQI4z2T7YSmC3Xp9uHB0jk6BgKh1nRLS0PIpfI/0QndX
UhcQaTpbvxXhu2wHUnZFBi6wxEM6yEIK7NvC8PBf7Nyk2kUkyf8mdd2X2qz/mBFA
7nB7bk63z1K8JhNrHttrrzEzTQJ71//CcBsbpJS8GZpBfPcvHLiksdX6WU651SEo
lrIu7vvcZmFyVwCD0+5B1m+eRh2e3lOr8HtsKpwJ6aSCiQSICTPCA+lWKs+X/6My
4OpZaZBwdpzg6mOHHAuMzIBI0qiSbASyHUVPx3/9ZInpXpEjzi88nEFIdp4IFtWS
HyP4NeqYQ3ceXCkwLLDzZ64CxFiP/NJ6JtWDKCwLeLowuylPIUDQkaECRy5bmUSJ
hYnuW19F0w4ci1XFrrztDij8oXpmgx2m6sVudZ+y4O6tOrOGeFDE7nyf/rObhy4c
5CsUEuFVLgeC+3K0Lt8DNex5NA/gc1X0YgLSK6e20EAZUQzfrEfE3GeIGBu3/wzu
TauPMM8Tm2ItMFCuZXVbOzlWEg6rD129OVyIchsod6x9GeCH/yADI30Fk9gpLeVk
cfDNAvfan8K/N85972wFDBBmxZpWGkeEHSEvF/eaIqSxaYdXB85O+xqxnulxMcHz
HinoDzFjCGyo6Yhn1vADswZqeGGMTVkw3PQQ3T9DY81W3jjSFEbwlwL5jDLgclIU
skrJKBh56uU2xzb8iBxrZWs+u87FsiM5JwmuhpzpiA0+pl1BdO4WIDQIfHMMAYpe
LKCLkmLqrwlqv5Wx4eHk2sNHQaN+rAiJz5OoSlNh6NZKtic7fSnWgIy1dR39impk
4FCjWbA7PniBHKAZKGF/Lnv1ojRJfL7Nj1ohSUQZEhmtAsDD+bG2vpzs5lUDdNbW
LxvlfkD4mXC3ht9cbP1LILSWECHi5HAJGSh9ZratF1Q/0LE4/J8wjancFQ118iDk
LdARgEU/D2idpOLkV72Y7Qoyby8Arqwk3HrZ/6kG+8eMGiB7YQuVdFLedezYTV2h
l23ezt413JtlPdEzE2o1f23VuE4lignwn7ASW9pUfrHWVRU2Ytc9PNjxm4fDvoCT
/tGiH9gd2uIQbl9j1t0srfVPg0cl9wphm+QbiTSNqoLYHX0gckbWFt+C6b1h3hUq
lHX73zYyPgcPK+n5GY2PyTepHvmoinRFnaxwp8TLBxyiyHJ4q/yMIZeoC0SXSf3a
KkEYMB82GDi3wHIuQPNpeb8ZcbzAIpQQhb7AD+PaTXR2Wrf3HB394ZvFiYna+lvX
9CSPOGRpeSFSqGvD1n5pZDMLtnlhyBiau/+PL3a5HAiNDx7ARSFwELG+fMeBnzA6
adv/rKOkN6QY6T5Na3ZlahhPgXX09syv81mGW+mR1xv7AinnU3bqxy6YwWkhnFu+
tnOREH3jrUGOiLzG/4PLepTHMH6JJHVD2lubUvQTRYk7NRuZ+ZBTdkDAY0B5Kwm2
bskPF5Kx2DJl/VmSVL4uh77mGLbo4Va5rOHgCNZIcNijq+sEtefA7QvZ8hzuthRi
4B8IwwVD9RIbESPugvdLMZBxxF/YhbnK2XE04Jrih2QUJytgiV2uq8r1Bh8l0RUt
e3aF0rnJ2MIS0v1w35a2NPEXEqOBUoCcjWGvElD66gm1z6asxkig+fuWkX2FehGV
06I8/KAtMGZbksoA8CNfPmgWCWEXZigY1QAJsiCmt+rol8AxA3hCaLaqClJiAala
ap8LQnm2DCeziCbWy6CbsDlTEgIv/c+XzQWrcR+bRsVgc8BhTfbMPeZ7sYAdjoy0
pA4xZh/t5uHSAbgwqLtb99AAvOo/U24Hl0NM4/E4A6wiv6diHHQgDSVo76g2Muo8
Y0beZuiJQB5qDMn0SiJHTfTFtJ0B58QttrCUOrrH+qj6l8t8Rf+5Cf8B0Sho95zb
ZibbqIbzbZKMZRAvO8oIvrGqepjvJCfFw0tOgktg9vVDgsvZdP7HbbTiIKMg4MCW
+7xnD3uXtG1cvc5aAFEOdMyrGktOVZ2UHBPH0DBe7roFTwP9L1aGc01VcayrUCZx
qDs4FlXWpHn3q15D2LPyU+r2vtNL1FyNzV4+E6Aje31fmK2BfqtmMjGH5A0UInRg
uv9aE8CepdmVhjDOfHnK/f3eVu5xOhHK7Vjh2aIs5DH2SoPlo+7Yns1HivWjavXZ
QPWdFt7wEHiwHOkVQ+l0lmj2BkDqW9WBD2qtiO1iRvn/usYEPBAnWr/REaQTYVQH
soYUxLK+mHcvSKSA9cGqrjQtzsk9+2U2+QTSIBq02TGcqBsbbW4UoBVtC9pvIXSq
BM9Ck5l8S5A8j0OVJZELT3jkTHkH4S2pR4LlQZXTj5OdCXqVhCwDKlez4q6zscvD
jtwXi5YhE7dgkLBMBWb1ubFtzk86iQzo58eFIed53J7D/sXgZZi6cf8YYA/tQtgZ
nSVtJHKimtrH8J015JzhcwJc2viQaT7GlmRoIpefqBaxd0ssbeIHciajUqI07Dbl
lGPIqvicZ7Ao2aKtm8IfzTW4XVlTGQOg7RUMdgvjBSHdBpdYmQRA3Lp98M6KEf45
O3UjK8YnuxZvW09aVS3/PBvTP2jMzkwxqB7UqkGATZXlDjUU2tYrWHRhnKnXxJcX
XLQ74yMCLzC5O7ZztnCIQUHSbO7hW4NE2OrA573DMhiKLbm2Py0Pt+KV79Ag1GXl
DGHWR8nmdyKd4qDb46x/EGdmAOqv42XA/ySr/SeEpjirTryuvXDUXFTWfjPEOdWE
NKjtXdpJn9fL3aMwUva/2iYSgDp9xaDdEXMG4DMe+I5z7dos3HGbEQ+HpUfku9iQ
kGbHiqDiotaoT9h5oJZeptCblSQk818AwBYnrvYuSliBjgr2h4UzaSCxOXgqjpIj
oSgK7MjCLmt3allFfjIg3wjrifysugyQrnRw5zuTLwBHQtUcbnQhmJczTHBhNeG9
0xVCp6jWQsyRsB6w14XrR491UDE8apnEHPqDmdrML3dLmnfIz5FYahAKoJYTwOi+
g8eJveMI5NWUnHdbWx+QZ5DF3vHXk21oqhEIFhn5N1z6Tq7qswjCYEqBydjr/sC3
UvhAQOVUcZs2rh6WowXMYvc6sKQbdjbOPicNbDnr2O/4ZoI/8HzPBtYaydfwhPKx
OI9rIum8/5PLv3RzNi6kFjvhr0XgZqiEYr9Oo16ioz4rBM92Xk9ZqeRXeSVwaMmj
DxGaoWXrWLHaMAqmjit/XV4vA38PoyYIFTQI4oYv21fdduzLLVC3F/+w84+pZunW
HEs/QMDjAD1JMbSLDGtdkzPoE8TpJRpylZ1kD3OGFwwTD4gni8pz1lXT8FVP+ZL/
hHGKnDplGQ1/ImO1uu/LqjPJWtTdss/sonyBLWFLuuVPkoQ3Lt3D1Bjxt2Nd6mtj
qwmZCkblllR7W/1LAE4uy0Rg400cckIwSpR8DULNvoWPrKbUEEUqAmRQ4s7hUTSi
f3TchLYlzvuHHj+OqINEZbwHHy4+Ijs9prmfzeT0ajzzwpicgljKu11/2az3vCQV
bh9uHUsktdN9ojm4aJz6V0+kT8uiZIfTGrtWOGvTgMqjcf1pWdt+aHjkrBg6wvQZ
wQ0kaatcd3iVgEUnwTbhKXmkGr1jfoSmgPZ3hCSYA5H+9HRb0vV4M2e+Rd/atsk7
9BvrdeWphHcEIss/ub9/EUOAEAAnvWfierbXJYjVauJkxnT6h6fs4ACcnov0hCfl
UvEhq5GOQskwNZyWnj8qWogKDmAzbpK+0OpRI7RSOJ/i4AVTMAJlnRcFGFILs1SL
k6O9b5MyCajAzbUYvwPLyTtheyx0VwWggjQBMo+0Ozlev2dVJgQ1WSEWSV7SwwIe
bWPWpb9afZ4ASuMbVLwIL149rwDyvuxh9HviRrKBieTqRMUrgRlv7iCXMkxPhcMy
/JyDPCwCIvE+ugfMzYI2pSaPzu0uW+47XJVh4uN4pJZxnJbIGG2XLyJENmchHEUb
kmVleic40r6KonH18UsZCAPfYp/TcQTMoCdyiN2MFokwCbT9WLpyju/lRDY3EHFM
xd4NuQlqDxz2i//av37egfNVAb6sH8nviqm08fL1bxu+s7/z03J9OQQGCEkZoxLe
X8x6DJTLFT/IqByNZEy30km+3BTZfmWqdONdX7IvFWI9HhnJ0vuQVcymMnj0ImZe
KRVey2L5LnosQ/4AO2BkTKC3nJgYWpLJ2c0CZD4ukLkfGpOpZPlJzqotZ9hxI28h
VLL6El1+Ug+JaBVXEgk4s0n99rXyVTzJ4LG0IJr6JAnw7EUUCe31nTF9U7q5jlNr
+mcS/zVNssqPBodCCYyx68Ig7wiLjOfuD/fwdNQRnf8c7KRnf9T2w0tRMZwEg/IY
5wZVX1UsF1fGqv1mEyV6HL7FAepz1JxRrZLFI1qWhwd56hKY2D3Egnk9bAGW8oao
lO+F/ot4S6eYhXIrcbh7bch7/TZR10s6HAsMVfCEKE7h1avTSw2GZmhE1AKybfLJ
BkOtB3VPuC6Wj1RfPesIMq4N1yDLIoLMx1Od5i/q29kp156JSBgKQlNbhxXjUasM
wNErKki4T1N/eNQ9J+3u5HkIMOZ4914JOul7a/AfOAEjPbRYXrhhbSxdELbRWeyp
byJZ++Z+qb2t0cLvkZDxOhQ2/qlfCWxxXjA3L4seGvId2tZDpk9GXlA0LaSB8VTC
Nvl4DLcoC8VM+QE29evNAL0zK1vzjJZKIMzGuw8saNI/ZJauVM0hwsGvi1XANpO2
/xYUSXTRT0ZDhHVr9WORe6A9Kz8EwOcdShvZmfrHJV58IwiDdbkk3BwyvlI56i5K
P8W/EdfIDxNDruuFqIT++weWEquhKx+G+5YZD5Ya6PvUFqWLH/u+1Z+If62jibZJ
okGSNH6Xad0nK7SGGyoe0zdB0pcSNUIUFbLLoVeltzle6dBIWPDaaX45t3hqOH3D
XwAjJTY7Qa1be/+zuKTS+9Hl8j06IC4zQwJyDYc91qyd+dBwshaUHpICdId8YkVe
ALqBwXnLc1EfyVU/zUfbGjiq1f6o62RKIIl7HazTo0t2odqrh43okpzyPsO3+rA2
SSnkG297lEF+CFVMlS20TI8vNhM6Rz5GZCGjD04dZAK9FSk4NuC45M9kZRdtPye8
sNA0MXq9Q+ebvbdfQLW1Zk16yfWy9A5QKwmsUjuFeKuZyOqrvPr6SGJQFzQHPcUO
BJpiCWv1g8ef+edJUsi4zBMyBoj9SB388ynhO2k7CJ5RFjWESb723+WoD8GqVnpR
jzQSHoBlesJVhsymn7OdL5gPvjHvq4A/hiN3wtSuV/WWrJH5JINrthjxgNEy0AFI
FTySUfnK7uvknzKfrGCf2LofRyZJTfakDAZdmvl81Kb3i3BtZne0wASzP1QhrNis
xPXWq0SULaOpv13IldQYczXeHJlJ0aauiS07S43xEOQuktgocrmeyrbrqq+iDYSE
fVaFABSBIPqzz2Csc8j+b6yidjTgGRHMKUXiV6FE3hG4HzQeHYWndv2T/JXAwCtb
b4oUzfGM0XkJyv/Pb13b5Xk6EtBBF9NZXyRL1Yu64l7ORC7qYDhg6aIeUsS9eH6u
lEfY+q5N1agBhrqhn9yLx3GEA5DT0B7tAG1sBpXzT8uKT8SqQqG+6Zyy1qs5p+oZ
zXQuZob32vJhfL0HghgFwK07itQ4HCR4+Xrg+CoRwsUCT6SS3JnrpVtomTPhPiOD
am2iu5UCK5SOFj19WOgfsvkxVmN5bXokTVlwPqnHN65LlhCxFJO21ZDe1f2RhQyS
6+X/ZEWMxMe6dzilap0wFl+C7fXAXScvrQbPqvsxplXlefZv+Sm1uQ5QQ16ct8EZ
X2dCBRYYAQeuXhv1pQFTRw+tSOfSEKqlvyQy0T8Pa0jIvN+8oMJqjIIOeHPhcq94
O6qPjx7jKJZJ5KMG3c4V+uya+m6D8fxuHkk2TElr+2ZVeMzN1uVQXRIgb7XP9FKm
SGYt9PqMcfQYbZJ4AOD8kA7NEVUH8g6eugy9OT9FsRQVqiBRExH4Tqkvo9GYC61s
04Wd1PLyyJp1Sl6Rn+b7gIzQqWsnjFwAQdNNITs1Z0FtFhznvmL1Mct48kCRUg7P
hz0Qd/RUM6oxaKlQQlydoMxKhfFFI67WCDoJB03dxw6OgkkVfHP2/d1NTVlbrWJ6
WnqMJ1Jf/Y5XF9d8GHaKt+2B+2ZMaT9KG4M4jPNTKlAdrMNMO8CCCbSbMjZ8Z3F9
CAyQROJPmFRmHxt+hLRR0AKHjaOEEQapbIWnhWNo+T9Q6CgIK7QcbOkQwevmg15u
rEcF+4xwXAG1oV8KkAYDj43qyRvkpeJxs+BoBIB7gi8h6HNBqaWd5qwOMjMDYJhD
pRokYezIiobOqaPGZnnwgqlaxpt+7oIiMR+DQiAA5czyY+M1VZ4/VVgZOtEdd4Z6
mN4DwLrvuYz2VI87o6JU9PP7KpWDLKJFP5IckCm6zB2iVr8tL0W/KzF0hh5clpUg
+9wa1FeNsW7mQyIbnE8DQbmOc5Y9uP82sWcwudCduhZSpuDRq1XuPqVyRXKkSBBU
/OnZO8QRzWNj/gVqm3FhmMDjkZKlL1ZQcoypJ9NDhMWYp0L7GHyw0jCKUBQ7ppfx
trYafcjud8Vc+ccXZlMIADxJHg6FzkW8LdW5wFHlGIsfLEJSBAFSqjxcoHlfLne8
enImPdW2TNLyr0bm0RsYVQxnVpzyhJ3UDxir+B3uIkCWw9xhSM5QsQtkVPjB33df
vdno3lnNPFA35bHbiddCYerro7JGbTmvnCSZv9TF3gSMak6h3rPEpNuFzu+Gr1Iv
dK87vOqz2vhidY35mlrt6rNDNMQ2OhEljHDAG9T92xcPF/Eiyn4kziRk35GJgIhp
t+hlJC/XhofDSWUFMlMeHGHKWpj+xLexZEHPOWtCPMLYL64Bu6tyiYajJ2Gj2hkW
NSZTPuEUYJG2kxY7q0JnoAnq4yLeX+lYXjIU6GKS10585it9lX3dtTPcggrvoAsV
nOYdvC391ZX5fE7WoHO3iJGTFVw3umAT79SNMbt3TNWrxrW1luk8/1xXeXzC3otb
bHfeWeMWTjoFoTSdz6CYwHrrvvoxXCpvY1ERXgjs+gw55GAkwFK1OIG4vfsvQoOj
kmPgJQZHQp6FisYCr99bGQXx/d+Ad/9NnFqoLSPJAEsw4US3aUdCmfUdWMyGeOu7
FGC0Y1i9gW96FDczKAEGJayojxtdaDznn7Tr4bqcvEFLlkBSN5rkxlW0OBIWVEn+
HhgNNy3EXw4mCcF+z7995r/CqLsk8hl4sl3ruMGWa1cWSwFah+LfsG61AEI/MH0T
3hRw+cfHz63xiRBmv9CsrDPZxOtsRf1fvbvZzD788vK+IS6a6WoW2PSYkzkF05sJ
9DoB3Py9qcgjv12MrW4g3n9fQSO74oV7auUG4eIc8XgFqyKgAr42mBDbxBSgUMXG
9fsKWcrNCt8nS0ZDPP+56JzFakXgIcorZXV3gZJcLUrzpPQ0suRyIMi2nQYbKuOH
2t6IwntQH3BFA5A3W3bt/l7X0Ua7M7BqaM0ljmDGDCbeTgoBlhgPc1mTKFVhwI2K
jUgcbvPbFjg6IUSq9zUP2hCAshApjBMymOuF+5dn8027tv9aK+c3GngLBmbN09Mu
xzv4tlQojJiN9MtfxFLFGTIVUnajadnQ0vB0VbcqGfIaxH9KN0jpBCf2BjAag1ph
YRn7MaSYtAbkMV7pgrUTglhaTCVX6ClfwlX51jM1q5cS718RID9jSoUfZgEsOLk+
ABcmFNZ3WQIdpj1LiKGF7k8G69k/H38c+byo5GX8dZlSqHwG0hBZP/33l/jy2hDo
KE2AOPMq7lTbjjxiBhRKeh1HqaAfkeIKB2f9LU1mj6j7WbY4ZzmM4go8K8Jrjrk/
nYyCDRK2ajNgNtwJOyG7CK1sLDhGLvos0oJRpi7ezJWYobjR7Td3KvA963mzo50W
lhKyKlLDBMRq2gILB4Cu2k9ZQQdZIk3QxWzO6FVdzIppHYYhDzFmU8pmBa18PrHu
v/FUgWS+0QmthMHEAzoQHCFrg01REcU7xMDnxXoG6ysrE09w/31FzyV1fnPxW6as
0J77ZxKzVS/gGxz1n0oB2nO8G1ilVvY9DppdYdDSMg7a7fExsfp9Nhp96YEHighY
I68bfL89/68CO2O3+yGe0iV/RpjubEerfgLEeAJzlksD5DNZvA4JmEvERUlVSMzS
X1UuuAYlgKdFEr3K5n6sJuqKXmjkD3C9UJ82TSDNZzwmHlvGu2/EpOiSxuAGIADX
qnBxQ57wf7Zp3+oCzUdDxjGbOQqZK40tz6lYHdTSGR/LTq7OKHz0OBm1DSL+tpOC
xtAzQmdRH9h6Or2y15pA4kHz2WBstPev6HomrJ2yhEGY76lBq0wJC3mzpoJNslmr
F/0j8Mz1JqKYUP85/04G61gSpBpSRDYVaTff780RD0lAckUSdZgkpWaO7m1lRB5s
jARNGZd9K9ifFpMHXbyv0cuhP7vvVoksklN1w48nw+1pXPYDUh0/4HKZZ5UmwqJo
U5Za4YW4XGoXJd3NXyeeiiP3CV53Yrkxu7zjP5EHuqt43nRqNC0H66fZAPQKnyKS
VutfZS5VjQ0wC58QxrvBW4VhPrrMd+JXQoKPqW7+AAXXM59kd8j6IG05ITCZMTUl
npc/dMw3mVI2ked0i+vGIRw+EFqTgSvqQz1R1swYDZoSGwkQchSPCIVtMXZyDTJW
MoF2lH9nJsGlmyIGnSXZTq+qW8dlxM+4phIBme9U3plOchv5f5iEvExEreVgvhJZ
ImcV5SGEH2fjf4itdK75VKlLjOsZbOw8PhDr52YTtRsE6hqcWOjNYSwXW9NhT1j0
Rd035a0JTiO838vH32zuAH18oJDeuloxBXKBVm0Sp9l+BKpmRsEYVioqJH6TscNI
5BSxbuRvk7ri4ZVesnlKdnTDNZ3P1y+eIo/bernMAVb5RmPdHcKB9ZRKsHQIFfU1
ZWK2YZlbDk0BVAOp30fgFWMyKJc9Qvm+C3L89NRdS5v6be/IoVPRgB+WyYJFkzPx
Wz3+0HjMTxB00/yOz593YwTxsY+IwkDn+QaviEA6Osf9mz8yQMnkEiv+JN5vg6Mn
S+nmemwG4hLOlkX5FfMhbMBId0ejBW8iBMGOm/0YylkZadv+ZwmSCeX5KHdp0s3b
Vmh3qonCmnRW+T9vWVOTibyD3uTcCEj0TrataTvw30iKa5eLjPjVu+4A0Xlih6Ez
HAKQf+wgq0rACFq6YeQ8haZ6hMvf5CDuvTKaBeeEOncAkvsH6Q6YKpPhBy0a0nGF
FtgS0MjikQVRRpLRElXBvj63UFBBjLIIpK4EIJBE8vA6QeLVGtACknDPDkztcTjB
rXWmXvZTr2FQ/WJckrHBb0+I5kCwJ+pEu9cVu4LHR4z0ZOthPFwrBgiGnfQ7EMtI
ENqlibKS6lWvuotr1ynud0b6QZEaH7LkY1p0YHTtqyIOu7Bxxt98WI4bAluyyPkK
4jQnJa/Au2p90snsmi/PCOMF/MP4uJjGz+N6ZzDIrEmvB7KnLvWpxtcFXEtidrsc
T6ECc7xBYARRhv8TyEHFTyqOZ4S5zN4p1chkiY3vfqZu53MsPEg3UmYg/GN0mq0p
h/Sbcm2PF/+OeeBbQc7cNxjM/+SFMaVROBSTkRbsj5EkleUkne1BSUj0pkFdkVE2
JeTdo5lvSIFadSxiXOlKlm8n7Yrwh0UP5YJC8GyteIQsv5phd937wNMEOaH9B223
/Z/yv1Xnqx6Etb9FAnOiGIgaotyQzW4CG9kbS/9cJ7vTTeCla8amTml5ANrDIj15
GqrJJ3cdBGMsEbpeVLqAQUnbHm28FT8h0g8JhApb47gUd6/Fu6HZdDo9D+020pHf
mdB+p8zO87cqQOizNqziZocaErd0MqIe8t10ZOr6lrMtMvivvKHtsrTZZkl7R40j
WsTzykyDoJgiaHTW62+fVIuPEdzcwH2ezVFj93rQ27lc8ToY4vncvUl7vvhyRdco
sl4cpC8VELPXDdd0QL7XOZpCEb+MLQAchXX9NhNFUVEEAIXJCO+mM1b7KlsGJnqL
Xu9Qx+Z/ZMXzlYiMokKPtjg+ixRwg4nsZBMJtDUjZ4JFj77Bb7/pgo7XppnnS+UL
bjtyG8ZP/q3dCkyyQ3klAPblfirtksKMB3HU6UOHl1cWxJTuck20YmQYD7LGJ54F
XgtlimhbHwhD2PzNKbpQgZtgjDFyG/8p9lXq0zHucC+ON0fB7Lu5znGLpEeBjKwQ
027XKJFuPzjtse5F6N4/+FrmMTUVsoRgEUkVF4HE019AB1g4NO+votdwKieZJYA6
1XOM3q7Lw7XpoYmEY1jS24aefQauCqdDS0vhS4Lq2L9wVLMAI3NGV+UbgV07/5x5
ndFDlxLwo+dpWuhbDdbf/KDnzL7qQkWLkJv1M156Zzz9LEDleDWX6bWpQnCgs+mz
9S8MLnUiotQwG5hXHXJkg8512QYxC3OzC10PRTAzQV5fakabtwMla5hJGMTZKGtg
lNxrHT+gdqQS7kTlKjue35Fw8zw6iF5SWgSlwGu4De1PgZ5eKZjt7kXIxlnoa0jJ
B0m6lu+HQX74g2C1QOusgkVKPIaOR6Wf/GwFF+QWvH3JrksBTxLU21nEUaGGqhQJ
E8xHAmRPlamu2yew2q1WFUEKVDMCpS4rj9SxDNslTR5X5OOFuAcm32SD3mxQR58H
OLS+RUcfTTCZZT9yIRA/HnuvhfN01LFP71N/KJ0borhvaGBmusx0rjKijUObnW4o
0UiNyoPw8enOdT4MO6mchdJeVXsnAS40FbT99Tslx/GfilTY/EAaXUkxQ+jDcAko
kiqJk0L+Uxiv5sroPBLVjY0KtSce5yMu9BFk91e0vop4d7VLfnHxo6hgpT+l/n+9
tiUjhOQI5KYsRp6ZmIjzOOCiQsutFpDYXQgqij4jTgbr0+pzDoYfjg9gBxWF7mCz
TlW5eRfLfOXIaYyj00QFtPoVyhK2cTsFFlPuIV5XALU2V5J63En+d91tJETI7ct5
i1giU6/2AUhuJwsVcefs4wo50PY0JOFjCoG9lT1RiWWq8H2aFRyI9zGawTKHh6tF
v9xxFakZDwcwon9XPKnOls8HqjxmTLDynrPtZsYQron6kTbf/LfVUET3sm+tiMGy
W2PN/iuR+9byhT50x8HANHDPlCVtkXd/E2sc09YOCbQUUchBkpiQM3YRx6r8Y72D
7Zwq0W7IdFi4oY2hmn12NmUw1vf5YJjjjmlSvcl6cQRF/nyG7rEPTnyOLdxn0IBQ
b/jyADPolP8QMDjBlSi/NvvQmoJdX5zuKddods3itcNdyks1w0V48WD+3NhP9Z94
TQslfGfaUD7Q+SfWNnv5PREm5MfEVI2mL+EEFyuTgCaaHpQm1i4aNfinjReCEU3T
psdbsMBPAhibcMOX3T3J1yhY7Oi0bIRO9K6nNmHqoaN8JRel7TLZMzgqhg4FymQA
QLJ4/dGFYdRiM+thqFuCVTwYeLVKEYEXskrYLBoGLoHXUN3YXe7YVmFoLdgK2i+U
9U/Ta4z9jATE3fm6rRVLePMebPJW5guGKLgr83PlwtCgbXfkt4DOciiL8pNTtjT9
wN8b1p3ZdQmgzyNyOCAf1cKeb/7wYsewgO58Djomp2K586lpr9pqPnFAvcSad1HW
IZWdbiNxFQLLtC9bB+qGMDxHWZSB+g/ZkgHjA7qeA09+JL6cyHKxG/4Vm+8iPTcC
ZSEiugQddpWdDGkd0NtyRuA6oVrgEAnlzXZq4kG4l6oMpx4h8tRPGA2eGfpqV8MT
gt0gGttHVTj/a7r37Y9vqHxx34hAx/L1K7N7AAy4oZ0aYy0Qhp7Wkl99V4nqbNj7
s9QIfn7U1ZZ2gDC2hr2To9oh2MS90r68sOFWTjYCl8Jim8qS+CijLVWDoAz+6UjG
aQ62k7tkJet6xSeP/PFCJhXwGQgrkkUb4XwvwAlCbVayAAoRvvsGzNK0BIYRqwT0
iQuOc2tZJRmZ0xrFxkRctFCwG/zXS3F5h50iFI9Y/Zi3g9vBVq8lSYEr023+3nij
b1h6+scRkPzkzEfbQ+RfD15ZfKsWjldkfOwQPtNBMAkYf1gLbwm28ke5PU1J65rc
JQnMOpYZD79lOnvPO7Ai5bFg3qcjBcTTrQpyAai0Zb41SwzCylHPVANdz0oxnvWb
3p1nGib5Cm/wnRTFB685n6YiGXGe3o/XE5BcuAN1zn0/yrAXwh+opalOFTmihSCV
rIe+nv2XrGap+YTyWDLhUZknIXruTUuFdJ0vGkxm6kRUYTrcQ1b4IRjIL4hcBjEH
xTrXeZaReoXnQmbnCrIRol0rcXYkIYBbeTt3dOH0+6YGpSorMPQyYMRxxV9k5pry
sa7qj3zrMUbhRuO100fO9Vl1rmJ9EOVlTF5PoraqtgzIAMne5aLDMXlhyh3T3K6F
RhOwilbi33KnpzZ1HcFNh6GKhgCzApUXceyVCT/lnKa9wq4E5rznzlWmkdVb6dVM
PyM1QW8JL0Vto1dEcdm1EaQr4Z70jeXzow4K4zPd2wOFwVgLneNCVryV2mA8u5tZ
iLZ2x3LWcIkxwH0X/4t6Na56JtWhWJk/Uwc8t+Q54nRatM5jObXrHv6Mj4BWSfqR
H6tkJ5iZEkYaNB9p26sZscW9jWUvB0lfQQimom+x5osuXDZqf8O2Zn80aIiJYxKM
oCmRvTxbvN68iyd+16RaGrj7L4+Pp5XlouokDPbIynvYFLKxiwfhTXz+ClWb/LJc
pxJiTlcY5mejGDbDadmEY3/uiPuzFbzIJtg+KHsl1apVmMP595qvbUwN+u4i7HL1
WQxgC8dDaBoiay6k2Jr+TbkbURDypOpwpbzcY+i3ipD+hK3INlTUxiKdLsI2BSbt
/a+CxLfihafa6ziIncceb9LRUsEJhCSqo0bOhMMv9wPR/JAFu4SZSXgrDlhhZkoR
O9WGeCCrOTDMtJ7df/w23Q0tL6xG4aEDiyWi23jfKxuZ62hpb7bWyCSGDFWBQZ2w
2fwOgYVHyl7y4A8HiYZEABsTd5Wxoh2dLhRklX1mGOb549sAPMqv4zGMqw5N02XA
g/TVkVujz/dg4PcwZCuY3Yx2mLYGF+ZMoh9sXen9KyMKNugNhJP8CjYxgejMpBCI
zgG9nh/6XwZGsgM/m/If07JN7WYsjeGx5USgRWUdqyxc84fa0boKQEuBB6ek/HLC
qxSiPhkejg4cHzO411oPi2kBStsAIABIaY+YtT5v/pk/g0NIzYqTZGVk1R6cmvou
s8tZkoAh+VZ2DzgIWGHB6AAoE5GoaQol3QJpIoMeNRVCj/SiYtjMBPNXOP69gGYX
7Wpnq8BlzNkdVXkjX0avo2GNX/zgBOA8v3i8kd/OmCeS1Il4zGN3kKAUsxVJIgpG
OIRdFCQiIrAmhJXdWpDYlyOar+S8d57SndcbkRuHQKm8no0sNfbkhXCRbkp+l8br
LVukKeH40YwVsgcQp+UYfe3rCFuGikcvFZE9pMzf+u9Mq2G/CbuB1nKLUGRtaBcS
wUgusJXQ3AaEqclh9pTkH3ejpThnQPyWGNUrFE/NJ2UaiNMfrwUjpD7wE7nFirbt
tDkDtu8FyyHcsEJ6vAqRHHH7vuerUFASe/xmJhEZVwWg4PdFpXnnF8NliY3hONXA
E379vmJf7Q6JwccxMt6DyvYaZldWXmPQ/kvw3h+0vzCZyFYPkEOAzUXPVECQFEUe
fgEUwK8ImtLNUGOlCaXgj0kdDOJJn6Pe0uePLIujYm21yD7EG4X2VdlgaWZJ4a5T
vU1HVrRp42yGe6z6DIBHHlU/GhD8n0wJvu34aQDRPESs7lQbn7xDXoJv/sd5+yIQ
ISV9T2SNbv7fsgzvCAuw8xaQpkJTEYY+eG9tbMx8B31tOjeOWr9olFQjab4qYgYT
LvtS/ytvdj5MijYgWinEkyp/B8eh3DuGwSdA/438OEif4f1YMUirPxJsMNf+/kE2
4bdpZWzaZEYBabqeXUW538gO3MIwgSh8EJWodGRqR0KBKRySp1B3qPxGCecWoNHb
qPwcgwE9D6H+ML1sWpls7prpvzT3VTwiqwpfM/bcMJjE6irDkk6BAumfT3rYFued
rMKANLranCfS3uIkFN1IHBeVWy+cA2wNi9Fh86Doww1ZRSNN1Urt/BUqPdZndPaw
mXxeVCje0q05V/6tEmJtFzqxkKCXwoMO38+Ukipl/1cYgkZvUgiHitYlchJJHwKk
pSS0lrqrOJtaGn2qtyyl00veYxn1F/2FmwHORzLQVjvR9Y3sg/hZvzQsBU1h4sUf
aTQyCaKaFk5V1WCP8Sli/YQebbQn34bcptCT0rWpjE0oIxS2dmqFBBVIxftOaedb
QfAoO5EMqcHKW2mtN1TwdhOoUiV78MTYHy1IdH2zgMbj0yjDSU4Rqk0kA6nVVkZ1
e7BfIWekZUf/L0CDOYx7VO0kD9EVOvYBxCX2LYOy+w9wDBoNwIZbBLrLUlGzEsmk
cudUqpf/ia2Hq0lpT9Dr8JO7jcq1njhEuOr/sC64C5O2PPP+OFT27a9flPm/CMHn
sFW5OOCs4trP/wIWfmblocjeB+fi0y6m7c9uvSJi4kqvHSwd7XY9Qr+8V5Nstf5C
wcF3bO+/Ibd832M3iWwL88DEvhrKHla5txipe+NNMcHWQEuFl2/VbqBloXV220Gx
Wrh1usFpF3dB3F4DK+Y78FKri8hfY20/eTRaSRH01F9Guiewwdf9LxIu9SDZ9h+Q
XhLpWL2LjkCyXAu8gJ2Tgvs8+rQDcQmHqnH+USLOTxge2woYVrKoh+V0aLbiicoj
SiYt9dmyQKY5VIzhUm8hvqSNWDT62rZ6ixtHtSwcWllR298Np19vF4Op0J2cPVAm
nR2MLZLKs3PoiVVGGKzgJoXYHQfUyXJKa5WubigbiFd2Ud/1SFQJTCG0mM+E5qpT
DtuyrdFsuoCJFIDdL9Xyl4i5IdsxSmEMbeagVfKIte7mfmYU81CBenHZWFJqUQn6
bTUBfHmEWKncX9nbDAp82hfjf8NQCs5by1n3RD0XBWkKiHsj+IuIh66n2GqgjAeo
TB2FMzHNlL2WBphq698eC6XbBu5BPwCac+YlC7IQAofur148JsUn71Ln3J8xOQsA
K6q17ux+hzioOP+18p1Oes9FYaPCNNWqWJKeDAZhB/xXkVnT4n5P2YQDy1kXVPgo
V+lf2f3nsCHQjRQsEqpy4L065YIY4Ka1KYZcW9UHz9OCaHE0NZTeX+EKdSzKI0vQ
etmRh8DCKkQeKoR5CM6jtW0GXJBN6yyY9Dx2rGE3S47H9hh/Frbf7FGoK+kiwiHF
KTRTQOpnZ65o330vRAe/iqWBDiR97km/Xq9oIyC8yB1Q/DoKy0GMHIFulsAUebfk
eUEWGTN2lAR5fNwbmy/vnbl4xWK3w9AKQ1YF7GeJX+4xKffBwgc3yam3gB7M9bbI
mrAiDtxqNKQC6LD+d21RtEZ8v6uThKYPeD7x6WdjiBAZGvo8y86LbrOnBpSxSFN6
TuqtsijJj+URMU5KGESL+xQShasFJLWyJ37Gh+A9HsV1oAzOJsVEwwROWhtSSjXj
V5PpjbqLtX74liqrySvQJhQWHu8fmA+4l1mQLXZbO3ez01hx4l8ZMQwB57VKcoFb
um0ts1YAiacXbgwyIj5L3iWPA37J0XAdX2qJ+amDlzpVApP7VyeTQ8MYV5HomI82
0/Z1B6x4uMidQlYCa8zS5tOUhUT9ThAD8UjXGSQHk/5RYM2M6M7dycVZoKmn4uei
8OZop87sPsvcI8dWl7PSMcWW0/rdtmTngNYorClfyaCjpkbHFl/dvTH9FFVBSFq4
ufR2GC9mN/o6769REqJK2gckI3/F5oYV7p2sgjxun0rAjAsnPJ2rGqPt3tNLnukB
WZgbQvDoiw39FFdToEbINPYlTB2CA906WuR6rFeBThWPgzv+6IlMIwqxgl8r2CWH
sSF8Bk96XiPFbAL6LNpcSrWkxyXq6WNgvuB5nIYHV+iz+IVczDY6KmSKvmQIyFCb
2RR+4L/KHkP0bP/do7OP6WiWUFmtMRnhPsuRfhovIYjnQ6HIB2htQhkfNQ9GABL2
j5L5E3qBi8WTPevc0SzvHONXXktBttGwJmqx9ZItdGCM08w1vZIG4IOwZkRdoJFu
XXim/Aa0BecMtZYvw2TdDTBt7A0Ex8/FK2fw1LIrYtfyoGeNIHmszj9bWqZBybmi
V11r8xDbLfewL9EhP3gSxjMj5vyo5HbxW4BogyCx5FJKHgAVnmXHEKO/97r0r1wV
rXZeGcbrWDZ/VM0m6leF449S4ObvKVbyns337yPmCt2uev1ssNzrQceDdqtpDavO
XHnFdVWa/blhQ8cKiGHbWywwY9gbZgVG4Lgc+brm5zhsPqgIDiE3TOQCKB8ZGffo
gkrseOjtfKCv2mjHmtbq+psOPbe/SDRm/S81bQlhC9YmuaiZ6Qd8d86qnHfEvkWU
eeHY9iK1RKia2LbwOOv33+iFSqvk+cwNsdipvVmrITwVdaGgjExO/M37bNHm7ASh
SxjHrf/Gmqn1rpkzDcUp2UAQUHs/becQ+CU0MzNPX8SECyJevCn1YQ+2Bec6Jm4w
Hx2AW+qlEQi0jd5ZBWtSQLiUeikHS2G5zlSP50xfUSABQvSSd6TyBNSa7k7XM7mX
WysO1vfTQcM1ygRik6Knd3opFa/GrnyNZzGUSqv/XUjvgp8qKGA/Xw+wUSEIezlT
qqgvcFlpmdmVxGiD4D0qJZP+qL0PLNHBRAEFaSKUyngqEBQ5O4mdggqp36gjWpPi
Mv/2Q717uM+7YHEIx3PGhDGbzwX4evQ4QS6ueG7ScCsxI80G6dnNwGUXP4l7r5h7
stle2zNvrtjxOZWn7r708VuA+xjLQhjbncaLNmW9bLrW2QGdxx8XuIwpynKAQ8Uw
pQY0/2Aofg0DlvPMe7d12aq3C3mMfedMW15EQciQkn5TVoDWD/nUleinSby6vFEr
mf8YFN5Z27ywxzTdVwkfjmGwScLC0PA1/jdSIddcFjI+0HZfvq2D4A/VCsg7yDBV
Z6S9M7VyXcYDwQCd9LGk6UDWQY4XF1EPX+bCN6/uVCFtUtXx10ifTzFc8i7ztcYS
nU4LS4Nn1FOGHEQfhujN9eA1SHr9taZnxrXEq+TgYJMd/UN6ce0QXboYFBhzEQ5G
RGIPtc0AfSFkpHdwV0QV2jOEsHp06CA9Zn/L8aLEj/aRxr9vHRRb+R/cRupDLHJm
22uZSzcWdQqGUVR2HV3IEtGx4QXgxN71bX7dmHWQo5KkwZNm1Z3KZv61cpqFKwHI
4W0KF4BiYtfO3Ob78Btf39r7+0dKN2zYbQR+GT8ovMFcATPD5xaO5MnkjNND2BMk
adk8eX3N6vyqQpWbOPNVMu3jYEgA7alGMdLxUJ0ed1wGZu/ySyhQ6bjE7NzKsSHw
AANDslE3CgLUWYhk7NCtK6GA54yzYsjcDEtcAFKYfY9EhjZfeDS49ykx9qupSVI0
kHINrIZqgUyoOhtSs8kSrDyIx2vh79HkZzV/DZpU5LD2H1X3E+ApT0eFVO9hwWQ4
h871gYyo9ac9jVQvXbfsBKnP+k8JBCfWo95T49SLjpxQZxDPmWBwwEAeu5/qZaAD
qu51L4G9WC/k4yF230D7BPzO6DQtsUKa3poSqXCFjwj60hwO/ngb72e0Y3Wt6/kl
Zij/XTm5xyd9Nj7SXwtdBSvSmN+BxZPOe458OB186Ep2KZMaQggLw0XjxZoLXRxf
Y4L8PXJ7RsmlI+RCPYpi4Ut3WaN1sreggbOSl/psAeulWsOxKg2FB2BMKAexqUUO
OH32ka/yBTmbnHjjIoAf12VP0Xw/4dBHk6S7W7IT5y/oRuwj1ODxNdUPM1IKrAj7
7vD4ji3ZG11o3v2KSAKTnIpyKrT6sJ5GzR40De9RrvvX9ueNQH0KHB7kfx0sD832
s7CoNzPWJ1xAjR7VczWKM1c2/WKQe/Tbyy8HOm6E+Cvwl8kLm9DXxNwTvfae1z5M
nUvUAJRBibYmNV38R9FR+oQ1zR1LQszTROIvVmM0g62J+A8Q5O/pA9AsW2wOiAFt
NKrAL+Cont5SS95LvTpZVxe9hlUtKoq2geou9BB2QCQpZMWPctY7gGelJq6sN6HT
G9NzaUfHVNlwJAoMCDVKp+6YfbtmEt7oJurwhYgluRq9rkxVOwWAmsReLaL58BCo
s10LlD8jNzWDRwpogthDv6qc+F0Tg0T3flkhbS+F3Fvl7aZuv/2v0uTQZbRnem2A
xTCz2/Zk0BMwBzn4K7gW9jFvNwwaoveMuxkBO4aEEcW79efugEHw5eULtBfH6KT0
2R9//u5VidFMTGZ4s3d2v0abrbrcqNsiS68dWKKzj8ZvyhiEgcg5LpMNxn731tx0
IvA3EK39AORrIzyidVqyT0EO7U4D2n7pd5JmOgC6kGp9K8kYM+Sl8Zsy9nJBbMYr
gStQUtWps63TMB6aAiHLpDvgif1egCCYq5WFUjUkRPOKwNJV4kTgFf1bfIK9Kf/o
T5dWgiSp9X6gmVc6qb+3I4zRsHKBDXi76qoojgzD6nZ+kjnWzQgHABWxTOg8QbYD
N9TPom2w99miAzdMZ2S7H1XW953UXIb1dReuavurDdXWBmHZsq+1d5xok3EqWSMV
Yi7rhSk9n5t7TKdbls+Vk9MUPz9MGpV2w7VZQINfVhatQlZ0rrd9OM8w4/ZRovac
9XNKNEDvoi72R4jqq4V5txQK9RRTstm/9f0J0nY9es7eycYV6Yxo69I6lns91clH
XafzFJiEEdEk2g31CSXTwbYAwj/RQZVoEe7RQAsnPZaE7MAAzarA/0P2evyYZPaT
nV1qER8X18rJEXkLPhKRQYDaTk5u6wOdU9kDcb0uQ+cBU6tUf2/XcHYNapHWFs6W
hE9epRLB3YF6me18O6xfY4ndoUe6Z/LGZxD4h+Hh4nQb4QKPPLs+NHfea+jal2zU
XlmhsMr9QyElHga1h5D22OBCCnoVbkyYW4bsigwn9ZDfkKQ+he4ns7v4oe6l49q4
hO/4bIQmGoZuirbdQLUdmgGi6ZotJADSAK7y4V/FpT31EkoTAs1X4CC8ES11lNSx
LjmVv+MzDkf3a4PbrubaKFj3foWS7ZXJJ7/CiUIW58Sqiik8E1uAqGqALhcSP4Wn
wygU0+mrI7U/3+XZ25yON0TeeMkRBW7ygBNOPyrAGrNVsb7aOy7VmMQ+T0CBSlj2
1Cd9i0ZmDZzaN8ttd0Ia+NhkoASXdf03ZUgPpLSw98eSYbG6XGfL397MlImsmXt/
P32szERD3FBntkh5cTqq8SQTbMwSenn+B9jHk5YyH2r5dYgbA2Rk8GcIWbQQ8Dmk
Q5g6V+6fbo1nccV+Z8OZQPY8PDoqAHTvSpddGG13C8bvS0Y31qWVOBdi3TWaOkNt
r4sh32vBOoJ1VJ53udx2Gh/RQUFbMuLbaLabJUE10Zc+YSZ9ZtCM3uULTuVNrLi1
rKvW958jwhO5Z8ojxf3H6GmmioH7lofGkDtMWFfCkxf6B6ZId08385YpDT+/kXv5
H/toXXMyl+eLolUtBllIW0oifXxPsBUWMs/jXez9G00bMdP29dQax339ixN4HWgQ
sdrGQoxukEaylHtGHVZagDNys06nEVnzRksXhCZYfT/TSDPzOHAlAdHlZ9qqaHYv
/rVXf/kcIVLBfWzbxdnmrCNsRf6Eqqt+ifHjh0XVDK2Cm5fZLykB8z5Lg9fwS6MC
LZqJDOl4b6rnEvAqjMIkGS8W7BaYVu5naeMd/1OyronFKADyN8eM8+HsSEfZHZlu
P8/ybOyRZxYpoPyqXQIwzabjRDJPIBCNOGrwDOAWK3z38D/YMVlSaZ2oe1gqaFIE
5Yi5FO1svCgma+qJLY4tJhRZHKNU5XT8uXw/6u74bVzI3ZV+CkwgnAJVGqCjoMG2
NGmsS1h3DD6aeRp10s9bRuicRwtWEuBUOP52zz6W8ScsVFGLhh2K8dCpKM9hrd5l
Tm7HAu9sbxBMUJ2XreN5Ah4Xw1gO97pEA4H1kt/Net6D150cc6Ql8Lky7ATORZRi
mi6NwLYF9ogbq7GhMcvPVnQF30ZD5ZO75D9+habMMSWatCs8zsgG+bwZxcbaV1CB
MV/bXpHYZ8+6OwfuKlf4mv8HUeZsxf9ro5V648RV03kGow8/Ojw3Y3zHxD+wiDmK
bXlRZ3ZeyASapHfRgEE1fn2MAtfeMUtQ0XVnOLNy13w00QbfZvFVSlQez5SDYgDy
EaiBofbpDVdLy0F8DkFxKsuH8exkTo0i0ZITmqWBfVq57Don+sERTE3pGqIrFpDM
zvFh816OMemWFSz8hGPsZYd2rJifrEtC4sRqMun+7jhapA16/gG1ld0nra/l0r96
wd7tXt/ztqTjH4N/yDiZdeDBe1kc/KN19zgwdsc9Cr50Q3WS+0livhRepki/vdET
e2z8SiQp1iQFCsP+MZeFnn9WrmwJspP4dPRP9WOtM10JgkSeqpatV9j2jSxBj7Gf
lhku0FInvmH9rOZX2MK95GXriAfFcPN6ElWQgXyMJrKDPjXMOhFSg//XpuYOkVVd
9EXwGJqZ4J6fxp+ELSz/CJjBRoyPeeA1JHB8fEjhxkkq6hOfZQicUD6WMMUSiuCC
DEgxdewPSxmMcuOvSeAyxwCMt7I/CPJ0FIiKbOdvqVDTy8CFPpfYcO+5wsRTFdtM
vqdZ6YAgTKds3tEYI+MSps6og0ZjUHERgi+1O3ygT8X8lrKSHqQz8+vs5MuqxZxJ
lTrWUzhRbL1b0AeDzsHH9n53NzoOogKdA0etXw9E20tQ7S7/GwYhYO+rGQlA2H/s
XqqyxK0Kj6XrGsRwt7Qot01GjfwL14upDRaWd81pN3RLBGfChn13rteojlz6nxWm
HVx1CDla25AWLiTpnTkYbqOrCP4cg3De5QrDN84XP/r8hke6bBNWQZrlAKpDogbQ
VNUjIY9S1kVgu588jSpaogNBH3xtl74F4biRH1qigJsynpvg4eftZmvnB2VG9oEP
RzvkE9nB5x6IY7aQFXxYD4/KfZMg9dPNEMcuHka3FR/ApN4vuUFreIr/rgfvmQMm
sofY3OWRhaixx/jrSgeXwW27F8dGogvOinj/xfkakdNrTIeNRnoir5QN52lQDJjh
XS3STtQWAd/WaW/vwUVWvMdQu6HKpgdeIPpSECQSuBa20PoPvIsqB1fyuwQZCzUE
zO3NscI9779un7cUfaMfBA/lQCa/NKcEHfExSYXjX3zqGK3JcaK2lXhwFrI4Kssp
qRVYnJ47lAaFkdZhBqUb8Lz3UnrLO40GTI8Eg+v5gslFo70s7LKv0FFAmqFPchL3
EBAwKP9Gywgmi27Oda4uKF8Tpcji+VOb9U2SLqEgPgE84ygdGY7LZ5ZhC2TTQ9Js
/a5fg4LoGhAy1hbA520ch9+Fs4OPm75x6MkCGB1vtxxsbCD3i86MxBMydoXIyPr4
0nof5zW7AfyldPG4REoFx475x8Scj1f2J2QSAEYUgPY8ombzZEg0Is3AhRHreJgl
K2DVEaU438nw5+b29T5+2D+FyTnaGtpIAYHEe5rl5iBIce8aFdg0PxdKKvvfK5zC
pVnisrtK/5yu/FCtCCMrmtRUS7pobkxMYSMUSP8Ud7sbujaFw6fpTlc+wD5nEi2D
jGmzLNdm6dnYK0mVNgn9OLho0DdvTBSoQS1h+KEQ2zre6w7MlLtUo0zCl27Wnnoi
L3va2oolUzJW3NoJUCpmfffJz6Op/Grn0GF4jC4JqG6aN2YR5FnpTLkINjCgtwt/
Wo0wRY69W460GJ8cefjfabITyIcSe3aFptepwnnFBbJ/VzZmw7asAlKnk6N5gfh2
IzszR8gYO59m2Kfiuj0sLTyILlUNS1PiSnRGLbxrpHdsefcxKD0jKfhQHQVWJIkH
19or+fxqt2XTnSUtWx+VOMTFDFOlXXmhQ9gWlK/RHd90uE19KCKvCkmwMuO7ei7S
DUtIfjFY5G51GmnO69PygqerkQK49nEPH3sVMvy7/+pzCpOLZnHqBcmp9xp+qpFo
6aBfIAQIJYqXvrfxhaRExov5w4Ecigo1vcuuHFN4fZDEdOKgedhNGYAqEc/xgwcM
rGg0dMX6TcLkHP8kbmy/5WqrzOf7q9WWkwOQ4Cakk5KFGIOMgq5Sj0WTN5+whlJi
Rx3hD6XAWODTWYFC5F4ecxkpT4TFL7ZkCFwoOXHOFyHiRHF2SncTAhgKB564knZd
I15aKso7WDjbkVXATu01beddh84dhoQk5Df+3WgJxpyx18QN4WwNF6CFOzEvAFU+
eD/L3e/GuheR23Sic1jwXeD1gc+rvVdu+DywHo94sLKbJ1mu8a65LYG64+6cP/CM
wli+hkvzE3ZtfijP24kdIRhfOhl00ydO5dKFs0uQ1i/57jDXdt13uvX6KJ8AZIn9
kiPOBqM8VWGZYo9vL4EwR1l1dxEPxCiC/pe2Nh/p+a6kUqYvV8QY432838G2GD2q
w+nWhaFqM5cUVfBOjeREiBwipHlmrht7SY7OTati0EvYCLbfsGbKlgT4VBbNaAUV
AgyT1ONUSjiwklr0v3Cs+sUhp2WnOVuWuk7vdzoqujZ0HqAkHrQBfNynfl0t2Jic
qfA+OxhYvDYw4dUD/7PQpxF/lqzPnGsi0WeSBQVGhP/9Q63rX2oGrjP4KUlB5z/v
33/nq3xe0qng/qOXg0hTPouFRlsbU+CinOL9yDsuShb7dqw0ByzstHAnYgHtlPJ6
RA+KsTZNjD4Dvw6fSCv4Q3gOJmFuxdyzFu4YgRBEWsxmfO6CKSPm89w4oYjMRRpu
NGp6ey3KtRnGuUk5SyittH1wBWPk+yuNWM+2Obu4xdNdnj5+La8bdWFUDUrvBGZx
hFd3sxtIpcow9rKgTS2dutRX/K0X3vKPlPAWBr6AEki5qgGnfN4JDOij8WZ7cs65
81eMnOb767IgYYlWz7Rl81UF5GO7FRiZrOnRMXXX08Hw4DQ5zjzEA4Q+4MRnRcRj
eX/JCLBW0cAiHtI2AHVumBA/2BPrZXidjb2CkvcLuhaoMr0qIsppZC1E4yJhSntw
axzhELP+/KKIcgy6kjOpU8usYTKbfBUFGZR+7CF1+rZPRdR54RMie8lXeS1Skn00
UAOPvhAFCTaapAujjZ3PLO/HugA30b7RH6wAhHyx2EaNbhtoOSgpKqDHX4AUnRYu
kQ+Wir4vkU6Y3xsKT9CBT2rPUFXn5VmMBCmWPrqMc6qFauhu7Sw7Gu69qRKMMv2J
4CvjURQDGj4Iic1rjcQiHjW3I9O/nZslmpvHzhtLOmQOoIoj4gdOlYHOjvJKNr9R
ww1o42Ry/UAq8QCTJzOtSasu+3wracYEp81iEcgjnjSjchKNDLyafBnf1QDORUDq
doRWdOx+U0VpV4DV4NmWe6UQQNkgHfBrCBizOQ8VaZDkpFcsoH9Oi2hsiO6oUhv8
a5gDm1jeFx9eVakFEkURXExS5LOC1GEt8o91AB4kUO+66PJASpAkZOhhG3mD1s71
aoWj7BL4hCMG3Ul6iFypQO+wrdMvyNy11ymgQ0MBtSrsQZwSA3r4gJU3RPfVBShi
ju/v/xAkAoUn2vfzWPYkMQG718ShNZ4twhtQ5do7uzJ/y4QaYn0yfJc8+Oxn8N6V
h59hlqRUvljq5c2pZoe6NgNrl48+Aqv7ZQHfXi7QYRspo1bpy6c0/433hHc0V/mY
mJMmmRYhjzfiDcGz0dify7Ckw1XbYptcHezpPXRHOt50z+LeLNeddx9Pcw+4y4vp
fkZQuKAvqafv5v0+enolJs02dDAVHj3Vxce8eTOf8573XkosJ8B+m7tI0L/4IsA0
kbyR65PTMPFFt/8oFRQ/Cs3eYwEw+s7Z9B5kfIimOL9tAVMU4LTRdIIodbIun1uD
slSCNkyEBKa5cMTLTJzTfH9MEzKIPb1vfNy22monnCetqsiLdWQ7gtLHfiQDIW31
52GwwVWbLk9B6Lu/A/I/JUCOlrVmF6DCxEIsBoDWgbrOSOMqDWouOUenQbnrrSMy
Y+DGkCDBqNkIBeFwZRCO+P+nlmWPef9v8e5Pdyq9eDNTMEWoD0LgOzyMOG0fQ3xM
ld8KOxENY12j33dxje7/ul+JLUssZ/Hh+xATr75YPvw9gU8BJ/wLJNdWtb72pPuH
zH7Ttwr2X+8hxZk2Re6xfQxiruAN7DxnBD6CbSqEw0CPXR9/HgHxEsuFu+EEneTD
O2QztT5X5nLtAG2kpouh80/0cOmOF4Hs/5Hp6OSmr1mMPff5n2/XBQ8EB5R/GsBN
beFonXq9PKfda/DMmd8i5KmG4a1lQnX4b5R0I2orV7nhC/IdO/h3NMF7fIC5ltMU
3h7ztL/Ixp4Rn7uHlWIXgKZZPCbG7IaPUeyzFw7RZPQ+wYag5lmlpiffBE/Xxdxf
lbpRuxJkrDUwqfhRg919WAtws635u92GolKFPlzTl4bYjHJ6K5uUMvSVwnP1S06D
8eOtUzCfBQ6s0Zx3Zz2XrnBm+ajjBf63d2hGF10Jz2ipjRMcIZH7Ow7nUkvpR7xD
t7fun1PHKVThrNKWwyCYq2RL1JLqRNdunWgID1E5MW8O5CGkig2p3d0Nq2vAkGEj
fBMUc9FFn/AfpR12fUvFC5WnU76mIcmGT6axHhSKjaio9GfOzzO2v0kxW9xymDpU
IJg8Slh6tTNdF1dZyV4W2dx0cnaUq1T2f1sJ5RMjDT2yiUzFYrnAPi9wTo8T9EIA
Rd9B4PCpyFk9oNdjYaZU1vKXFM9ue1yQjjqq4uex5Jh9J/J5gaVbggg06pPy9DBq
lH8b3QqTOA5vc44MUY5lsuTxLFpxTr2m8Z2KYXaa60wkqnJlcyj4Ari3kATWl26x
QlcXw8rZ/V7hljUzn7RHfaZnUgEx1qXRQyj+S0rcHcvXPeft2GbINJcAviQBN23d
BXtNCix9jTbrXgk/ZW+t+mdNUnaNDvipSapvLY+xHGKTpZn4cQcZNUutlHBnx5lL
NEahHoefVwlLLmI+qg7HXb665kDawnPwkBLEzoMiDGgut41xCHC/L/W3rGSMNP6T
qTxs4esv6CvXcIYekFMePf3DXqr9C5rEAIxmM9kEmk7x9Z05jBqkFYxf/SGqedZL
tRCxbo/SSTYFxJ5RBRwXahNjaLkg1gQ6ccJAC6eL4YfwCX61aBFo2JnsMYXMkM4G
KNOK/fG/9OTVSuoxBnHkxO4ogll+ojLjn0qxAgW+UBo2seXWR8Yju60xayjmOCsK
pNmf45IUbEIFMHkIR8rR72omCoXx+OO4MmGLWbj4Hy8Q3wWrQs3h4qjDzlq9Dx9c
UPf7S0DFpVPtgXbP075zKHTSMgpjHSDfLAWcKE3w08EKTXGJvJs6hWlIyzBh5w4O
YTDseMJ+1CZsN4Zy4XsqgHieM/ju+NiJTLlL0TlcvOewO11uUFFTWR5zWjvq41ad
w1vxTMHY87BXUnMkfJkJRNTRHwImKgQ0E3h64H9LYhucUMiGx/6cLbW/PATVc2rf
w+oeMW99qLJcH+JTuy1a6QJMizwGU5FzpgESRiMXvio7+kzddFnog5+0G2/hAILs
20LFmxE32QTPPaUsdQ6KgkJnDrJfnjLOfij3SAqsltru1Z6yRiNd+O6iV90S7/+q
O1oB8mliBUdmhkBuRL5/FY9vjalFAne/+CrMEwhhr4ifBPkDTVcSoSfB+9w1NsDr
pEMsOjl7B7XHvpHRLmNY09elcBKyLVAtp9U1P2R1Gzx39EIHX+XGnGyJEiKty6qw
FozlToLFj72beEd7p5aHH896389EzdOYdcIRvGQ8xB6LoDwh2lrrNzpDn3GBypVH
B04fWciK8yDnw69ldeCGEXLU2/dyJftZ+CJLfXz51A4Q/epCxHP661UqmaOnAT5Z
wFOMuByvtcXvd3OpmK+PIJ3ghuVdTxL2l4URiqZ6yNrgNG7O7Laiy0L+XtS5/g+0
I1Zwe7CjrNrA5xH9+xLSURp32fcTvR/Tks9nVn7UyROPAMqoV2rNsRitaCgUkxqZ
xVoDl51uY5Dk8E0eXJxYr/c9VHvDFPjSXzwrj4GPiDcXM66hDjmN9FXegimvCnb/
xVUYUJ52djNkAc7p5xh+eVaNoDbtMRTfKYs5jh/CJSkj2T+GXRBGliVIu1sjyTpM
wYVODns2WCNUqbzoMDyfXA9a0vhRUv7k/9qTYwDzGUuhjaOA/hCmhTyX5QKy6y+u
4RWhj/ZXkIMJhHcusFTKtnsAAOIcbJ1jiLwkolamTGnbQK6MVC78I/W3DQcpEdkO
3upuUjJrbLc69YQNd1udaOfhDE1gHfXYOVdtI6g8cQ7zyJQrd00rGCq45OirB98X
TGO/WA7gApiw2lUDxR6sfGTAY/B90M8vKPxCPh4MbTgL60cifBeT1udVHvyDAyB/
7/kRVQLC5g/8mX7fEHSQluN1OwekoC2GzlwDh0qdy04AF7DzZahJqM940NPmPQ8P
ada2CeOpa4ekqvAs0wSAFdppCxJMqlzc4SiuEi1xFGaUSeItAiToQEX8ew+lHFrm
96jFO6YMwvvKOcDBHJ7wvZJTjGYjuFtUxiNfa5a1jDg6UW2e/YDjL+xYA6g11S5k
sUNCNNJCeYPvX5Rrzq4Q5McLjBU19KFU18gRPZR3XpXEQk+aeVDxdGQUiQ5ycaIc
4TtZa3jcdKhWco9bqn97EhLaForom6uIP7OFJaCw5mxELukRBCsmM8p7Iok8qiQh
iKb8S6dUiH6q1mjqQDVfwghBAbwl51LkSk6JbFOHTB5r7iSAfbOuXgAldMmcra4x
V60SJmcaVFn5Vh/d1K0SFb+XknGElWrVxHWYvG5YmsLzHzdRkdh+G3LJRwYZN60R
fpePAL2wFIUe210/e0LjKwAaEhrJvdiZu3RyUXH0BqHvcOg5h3AgVUwqmqU1p9zi
DLHjzXk37pX0KSCmomCfQXdXW6N15cwgjYGSXCArc1q13Du1eKVfiwOAKMMRq4uO
G7ffcEMWfTVpZKch/iESauSMs155RKOr6eccb3J0Udr1aLejI5DBhQehpBHkVyk+
aZNGVrTnW1VgBQXO7MDJx36atwE9XkUhZgqn0jPt1Uq1NebC+qG2X/PZiGPNR+wU
F3pTGfADR4pll/2x/72i3d1o0iU+GP9HBvgktcYz22UF0q7LhaPQyPFHZ5Q5mhCV
JTt2pImpBjNZnvh/IaCIi957PkURiz462egX9SpOxwTUTvNfxrTHkLj9OmFlBMF3
jXr2q5Tfi1bs5fcdX5fHmezehstlJYYTm5K4WEHRcDET2qQf3k9LvtPwgfkg+5F2
Jy+BuW/hSbadcY84R9QIpMIXq5thwT+GRZznAQ3X/WazYHmOdc0oJzbl7DhmsNcv
OLyK78hdHJgF7UO37dGDP8185NGx59unjBChgD/oqM35fUz3Hmos84MwhdsCHak+
0vYQB3709KcyGYBsKY22nw15IIk0zCpXTmB0kpoEM8xFDwdDeCyj8olJc4hIHbfI
P60vv9VJxq+doaCWpc9gUe8Cq983+6Ym1iMNclTm5zXv5ZS0tVqTdQsSoeeJdOFC
t93LlUvuWMkMfYyin6tRM0LfgCA74YCEiWWGI0LnhQjShcJ0LOOUFlosr+7QhZ56
KfgTa4Ck1Pz95Nglc9h3ivh4pLJXOGxrBd7OJ2QYdx9W5oXcBq3w70liXNC0oKBf
0nx3hLNp6AMNZOZ7QYtb/F81GAUVfpiJItsfMDhYZgsDN3We/xRmFB7Lk4ekrlhr
7a8ZXFQS2NvfUENTJwXxD2+oHWIiKC1MZzcs0wTwC3vdOGZBzHkEocch7wqUoO/K
4yFYxc7pL9QflKIG1rdThUbrgApGb9RmLbPbq9wpKZ11GsjZw5q+yBLc8mWoW+xN
szAYIHB6dCUMj5fYKWLyvPcsGavea4bEJkeoUgJu5cKIva2zdMZtnhcrVKlGVYbp
v64kYCX0ADrjOvBhWdQqQqiEfXeE/JE5Wb6Xcys/hrwB+hgElTw9474kdV4c6gox
VBt9gvsO1EQHp1VVlNMEq8pNHIqX92ditqAJ2hmw6YhnRWOml98iHzazx6RAk6C8
CvXHGk56dVOcXF+YEFI395saxA8DP8Kmt2B9wiEPwdX5DpM0TZh+wAocHC6ti73R
xb7ijhzjKfcQKoVSe5s1fDBswEgHPLe6jRQyLbmbhlrlVyu5+LfOkbYhiy+h7Djd
x+LAlB0LNS7s77hrjMw8BD/u5KSC98ABaQDb99+v0ZhfbU6OhFIHRVE/pJ+2sgGc
Vb+3WAvu1fRtQ0eRetDxwdpQSd3gju/LInzyWBXuGaRZRvz4FSwmZDxNvpqP/sw5
2BPm4gmbE+GSEtKT/LgaR8ybe6RWiX6EGUaWRitUoxjKf6nVH5bDrM8hvie6k9re
KlitWXidOcKSFSqReCmzQCgLLVy2xuqg8cyeYlW4pW1Q/uCSmxLFJ5hc8DJLrD1S
BydSolE2T716XKa2J5q4kHL6tOwn4ZITZYwC9VUwlICBUvEtGMk6kuy2hZGNVTzR
8ItyWFFeJCSMkTT9u/N0a67M9Pv7gJ1xeK5/f1DCwtaYz92xMlle++YlUtf1KIrU
6BzgnlEf3c4bJ1gEzyXA/gfxsqiMWAbeq9reS7XGkULThTEGHpDjDCwfJDjMlKA7
ad8oJGGVFfhzj5cu7cvsd18LOaobn12DYzaOTM32RSD5Zhzjcb4yFvNi7FX7vcyX
/8nG0O/KtedNNReeco46nPiPUAbMYplIClYEJRYYfcCDdANHleZ/DIU9JR4y+uXt
HC/5dO2aKUSlDj5K8VO+mYp5olHwCUIcEEopiA1rNxc8MSnBh1ocjGnOpgKnLgq+
z0dtS3ZujsLB9h+Ed8AxHO0VHliRG+uoKqUa3dyJIRTEG+Vpyh3yRvWwUwB+NArq
9gLEL1GS97oYUUPjSFH7It3bkbbkSk0JNrpbRrLQSZBg0xJwGiGLT5PWeuB1ji1u
nca0jfR49qBTlZccQ8cvHbxshJjGCbZTC2P00fcJ8feX2uTvuK+OrXY5Q0GiheWX
RW91z06+vMb4GoToam7E+N2kilHs65wtq8zwBs6OxLWoEFuyY/ch4ZAZ+IqCA2+I
Rb+suI4L13XQkDnEnHcbatjmm1T1NnUwY97fwDDLO+7jUQasLIAsajph3XYMgIuK
TjsvJ8+/mL+74nu6q9o7/XgxaeUA0I93YQ2Ufy3KPn095Zc4YTX5tyn6QsO0LPnh
ek6NShTLoJMaq0DWGm9arl8qUn3YZskoY+wiTfxzshfNytKgGta4HUaMsP5bi8H7
g7KdBwsQu79CQSSyPob2rxgWjZZ+vwuU7BG7/4rxfjHJ7lzJ1uX34QECG/cvTaEe
MbqU/Gxqhy2N+wIiuGE7/3k8T/3KicMtzjUpoyaDi0z1JaSyAuJO2E9fXgTKb3tV
UlZc/oPyVdTlLm1YGsDkICwqqt+6mzNFCfxvdLIVx+NPXAXxRerqxrOp/NoFpPVT
PSEOCao5CFmLL0tjBm9n8kPCRZpXH4Ev+VBQPTVz5uQZoLlMh4Vmkpjs0SjcJ/+k
ITuTAvjDQSN1uDrvJ0RXHa5i8su/SFq8ys9YlTouGW4QhVWCmyHLAHzmghUelGO1
knkwJ7fYOUxVEjCwEWbc5Z2BRf4h7nWJQqfTxQ94h2iFHu22H2gjg38LL+s8KzM/
rrGoh2nykbwUrWVvZijlV8wgwGE0roylzGPm2Tq3aea0rrMUHQtkhf4U7aE+RXUx
lRg8aVrdVFa4n+nUbCggKVoI1KcdeL72FXni9fQBMeb7Ypi7wyNftBbAd74nIICv
8BXZ55IYdAIW2hNlYJQ24bKsQ4Pz/Rk3bly2I3qfuUwgb/PWwdNw3f1z9/o0UL/s
iZF21oEySWtLNz3PTEQifuuWniep10mPklVN0UJXG10kGIwkn/Xf34J6SlObWFZy
KPH8HSNDz+9iS1JbDNzsZPEfvyQKjBxeVK75lsfZPqntbw6AlPpEbYpdZf1MJW12
agy3ttHx1c6/6zC9DGvM80t8++rldkVGfPNgDq+TnDlw2xh2AootmKWj9BZ5JxoU
aw5rAqy+jB6oYOXmXl6StOoE4VlOl0EerF3SrgMleKAGyA8fmFUgumyEQcElkktS
aWW6QdtKXvkeGo2eEloMuoWCwuyMYeBUW9c9HDahqAEhDxOKq7EoIHdBmSq5xSZx
OIFSU9vtFju6/rUXiI85SCqPUC/rviIz8BZ6X1cafmjYSHc5gxLQHlMdV7zd09lF
uI6LPS8A1xzzVnpojkH7yb6LYLP8OMk0XAqpdQQCWbhynfk9XX/HYFr1osJXpdLz
BSQVlivRwoZJNsEQMx60mNxjBtwZgiQ14g79LpGD0SfsPf5K2u33ixokSPZ96sKH
u7EkmFHSEDw8rOWbxsJW6VEUmTCvjF8laOzVj6K8AVdoED+P9ED5EcNAfxJZHVil
mqgZZESi2tIPjw40ECQX7rzN+bbQfsw5qx2Pe+KGRw5UUoWw/z7NsWX5UdVG2cfu
t/yTQas6gC6fF3Jf5+WlvLL6gh4BDI0NNHl70xVrDCabrWI/HARWjwe9sujMKz8Y
ZR51Qi2XyLCyRcbHSP7EBykmG/D5TMRiIEjBbP0wtc3O5rFjemGTTUxkXfZK8L5G
WkMh+3qHrmNSNBuGabSz9phzF9WsObgFS4giEIiay2ESR/TgW6YSvgdSrBc81JD/
K3chLg/EZz0ot4XVVMmHEMAyaIaZhw9i58Ao2JIXeB3hdmSJguYZI0oA66WtoRNF
CsTVk+Amug7DGPJ4D1JjhRE5tDtUn3R+Ud/YoH/v2ZpuHYdNI415ZQpljpF7Rk0T
qewhqMeZes/h6CFuzQ8Ghtu3BPHnhVF6WEceT6d+2yHJkwhWSzC4TTy9eQ3fmsH4
ZmSFWXqyzR+78shFgQlroJXAngv3n0w+1YNuFIuKXcX2d5iA6kBl2a/i4A/LT7CY
hnk7Gc9FEkBU03eYDIldS8K/lSwKnp0AYYXYriWPEA+abEuTbbxmaZ8XKJI+DmUy
8CU/iwjMVpebFM4IXtQ8Q7h/t+rTx584ij8XlgNifQZwcLl9uvwhhJgeXHRZPG3Q
5rA1buEccwjA6H2m//HrSN/0+DDfiIPe33CnPXhA7YAPy4RfmAx11kd5jCwpxgXn
krqBbga3svDXJ46QIQ6Gev+j7crShERMa4Ctz82qbN+zuxS3n7eYwjVycHWL31wY
5HWn+9NIa8hoDYg0SZfLllclndv4TEF8cJu0RvjElQsTfcGJVDopkDvhMr3jMjMk
t3CmN93++3mfj535E29DfGuRVsGw6y6ieqFhVVa+hhNockxoDJaw4I62DwkCq71j
fMc3SyPae0H/590tsKcIfywroxCVbD1GTXOj2axagnGqd1uSqDx+64KWe2zP96PY
rXG0FPrqp1moI+FpxbxqisfnSQl/KHs/WzURBVYI0pgSC6cjXAjYtBY3FVASupzL
NCFlJLCpNLIW1vv9Z2kPMLwtvKHIVArx47QYBXwXfR796kBDRrDJ4j5KKcOHYfIk
E9hh2UIkI4CJqecnDjf+VFwrmRryOdcZsn0Rox3PVPGR4Qs2nZO2fTRTleuIzm7+
uDhOHiIOreXR5KE5Mz1vfGmJTY8nLLI8gjOTCIbCZ1bDmiyMWc0a1esaVXzmWrCt
A6F6c5sztwSZv8zCvObWqH6XyH114oumd3zxm/e70IbWIoO5M88ylc9FLNgYhnN2
yyjVzAVaj9B9ToDYqJENE9HjZD70MhZpffxZKjR4OrC6Z1+CIoTy3ninYl+89v/6
sO7+uomqoFCOICjkDQd/TXrXrOqhZsmKlWNHfT11Vl56blQW3v4Nx6jidnylxNXU
oqkyOLVsTqCf74W/S2XyMpYMrty2qCrIZxlRSQ3gQiXdD/IhJvLpjhRSBrtEDXzD
Pou5ucjI3K2xaPkyTCUDLnV9Z4+DPDiNnsajIZUj49b8qe7ZOL0tZKTTqPzthoHw
H1RbR5crW8TvjIoRUkORE/ppL5eo9ug8B+jsU5XBjknhyQjPpn4EYqfZBqjueQlC
NkUKN8DIdHS8+K2c0wvub3BRpcuZHv/CpiqRNGIj9ToYie19hinrtZ+f8Y/Pm+Hn
iwfWhYH2dt7ImTvBHr/pd9nKN3M46FAc3JbqyMWyoCma4pUtN+4qZstReGO/rESO
zGX5Xg0ujmWDzsJpX8Q9FXFaQa/22xNyxbqMrkAz/plYuDOSQ7cJg76XpIqOZ0mX
GQMl8eQekyE2CdUDg0Qxal6lB6q01Y0DoCpQlF+BWppmSC4kdkF45U+rceKMBtML
XvogKhbM8zCzxH8EaH8D+Ls3DJKoFBPsy45LmqaFKshEfKDTLJyPpYwk5A/i0cUQ
/DhKUYqz0fO3+xzqJNZbpn22LVlUjosse1joTb1cMDol0YoaaIkbhfu4RAqlu/1D
VfFTal5jt05mJ/js9fXRR1GDLEUmQRlT/XJTvS2WZIHE3fbLlzTfN/rQp6JJ31s0
NzFPC6CwxkFzzrog7olKE8oQA3rqPK2ZyZ6ErJa2OVd24FWPfQQ3OTYDqFbLZQtN
Lfak6B950yA/DZxvrg+r6mJGkK5qRQOGGI7h1rWAHLWlJ/BQmu91EpJmWTl3NexU
/1Spn4tZqIkWFwwaf6LmGnKp9vW0ZlRr9OKEdi6oxJIh0CLsPy1DXbhPrYg+oV3c
EsarSHeyMddwwxdZ+YtuAvPREy4TWPZRaxh7LdAxNXqCWAweUdo0rjLV5h9jI3dv
qRrYR3A3ls39Wi/4/NjmE0vEMrPZtsPJcT2M93n4k3SaXcASqQZlJ8MjS5vVo/n+
EUPuwv06m4DXVqwcnXPfhu/VNEOYgPAX8vELGSH8ZiPigJbZlO+kRPE+0l4DcQ4G
rzVZGGfh8lHkM8TGZsLJdybQx3lmJ2zHiIgN0yw5fVsRQhWXCk/noF1iqL9ObI1+
YxoWi3poU0I+Qy0NHXxKHwS6OKnViiUr+aq+uGKruPWxgtmbL89bpppKBVSoYGGo
lMPo6u1/qzbY9bi2uAE+YbA9dQ490nVpJslmnJOdGFPYyhaQz+Tgf6auRgjhenef
axymsptU3pkOxzXti3vnv2fEbYFfgLeV+aYBQZDTo3oYhmA/w9n5j+SexgsQ2zy8
nY8182eDYq+lB2X5s0aYzQHtr+qizQlJk1u+ekhIsrUW71Ff/FBhT53AOgolYctb
WvsZSBotzan0u6Bqm6VlBpO5YhIP/K6pu5VACdfCKYtp7MVSAQIiMAFqOwrZhzj1
MpgjZNoapgHfX/2Bj4U0zkNg6Yswxr7BjvL05WiD32tQaE/ZYCbzh8W2rLJwYyPo
KnVJI2l3TJKDRBqECkvoeAzkMIk+7CD1lQF5C2jmHXQ+AYUi36P95fqDFsW/tVKh
odJWX9Qh3bN4TEVle0KNMrt/bjdWP12NyDDK0wIysqJb6+JrUaxduxAUpqlYUT4G
Pm4b2BtnQbT5FnR9nLjart1NmmR3U6uV3awQCiefCoUrbyi+ZKTfYegwWKmfAETs
qlpQ3KxDuIOJn4CZQyQSIXsW72IDuqGZVVxUgbQiMA80QHtZq6JwWHldYNrndCmf
npIj/ffOtXdstdsVrkiIzSiwGHu25olmN/vt3MOvlmqY4P3eaioZ4oOsalU8IIVg
aquGsfDpet8Ng/CBryN/HZZQW9HZZiYxw8rZgj/6u7UJ+tnpU8ELThdL0ua6yBij
sAuXWfvfY3Z/90tqw63dJwIJK/1h27/Mqmc2XxM1N1n9GX40d1KlYRCHSQ+z7dDJ
RX6c26REae2rm5i/p62A+1vkY+4OfmN8WBYBmLDjgTktytuF76u5HvDXMyOSjl1g
JVyH/Mg/8aQDBqMt7Xwrbm8ZQiOfqHDYvUnsfFvFTMMvnPCe7Tv7WLjrOMZlBQWF
Ju3arU9t5y7t9XTuzcWlf9+AnbF04kLso/mj9+UBLqllap5E/cs2JvoJznOH5JWc
L+fDt8Njp9QkMT2qzp0qVHQ5SaZxK7udHgpkP7jrGJUTgatifx95JaAXXpHkXLGp
bJTRJG9PxmFSQqRj48+KJ7SbJbVv/lncDQH8cImyglWpuASCub2Zmoc6P9b5OiJc
Rpdf2KAuICspGlScUrW9OcDPvdkeKqkfM4VNCZtkHQD3w7d2Qsqev09VVR99d2Fn
oZsTd8HZs5yUMHCJZM4hQDKHDMhvKUofYFR8EnNwYX+ONd6Gkk8mLJBZoQ1yG+3A
td4G4LgXj5sDa94QWWwiNy67p4kvRUpnKTIUkbcF5P1XYeuMMcHGGhAht3FzRzXk
PIFbctW4NGRT7xXPyU2kK38uUgJxHs+MuBGhY7jz69niXEB7SNu8C3Gg2ZWo+YdG
aPdXhLXEvC8My+kn21uatEF+htR6DqNC3hKco6eWlLMv/dESZzImrLqNCDiT53ez
aLNjK+jg5cuBTwy/6dQojPT8F9Ux9QrsA3HDr6H+FJe/raUk4H4Zs4i15/o8nER7
iXdDxUJjqC0Q8UmGy5+gIObw0izb4bS60b5gMFNYGNoMvg2G3lUYP5aqjMDI9Mbh
PnDYEGXWeQ1TK57bgWH9I7o9FUj+zlX+UdGV/OmttN/0wot96YEsNLteLKc8XBqt
E/jcbMuD+0T6MwLmUhQg7QP6PCzvULJu1G+X+CrgOoAqUIK3mLKPlRUN8WTQ/hO3
kBS+rB3imJPLfYcB6/5GfKOkJyfNNAnxPjMbFarJ8JF+30d5gZ55MLetNRLnAIhn
bXJtw22sDW4Ocu6pwwW27ksfpmZ+XXAkrx3TnJRx3iEEQn06MEEwWjVASK/8GCbo
xdvRiCPSwX0m5Hv4B43bDbesMU/9onKER1tuCXlBQ1Fr4ToC2HlIUsoOaDresbRM
mU4T6xF51qBJ1olw/zsi6wbrGKXbaKB59wIU9ny4P6XuUHhGYuWxJNf+ZdYKXHqz
e5yWSNaqcav0sFaE2LuM3MVqDXsLVpzpUqVeE1jjEIDL00laX+Ukp1zqi5j+DSmq
Ny3BT6jMtUeuaDpHMavqw/yx4ckDOjivj/pmfQjqCeAdpA7TDdHbEBpY9AsUuGpj
7k42tlr6oE4rPsldtoh+2tt+sNv2pFimkrb8xW4Uu5kbSbldtZTWer006dtPUPCB
gecpU57Z/CXlaqI9ns6RcPwJm0FlHs0xouiV+J7gXRV/7I9d91FOF/JIU8drJYNU
WxQSTHzIOmx8j4m44g/F0mHVA3sgSPS5jdTl3HRjGNpz1+S2g29Dcw6CsSIqIT3/
sWN/QAVXUfghyfzJtckq1Tk5FrdEmz5oLFPWEDd5FLniwu8vUrdvyL2Uo8oChnJ6
l8uXGIjD+/CMKO1+hdHCYzIpA9nnOPm87fzx4w02JOKfVYOTmrzLO/bmsm00moj0
5nzZPzPgdp2I5W/P4QpMpCPUpAWRts9G5TQoKQMX1b8n1ot4XK+NS9Hqub3mGrac
QOna5PN0rOqnHszpiDSLHRY87J3lIxcEShJ3jF/LuqbC94DDNW1lJ2iTniJU2zpB
lG2ACOuvz3nmPlsmIg3vftQrDzJl7J3bDhbnxIKRgYnT/1efg6ycjTD5aU0XDF+J
NQ6mduVi9VLFnQwXGFZ9w5RN3mgitEaNX+doJitRX6H8+cKTr/cpt2WZHjx+rE5T
jxIFPHMpl4r8v+Yo66DWKZx5gPGKlFsUebUwUJ5kh9HyYcydBwfzN9kd4v5GQfPL
O9O2qxTjJ35C6LOF+mTP7OQ4t1vdyLTVd2Xb453ASysb5Lbs4+N6ZPgiG3zUZ97t
Ak6IK8vnFLajef0GzpZb7ZCPAX/B0mM1x5VupXy1oSzTO7+8MIWG+fxZPufINHho
PeRT77VPAnHXcS7WOGYtQk0o0Lsdv58OBKLXbT5zXgeyMOOHnNaBfztRp/Zg2cL4
K0I82vNal4Jnm0ZqU998l/Emnwh/Fhw89+NoBAy3n+kni6Yg0Hb5ELHxZNpBijfs
AT/aEHZLS9E+zIZzO0vmYmOw0eYTqyIfw/XfsnJOuzAjdWwvZyFW/Jgx90PmQ5x0
2EGe1uHEMHArOd9EYGdb2Ayrd8osNfmLBJ5HVDE5bl3YOmP8K6ArAeWr4YZA/08Y
6faftlQafxZx3nAbzFHqKVVfJHse4iR/CkAbMJFooJ+1zkHWrIYtoSeH3sh7ZGst
oIgQRf/JqBVia4tvVq0wfFnDtIuSai+OKBUthz+OR5udPFE7dfjSYdkIJ2iFIFoL
7PekYsTHCvqYSbjFVJNgFehj2svFcTjGISlOLT94dWTwoNEPSXk5myxd4d4zcnZ4
ct0prrguZMB3XKw7KfnK8OJWBzbT8vlLn3Ya63JGjkP0RaIblxHuhis2Q9ODYOMK
wfrMO1gyYXybKxAOciapiGqShlNv1+O8YbJo8kSrjUKMHn6hU37NXYsKU+idvACm
UEYk5KZs7OO3gLBefXkgvsple6pHHJ+GhqdhG+HcuVUDGUvsA0IE2oWAMWhsJCdG
czZLwekgLQb8tWDcEeJW/RNWyoc6yCcOg9MEUWZDCYDv/DBNDMaVfHwtLy4G9FZK
u9tpLt6qPn6Lp+mgOsK5DMhWPJtOfckZmjY80+qGr9DIs6u2Vkf5nw9kUUJ3PA1M
yBuIhFzO/EiTSy4pNt/S94zjeXh3wkENXFwsQvsCD8PLs/8+bVJEvMFASxL52sBz
SpsOzCH24n4txEVsJ6WhPlu2fqAo79iGuWkvwwfuI+WUgYmTpIgGieapCyKo8B9S
Xee+sO0rTbxIT9Hrsm7UxR4oP6Wrk+rFKS/olyDbutAeIvaSmolBWSP7SQfyY4NP
I05LiHLZ+7J+nGg2mRLISFeV6hDbbiu8HL+7iqXBFnYdoz72NRvEHpn8adVptP5m
HC7akQABM/W6yIza6c0fWVT8tFmLjZwHh2NaJ/ZTr/tmxFg0fTvV3AI3J6UTjyMc
ENK99gmvsmOapq5QauczKRRMsXZbLJsjVQ17tnB4/aa8LYYP3kJFcMB/dzViJDdO
dxijHuJY5haXuwM70GeRJhopx4f1uJYAcZogeC0qatKfg5YsDo6iFd1bDF7ELEo6
it/GL1v970DJpbxaiIHzxM+8rO3obwDYWNFxfx0SSmEG1vwUHewfqROaGBrpyQsa
KsQI2eFUNhym9ZWjRbvWiLUPGPWJgXRqqAHH+yWTUL0xLvihfyJvQF3ujgga9WAt
HUHz4yXiKjAurAgkXeONl+9qawuA4WLZATVZ+nbyCQudZyrfIDmbVUSmC88Xz3DN
Rs8K58CZ/7XIbB8VbWsPoDph3j4KmrHppfQUjtNkv73b3JwsuugdeVOzNndv30aB
Q+PKNYcIMdkTG7GS0V41vCQCRKHXKW6CkwLpykrB9sqrN+T99AAW5RS+PxDGaXMk
0CnQ6ZHhZdWj1/+FI5628Bc4pFM79ZXt6EOUAKNkjL2ERC7WmlpsRCxSOT/Fr8Uu
F3nMIsq9QiHrk5Y2ruNUaMR36aXbhH1yQ1gdV7bpOKS85vI5vv7qEtzfPsXsOTNf
hW4lKXr9MXuNBJ0A93HOJ6oEDjiYCTSjTF4yZ19bYkr4JtlSycRdv3bmNxiEnpnY
XsRlDq7gTjega625Op8rXjUI8IcBrW/1XIHYj6Z2YtLY3e5ntUOTocVUpJUwOr+M
N6GNeR0eayj5EDZWMXXuDB/tdqWsDA+IZgdDK+jeRs2GSPmzSM0BXmccDJU+KpLO
TkVan60UhQ6Ols9befieWuKRu82xMDNf9THTikX8jSp1xtFLtIsUIZ1jCvrppvCV
uo2OpzRmaajBLRWfd2YXPhJKMdRI8y8Cv+l+mKLNudEKfGT8Sd29PLZs6U2GGkVi
bnwMXfRCUJOZbL5Bm+J1Aml855fz+k3a8TzDj6FWimfFTfit9pgfx3DCsfdcLWP1
YhyiT7MKsynSfjiNh8gJNibyBrR532m6t/QdfqnND21npFestKARWrRj/vSt6dzt
a04yaM55LhCQluspZ76Jx3Up7QGOySUoYuf0mb30AbGfV4dtXv8e8NI3gBDdNziw
NuAG1hzeZIjSwrBF7dJP+gQFQI7ZV+AwYd1ac7c8z3lgBei85vRRPWzwWJCfwAIO
AudzFLj1BXcYEPtnctY+P8EgiuD/jN9IZatnU/S3DurlbXSfNU3c9RZlUuXwMDne
zv3i70bVtkOyoZvlzIWsUdvhJ3Y5uDlZ8S8dVZ334YfjpLIAVW7UpJRsUTaT9iE3
xKXyCaF1pjNGXwevNBnqqrcUURQ9aLfpmL48zuiuRZiIoN4f8Pn28T9LKSrgPHkT
iusxJNaMh0cpl9u/Ny+V2rZPeYTegM2cmpa0xerh81nygF9dr0Cc/uTKKlxrsc9f
3XvZsHacq+R3RgjhU+m3syFM3C54D+N6a2HWYv8nzmBa+Hd7/JoNQcKIAEys92Xw
swyOGmCOggmdas1cU4qPoKqt6Abc8l0flMh2bMmurBhDDN2Agkye6mKPxiiVgAA3
tBh9P4p+n1/p1PG0fxCwyLN0wTDwzWynEZhaaQB1AJhzX3QDpA/WMqoIlD2ZMrg1
JVLGgezsLc/ZZpCj5swnEDF3jKpsTNfbjR8HT8d3FpUnGiqQQpS4dIWerp2TY17e
eY40a8yyJ+/5XDygs2J6bnqeIv1PF2mvltGGGRG7xKQu3n/CZXpWpRl9Dg6RHshe
YP5gQe89OhilLpcjTr9ueJzwP/3xd+uxbR9+BXv9fXOQceNjHdmu7r/+qjB1r33T
KDnI2bj4edY5tummCjQQpUKTfdaVTNjWRMJbpXBVd+VlZzuuqADcHZGO98P228x2
iAiAXaGRvcBBxGuNSOlVUPzKKLqLR0uzVfB5f/etZlf6Du6N7InXO6WFNVpHyPPA
KYQnlrq63B0YwyosIANzllSKl13Uzvn0v8O2h9+cvvu/ajEbUpBNs7is0k3E6Qm+
+9l/Wtk9M4JlKfrBlj4RKHE7I15yQnHXjtB9gLt6UwEONJ9+g4/0PEMDG76aM4ww
G6NUXzKNKTwq44/xxxqswaahPLOZWn7ZZBXFqMAwfAR3kwZHu1TxxJKX2br/rlbb
k0T4F62xwW9e4WhDMg1XJcdpwzK4dwwAF67ziN9E5b4Bq5xEmFXU5/nrKTQJwn8W
EhoHFWqQKM/Xu1LB/0VWWHfWnVdLNjU9dSS/LizCy31GIZgpXNu5/Qj10cLRJg0X
xGF8oS5SXiPa3h52c7IurjkcX5MfCqhHQcMmf4YgScEwK7H4dM1MQYYKvcYs4Uss
gKLu92XUmWoqXMWzEUXsPCvo6kLPc7EbioBlvZ/YNBKKiNgNC/ImRtzvGvwcGtvW
+DU6YYITrGnoqaBP5NkQmi1mp0lqg6B1HhgtJtVb/OCpmhlbERJZmtTrtLsAo2g1
V3JJO+nwhX/rwZGvlyFDJ087taOHavPYe+WsBOq6l/wBUSBvoVX1UWXFUXnPD5Hu
V8XEewU9KWBms6+msuhXGqEPd2FqO+NO2W9It3KY8mLh/RATehZ0lhhz7hRSBjId
33ehx5JwscJSy5H4+GYkf3TvAi6rh/oTIY8pEtwD/7lIVOOO+BVEtq4lwKOM97c2
mCokjyecQLubE8xh8I2g3M5y3sZ2o1FTtzWxnhZLjly+F4CoKZo35tuQN5cYqrCW
Z7us68bVAn7+gYvWxkeH8FyRto7WBTyGcjRsixoos3LKxjH9tWxuRgWfgufJGZRp
iKi27RAYDHcCSZf/jl/GuYLm2rmjsCcgn6FvHRgPQ3gKk6hEuLTpt74Y72ZSFq8c
2ztCdVw9hJD6Ni8dxK35kkzm1GlXTqblzPR3hPyo4ySgbZeeqtkZAtqxiigWi7SL
PPlYvELU38hhVotZXZKBMMY1uTBLGydr5PC2Y1PcjDdzudRM759hruYzyFshmrLM
5AOutw/i1KKiL3LM6BFqq0vsj6ODzcSs7VcEnuEekXwmPnjM/imIWB3nIg+BCXA5
WSn/qoFdeIrmyAHT4hRGUP4CP2RLgQpWyPivXcm9IKzQolXO8IJZpAd9QkzsGNDP
lpsdroBapUS2rOVgdB19kA2aV+LgJOeZ1eUyRVFFVCaSCVZD9NOZd7sBF3RyJJY8
4agAimAf8Llc7iAFKbKinC3i6jlZLrQGBq6fonayaUlDvVKvkHOw88HmmHyU+Pp7
NmFIZRSlv5qVnF2CHumvEMujGm2sAekzBuYEcHTEKHzCP+lnde2tdmOhR0wBBJ7B
RrMmFyH2ToV3QamdxGl4xLVAnbP7A0KB8Uqt3SGr/8Er2deZGQW3XwEaByPo+aL/
0QcuBAN4gqUAa5DY2glGJqGZ+tLSTRC9R5eic8JpXY/NE4N8ITK+se0hUShQS6eR
3Tln1Vq21mKrHCmoZcqwyF01NzbWDfcASdvgLQW0eoueF+qauwMfbllJEraBM1aZ
OOmD+5Mae9BnQp1y9bRORiiiMFYX8Bmi2/V3ImtQGZJ3/I+uqXENERkcYtQ8pZQa
keVs8C4azqszFLBPmn21Kd/XplPgFjFX3kpUJ4itEqkDxRiThX5u6gMkTtDDiA1m
VUBzrN1KOHs8cX+Ax7eDrqddeW+SsBPKM6aQRSyeoMVMTGqTbfEZjHV7f/nbBRrx
pZ9vn5ySc33sF1OwA+2FiRlAumNjfYqk0XEG67PtS/ZAXdgeSvekB9xhoKs+M/ok
I7S1IFbuedM41vYKcR8Mnqu2B8FuOXED3XwcW62S9T0905lmkVtdz1VjQ+CiO8hH
v6dUxNxudZoGi1TW1fKv2t3dQrnVdFPS8zSdQsgl533FkzDMn6kUWcP5DuWxztap
zaWNMhYELBB4yrAA/wucJNek1fN2q3Hxc+jld/m7IvIe/zxacrT7xBvgBIvnsYmq
BVcO9R+D6RH5fSr8wOyLeYo6oQ1MMcCm2C7LIb4P4xucnye7Sly95fWW5In6k/Wz
Pc0txauytiV9JAO2o1BjFxQatbK1cerizNBP2uJowaejzHUpliE87YGrlu44cYvB
mVrnhvkeUuBpsYBY7w6htrm4F5CBBq3Du06uLxZBeOPcdy4+lIxA1Lo5r1/62BKq
W6yPMQaAG4sYzjTh5xF33ywBS43EkZ0JFvClWI0MVXYnZag4qtcaCo62nCX/1bku
cx4CdSx+ezdwkH8NqkeNrZAiGxvWRyPtM3QSWi/J21d0tL83Vuw+kgeuj/GZsuMT
TMcNnxkPPk2ejg6txrVRh8ukc6/mAaBLGc52DKGxTPpYtiXTTv9vJi7+UGUUThFQ
ZTo5HzKkHd4yBiwRM9UbSMApGg4bpOErjRCCajqPsydK3ohIyAy9bycQUBIlAuRD
HorB+jR1UgEgw8TR6mOJ/RrVsoRyRREjyl+q3jmVT/hwfu9KFRzPoxF4iCAXdTQj
4pLEgR7qPFUc7z3BjkWebGw8XEeGO4B242prJpcxWOyW7VAEkJMONODlyP0MpXG0
w2WQsluEwsRka1zX96jAyc3qAEy4PftSc3YDQ61ihmASnUE2UkDHdRYOwDDPjIvG
YRrS+NTBl/4TTijMDD6GYfSGvekN8AuP9L5/7i2oYTZYFdtvBQCWTRVSO66bKhAN
0FEo9oJ0Q5UNWa+YWqbfLqMRRkWgmg8GjThPlHwu964a381/bA4jQ3croorl9Qsn
TYHMfwGDwIjI9rGhNOs0jNcNtsuncIN6isVaKZdze0wYykMD4+AuRUeIRvSJvV0J
Oj/ovUvNiFxnq8ti7G2FmdDmzBfkan3pZQyb/KckL2LfsZuKO8gN0n5vmu6Q0/MD
bbyfV4fdjSd5Lm2ho2qHK8ORi+XpuDFLj1LYWCyzeJ3lPyp7O1OBS7uWPVpqv0Ok
KeD3dI08j5QAPPHIWMfxFynNwwF2E8SQd5XIj1Kbnf4t+8GCuh8deRlU8goj6qB3
72q8tnXUv0IXLbC0ONNn3BrcA8ENgHdZnknF2KCf+UfLxGImUzVtvzRPliLHvKHy
wyDBWOxyriBwXNQsD3SAVGE4sSRA7klsiZEKTjTLSTc2bv384R3KgeUl3IM7TZaU
3ooGoAMBCZCfawTJaMCr+IscSfdPG0FcWkUeDUjAlmOKNcRbwQ3YfhzOUV7bHmY9
q7gM4z99DtfamRRsj5vckOpfAI7IDqn0xIPWFIwiT/VcZ/rMXydnHd9xDsK3IKcc
r/f8DZpaaAJ2YMpTCqoJMu/203chj61/jrYfd9nKhZmGlc+kf7MxwOk2gak0/8Vt
+dDUJiHzG9jwEMFVDAFEr3M2MyIUOsUYYpbJW926TS1xIxV1L/zJxwmltoWWtkgL
yeyq+V4+hQwHJtIOvwBXhN4wNRIU92ZMHxuSV0VEq74vDo1A9GMqefda/1DwbpFH
a5rtXWU9dGWPNuBHbT2NWlpKyWA3M2NZCttszYX2bTQrlgQKl0Wb869k+6nc0RGX
bEOWq1dFyCK+e4ad2l1DtFu7WZ5PW9/TZMssTikw+rA+eFD0pncC1neTlbriIm8f
4gQ4P15scBaTf107bhcg5vsleeR9ninsbLPyeZTlF4j6OAizxxjh8AP+5s6GcbJC
1RECaHAHaOUJuHeSrWvS5IqIQEcurZ/9H9IrQbPBXbxy24FeBW4KTT5kofocDa4i
pLGlFVzhhKvT/tJ8/BK74xfd14BUq/k6bsLNE8+Z8dTSGOOzmq4mPqGNrp6Ge1Df
HKVmHCVD1Wf6hnYhpEbWFpeHSkTRGPCCQaCCM670GaRHsSUT5fuE3ib7nrOMcNu2
xansk4603gCQP1+bnWB2ORn7O3mXmjBJl6/QFGL/LReORAtZ2pMzRR5lGa02iSxI
Ab1vBtSk0g6JxU+a1k/F+ss4J5HsHLh9pam8jVfNxbb1P9/xhPNf3sigWGtncfvq
GvR/f5LEb4QAPfwtn87B+1wHJn7GNlWtjxv+T/Y5+n4lrDr+N262z6JJD3i7Mr+v
WZ2DaZIKt6rPly8OQZetQcrqA6u6AcnFKE0dNtslbcyucMX6csYDo5waCM7/E9SK
BkD/hQtnazuL74CTRb8VbC+n4hAMnuTwmEXukHdAvp8AfciReIYNhaArqInpBQ3E
ar/R3XR9s0BDlpkzmHu9tKA92lWIcP/hqm3ZfXH2pZeVU43LB+GYPqaefi0H/YCo
nxpJOi5yy89enykdhXqXWDzKZZSKB+JXoPBnmFoy4RJtHtYMdLU4vWEAgvdG3FW2
TEU0WrlF7qwbH8iUuA6ZRiqse3OIM9iPh6XeCpXyXrW4n4z3VDl4ncCBcshtFcw7
gSWGZrT4JELNcmVD1IzFqbcu7AC1RauMzhKa7a+r9N6T7dosjuiAA5mJlyMcTTec
Iz3ff2YcUrH1I0sSGR4OwN8jPPEiOwGajx8xp9IBn+zYJyb5XYbafWq201ZhHf17
KExRGFpqnbRU2sMW3JMQOiaEUS59PNdtvXXR4I9abr2I0tvXEqJum8el28QbAOXB
Qs9vrQ3bQ6uu3p63h68F1fCGYfKxyKEdrgZ4NYFYUnrEzN2jzFWfj0A6zkwcZJ7Y
G/IriZBZ7tFY5WjKYdBNnNRVLrj9x5aIdbFCYygZb4B0VcR6wzj8XJOh05BD2sBa
tyDud8kpkinIr4p7Rp0c+oT25FvtPfcSnhPGwQenSDoTZAUXqXeYbPRz9KNtWNt7
9eavp0bvKU3UbajKk/Q2kEwefLTvdvSj4IK22lp/awQfUct6k3VJhXNcVTG29KPC
4TF6l5EpRlfrpiTvPtHfSqCJvAPJziydKi9XXttltJcHdHZj1N79TyBXVADKGo2L
6xvzmiHniZbuq8pI2LTrcT1SNud+87k4BD/VSqPeBlbXdR7JTpcC/dNGOrW4qVFd
VzxMZQQwq31vLfc1osRCf9Nfj6ZvrZun3RRQYmmirSAmV+Sx4OkRoDPRD6q3R9rd
fJKxRH4w8Qw2XwYihajvLCghaRzrm35MHHFuqrad7TEjUG3qJ7CFY22GSEYbTKmv
4iSCads6aReOicbdgvuz/xuBYIokkc4Y542cB+PfNvhTE6/XObtT/KoRo2r4PsS1
+/qU3oYl2pM70lTY7dj0s91IjlKgij86Ac3L6cgRBxORr4AptZ8vSS8CIPz4Tjxt
iS5pZcHQdQvQVPEJLVyCDRaR4PEIR7nphSj8kI8oNvWoxW+xO2+qq9ydrsAVYk6+
SlRdGdJLWQbrBMAhUFabCjribqfgkTcbwi1+pGuvi1L/e7AzN3AIhgKjmOd22olr
lA1LLQyhAOLVqSXFoPVZlRvgRIVFwaNM027ninlt76d/MvJndqoQlJ0nOePzjYu3
YBOGCmjPxQejEvVl2bM02TkFVq5gdzPgXUc83+J9uzLfEelZadKc0nl4fcEK1wwx
eFEo6QlVFTJqEdmcWY5ReE71VcKtbwOEy5mDSisLJ86JV4swqs811SaA3P9dEYj8
kBGr/kN4gRZQoo3dLvypPFM4MRhwWeK/4IpUdiWSopLisM/yKDGeFaeS967o1E9Y
wwXBEzoF3Q3d/fKDFKcvF9t81MFziyWQjgDqWUY2TlBuksGVnSVwcuZGxHpowzOI
0Fj8DUJJqycnlH9IMPALKGNkleeiFxJQnFCWBozabcfVXDq2w339nCxtZOz6eJ10
Z9+IwsRtjOyOX8mBHTPmXebvq1CMAQ6n2dUdLZWwuUiSOXloDsIXUjYx1/z14Tls
71FmxIVTvPfr1qktlmn4ednKEA1my+koWBKdd96V2dCeDSuOjy2H/hcKFOFiTJM6
UY0iqhfVq9oxhD1uLyWX3BwfTkj9jgLhzQHN2fErA33JftfVMGa/eJscBAY6pAvf
RNEovlvreL2JHD4wmO8+Z8IjeAUOGLbzl0jYVAIR1mIvrpEHNU33X7/2G+Vs7wbz
Z1FedHRHAQRJqO4JGoMOIS8TRqjVYKoj+26eDke5c24ueggVF2ognL0bU/lsxOQq
ycM6d0RBM4y1bcKbJe7mRtFHpms6YoM0kqNx3K8O7Y4YhBv8ApgJ35bcoquXWjt9
aueR8zh/YQP64LiyJspZLjPYIIQYmHsDAoMJxaEH69t0/INQj9igU9ps9IJemSkq
ndvmhH1tFLJ7Wp2GPmiwot32AyGOPEkAH5hxLMOclEtiC5xKONs68WfbTnPzaVxg
UBJzqh4J68HuLa6Y7C1G5o60cySTNWMIcYSkvOuQBwhGA6Bw4g7dC42RUYfJJ8ub
bdHgNe7sOJlQC7MTl1u7Gt3UhXQT6od7+SIAAqPYYwqhSUyKRNo7hnTHoeNW9lIl
o0zJf9uKZrsQy77jHAb8GxwIkbtewekq/37kZKBOrlNETENOWPMogQYBHxepyV6p
Y1xGuhhm3yHG0Wvg06ru/xBtstAb7GtCtHeP2YyVabJydzhJCvHt+QENRGzoa5Cc
Yc1eHskAmU/wGbp9kXS68L5Qfq2N1HN/Iip5/x+6Zdr/zu4vnfqk15s2evkVCsvN
m4X0z2RxpNGYywm0Ov2UeMTSr1ackVoS6qLDU19WeCUYkkajkH0L4sW1LcQiTmZs
dNEMXOa27k9N7VXGoQOs1QfYx4JrKhDd6Zfpjyo7bJ4NxGO5nWq4Ugi/hKSJLSm8
jEJrzea2e4/UEDKhS4bcqrajTJNjm35Xe4qs05WPexLgL47ew5vCrOAlhYSN/Wo0
2GPEz+1K+axschbAJWayuB3F4NRfu/jF1prFMy/8DuZLQ4vBVWSKm3Vt54TlfKSr
zLeBAWzVuXqMijagJkhpyX0yW+2ZBIBE4qXf9KahtExS6Geo4Rj7xMpE8tuLnXio
p4ybfi7UrN0ikFKQFyOjv3xhfS7GVkO6a1qh6pSVug5mHG2It6xFu31cNipx3jFu
gqpkZWM3jEzuAvAXK9IJvlPPY0ofNmprnR5euk2RIvzbd5DX9sbugzHUbewKR1Pp
ghCFsXzkc+5irXj1oOeZ6SdQMU8DoE3uxuNGqKNN1V4vuJydiwBUg17iQHNKE+Us
N7aFNMhNk9ADuOFEyYNmSyEO+zCeeJ+ppk4BR0xxq/STthY0D22SKXhFoVY1yzqp
R5DjLtINw0oybalL+ioGxMLnahyMSW36Ld7ZI/riqqXNPzwk1LLn571xjPQU3oBP
E7iJ9rLeA6vjiY9w8BxkmwtsJMER6hEADTUbEUKRKyYfa+mb0uxwv8IiF2aWWD8a
1ilV+dBip+WXaXtmOup1dIdhz+I9ulw1UK+7YwETS81rFYnOszt6hLjtFu04bXvm
0L+5GUYAgU3m1PabINoEsxcgA+dKnFvOGHthrFbiv5iX8YwudpeeduP6BazSvQ0d
raHoO9Ou4rFNRSD03IdJuIEQLsT+5uZ6YxBGU5dBgl0SDm/MftVYRVgFXrq4gmvv
uFHI6ejkh+HvxeZgP1GjfOGmjUruGbx+akxHt9vj1+ihKYF6+weeaF4YtwgkugHn
JhAlFuodiNapMGXVJWjN9qJvmC8Y2xLJbvNPj8Hp7Vg7JwNDnnW5p9HdK230skYx
YY8ozeYZCBY3ZxZJ9Z4rmCb6giyd5UaQC5JnPr2j9HxJbqj2bSa+Pgk5EU2xFt3l
pkxlLz99kaxGpUPcVybbKyzvMpOzU8XT10YmknVVK9Y+o2gP9prqskZcalBHv3Bo
BsVjMxGVXYdB5BnThTo1Gd63DZ89Vog5qIyb3fK/gTxmeXzkXPf9yHjcCfjwFHoj
o6xA0FqgFJWTSm7PQZZUh3Pj1QlUfl+8NbXudLypW2LXFkxuehH8ZKiPI1hPVPq7
gE6Mt7PAen52cdf1qj2RLsKqyx5U0lonxvcBvUGKhtAxP6oBoUrfMAPyBBbgYyK2
fcr7pQHMBuA77ZDaZQAWy5v+XsojbkmfYTouulvMfJoIc2ZDDHzxSHQ9iX/evSMM
t128TKA4Y6O1bUWLQTjCxHpHtrCrpFeNoHjKhH0pTvNrVlGGOBz9Hi9DZe2Oijcd
5J5IqchT9tNS4nwbTOSz/yVAW0pLFoSUUkzBXmxbyTyG2cAHUEpgvInsWCN/PnO1
XcVjzDOeKoDRX5xR9gTt+7SGkwj4UN2r7Rh6N4MjSvCFrgV5rTTNbEXxsjWatTB/
2oXYZVGR1iBhRaZFIiI6QSC91+tbpykb68sh0EMs2rIf8OmTDFW+0cjdWUd4raQf
1lFB3+APMWloXVnKeLExA1udDVja/4Va2oU/FF+z+tZDg56dCGbbNoYOvW8/khtW
+qKgw8TZrO/n6fkycp4nvI9aMffAoZd02/F+73vLpHE7f4ORyzLgor0sdjuVplrX
iVm72v0MmCGyUkK9CnoESJCHcDskbXZtGkw5jC3rHRIieIId+9CXICL9l25XO+gW
bCbdIMoRXkNHRmQ5muXj5hOUpuTvqMBLVxr17mPgvVvY0hXFAEfKVeEIaQWuKvjh
e+bZvLb3DzN7WPh+OUXk4paNRIdqHB/oxvt/3UcxZ+fEZGe1GrdM51toivVQvoXi
JzJSKFbNcZq/mOYTJELGnyIDDFnJdtJuMcZYUBOwv8e39n2FG4rMJJ6FUXjrYEm6
7G6dTFztBCj5vw8ASiixTpM2hFrd2nQ1NzmGbWSX0Uo7paJO9sh8nd5m5WpMW3X0
7b5jkUBzcjhv+TqswHkHkdBRORtimVzLSF9p6BiZmmOroVUNp81FM0jhBhjW9jj1
tPiv8AAgBuFLMmu0cVDnE5Vw+K/hvg4F6Wah00SsmlOXzC3/czDxajgOFXxm28uh
lgfa7wqo3RYslMWZsJ055XPHq5IvfG96KIXsnut6RS8VYEqAo1Vtk3n2DFMCz/WU
lKu4SBTdpIonR9W4CcJuXIAv07LvSI8Hvw+FzSIwO8GxobCq3QpcUPt+JRZUN0pF
NC3DkSuxuJxwKkOmhoG+r3AnHf1Cq/cUowqXRnir+8VChOTrFYfQXpLmDYpoNQTf
X5NtGvTZIB9zGxfFJtyr1dDi53caN1HbxrSUUyjLXMKy3X2clPJY3ZpY1Jl0ZajD
Yb4bqA/uKMk9QBiK8Nb/t4MnriWTQlWrKc0GwIv6KECysB1ggWoSUP8+Ecog38Wf
D9OZkN3u6wEZriVl8LwZmJfXfBMNiz0GD4whiqO+IW8NORsULdH36JqsGTqmr94n
AYi0i1T8Q1GBtG2ixNimxJdc7gbpqbDFqVn1hjlGsr7zzPgECMf1JDTnDGmG7vJ5
x90+275D/OvtII4GKOAeGerrYhRqCHW5Jr8QThLq3NB9Uxd3CHGYlubfNetSvEzo
97BckwbIa5RcIerr0CeZCQzY9osZhc7LSbsqjib5ACl++oxwmlNl0UKnhoOshEJy
/84pytz0QiWX8hOTCXDp35uLrDtrXJwcJUVUp47Zzy+oPSg/Nv6mF1QrQQwJ3hZq
mLMw+strIx96c5bd0qxUKsD779qPCGdDgZ8RTWHJWMyJpdO45fP5SulJ3jhyMs+O
EAh+5FWCamULo1ISpRroTpHcupfMxX6kDtHu68os4K97rWWk1MsOFi5e7shTIqVP
XZ81pw9U4vDwcus2pIXCBnz9FcwoJfvcyXf9rL5vF3G2fYCJ9DfyomI3nVzlmBlO
et8kxeMIMjiY9llmAIfxkrcQS4VEQ5/CFi4av7utPkSWqafQXeotqqzkXTf+vLts
5CCA4wtAn7ifN2gKqMFEi7H9/2DF/mXFbWeYw9A72WoZj6heThag1bUcNkrE7/bO
BNRRda5c23YBVN7jXbdx8A/XphLK9BILYF9C/fclAC4ZRyk3kF6Dx/luxdDYR/B6
pZ4gSSApOz2qGHeFCHPJTDV8FmYrhoTQ67PDsmnNEYnB8AT2RE3Bxi5EJFexU6qq
Ae+zgAL9QnveVu/xt8HKlJteEtJohgJ+SOWR0dNjrb2HD+fQRYp9Ox4dov4wr+8J
+LiH7j3TQeAEdDAjMGDSS1q9e7ehZNjARr2R9wl78mz7v9iH9wzFeG9VsTzfjMJk
o0XXign4oBZCSMc+wkBQUwNpip0xUkz6cmdew8qmCJRtGQVu7or/MYyeGQmQ4ytH
fuFEmAaqtr6/P2J38Y+tosj1Kdmm7ohTCEuOEVX6gmVmdlUVi+L82d/TEQrjYH0W
pu4xu2NiBzxKIGtYjo6dx6E6HDPYJUQWMzTYOWnKM4BLsKFUb/HpPIq9N+zauEHn
eh/VrFxYyBTMbQjf6waJk54DACWUrWhWFwhuaLTPNzFmIUAMDqhGPqd8OmZBjvi6
xuWG576gWryX7cpGoBbfH6D9mdrpn90i1zjvCjfaPadVJSgfIE4Dny1wMThOQ0mU
pdl6RIRpiGkWobxopTFuLRzYFS8nycEKRoJL+8hWTTbE5i5tEmDLaqpEeSPgc/dO
GmqbILx9DbfDzmVaY/a4o23fwPY1HYMSg0dmZwDxsMO+FMzgRhNc39Ihz+Bb1pAA
1dRxDnszRJKSMz6IUqP83A12kWgBRpAK13+bNwWR38TmD/solVj1zjkJE+YGQd/M
XayYPDhYGevVvXqc6RCIwRwGFn4rhMj6Z6ndPjdAvWoyLCXVFgd1nDEfHNYvc0Dq
9HSq0k2t5jg8Ghi0YFMXihM5S+80XPbWHCxAPRbyfbgFP+jxjtS6pzqzSb9WGJ7i
xYIKLydb1dny6jAshfi4DgJqLIXCzd85/FgR3Aijr3PC3EmzoLQeXkZj6xB0ViS0
lZoToYPogKGZEmR1RN+hXfu7l5ZceChM+fBdyATFpXU/qA6wgxKfNoIoXuu6vO2w
oXa3TInoldsP3/uXqbM6h7WIN4WO0cQd7Z1BIkoxo4yKJJXwr+VWNRLi9RSmDaZE
qkvgVshVJnKDqB69CtW6nrNUffXZcjhlwmmsEcUYIrK2KWq97VHvOToQYFSRCFnV
nye1K5fe432aaDC0I78AtmRgUI4jPk8FbCiEdTpAb3U6X02eRE2WLTTC+95YKwfb
KXol6ppKFGcSYqF6LdwSPN2+dBBz+Vy04gj98FBa+aKbx1W3LVEP96yCC36IRPtn
PG2Y58nGTVPA1rdSyE3NQ8Zyg+6mUdb4zxPpQAcOz4OpuyfRMahyjLQoJnVUlAm6
F+EC7OHNUCcWfsWBxnIB0fjky4fkiMVuiDrVgkGMuPM2b3C8mQ4MGTO9aVUGiEqQ
AtYxoAMAQAZgbYTe+kdRBREZaoiwrSI+Z3oz7TjG4XuPB19hUBqa23bT1zrx3b2W
i0+f4T+5Ujo5DNbgKThaRx/eQFPO7OzrW4ro6iH8/EqZbfOh87/PGE7m0cEPwFJp
nRJa7ktYtOM4nwn64/2BmW0Mmt+IvSn2xugmeJZuUcvhOEW1/Y8u7wUzCjYUK7HW
eCaqz0J8s5sTzehMjnpY9yE29O8bj4Otw1nDWRgsE0sGAHqxGGAHeAIzCM69z27T
2BRrtSNDF0lQx+rtZnzohqjbinrbdNKqxdVM5MnHT0/Rtu2Za9b6Tc9lozemdlfa
S0hUayvwpQIPjLYZaNqQSz97ki/wiGhXKi9chnPLDhlwKfDuhJlTg7y5/kbqMaSy
m5+e8Bl/HlCvrUL3tE2jmbZ553SsBiX2ytdxJ2UDRkj7u9mQGIh9eVE0M1D2VUEA
eOWtoYn61GuqLToonx8bGRxOhPxzVcCpKKAFIRNEpwFUi1ufqi78E+qtos3dw+LC
uAMOBo0neQPZH56yxy8woMv2pOe148hC0FIVhw5TYeRQ82McoQYXWp0AwhLOVxvl
N50KLAypi1+Lwy8jQKIU6/c3QKrdTzV1bdA8xbEh6C84KrT9odkWsByqGfxonBOi
5EGC07QpcAZ3oB392pAc3v94ifNhpMsvnDo/z9AyCYQ/aStwMTx+ZsZbXpW/u1jN
16ogbtNQlfQ28AKyzaBZPp/4y2ResjJ5xtZ2s1JWsIxVqmDIrK8UvGbeMdMXLKdW
ghA4S9Bi1sGSOQgYblQADOYXtKX8UeoLINTE3LfusrLxoDoNPYBc+8/VZvXLSQbx
5e5rRHgVqL+Ooom70vhJbJzD6z+KSIXks5pm+02ahj8InUsG111c2nZiRqxCiTOK
hD1npIiajp3633THcmOwF+ZhYAnj19EJ+sp4ZINjQYxcBcLEYb8vWIa6xRhtfXAU
557rDeZqVfJBZ6z4n4mlKm9FhdoBj8k5FUVZsymWGgmsKQ+bg8r2+pTCt1+7ribW
iLrInuYGxHyibQKLxKbvWBeUk1lJxVhT1ftPPiq+iBhAr/ppQwN1orRu+jqVDJSO
WuTaJATyjmYAtKrkMZUIdwh+2zj5DQQazaxHydWNAxBxwaWNG+ctqNfhbHguS64t
HmUr3dNWkXkbof7HX6utE0CcxGGWlT0kbJTwrv4JsQnG4cnkF3dw0p6BJ2Dz6BtA
QJqiCvzDwKUmoTUkRxfrtEvSafnHR7rjL7j4zQ7Np0t7Yp9uYkD8JEuR6Sn/3dba
duOf0+98vhihcuvlvfYBTM7+6nF93yhds8/e2HZIrvMYR5NjUxN4yDQStzbz4p+B
jkL7abH1xK7CdrB8YWIv2tvpzEMY9C4/6FUvCEaGR0SZkqF1NyyJClrjV8MBa3pN
8/3kztxL8fsIVO7Of2at/9qkCXiSQZq/GFPeWH1v18uTsZZUZ+AhgJsD6yezZ1mN
qKogLx3if3VST3ZXMKutHVcCJp2bLhvRhh1WT/lpQViUxgI4zXg+ZMRN7cw61Mot
lFG1VZaWhvT7LeuCBKVnd1OPI3Xjg7v0W/hJGBYhmBW6SK9dtQrg7jMfbT5VxGrS
JIr5v+uRVCQpamBK467iy4WRt6JklIBXW2H3VzBTWc1JXvdyA1K7sesh8/iKGZCi
0ksXHupSB0n7BsDc74YhmsCb3GFsSmsXGB7zXfufC69BTIYOTECiXXw171HVDz4p
T5FclEg1RRe/rJTU9sYS36hc8W0VTy27w8eG0l1gMInRCaddXAGh795tlcSkgOJF
DTUXLPa4k4iKqiwZP4iiCDXKZVuZfCpoRwV3+KDhcg2OWX0vSaTtsKIwARYYMXBA
7ODjrgDaeayjycuW/c6Y9XPPKUSck1hpgpqW+ck30IEO9anjnp37f56FomvDNO7h
zkKeQFTHy2uKn88LcqVCynQgZTtDLRd5PJBTHpfXCv3c11NB4G5SFdBEgju6m8R7
AZn4BeLSEg7Npckt057FB/au81vG3yYZ4jK8ms7ZVv6T9aafTxEBsx736qmyKM+i
c6W59vbUbsInI/vfEgzqsSH8AS1qdbZi8ZlTR1rQwXNjccVVmH6dsFGnU2TS7rLW
vABVatCygrIjvlBc0SstHkZMrvW7Y3uO5WpN18MPudtjZz6awATxUCVRY5QYPsy+
u1BOTi95gH1OPErXv41UzSSPemmXp2nYdvyFFDwregK34A4ZG6t3ILF91cZD1Y+g
zUzutuhM72JTFS7mA/tGvPzBBby0eect1CvivuFMnsqX2oGQDIVI6zV6nG4AAWrH
4pLGYJJzCiuGJSDOnNmn/kQIsOjsAewB0/eKisLmVKbgsvY5heaciQib/ZhbBgCC
/ydsM63t38g1gs7mIRCXqsbTz48cAWT9b1rWJUrHhn0A/3Tk6JvwU4rKuzMoYblv
jiVuXff+xGGK/is7sdkMujKEsUZcdtm82Gf74zebYnsfpLk6+8kASkpopffAOPpu
8ExqZ6J/dOnKMNiBhwLXhULRdF4PT9PUXfdySnuMCXk9hRjPX/tCdxcubvQkuKk4
CN8qIaPPXKYCzWOa7pwFkOYaGTx/r7QZyE90d2xahKCn8Jr2yAqCT7adzfUpn8/A
e4tsYrxlUXsC4kw6lvLm8zeDG0sIRv5xX7wwDbetHlxrrHYVlOXKmE6J/467fSLv
Hw07h09C5hvxTenDAnn8zNVOii7dEAQVqMn0O5WYOzMsY4GtFn8c8/+o1qpBrfwY
x/dk6jHl0y3xHyqtOoTftn4CR5ssUraeYoGEbEWSqpO/tSHvN7oA/4XAoJB1+lFn
e8GAIzDZLcIR6cJyN92me2XVIFA9mo9KbTo6A787QMHI9zuqGT7I2xgbq8w8ntp1
ebXMyFe7+hfbr5xPfyYbjWkzztBqM2L78+hStwDycJWVPoprc0HlJZHtviNjf4Tk
sLFS+mZG7vy8NR1W5TxirqCSqOOlpaQvanNKho/VbTjC0P+Kyfg2ujbSkACjZrjt
n94yMYdnttwCKdJQEViTwsveeTYgtH3AoHGRFgrUZEtpVLVtBEUvJJheaH694dAG
eGpboy2xy4OV3CruwbaP0J1eyYDum8TrkTYGf5P/0DPBKWCA+tuG5J4D2BhjIafV
Fk/mEpxxKO3tu6JUMBiTz1n/LXWC77coDmYFQXSWylX+oARMMjk4o4+P9KKdxfZu
leB0/w31Ghf+4xTkD0+PKfExPiSk4CkjWxdLBgSYMzzhVQahfPiPYcAm9no7PGCU
MKH4so+iZgCrIujQZSiiRE23QuUtFg0oN7Yq6hP+5voInuISc1FrV4iizkFwv+/E
GFfptYam3BeTJZSP3PxR6KUZE/vvU4R1wPfpwf11VeWxa/Am0JK8xRIJcoQot0gv
tpziRkhrqByiZkn45w+WdJ8q9676QQ3Xg5nF2CZdX0r+MWzuSSI0lV+5EeLDfv25
Rl12aat95/JSub3kTcG51RiW34Y/KAdDhafwHTfHna9V333I3X0LUVRfA9GWXnG6
NxuL04RdHdXB8tVwyHbNBPEfqYz5i0lcRnu0FQ1Wbb5rbzBPKBDNTwn701SeJ96C
TmTmG7ZXpXW3krDG3U9OnFMjGTPaoKEqbbzrY1TyfWmtNIYssPGEloYhRKxcTati
cLzgJx1UDSVv0x6B3pV1sqHrUyfGNQWC4p+Rtc/LAMMoG7fxAkkNQ4LBKWKm+BHu
YiDZgNm8EPCrSjjJqL2huDYF8ybD9yPZFDSCGV0z7Eae387nIcNlvtciU4XiNJ19
oY2Efpal058C1LZag1G8ruVEPzl2Sf3GWKt9oBQKpijuccA6X8ErqwMnwApmrE98
lUwsYEMnW4KzlWmh8blFk5K4zeNWHkDIPGSG2Te65Gn/bxMrtdtBCwKjSxXLHMgY
iqCxOC4DtHdmSbpuwKuNPxiFULwlXxfrjXA+QU31gJb/KA5ow8C4gYRhZ8TADgVH
39Clus2C81ctVBwF1hZbDvssm8eb0zDLw/WX6R/Yyy3LHkt5+yRIOWrKOpYXgCRW
/JiurbXze4fJADGPu11F0BYCwpPR5PTAYI80vlMfJFlxlukGS3Dc7D9IgIjBgj+t
hL0DQPXEDm8quQaz//8qeyKBuWNhpHTwKXt7yceiYtJH4J0SOJ5O7uQkmtRJdqAv
s4M3rDEn58SmOMCkL/oMXWdT+Igww8u6OAPYGCtuVyW6TRHUVimln5McyRt6IHsG
IaEim1gqjiCKwH6PD66Mc+GeTb/fpozxLVXUxUk2O6y0X4d3BSrOE98Rs3vu9H8t
Xdyu6LRh0j6KJAgCEm8veVQJcg3/4aj1zbpckM+iroPqtmCGdTwKW/Y82t+6sNgS
mXNNqRA2RrsMpAyVpFcsxTmpqt5Mb2TSHYWw4/pH3tOpQEAPOZYlar8FA70lYJoP
ALZSQcoAkQkgHCPJDmUjV3l8P6QrVeRhC7CIrYAoORHj1JDNxbgT0S8OWJB3CHaQ
Tk1/ELCgY8P+P4gupHs7kYMDE8Uq8JkjqCOA74oQz6u7qpcJbQQcDSr9GOT3dVn7
iFr6xi4S9JhcREBvHZfmXmxDaK1xz2oyLYqh2S/RP+H2BqcS5KhMG0LUnh5yo1ZE
UpN2kngnOx+lQ2zaT7cAdVr+Mq5xn0oDnS1/PJ2coMGQjSyDvu81om59ytsSGS1c
OjCHgaANZ9wj0w3LmzRQuyMXuXCCLn6B4H1Z25+J8mfGoq/swoUaN0TMLJuA/XFh
qLLKRxJdnheFvbuMWLVqetnjPXtGztlyq7vgFZMChlw6AmtqqJAP7pjMKZOWfhds
otAYH7hCp7m7z0yJASEvRe0UaQzLcRb1wWGhgGq6hI6b7XsrT+oVBWiNDktiRLoC
X1WGJhsSxbZ3Lxgwhr2BgnKvZBNaQwLq3w1a98FnFLzomonVhwd2YW6L17OgT7oa
a70wPKsa+R3BV6ZfFDAcyLtMyslOqXMsKXTOA/Ocj2PfCekb9junIGYgoOiT6ims
ujOCpi8E+NduqtUl901/XiJHRZdlyYXUuzHTA3znWDU/PeuAkbpHSgrMWwx5U2gi
S+Kc7sEYfpB5Jcm/vd6cONo7jLyoOgIqAsx79Ltr4H+tqDj7n0m7b5V8R6FafL+6
fD+xItoW3eApfDV9lh4DF/k58D52En6PmgyUmjCtylHnBoINDoNll2joOdNj/CBz
dB+kz5sJ4F9azbjGfuaOBy6RauW4PhCFH3l8gWhr0OIoGQj7RDdrGyXx90gT5nDM
pX32HmBDC28tnXlxDxa4uBOaS8ltWm6jXs0IzR/E8Qtz1L6dXHp+hAoRDJUCovfI
1/Cb3fHTfwrBGQJvOu+a0s2oBiPJ0YlY9KtHNScNfUyyJ7PSoaYnPkFtFQtuXTtS
sX+VVp2HyKrvy4xeRSXywq2U0LLyQlW6UWV4R73yfp75OflP57eLJcSQLqdKQqRF
AU57aXrFwZb28+PdLUXAb5dhn/IBF/PBagv3grsGKJs4/sF0YYvcr/LXV31eXyUb
gRvefDKdmTrIZwDTYTgitgpwihMvSTSAaaItjNSjBC2Rq5NVRMuYHIH1ha8uGaZb
XAJr1+/r2ik3PLTB4GqOjK/EKN/KUBY11GIx9LhiSJ4Y70W+z7bLkLNXYd6PRWiv
xisiV2e+CcBZZ0dqMEW6yTfJ/Aishz+JJ/CC3olo5Z5af0L0X/nTUvubVqBQr+LS
o4NUdNtCH2zB1SQjasjhsjh/3aGfvOo8fcykGrBTIt6XqNxA8y83mP8x6NrUEkld
ORHL5NGf3/NIZ5EwZKHa5/9znYU7/XPTDibgk2j7i/AIDUnadhODe3yjVYybC8Ho
O5D8QG5gxXWPqHS9nTgg9TwzUcLJhxyMtV+XeWn7akTXmnUbAmoA7buVhRDeJuji
tiVi0+qD22bKUDjdHjxrPTKmlBE0o3pWfuYblPxM/9p1xrhafGT27+wi/S8h/Rae
whO+irYv8qQtoJMisECLBO+yS4cG0YBz/nvhvXlqwcA/feqVaz/sSS12m7K2b3IA
syUlqIqwpjf3VneOsKQjY4DfzwbXdzlvp7lacg67ea3BVPxuGm+F8KSLzswIg3RP
pv/twag3bbtYJzB7wkUGPTRFsOWLmu1fU79J1A68rkX8UrBgFta5TYGeatZ/eXMS
FN7swc3JyXE4lYgV7vbdI19mKIqrKVdvxDO8On7k/zGFQAE1BeXPGI27g2l5KFzF
Z1i25XnfdYlKPV9RCpKL/f0HLFPkzBM1KW5A2rc1edYN3wiGbdpvJngvOAy6txqd
pXWTY7v2C9iVI5/3mvNvMh4WaX4QqYUJGyscrFF7pM4KxSa3gLzUGk0HFh/ndqJ2
tf5dNOyGd9M73rFrINTo78VWEnS5YHLIewXKMIv391+DCOqKZlsHIj/zVlfvAiMP
TQz1TkLGtUWqM0V0Q2tLBIDayhzYaIqOjGEVaAPzE2YK4atLV9xLX/5oIne/MvaZ
M0IjXQcxP8QnTfcLJYekZo4ctfg3V2fd86b7eF5zj7dB/bedAbuvaMMOroHD2j4X
szr1qHvZMFiSRFHtM4UKOpMu89M9rTiNXf2B1fVqAmqN1mdMHn0Wdtj0ZgGuVhGQ
4KxvVkRmPRvGxA7EIXpgQwiIULzao1O9FN6C7mNC5JFWezM2qrwrUcWh5BHM33EB
O6eiu/qvlLKA+fuuMgAxl2xQjes1LxJ8Iw+A8+/2NY59DBiI2zRzAEckgDUv47GC
Tb8bzFYGL1DcSqFmch6Sr6t1yITWJ/rIIuTw+TSBPhhWxyajxtZIk07ovJdyOIlC
NLuYC5JLpNUiw0L3L7PVeePN33J0iM8r5W5b0LVrjAL9ehOkc+PHMf+z21aFmaxO
2qWpsW0Ul6bcz1pjQJdC0c/hsqBQMp6kKS+BvtoMHxWz46k9A8VeZTg4YnJJhR8o
WutLhnYIzO8yhVdkJK04ElvYc86VPNnLtSaaqmVsgJxJ6/4BuF0xSn77TRE26e4H
BMS3D9MofmWZW1LG+029FUg5+WrJ3bxV/Mjyo3MJj4KHjoQXMpCkx6WskpYnh0lf
DgV4gdRb7lWc/19U+rF9RL8Vw7gU6rj6dRY0Osu9LcYGNsG86H8ms9zwxqmWvRic
FVWdWCvaOjzBf6JBwwv7pI6CnD3kQEotAliZIXAiAvxqNxcIaAjNYmgbN74FAeKx
w3RYbF51ACUXvdDW2+UdrnYpVm/a2kLro17UN8AWzWxdgNQk3xbakznX9q1ce0jY
ASyn/Ts57yGc7XUTr9aD/GPnxvhuUVavA+xPQtqnCinEuegdsnPDf3OXSgnYv3lB
vWPTTZHS08IQM03R6d0Oqu3g5dR+HCK1RQ7cwYkqI32CyhZliYYPxw4czijjOgds
4cOmQzjrQN4CV/VsvIO7t5C0w3U/lLz2GoNSzyS9RZoLnZTJh2qTEsUOQmUiJuXQ
opbOS5sHc84bAwRrkY/eUMi9jao4nwqAiXOCsArgatsntBZMDW/dFmFSHGiLsJwK
bet0z4Me3ZSgpi8QswQ74un7R4WSsBMdCHv3UrBElmT4lr+H+83I6BhvmLcCPrVf
JeXfIlfMvkvIrw8xB2YdjKofaoZet7G6tAP9dX646UKgjhdgviQeiiEhKhfc+egc
xcW2cE/X7VkHdz61Ex8jSRvpiUeL4sqPOUlRnMyieYaeQoHjlThEGd6FWd9m7jP2
wCVO8QQHsozltI05u6HqWAajYef4+eEanOJy9sds0bPbojE8AEknDtVi6NlGJ2xV
k1+Kn+PDj0+ICNQf5Q5+Jm0NCVXPcz/J1aeAQ6PmM3upT8ghbUp9IvMPpUvd/UrI
BKdwPeBcsPZsqsU5IVIkEeAokj1BwoQ3jBi1r1BL+AMZemSCIyQl680PngJ3Zjuo
gvPrisjluGQ2zmGtUGRsd+eV884bmFpwM+UJHkO6HVSyhzQlAOTea0rqPhs9OODr
moq/U2kjD4+79/EU+cHB9GPGeucUlKsj2i45SAZAzwC13pL9DKOiFMMSYtZ/uEes
xXQCBWsA7QX/jy9Gz3gSbW2xL9Np3Nk198gjWOJcaViGNBvZGMxzWf3WADmQSlPp
be9oIxAzApzJwAMiWbTpIa9gVO1YvVlVYO49WPFizptZfzTKV4SumnAJIQHL9FhZ
ICEDacWEqX2n5q/9RmdB+m/UQqMhzHA8o8SNLHoZRZ8qirJjtswFjjCMmmzuJiug
au8ZMxSbqKeonN/MVNbqXlChAujEv/VBB/k40tMEO5p6A14A2CHgW1BQ2r9jFxYW
2A4+u5prtvnNISJCXdvEV5kHho34ZEiNtZe8kRXBbAn9+vveCjqRbQ27RtS/Qi71
cMn3szggtEM+MYiqYIr+mcntcfpbhVlCjckLU5Zpw/zRm3HAfvgJiaJv5P+aOsF0
9it32k3cH71J6AK7XHdGFP0Aok6vZYWCtft2H7zrqGRbvp1O86ifYTJte4VmYTJ4
mPZnNt/8A/as3JHsLTGuXKui1l9Vio1utr4eqYyD0EmVC5KAL6xwpcv+Skt/khRs
p0Ff+8lWWSebfAu2Y19Eon9/BEd+8rwFwXL+00WaHutzhGcPPeJv0KabX4bBiVcH
T/HVjZt6nUek2FmZU1MhBv+axERnrsVF1s2ZRck/krdbYKuICtzCqzHem3vppJKi
Nk6TdkFGUODDpvAgL3neP5iiU/jqOeBFcMPGN6W5kVbTGKOavrfu28TC1GmZ6nIG
ajZEwWm4WTpX3kzXPTGCzYYvdiNlZ0le/fPDYC14/Dm99C+/0EhTx9/adVZdfzom
RPdo7IxV1hjzggcJHL9Ity/30Dyf/cU7xPzlnB4RQnZFlRMb6iserPDZuEdsAxVE
MTmWgKZSGLLdUJxmGDEjpibL8vO88mJZMkuHrBvukrq4/CGx86XFbRRG8VeqkmBx
JRPEyBSavDmfQLIXD+6kTHLLjU5hQu3CbJlUoM6DAhdC2MEIfFgwEp+1cZ/6tIOD
g2klYlXZS9f27MftjH0il0tFUuJ374BeWQmVPs174hJTexgttNg7LV5mr4evbFP4
0fcIeGfTaQ0g/aa1IcwHMxTQjHxqvu95yB9E51vta7bnQMfEdyJpjV+6fEQiq1Gm
PcbzJuuiEcSKrkwYrzCfV1UiLtDJU2/I69n+6c9h192q1mAjDbzCCmr1U88l6Cr+
6slQ7kSF+AveqlT+BnOjCciLbm+kSdCU/CaDWdvc6lv8nLf4L91VsrctLyey1v9r
MJ6MYhVQsP5O3Z/K4VElun8NTYzAsxTapM0sQEOOe9KTklYJnRK3hQvpLqTF/kXR
RKJfdPiM+CJO1auBmqfv3SGZcyYx7fJVJPSpoGct0eyiJF1xCwqdaPD05CM/HyAn
Sy/OF4a144MKBKacRlKGtTHhu1cMQKCFdEqyTszXjsjWIATejblfQ2h/M4tenrJo
gSI9utYjyC6fmSx+Ap7VkG4TiZJvs2SUou+gu/PefCb1fSl+dyzJYrS07RHOZcoe
3TlHJplhljJzK0jXBDo82O47GIPHpo0oU5gK1FNFCQFEy04CQsAdQL8sDGHMI2Qk
iFGDyVnXrvk096S2fZE/238MiCS1GsndoJUivyGVDGS0OyPjuSguxXHMPlpoITlX
lClaSe4yQfxbcWmf/vRlxocJ5Jew2qs9xrDPAxGK/zV+PuKx24Rt4Nd6rciYZrVq
zqN3cWtYS91KcNnFL01yLIdLQdg6TwiCXi2zvjHJUrtNyp4R9XEMvYxZQ4xoOJ/+
5VL1zgOYLiR0Nby1VsbaRgnBdjeKPReX2dMc43dwZ9C1dQd5qy2+RwoEiaYHuYWw
0x0N3gPWFCnndvFBoth0oxeVlFVa60IvSbJi6wTYYtYrKyxQ57ckfZfX2D3uPmev
xKEbS3v8xO4TnfOoZQoTVLiqaXGj8CIsRC77XjzI2m6H94mVAx6IPA8Fk7PCs7hj
0YFtV9ZmUHM/dSvB8tDaYuo/EFY4A3IKsNdeMGVRysXtkGARutsZBixn51FUUlI5
p144V5vOe4V3TTV6y6hQ3/ip1rEuBr5KCih+wB13Q0SkwQM7E8LSuV9rushC1DSC
42CuYG6iI7Eugb1fdE5pxxtFDko8RpDiELFPQR855wHuCCJ98lYDA6P1B5AxOXW0
soRau7AKWodm9oB8cP3Vfo31edhglWTaPXwuQlKWgqwZ5o815p1GRl4KCslKiYsh
Uap0in7EzSPj8BUl4hI2v+J06DJfXDzNjNvArDt5SNADoU0tD4gxD4vIHEyIjSZ+
E/439eqJOCKsgFwE8bsfNXfRYFW8cswmU5A/A0udi2vwowIiDuKgAMhN8SFGJLPx
84WhE64aItCcJxgnLP95X/3Y5yK/AZPiFeR66TQGcPjF9cNQYOcrd1lfkxd4efWM
bxHkmk67l5keiZX9WgQa74ZdLctXWVjqIQTsm5UkdhbXoNv5Av7jxWMG2P3us4EL
4IHdofZ30sc2iE30yqIFmdOHQwqlxBQ/rPmxR1tLIb7QYlqVLypG83yLO2uDjv1+
1ksA10cn2txegIHx47gNO/1TiSYmTJQxnldCUf+JUum4f/s4OKZrgRM4NXTG4lch
8rOpReO3VEw37gMZSOxKDN1wqxXwmK9BWHcVdA3jvF43Z1MazZs+Qju6Rfy2TKMd
Q/YH6NItJCznAUmPd3++MSU0wHKtzjDBZ13rMqjN1tmBffugsPbN2qv6fc15vX0l
LhsG+Ldf3CXtBldKIao2pe1nwsS3+wDS5ScPBZeDoOtvZexbzMWsBACWmZZnil6v
ekXotAGc9U5KpsHBw5NBtHuGUk+42Us2uzRHJqhDDK9bJWxMIqg1xecOyF3pztk5
+1g0X4a4YG7TihI4CMQGvgyZBLql23ECiDtlMstpt+ROsuAjQVmurBPuOJ4CdJho
PcUge74HPBrUzE0x5Jyd2UCE4TTDwgup0TWJTnI74e49BbM7anK6BB7NBcHPvNbZ
d0KpU6YZa+g7TBqbsYZcUAmMQ4ip2mI5Y8CyxdcPzfmasuknKXsCM7Ii7yq1No6y
ygcPGs/fFyPdiARVbHqcfIKnDzuv1UwjOj9ibPzPIIhtrkvswUmhhnECYS4pGITq
Jw52bYzm/dcrcuhzh2TY4N+PZDqm1KHFynL8obxj+0V6II6eiE5CCKSpFHEKBkhh
Gv6FsW1AkahQUP7K9J+Ood60VWgZFSBQc+B+bA1g2A5aV1rBpOawRl+pU4e2I7w7
BDTFZ/+WfokS1i1vwm/CpCMnbmkW1L68QoiH0JXMrl9Brt5u3X2r9jAYf/LQBD3V
B54fzZi9TXfhe6hkenkqTMHrRf+QPkyMK34O2diOt7ArxAu3quVMZa+DwsEnxtIx
6A1DDPonTWRLYSg9xTr0rQwNMHYRijL4JrvwjCzx5FFGmnWpna4fzf5meg97nsbU
f+ZnaUnWW9rj8LfpRtP8aqTgodUy98LK4d92OtjDk4X78HD3J7rM3Dkc9K30Xud0
d5xOnvkKHudtrRfcMZpcmrCqj1u2PwwAcwRf82KgwTbOIhUqjkJs03VimKoikvX0
mdhste7FRNDCabc0mHT7hWhbdjmmHZToCuVjRaPIIKM7wOUdSZkUJgimdqvsy0K7
7dL4wgWASR2ROj9M/UFxL3uLUUeCS12MUVkvHByfyhFpaDvpLkwYhNPHMeOe7mzN
d1NTF8XGf2IGJw8YgVJ43eHMRd2kqDIEECU/wLm8/L5emnZiEtF0JkgrnsRPKYQu
s4jDx86rh7qHr765FMONY9e+zMkygfnpm+L20xbE/LorZwviBDtGcUem2GyFxvlF
o9FCHKUSpksOmVfkp/3J6k4Wqg32iigZ2jMXkSvzu/hCPZDry6cxbwLlA7dFpK3R
NfAnwCLLeMWjYfBymkx/rEdktL8zByCGBzE1zmA3SO7P+E6lscQPiGY8VqSBw7Hq
S4ZZh3+yW9G6OHpdzgKfMsxrWF3qEMlN1ssaWG5aVXAT3CBI5itEz6AZBYrg2d3s
jgWFHPRTJ4C2grYVClVlRPfH9+QG3UxZ9x6k6Z0Cxw4qbfnvQz7emIT2yWD9qjPP
Qjy1vUD74hou7g0TLBd4g0I5v04yw6QbfD0PBg4rMRdPkYIluOXApVRsOHhxSUfh
3SLOhQ3Z5tYCGkBj+E8oZwSULDaTjNuACEw/VwycLrgVDrgX5/18jLo7J5lL2UmG
B0UU5AMzAY0POTMzdqC4j0ch92qq81wZT93qGiMsTxLLjzgmJ5FgZRvORXXIBnxs
jBjN2TZQSyK37SOtqXgYhkR4QhUz/J9dJ5JgFhsJUNbNsHeDyJ7rh0+CDJBeAKK9
n/Sv7s1dpStvhApV5XTyCI2HAArV5EEpnJqNwrjCkGB9vEKdaY2KcLXxVzbMTCeO
7Y+l38ky+Btn8FeH8MTLMGm2axWcIMx4AALafJ/5iNOuvAdq9qrgnJ/E6r3AfvRl
z48aIpeXtcF21TnlaL1G5W71NxJ4V+CMbA7fB/Uo2H/ltemzRsox/GgODkIw3JyW
3LCBnH6kF3ALfKhsw/KiLyL77Fm8AoRZDh/QcwWqiLjcsdIGZZwkEy8ZuFdsv1FM
wq12H5uR8w3MqXEF8CBOTGGLo2oX/0mX6fB8gcV1m1JmibkDntCPiHuV7Ov1lyJQ
YOOI/OOg5JTrP8HmiDu7RlOiGrqxu6GdojdY2BNSx5gn0tkRv1Z1zY4mio+q00Oz
ZyxOcOLFJ+Jcwq/wJu42dOP8MA+FqbKjQtwZYhtJf8BZNEGCnG7o8Yh/uYgIQT8O
yCBXL2W5XjcjqxBU59dKdpWEfvUh61P0sNChLZfX0m7p15fqIxti5NQAErYqcMkE
gz4LhQTFUTPB/0iQzGR5QQGIvR7yEaia1cASCqUeJdugZ+UDZnAbAc30n4FxeNrF
vTMg/ftjwErXVGpN81kZEqIrNP7bvnjfXqoiu1/eQBbCYt1qqaUD1qlzb2LStb9A
/k1rdFp/ialJ+RZ5U6wiZ8Kgz9KAQKzu0NA1ZSp/XVTyRLBpoJEu26/5ukYwDRkW
nAPle///Hc/zNKsfb+wk6l8VuIb1X+FYMRwmfjybrb8EkJEMtrtw5CI55Yt+BUo8
jRTRhmA6UjUj7nSfHwcud0HRC75mmai1rJFf7RdeYoY7GJq+etKbmEJMexzxFyg5
uM+rAriubdBbyzvW+L4V3Wh/HE8j+im1sgH4C+k6DDI+NEBLLgdKVU957Y87/7k3
jXu3FU/v02ikhnQYCklwyfak8GBDx90eaNdITpQn5Sv9prk3DgUXoScXLkAXvcNv
SRGa8aKXEGs4ZB9tFvUcCqmC/eZeHUXUdMd5j+C5xA9SzEBdJMhkcTVpwBEM7hJo
EjzmYM7akC6TLTnXBS2wyZJYHPg9bBAIimIv0fVOs+W6ILDnz4jd8m/UbYOTs8w8
rnKtbulTZqwRdMe/LDLUW8N8oUYrv4XpSyDBOUWoYjbYC+Emac/pphja/iV5FirB
CXsqNTjqbkN7PcU1K8cEukhocqq9Sr3Ns7KnKle/wFuB/g50l2addQ0gIIEeRbwW
i9RjeZGmNmSbTYj6LP14xUy4/7eNeHfNchj71WuOoZLs3a4Bapebcr3gBplhMtBz
n3DgasjeFIQmh9GRQFr0RTHeuIr6fTBJqTaDtUUEsZufrf2ZYd41NfHUpbVqCQN6
68YwyLMg0KZrYc6M5s3oA0RVJxJrOx2//s8Pm2+pAR36zd9mloHDdkLFe8tGO4T3
+ezOE+ziI8nJj0JQvhP97iFJ0z+g6dxkiDG06SMBn4jNBsWxNtxvVniJxUpk4naA
LjG2KMEGPUiftlpl1OJTl96ejtE/ZHNdRvUeCaz4KQM1UNlgz3GTquRzg688J+Ox
3JFz+K2rbaZ5wSmrUHd2Cwdn89fNOc+KDuGxL5LWJYF+NjS/fUF3ISbmCbl+I1Ux
8AtyyhiShXDr/wHOj3WAwEg5j7UYViWMZY42SyvJZ0mp9tHgzntd3tjdUZM4RqRE
4I+XaUSvP82NY6EoZV4/NnGQxCG5xinEMhUlsNcs40nIsdQ/2VVU2JND6N61qtyI
B7PzRDVoMYUloWCptrMvithd7qgbf3VnopQ5Dp2u01hDwcs4qv4RyS1OEOdkG3pY
cw3rwhkowLEPJUWhBODwhMe9UjBX+Iub3CwU2ThaNs8rMcCXEF5gbKIun0WIG4A6
QdA5UFQpUvez4Apa2BDED1rC+9Bjj3fV/qJ5Ih5BAittQQcKStoe5PDyitIKrLiV
/QIddCao908ZxALqxWO1Sv4o+cRDzV5OtAKHjWdtRVwamHLGK4cGvY8dvZWiZwhi
SE4zxalyb4ePjduPerXVKYwKUivi8yOPSZgKl7Upm+Dh7KKuiwlYCJNBTUuR2osb
XxnKbWBH/Q2Yu9yLhoPmLKmoVBnHki7rTlsEJ8jm5EKj2Qy2RSPMY0G/zPlfvH+G
Vjh2YePShdj3B7z0pQVmYJBoaxWpq03TCx51N4ysnWPfkF04tVwr513LMnZx4wdx
IGjVPEH6GAJaKrskjIozcBnJc9zrjpMtjrmvpToX+1kCu7U4b3cxOpXcsY7NmYVS
CCnCd1HiIAvhFKzC/RP0m57dlxCGrLWgrsuuFVXt/Sab87l4PWsMhZLdy9GrlXh8
4cHQccDZ/lnUCAoeO6MX1vuVyIHZdAT58Oi9Ca3KEdy03o4lo/xon9myeMc1QSSr
Y9O53kHaLFyYX8p21o3VB08jANwx2vh4Yjs7qRdLKZjKYhuZJ5Ye3edV080ujGDe
L4KN5UdyVUEIS2J+hVp1ru84TZYzlZ+dj9Ekcg5ehW7D2M1YcBDTWYMNfYbXIjtI
KBS9/xY2VpyaNegeO3z/Q/z64W5bXq4XGmq9R8Ccz9J9+VvwXZQqL5IH8kkzO050
2eoUSseijtu/irVt+h23ILtJzeJlTJcEPR2zIXvutx15brD9oGiQsqv9Phc6Ce1+
I6WwGsZLkfF8maXcNCYx6whks5ccqO06x86zd1k9cN9GblYzBucuq/6NnI1ycREJ
e9Y05/yMe/WAjEw/3ok988pleG01dA5b7O5AQ8PVpUvxEJCqpKT2NQLcAdBxx8Hc
/bQDBxFRI/7dO1eXpzb11tc4zQXFn+wWsdSx4t7oUz9zbBsM+Ypb+1yAuXxcgQue
+YJdljUq/ffUK5KojIXbuUmZwF9xaW/OHen2yQEZnK2s8dLQjYoSiAQBtu4EQp5f
oXnVFl8Yh13nl4UUZ8v9Uy6crJ62cTwWotgQMPNiQ5JRYXP7ieQ7MDzOpY6KWm2w
FacpyhLGstt6ABF3XA2BSdrJ8x7Fvl97Vv9tNEDlaL3VDrr/oCRiB7brHN96I9Bj
hzvxNnChMw1EyTT7RCB4/20H2bQ1XXMBjiKsUN4yJT2mcoAGUBGlmvvVeZpS97An
498aQ6KoUxubZDWNfufQWpBRE0mrYOH58uUQgMPUqgYEq7hVPCWYaWUEBVVNqb4P
hvonqpqjhtndQNtz5xaraKtC3AhRciq4mAuisEtXByCXDVgilwOLL1vtqGLZkmDA
axhHpq+S23Y149pYA8R02gIsnAUQJc49wHyGmNmBTfoas84qLTFUey20bJdDm0Nl
jSMq9J8Jon58iyvdLTlvoAEf8kF/G2ascnSQrl0pv2ggHwP6lwLh7Zh6Y5SV2fNK
uU2UoVxuQpLqkSVb0ScmYG4yOKUHg7dZdRQNvKnPGL7zRXMxHXa2mWygM+x6U1xE
3SHhhnZSZLz7l8NFXp0jVdBFfUF+3Q9Jh2NRYjcSoRmIt1foFxAPS6Wprn5vQtRP
pyhGIWjIBcxDHZWZM6cf/OmKAbLvdrEbQPZ1a2EzpAXWuzxKlU6/k0TJHZADRcTI
1a+xxPxCNcUhdBB0Vo+7jx+IWXHDYncr9X2eoO72i95IEQ/593JRVZPjRapl5yus
Afo7JZZEGoDadwaIeAuMfJIbmqTblhJHPefO6ZO7M1Myau2FVMrauA+M5ZSnZ6vd
nMHSqWd58/nBsF/IU/63GZ7bZTY0PLF27AD2EizAh9ZKHAiOVs5cISHX0yT3ZXxr
HBObGFxa6In0+1TiEpMt9/yevM1D7zDqIWMPI0JY3XhiUyNvOKohWk8UKjjN/j2S
iRlaJW40emF+YAK92YvF5Qe+JDPcmrWm2aEUONcByDc1P9baPI7edFRvo5p2GXXx
7U0Jjpw6GuADZkyaVz5k2+8a0gQ6G93DsIvC7QiFagsvA25nSn9XbENF6gJBf4uH
TSau/0b8tWl8dxObdZ42sjjeMfvlc8enfpGSgUKOCbHXoLH9rLjlzXszUx7FA+yH
+tk/dElN00/drYfesTplytqNmlRVqoMw3wXiXwvUZ1k8P4z8hD6TTARZxjl77BvY
XW85eGn8OlD8lzVkqTfi4Ed0rrbbLrpS5qN3kEiNSnAV90W3WRT6v8Hww5LhyB6m
F9XOwtQP7f4lQsCJsCIt4pdC8iLCMsyUjXRdHkB7mxN5aLytLqeubTitOOWBndxR
KZcwvqbr3Ap0fAk4d9WrQRJnm/1z26mnyPYUSDJ6eg4qVAxzKB0Ye7ZKAKbMmOB1
ztpvxb8YCJdCYO99nVV47UhP6rDBoWrRyN4bwOAeW4rkSgzPy299AF6UORiv9/Wo
/H8DTIMkqD+8NgzUbLjqaJdWBNYuk7xvU+yqYjO7cKOCcZmp94+qb5wJXR8AZoB4
YNu1HEcTGnVJM2kLv36Af4kpkDqUz7uNI+GAh2kWcx9SaNmBsyubgrKDgofNbTxh
rvF3BXWWzsP71q4zvCCmZ3mWuboKI66hUWUqEgyYa2H17mK/HqraMgvEXdbldqRP
m3AwwH84HVvuEFU+edDICQ2bbUizofLIae45xWyUXmxVtyBlCM3MtFUHewhzsmAw
UqtIJkvQVmrx9tPOmEEepPYBUIK/4qcU4y3A3cuVvVUIJ5FOxF6sycTTTjTpQdt+
BgnDRsAug85gySxV2/YcUpLUOBwp/tkmsPCftuzCL6WJyg0J/ZpZ+v6gtGVqXLgA
0BRoImLctU387g0jZAI44+xoxaCfVPC8UhatSk7PYQlPADxIkXT5CUYuTId1yPmm
ZuXtw4c+m1f/4vyYLP/5ZrxVOKvCfYgfM+0EfIDI6hfTPX9oy0EghAziqUih7q+4
iD5v4OuRv3iO4F5/cNBi3g4zjSlRxp8lW/2XUhwSBuh2O7r1CTpL8kX5BFm7Doh2
WXvyFs0DcjGEkd9lPfOS95RLfbTz8keg/bZXyuqkJSItMdPKFEUHrw+OD5WjuVeE
YA6PvpMfr6BkCvqOwMC9K+4lp5sCAnyjnZbRrwl125DskFuQjmFzN6Tvli7Jh2na
Ybc6vlJfvf/ZhzwKJU/dk2PBuiyFB2uXV0EqrZ/I14TzyJD23GB5CVgloLGQSWuH
QzMMRbQPAyLYq+VS7+M7HFBZ54KQ9cKmFQ0R0emSweTLAoKqr2lV0z6ptJoZfFxR
ra5vGR/WR5TkV0LV/AfMfezyROxK7vgdTGz0MYukGZ6iPjD8XqN07FNwlftfr0q0
MwXJVL0Jh/TP518BVp7xdVO2xQxihShmQjU3iKqFPBsuMD3Jvuc9F8IQyjOy9P1l
QlFLIvP03+fjlqc5gdwFsjE0Hsvqr3Zwzcf+bK3nNEECX32FfPvsAKI6sAaKLbZL
T8NnHliqUT982Nub10jKgciKhsKmBFQm3LnzU49i3waJj9GQJtd7CVp+Z7ZYF/Ge
6i+pjFyYZsvLOPI7cRbkyBxaEt5xc812KNc4tUUIfd4z5P+KhDNPWrJXZ3w4GU0b
IwFuVAJxaDE3F2t0qJNA/xU0ICwwnJLdJDeuLzB+ZEvwxa6Drb9UmAnf0vUVujLW
uEpA13Q5GbhclS+Zj4QT05qF0QSVRoFKD4qrwt8NBRAntvfdDAcX6pu4MfcuUdYb
GCyNR78gphsfH8DVNvmHRCg4C8qTkc8tPB/lJkBecnW9Mdx4xS8aUP1jn38kGTg8
95YR5/PfL75iqivLij59kkJq1JOu6CFHRBHE/nqXopONtwq89B0wv5YdcKH1ztZd
NCsoPiJ3HZ2QXXN8jmGdr+uC6gvAgW+tUte0YXrTUu//bitWLjb6x+9kH5RflYqY
AVtr9SjBneOn9ksHCW+VVmEctw1ANm80driTbEsucPQDlzGYfzooO2p6ZNU+J9k6
gEIEdv9p4oIoPYaustP4cXaC10D3Pn1l2U0e01yuqr1wWXbE/xUg3QhgmkrYBR+Z
MuNzsn4KhQWiPZe06ngnQFNDaXSaEOzo4aPqvLNQAJFsDte3NglnCKseRP38pTyT
nEccLrvaXhvsJdPbkZ8LdJI6MuelHnkxn7ACXnqRCSD+EMWjDh2pK0/z817H+Itz
PZAWmX5LJk5YEPxUXzJrmoAZYoydP3TWpkyb7d1LPLqVgfDrn4fV/a2RLrn7SPdy
upN95xhMmYXmUNRvARrwuWrd7HVIJ5LTv+kWJLIH8yIBBVyryQH+Az8UigYFo63O
8LgHPSnqL2PRifjBrQLJBjKAZ+yEnNakalxoCD2zm7ebzo2lk/PGIrJrR3HWskBC
sUZa4Zd5tChKEzLqSG+eWX62VvZKtpRCCX7Aqd0VaOFZVOyU13LIEuqZ8MFjVP7X
v6AMNhB+VzqqCF4Hxg6bzSsXupXmBwRHn7A9Nw1nn4MLnQQwldorawcU2qMP6c1K
txhwNnrT7bg4Mwel8R5r6zYCMHzAEsj3AlrZqJlQteoO+XnlOXiDoIr8aP7YJMlp
YsNZFn1bF4ZKhYTHfNCJQseNglXiEbvp1ewQY6qpwSoWSGV/zXocvhiC/gbt8Bnn
NSseujUHuK+VJ4dwP7h/PtK3CIgNTXEiCTenl1g4HB8SNX13g+TgojXqKdNMbWxD
6+36YYP/7lkEiIze8KR31jjz0jQycxFMn+hExkY9n24IX0t7T1aiMNrS7pNPgOG4
kbeLsat2guyum5rN/WhQdkUeSJDNBjSQJN8xSWiYd2X2KrTv6rRRbndUmE5jNjRA
4WunIJNlPY44faJIfK0dQ0Uw945fdv6KFYC2RYbdTVBmN7Ue34J7x07MI9N8bZBm
CRnvIp30WF5otrK6yX+ChNTfcF39Fvkxu4rTbZsuZFwE9BCVrubLjw7Qam3enREm
Uzo6fCfiA+iihoeK+MGlJA/6muMz0v8UaM6KMC+PiD0iWR1Pn1lyLmdStK8OD21y
ev8IGC6X8f9CeEIAHVEy31ruS7SQfAwN/itH83hmjkz5m5ao1sBIndDSookn+56O
1aCF47WIUFu7XNQExYop8HglgQsgnzDSCZdpfSgjSYGBSpPY/niVJ9M2BBmCwLzl
eVc3clCNCmoP7V1eWUPdmcrcZz0Bfr3zcsUF7cyORELXCtlgTvtl5xrOMmdmUl5s
AH/sioXXTtInQArcJCmuB6ypeW2sYks5D44MZJpxwQ6jtgcKLfR6gigFZzdR6DCo
USh83i7fgzGNvHhjkp11/tCbdZcsQN2vQYI0GAm9xr5IxMNjY+AMYa8xk3cd1Oc+
yaEU/d/Cmv4ji44nWHIJHfoF255dFE+CcVT+nI2TtY1elxhUfZ+CGWHSgwH7Sayo
9dXwSzxpC4MCjCQTgfjJX54uWBU3FqVjSTcEofkg6tQReeq+h90PFDrzStiZoWOa
PMaoB074iTidwN2seVD+AEKuuKPkMuqPwmVaxDfh5bo8ejBtWjHLoqd/h+YWi4az
QPGflHH3rjzL7UbwCDP20lFVlj08IAo7BEb2R2Ym7AMaGCI2TQFkW/RDDTNonGdR
gWvyOCH/l06LS8cTZHEMG2Y4ZZ5PtZmcM0m9oVARDZo4ZfDXGNrAec6frhTFdDXO
IhxPlbAPrpJY4I2On8VguZKES5J5SlyrpVN15eCpsZqYsYTuaVF4abyczqvb9oH5
Gr6TrLbcy0w2fA5btRvCkT4HkzkCxslBR9C6/Wo3vrrZ0F7Vlk/JeBMEUh35MzE+
yKwFGpeDyVpoy/vSrEcVDZcdnIccWoRhWmNp0R/NQ+mHTR9UxLz1zAZtoQHAx7Ct
cTXZU0bF+dapziKPxOm/qIuHTfj5IBabDWpR3YOU2x5cSyqowDynXnQjFQ6hjMWY
0/jontZ7ilzbQ+3M+AysoZBVImKc5Fwd2hVfxkwkMGtOLcgxexdPVvkgTXy2dUjY
A8UoVPdEMxadq7+l8NOFsSSviIgqjd9IWHP3WIHEk2/7lyG/3TgZGquim70XlKO2
oGP0X00BoRGlqWMRRuUVjL+4WdRyK0y6iTiNzXcDdkhRHfKVvBYkHQ5Y3geG/qkz
G0PrO+kDLBZYAcOa1DU38G0do8eKoX3tbeMer8xOoc4/iRMekW7r1RzgRg7J1sQV
8FzAcS+Shfn35uok0fW4+zrgWeWKsOm5usspoTm5gjXIqs3421oVHKiZ0Ov66wav
5/7CHhroAdbLRJ77D+aGtx46neTy2r0zvo5vtqbFVFBoeI3p3xQzXNx7GR32NcDC
QLTjP4a27ZfMSagjJHyhSQw+hZQlXoJBEKaoDcSImPnxuOnyqb3cjhwO4YMaf7tQ
oV7r4GM95btYrWv3b9McY/oEdcDFev36BGupE5MYkAR0K8fk0SIhNR82q5TmJmvJ
CKKAwOdEcNMRgcRFCpn7/o/Vy3/NcODCxz6zNoItd2gOkZiWLoO1zdyBYt+X3GPB
WjWHwm+nJp6ijPRT3JaUl0vlJstuFwMYJLz/naklvLMJ9YNky5iQsKpUOy9SKDd1
+Nd/ujPAZOyVFeYFYYjhOF+5ZGfw9z/XNCiTH+w5HDH8kIrpsPtlP8uiOeLJIbfz
XYKjh8VdIGpIn03prlpwC+u9ncr9HDAeKmBG0TKp51/3PQSpDRenU63E2W0jj9hV
b7bykhmcHS1A6Jk27uyTbrlPs6hjhEsf3hTAhzCES8sJm39KnBVB45lshX4jtQ4H
Je2AwxYCmxZbymC+clX1RzTep0j9p3wNcr15/lCxrLNsh35BYpvzsylhErSFZxd9
yqSqhO1cUmIuOiX/9wjXwT2eRef/u/Gtn3Fot1UGSXdWarT+0B8Ui2MECaaW+XhD
N4aPcNbWU4fsa2/DX7jiN3f+aqcu7SI4Hclf0jdCQYnsiyyuy0fm63CUw1KpAIXL
Sst9J5QuxP4afc1jaBwz7ZRZjQfeBF8q3Aa8r3bLfUfqoAFtsHedmvyCJ422p0A9
sfnO3frpeQKUnnckvlxAEA6jD3mYMV7z7vE+Xv/yQYIM27Qqpt+aL8BNS63AZqq5
pXmbqYkh/bshyOc81R+WtzY1DWBBzj9omhnSqH4/w1rOCl0IxfbxSKTSnj+TuDHN
q4cpIFblhLKLK9FK2Cwi8l7Y0jPzK5jkQRHscLhfkYxAiu76Mkns2HnqsJpiW8sH
znbNBYCtzp6N9Zf/z4J+7XaOdjMa45eyq9oXBvGQ3gj/boofI0ndrutSzE0uxk5l
nFt50uWdF2n1N3jC9mKYiWz8q+0qxWiwpes8U/oEnAsgm++YzUd5WnwIM0+ns7Ze
EPsy/oTYizRdyIk4+4J0gZlj6Un2/ZQqS7/EkaSpBTDFsyGw196z1Jz5Nh8Qa53U
pTRENdHQVqbC1lahaTKz3H/WWdqvzVC/H0DoHlM5IVIlIh2nNzMw63QPrRokOnmp
ZAdDF6ajO6lLADwxmF+tAY8phYvU+grseB7nMuY0VxkKe8x9LuSKSv2dlpv4ijqP
Fqyv+8mQnzgyRLIWjNgv/tRaRToK5ozXXPyiRpNzdGp8f5MuGvfn6bSIWPLrsrZP
dSqL5Yo33r+AgtrKshOEko75zA9C+SqdLwUOv4WfZHsCBcmhwQ2mki++wLIzG6Vw
4Q9NxgcPFWCKQjZ4QC1GXaPBRhH5IGYj/FSjwS7IIYVyEh5RnmjVdfCc0Wursr5Z
hEPgYFYaUB+tFWEpRTZjC1U6bQ3yqxglvBTSZkFh+9t1eGhPtxcT080zhzacLybQ
SiClVRjVaaRbPx53e8dpFU8AzibXWHotQ0pyczQ+9JuUG9fqDGr4SU6INPOOIayM
y1ol1YTlwnPtkaT5ICpCmDVqqcRBwUn6QM1nBg/80bEQ0cSVag7PyNBTw+y8QWd8
WEnXpRONTT7CrzNUzcqoVXR+YzW214qszRMCuePZ2PxUYdyf8iCLaYCzba9uI0DU
dk/WUQNkDV5DSy6wlvkjJazgWO+ROfH4Fgc2v8S4OZl5A5C6K6lnvbDQL2OYIplk
AU6UDDdcv/UP04CovVyoUWnFdH2uO29Yh7VeNkXsNFB8UID3QlczZAOpUnWOaQxs
I0k1nkHNWrhFXk6gHE83WVdUxrtMFWqzrRTupBPCX2xyCLx/E266H4AqwdpZSQwC
yXgzu86xVsP0QWvuzeLjhFkcSLOvh8baMHJenP9xRP8l/I2rL/5Uqfu/1r3eLDep
iZHcu6887z239k+DnfYqaVLCwEFYpL4rIG0Pf2IUeHJiz2qks3pRcbTJ+1LzpyPf
HQqY4Yk9xXvLCmE3BCA36VL/ZDkJqRa130qk8dcN7vunubS7SBxNbgNFbOOD66YC
gDEkAGb187bWDqAcTpgAFRUrOKQTCLNYSQBev61jTsX1dARLZP/ij/8F0WWeTED1
pNz38Qh3sxzDcGBidhyOPDO696wzEvHd/pUGuI9X1frGM1VaBEb96FuTNy14XN6J
FC4zU/z55o/0zHVF9cvcZM4zM4Cof2qMQxQJ0ZiMdUoxA6xOTj3KtWTQ0FPVYhsK
LVP/8GLchTRSu3yo0EexMGS0/31Jf4QVwAzvuiCxaKXMFZQhMinX3otvR8UlHdKM
2q0cyJWtzgxjWg6YC8dTWTHXnCYYBQ3qxnIPAipO6Q37KySnaBpKlP4fXiR/feX7
Py1616Xr1XB5QzKoRnDf7Vb9CGWpqgCJ2ubjZTd9vSFxyCaT/UOQFNUAdLW4/Vjc
Kjxu92m4ekY7DvF92A6LQ0TfaD4NKcH/w/unAHls6LVL8/gPApA82CxnPPEq4VR/
wuujXsJYvCQZcJmKgyIKghBAI1DRg4CCsGNqQ1ZNEu0hfVwmwsDgeadmabo9xo7P
apps+ck2HXOR8b2tgfmPK3doW93XsBS7Q+RewfEhVO3WtoaQioSAShP+4GpsX+YT
eDu0AKl8BIhw2B+c0G0SSaDAv9zn6XM31+LquBi+o8mUsMf4nmHy9/u900PRnUtg
RuN6Zo0AeateNW9RRblf2E2j+cjTdCtoO+skwJUr8i8ctZBfRcZY2HYbvM8pjLcq
bhcrBBmA9PY1tYxtweT1QhdxHv1LL65bMFNELIuMTEvjm67jQTp9BQOiJ4wW10Pj
VTD20nYCOqg4Ykqvvx5ViXlwwD+HKMq50naHe/bfmr3RLBfxQh9VxToxYHE/ShH0
AaHFDqOUgTKmWB2DBG0I+3ka5JxLJ4U+UMgNeOYQL8wcTYM0GNr7IxlqnvriSqdR
bAZVEORosDY20cqeIxLmKbZiR8lvYRqwj1rLQ4ALQR0oi5CDN/w0Cm1i30tLf4bc
Nj26j7fcs4dEd2uXJo12z+mtqeYVmRtzWsGLdXtcrc1HxSutdhLoN+bffWUlsyFa
P9KfwCtwPQVmrlNDW6PqeqmNjnxsIfH+QquAFF0U8tG285SryV2XUBaztilbEfc1
Fli6wVtA9ZzekbD1hKXfjBcdAMwIiaXc/8rMc2yAdFx9aB9g98W4XVD5ot5lCPib
85JIiBXaUjNWK87uoKF2X/SHJ1H39eBI8pkJoQHqKwdLuGpUArWBaOD7LJh5cOsy
LIV057he2tNkhLp4gQuQVLd/fA3CN7Od24IkYcEEGPVFRheVtIhn59wErt/Pp8O8
YrsQWbR6fekzXtqrznPz/3JkN4P7AbURySI88FaHESObxO3/1lyydqLH2TcZVzJU
GUn2GteWes1aGYvLa+THgOQnd0vqAZywzeDVE8qzOXgSiAnWvYnGfaio066ye2cH
GYQasTX93OTESR5soBI4rppMTlimY9S28ZU8xApuC7QsWyCbjyT5lsqBc78dQqjp
pssCpKLXOQJ8QkUzbcGNPi7lGCnv5ZDOvPFInY6NK9TIK7YUU3W0GdtQzSZdTWSi
THNEd+YCxiaFue/m6b5lqScU8TYOw1AdGYjIu6iS/ijlRz+kbpGK0ZjN+EYHM1pT
RoF0RA+xbSfE8OT6901nW9hq6KKeEObB/lNz4K6LpOQW+6pjsTB/rRoV1JC2IAZE
KmFtTLafcu/t9Qv/nmFBBWnQ8e27PwEaNrIBXQEEGL+dx7GuMBmrmZU6K2HFiopD
8NGG0gJBwbY84emPTHQarS6ozWuqbDhjeHxX0LGBBO8VR8/EPERn78rP1N+5v9QP
vB7GVTK9V63bBM99jL821IR7Y50VajPXFWNUhs9hHLWgtPbXu9Cuv1D488MI5Oz7
f0S2zzZIU1NgCJQhI9FHb1doVr3W1yGod9Td6FEG3+22Vlpfbjh76leptBLH5quP
VSUThhlZA3tdgjWa3bPu8kRZepCv7GmXCVo6/zZfwjs75yhSu392L/gb6Fd92Heh
xlllnEWwO4r4BrxpRWYPC2I8h95mq7mUro+GxMg58O7OyisZJIVkS4D+jxS71wKq
KhYdbCi9QeAOIHsrQbewYn9E7dV4EuAPuGmS8Iv5V/mm32YH/wPCqJqQEKsu3924
i7lll7KzDgyTut5fmuxAbJEGlFoUVqgOLwkLfPuZ83F0dXRf3R0vhme5EaPvOZUW
uCbXeAvO0GYh2rMgRFdb3uRXXmRA+NP46GOrEBDLo0CIXZpkbqZdr+KKafo5Z+lc
MTixTyRlH4571eNDHHIZsFgedQUca8cXrbkKMZxhGQZAnb0sJnnsIspAwiX82vEy
q/Qz8oeiPni/hDwNGqC5+9FeeDdZ9EBCvstCBIXpFVA7Z7VNKQ+fpns921ig3r4u
X/OBk6UP6hz/3QHOUk0IYDsKSD3qZT+MU/p+d9mK62LF7jnVZPirPYiNUGY1YWpl
jMAEnt/ecfgyWeb6jWpxMSgeIJoYos9KHUedQS1yt74plraL4RRCMI8RcHhXiM1S
sStnOnwMIfOz2NQhNRPunOyErigUfVE+R4o8kqybQisuCUmUoGv1OLu4PK8+7O07
pHDyqz1ez6v+bSHVtBRJdr4oLxGu1weJZ2BzYvB5XpL02bXIE3kxghOUKY8IWrQg
WoUjMQd6HmnfM0T5GN+ou86Vfw/XsjLDDT2n0UERq6avQUUnJT8Wss+c5K0Q3YYq
jqMs2JcP45D/n8iErdyOqvfqnnblR7wKyLbcuzj6YnHXWwKzsAj40nSZ9GTTzo2O
HTDViaJvxaaQ77oeL56DV5iWnXP2Lo5NCZQPP0FNgqnWIhkKczyElQ+9fqD3qJXx
Ci3BN4sX9n3eUOhZgsDnnhK+vfpgd6NfiAS1pThiMjNLN8Wa5HbM+dZw8BakpF2w
h5PmcIHSTymAbNmq4aNQG2PVt68Wy4nw+zXZRgcsibLM2pNuE2YRCHv3qHWukjtk
HFQxhx/V76g3XUWE+4O10FoSTWcYdXOVNTbYpWJD2Mh+yyviSiveHSu1OjKrENHi
qD76toEQvqf50hGN8RZ+8Jp3xhTDEpVd0587CcUSbov5ohA/DrYtvu0VKgOmJQr9
1eyOvTdSylaY6TNg7PE7BVclNePyjAl0MrOE71sZvgCqdbMh0zqSRNbOKeO6D2PI
+y2UpBmoX8eqc3M0lmb/m//gy5jDB6nNO6t4kWAJQKU7z0iUNNcbViA5h/BXNfp5
pYc94vvQ2hPVJtB/uvSuptrNoBtOycgyUUELlBYHb67znJzH85SEkVLJENn8y27Y
aqLaiMlzEYJzl7/WyEAXV9r3KiLR3Ye6foBIeFsaYyROiHxMUOrGA/gIj6oTKTpd
4I18RvvbqVXeKDY1ipa1oYAXhF9z5tB9fSvZ1jjgZWBTrOBa+cetkmNeG9gQfPjY
9eDyWbWMHrtV51agTdlvjN/RRqlAG7jF6FtW1D4ytn7rccEO85iarplWwFFJOtR5
ryf+CnR7Iu2S44V/lB5cztls6XccQeHAVm/SDkYnTy2E+/jPk7d3JA3nKn7CCDMX
zCbjwZ8bVFDX03qsDFvK51D/pImLbpVMua61qMSOG7hnSucIMAi7DluqXbbcodlA
K6aBJ55YytjK+CuoaxfICABBZHrE2oYc+Ai/BjmLXYlK4Yjzn/iUGbhz/Ht/Ct/M
LzOprJxIQfK/6Yl6QTUuHihwMbPNMLdGEbk5KqXOddJRhhjjffyuotgK1UVRel75
Nxt9VFX3obtmjgKRoR/XlyMRzioEonvf1sctTE0KuLS+Lco94DuToFdDIN2HSkv/
h4lxtm9pkzUJaMFj+vJkB1ZTWZpv2HCCOGpGSr00z4kFiXmvVFwBXcE3xFIIzqbf
JPsQLiEBD3b3YP0tMiOtyKfDUkwrWiccnNqkz+VpYRi+IR0CJdXI1NyHGfr1WgZm
ooy5iZkWvgF3tzFoSaqRj0LSBwFRDVNoFb3K8td8w4Fs29DcMrHjcEvAMb93PGD5
bJIPwVv4YabrIWJGhd8v3rlKVVXnMaPEIIRzZbgxYagM+uqrPXblO2+IhmWaUb6S
jowSyz8mytag3WUdPAr3ycFNndYvNBLSiKkCrSmpi2AriZkGR6EPoqxbzgQER43L
5jhE8GBqfpCNV6g0Fzw0SRAWoXu3nN8a6zOm3tpil+90AFQT2Pxbm/TkjrD/hnHK
VZn7N7V7FGSlPAdVKlrMKXI3II2Cuz0vuGtl12Y9MaU8HYBx5MO1IVpbF5Gp8Rc5
xka2yjbYfijQXrbyk9QWIt5quO3yzIc+R222JVPyZ0IZPMSedbclg4TOfF3XYtX2
L/uY8VD0JMst3opwkDiiVvI957ZJM6nAseN1Wsc129PSXsGJ/AF706GYRuQMbkFD
fvFyf2L7F4QvNyEo5YerP9F3nKU+FIgl2N2tA2gE7xoTlzuDgPobFn4M4s3nEBMY
/lxLxMFhfExVo6abWOxESOKHPu/ORcGyXh2IhhzSV+UnkZN0e5FBycdBLIzjOriz
Gd+xgQFdXN/F+JLnfT/KXTDVKLcN3DBMl9EAu4hfKa77ziFvo6Xh6D9T8YwUwdEE
qffR8RIZfsllfqtzvT7fz8RUsscwUff0/EPtxUGgHfi/HQP6T44k3Wr0v9wMkYYq
h8JnbdnSZEJSNezyAu2Ye+YyXf+QttLefZ49anVfjrt9d/WqbsAQ9g2VM8xKY2Dz
OIdOchYzclOvd85Ijy/ILiigb/IjyKFhjeMgr3HovfvWtS0WnORVzoxMJ8EALSBk
ripDew79XRfK9wZhMhaAD6NH0gouRdVCf5dgL2HVGdYHnS1PFQIFXfNvHN5+PWcw
UjbPmDrbkrjSdD/dA/DfQD7la2X2ARWuQ7YjM1xChw3UtquhPsutQy1YXMEm0OWI
X+3SJG9fisiYaxqSljQ6pQIhh/eWYx4l1ygRUJ+PE14UTSNnjaYUFmRepCMyKDyf
32sqeeXSc8LNmuW/LfYeOj1YKCzyykB50pgGIAEsBjvJ1BhCW0BF6jXdXBHs+UCD
lYA8zr8HzVXn5WO48LAaaPZNlOx5qIwdFROFgkZI5NjavnWm3bBHGaYcwvBEIrEW
Y7r4saCymt24Zt1dsqLPIaLFGS1+ie6tdCylrFWWYjwFd8h4A/tyKI6Kl7yEHPiv
5EjVAVEF0RV+9yUoJeXeaE+FxW89+elMZ8PHtGNX4ngjvc9bWOKxOrOKxnXkXrPE
AeAf6360PiPk//hIl72pClR+/w7YOqAMmM7lT4fniDKCCuvuH7XBkGY0Y5GMzIW6
d2R3GeBV/LHrZMHnX+VEv2sfW5St/93ek/dw1ydSjDzvCee1wKy1lEYJYDrBHp7u
mUeBxC9X8qxFyfZzV/6U2XqHaLmxghA/0hvJZOkw3pjGhznDkboIldBq0eNy7qj+
biwZbBe/ITjoRKf2A1fdyHV/upGu9RMJPz3eIj9+mYHSdagOYVUaO9nRO1+bGXSU
BXZm+ytrjQO1KJrCwxemtTmaFSoSpgO5Kfk5IzncrJ0a0eJoF8cAJtHivVmF0kje
bmspxN/2aQk8H5/CvA1Q0+8ZEaZ5wkx2QMmJ6aaYVd9ol5aUwBdsbI+lULHLyVMJ
RIoNumQuJWjYE49/pm5xLYe03ttAodiTGmXoT/oNJCf6HYv52JzpPxjscfTGIYJ/
W9i4bFDz5Y+5Fk8HNWezGLX97H6ZPd6n/oeAdWYFcnRf4HFm5aCIdTw5NyWewr0X
UsxwY+kRmKDAwVYSZK8xW3Zc3VqdG4W1PKpcl0rb2JGIcq4j/TqhTeuJD8dAdRDH
kR8nbP4bbDFKlSOU5mVRyexSfcdWypxpfZkwZ4Vp2TqrB8nTeCmdDOf9gVcHmge2
Ry8Bqtjgh5ke0CdlHWh/dtJZAsBsOypjiKy78MwKluRNrw0z89w1eKd9wl4n8j9F
uJosy/SR5Tr9F/Ed+EZue9aGowgsBP3NsmQ0/A0BdoPh16DwSj5G4t7nuDjG9VmI
17siHZKsJ2nYOzRT7GWnr/6tZsmMR3+UHZu3lVUuC78CauRLaPbOLUEV6QduSAX4
xqmrpQ1CRJ7LVRZY7RhxnjH/Mq/9cM6O4EOGkXCct5KXzDow3k01g8Nc3KUhDNfV
HrQV97VbgTXg0moOHQcNr0zoOPi9R3XCw/Lpmlw4jPRocUHCn+8du7KuDEvbljql
AMkH+txOtnWOSrap02/QHGIa9Cx6JCtG4rx6qvCHzv+vLaSp/tgvU0u1shhpl98x
lnP4vdQ0q1uEhfSCBRVudn0ehjSQaeNCwm7Mfih3Pq/Z7DZ5NBlmaVkC5DUUBDkQ
F/LtHsuP1b/AoXd6+80oM+gPuP4+VVXPkxIZLKf2sagg8ffbHvhLdRhK5wWg84eb
qy3hrXljB7ma6qJGe/NDQ3JRuK2vH1OXZReVmxcwcpI9+WDHDutGnbnsnIEeBeew
m5XKfB8y+CwK2RNubPdwkt/x2VRHSn8x7eJBOQhnAR9L8zbR1RjKYp464gRaivAm
GGz0xsoKD1AkvsXasXflmujP3ILNRnEpsHwJpIGva6o8ozu+27Z8MZm/NVGMKfIx
adZLU6rQPlvpYeibMVnwuF7vtAo9ybTuW5Jq4AluRYN4S3U9oxkssIUEjjMc6Jj4
+CtM5NJDyIGTJRAQXXJwly4XMdMdE3e3uOK5NPsFrecTH1y3LBfdxNiVGJ+VqloJ
llSpBEFj3PCcJLf1Dkf3f55nyY2vlpt596uWl0zH20UZ8s7VCpdGoHu7pjO24t7f
ciYVmsXrK76h5+HP9gzG15AqlI9yHOvxG2y48I1xcQHwOuSUzqQ8M30vfq5if/wd
jFBuiqG2ZoVtWsMRGquNgltGyTe1V2Hvzbb41f1cWr88H9r3cy8AFW/59J9hX//m
X9oBja7COesL5zikeF+pc+iwRlYu2/8QHa74LNtDlCNil4nqjVXjjnU5F3mgkRBZ
HXGtboNKcuTplG4tHW7sk1i5PbqwSaDeQFdlcqa/5Zqjg0WZl2Y5dc4YI6kffmJp
CGMxCN+s9UBq3ohAkelm8FGZWPolTEYH39FIFFT5TITh22qL+mZieRMYNYIxQggT
IED3h63D/EKXrJO2sYvl7vJj9Le2s3G573io+mBjmNnXrLgdGHuaoymuWq4qNVCT
X0ZOZLhjZblqGZ3PZnBPvdP6SYAHg1UenUUeXKS1gLbglTeIHEaJ5bCbpjyPAEA5
nfGFNcHK55ActKpCDls62E8QhcR74/itk3AzLYDForVjGg1TqpfPigx6HGYKO1wn
jPH4u6zM9SqkC0IN6j+n2bAYppr60onRd7q9QeACTeHjaUh/Wffct9QclP4ILtYA
jMwoSppcvZkQWx0xkgjy9sCnmQYCiz1x6wGJLccq4L/+KAo//YG3PUm25Z5Zt5Hc
oCCILqwx6zO8Iu+0GXx/yg0UGbD3M/vuaFsajNQYIDips2Jk46ssimEbkQbjPDYC
PrszBeq8HXyCg5rcrag9QIilFJOsb4eZkyPcAoUPdwGXSaEPYsHz1FD1MqIFGrib
MT5iDme6+fDedpBz+yCTVirhwnwkV5H63ITX3BHEG2XjHr8yoIB9n1DSpaTSCHjU
zo+NezL/OPEvc4LJTdDjm8IG+uk9N/4o/Rr6cf/MOINgkWSHLBv7wzz/E8ITpyLO
P3J89oJOv3MpmGogYD0dWdreom+NN1SeHppVBFn+iCnuv4JZhMGaM4tYNxPAy20K
uWZoEHPrczpz+C1VfAfWtavbqb0uCkU69Ec6tRUkN9VLNZYtIMlH6HKdwTKKLWZe
cvzFy3BZECJ5fFPpQzapCivMzZCzl7EZE3hf6bXidKqa3opxJinj4zWZrfLcnCNK
FINd/4JJhtyhTgNi0MmafJb38ghmcwvwBtdUqHrKx5VlS4VqMWVPMldMJkl8Kwug
BwlZdI2a/CH4pwjrJ5NBTg2Ic9vVVcyNB2z48cIwiAP62RiqmIpbocVlFTLCJCCU
MV+Z4N2vLZX/rmwOyX8zzWbOAAdxe4/oa3Ils4sYHVrBzSoxZaFc1BLn4Q9zxykX
2UB3w2UAEHmf2EuB9ZlvB5H/1ZqkOKCemmHamXIvYp1RRfFmRkaH8iYk+ZmviVIn
d2AgXAzN0rpsW5J75WCKKnohl+kSRdzKo+4tB+4TBvtjGGsURzz61KwJTkO1y3UA
N6AmOUaMoUVM1Td9JgWeL/D+NqG1zcjpmHrwmlfVFoLWaU9phmtDaEF7WOBaRCBB
7607jH+pDh+hHxsy1YMxTnXHLuHIqSwc03o1B1bRJ9SGU2EEiPmK+oAlC/Aauiod
+qt8jTPIh7XFztGilszWAyk0COXSmSYbVM1IOQQRcwz218njE5EeMvARiSWPomw0
feW5wz8fsRAAP5ufSL9hVbsYrQHRV1VypRh0JLMuBGH7qBtPF3XLcPQw/I5G4LCE
u4grsjMXCKrlfxaW2tvTxrlmkYMCD+AKMNSV1N0j67HMsRbLa3eg4SEEFJV6LvTY
nc4giUKZCRrx7hDMRf2Yi4aWRyrqLsqIpDopJ6R42eEIUiQAeYp39CXrrVgWT63s
y0lwuwoPb3/KMkDW1mXgvZlVDWa9LyE76G42O7F1niO1cji5Gv1LLvM+fSKf5bEP
uP3BV990D7QyDSXrrySJtqA3Xx0bwJuIj/HaDg2zYQZnegoCX2/PXUAeZQnwTXog
cLbmkzfd8rrXEnY03ULiwz702GxMqCaufljC2FKST3s3SsUCGJIv16HVMi59LHkG
4eRo7xOpzhSc0xBB5PzUc5ysZK9L3U4qnkrMezxCKTosMnOE/DfAy1tWny0VpIeY
UL3CPyUhEfvMqva17GF/Hgt5ryIJ5ivmkLR+pFzXo3xS8FwULQq67p5u6gCo0rdO
WMZkKNhLB/v+r7QPQornAJ65MiDcezdHhlnXmEEcafi7TEp0rBwR8qGzUm9z4fF/
7IOL3P6Gr1KaWAK8W0tbKMZ11sOwrEmDfg5opawJvwr6Lmc6v4UaMACqqGXOIRC1
+L9CGCh4BS+QOzqq1WiGGQeP7p/WLGuUWYzZQV9Csi5A3SW5TrwO2TDk0znTaS56
pkgl6hEyU33x+62SLPnzqWNhuHwpJj536mAc2S1+U8zInj6vAxXNSFIlwgnwREzg
ZJZJZS06plTvSl+5QTuNupe/zE4NvXk9uXzmztFq0K5AmWUmFBW3sKg6d3XR1bBm
S+jxJrkYw7yazWkqkrB2oOdhXEylAdO4lBc5gBibgTJ+IknGoPe64UTeQTzE3rbb
YzCaQkFZD3b1xAKVE6FB9iFPMCncmPWksldUbZsOLK7RR37NHMg8+oyW7bW6avp0
HR/fXuU3a8lArp3NaDVWQEKTUqIBjSDT+YilYsE81NzyqT/C2h2wohqdq0C04Jim
lJ7l57/A/jqayh7memtO3GKfMDDGNWdTyg0u96pi8bzbx6/DN4Ud5eBTlEtBnoK3
1Nwy9BUCLae9+jYgw7w8UVQDjo3RrYAsH3XIp+aj9udNYg6BWanJU/+ay54mjJct
WabYosT4p6gZfMkx4Ff5geMjQR2jdUvV8gtlBBME7OpcFkFuQnW7mpaNVDN1HgFV
B1inFTIQtZ7cv0twN4jK/D00FMKZKYQpEWorLAsJXRxDmXAvy/et1XRHmbUqcCKp
SN2eF2jcB8i839bihcBmHy3WbOfGAUrbnHuQlJyAjo/pz9Q/3TYjT8v5cN2F1QIO
if12fqw0aHDFpF0WxQe6HD2I43FAPoUApchA8PMraSgitPecgsVKQNDcpn0IIKqv
qp6egvM3Xdb+BTA34GVqVEXlkWNKCymlEPX/Rn+r0AiGd2LjU+guP+lvE0CQvRcp
diAZ4HTpZnggnG/N1qJrMPo394TDJz3n21JCKISAZOh9J6ec5Fs4R34GTT/RTq3I
AiqJ49enqCnFagw11T/QWxTgJB8pfL6iDVzA3nVEvUS3dE7PSx+jibxDVDGCIIs1
F6y+ezrgNEi75nxgrxPDSQqeqFDPt4MVpn8/Hcrsbh4QYHsohv8cqirq3hSIIE6o
8bEnPUutlyPU+EXt/ufomhezLe/DHAsUdPi+96UxFUS8/wonkSIkprATH2MWcu0X
92k4z9ve8cnD/K/iKbCMHOJqBJ7PuxywVKmYSStRh22EiHgap717x629nM51wHW+
urngA+dhHxiVA9/+84U9FCWIWo5Sz1MkwC6IcTHIyEuLDlk3FdFZRcrvJ35d7aLm
sCAnL6BjExqSncME3k1CtKGD6UePfY6dIw88rbbw7iL/7N7KzUjXVWlmST3njHmB
9FRT5URiGl5GGAQgGsNgGWn9X2KujrcLgeQpczN4kGkQD6G3M+X4rjVKHr2QHWpi
h+DNv7rblaZU3qGUii/zi9GMkZr56jjsSZkzJ4nsUatFbJ1Wx4BdluYc2NzTWdQy
dy4BWhj5GDX/MzMxcgz5SSEAiWjR03okj4u+hFGVbuTYjoFD76kTWYNH/xNQUp2X
xy7KkQGg0hbPN35OTAzzzYU0KU+B3RIjam4Y2bdBk3r/TPgaelORAQXALDnMNrH5
wv/d/jFRyqakaKo1dJIbpk/pgfbslzzozNERXAbS+JcC45AcwjdoQfyR8HQJj26l
wZ+5npLpWFFuIYJKVYGr/F11sKxSzTaz3EMeFqO2Q9nTpSlkRAU/c+pANbp0nG3M
KO/1RKLc2FO6pS4EHUj+sSs+Nc+LlQCTIZJRilQirDdKyEdVxMbwO0pFYyKLKyLn
biL5wVt4MOqB/7yaEMgIBRvbE1b9D9KXoPj79CTXozNk5zwZNIOQGDWhMyeCPhqv
KgEZHqg5Dydk4RaQ/G0Y+7o3r2UeSwxh4lByfxlQMAO0hBOQWgQJ0JleYNfX9yOc
IdrZ2ii9YX/PXjpBGPto3BOXdBO1AYHdjVFK57O4ROPKX435ci1UGLe9uhcgWOfj
T7g+vjNfK6T+lfy16iKHpjGFpRzPljd0aSeQQl4rQ8fM8JexYK/Z/sjlvQN1GHd3
JR/Etb7qjsqWBOsis8CwuZO5NBbirfgFZ7Gqn4k12ZcmsdcvQ3cfi6UFI/bp+vnB
OCBxvdrTS1wULhj0/VXGXqtzZyreviyA9S5CJKOWJSuCQYZV9s5IaMbRl4JQk01O
465YniAr1Z7Vhs8djnTPo1X2J4i6a5UjO/GHT3hPV5kShRlpsmsMZ+m5kla0w3m2
anF7rrWBs6eGAYUuXzDYOeppVyWdZ2B4mtKWFByIF6AymkkjlFE8ycUktc/YNNWc
T1O5YVmHFhkFXYdCVud2Rh0MwYhrJhFyFVSQNPDPWst4rdYat38i/6PqRm//Euqd
loz7aqFH1rUBMx9n6iRZoPKtVXj4KBa5k2uQMFPW3NB3AuDQRQtHyxnSBuBWWLgh
oIz8AC6kMfPrscSzYxWW7XZzYk1DzSveVMu15w/tc+zSJvAePsvK7so+8nP0xg2v
5mTH+iplkcn15qXywmfuNAl9seAHNJw5OZAfEy0rImLLM8Wuk/DfTFYyk+CpDdqo
lWb0jFeZ/DG3DijV+f+4iKQYzZFw3n5A6iOY30TqssUCFwSHPtZjSr9yh40t4Sya
DIC2/Vere428Ycr+NXLy9Abh1s7iACki/8AAVjR/8lkG9kGeIwlZjFlWwpnPKM/c
aoYOC9BnzZgKT5DD4eliUVqdg8hCv86+TPm/z5sGDDUc0TGjI8cmsxHAnr7kP05u
umhAFKxsBhCiVFXRtxWmpAFmA5NZJpHU5UPM03POZ/T1rGSQ+czVChid/0ww1DPB
Apnp59N/6D1zfv5FKSQ2+PJpquamTPvUTwLpxY9czLh7Q81n9/rngtghAfnJrf2M
6CcOmRlsgxXSutEiNtfxXxiwuGM2teV7OZprMbW31sctNRY/lH7RUdn60gXmBsjP
Y7XK5y3DKNuV0m200GwAa4aUmqvLcKloqYZkqWEsYKfwqcScFZItJ0yHzfXc+dMC
ufMQ5bMy/TNhIsXye77CtO0g3BOmCqeBytLzgJrCipkJroIaHyx+Z6WFoGvU6AFp
dTT2AyS0knhxgjv8fZ5emXTd+EnB+qWXASLuNTB0WLMd+RsCo+OU8A83MfqPs6Kl
bKZzDljVwnB6w5RKUCa7oSv7iKXGKj/oXG+5znyvXObnlnXjp+Ji3KJfNjzfTWXv
7knIVa0Z1iOzkPdmTZ2IHNZSxadcNbDFbTU59mmvZqLRJ3WyJ64qptGP/XRKrlCm
hPgoeuzyalp92/9dTx4erq7d8hW66F3NndESV3QlLWbE72iKYLRngdbe52gskK8N
6OgamC58rhYa6ipvX5Epo9EFhy9AiXVr+2C/OyReE2dHry/VuSw7KDehNOpzZX3B
jJ7YZAEE8eq/CMZ/ZqYYdKrNGcDHi8CjJamT51Y8I2f+tZbhTYQI2b20YYcee8fB
6HzSuC6QvrWAVL7/BgnIjPMA6+PkZpcTkslXGTif1Dlc7C+4ROBA8FnE1kazWJqo
0Bb0pLnu0YPhNwGZ173fTQsvFHKeoY+G/PT3G14qsGmTZJi6lMdz26eNdp0cOndd
m0Lr6s/JyMEiPmV/eNHmnV9/DeuWTHWkwT/XLqCfRsccl3UNBr/GQ499pniyCM/f
dUrXq188FAnnRABxb6Xg+fE504JP+aQ/5KRO8YhSANbIX2Q5gOM2v3g/QEogCejc
VmK2BBSPhAyWLHZsQVC2LcJ0maqHwGfcUqK79UMSYsjyx5HCCeo0v8LLUvy1OawM
6ESJkrEdZTpUw6aSD16bKA86SapXa+UvH0myLH0zUPenJwMUbIIeyW+8OessVJFe
B/JxfTSM9zow981C1CATt1wxQpZNSVLON5a9nOzXQ/5GAKbVQcEo8ONDfhZr07Fg
lqCy4FaaRedviODjKWtbg09ZSxcXbiBupEwEzHo0cg4CrHKDDs6heX+9zyvXxzka
8BR91kxN9ywYD9KFc1zy3iZ9EfIq9oVsyejkc5ERV+4ttgdVJNnJRFdIUzcax0z/
g+RAPKqJkYHbFSNDARTqCdTgmR4oRG1V2wMH1Ng0fA7Yx6EYymyp0Udw4e0gK0Hc
FUdXFMruyZPgucpprJieND1uywMCp2B9k2fSY6+szVGPoC8i8Mff9kDRd91FO2Yq
fXUFDLox+JluVTughhqCWL7BN5QWhqhQ4Z8iZ0K4Pe+A1RaHc8cgQ6jjnmrlTyZV
mOb5hT1uoJ19JH6Zi6JwS9iWNk+F2VRQD0cn7iMrh8h7FsIDH2lakCeEENlDXduG
aKqvqqJdAChH3aIsb/7HxehRKaqEoWKa5wWtRwzyaeqASuDfGZez65ueeVcq7Z8e
dNdnApsdAF8Lt7JwoEi0J5m1+8adX4YMMT/1+XAi54Vfjw3FF3rtNUbEEEnZv/6O
l19J3NfNVdNtg9L36puMszCTrcaTNACdovJgALJyVpZCJZ4S8B5lvj3zp1EkT2NG
KU+iGWk8k96yfdsy7ylibEC33tyl8cQ9kThQiBZr/QBbjYmCIgH5KgtGDoeo+6Q2
Bky+ctSenjCjFFpTl+19q/7M8+1fcPbU4C+42QW3AKRZ+QgNoRar3WdDHJQ6sxSH
6TNgknW2ZtuZ8ju39fxAUZqhVJbENHwCv3mD6chgzRGIV0u1nqua1hfF6gYWLgPe
F1x2oR9F+tiWPiqbPN3c2mHxaH5LWoIRPpIaAkVasUHSl7kMx1Ph3rroSOydgsx9
zWD26uwBv/7uS1Rgo/pA4aed4k+yzCJkQgI/nMjstNhQ+OE6NhkuqQMrroD0T+Ct
tDXxMjFjjZG6/68Naj5fnMuBar4yVDlzr1ZjdnL+kTCd2Ogi3S6Ta8Vg+lbcs8DA
fX76hbQEEQY7GYkaAfIusuJoBUeeUlgTd6GHZ87sCg6KJ+u+CuEvIR0OGePd15ji
VDygBZh6Z0RDh3oVdsrYkb6Nb7pF3JWMqt9JAmOEqGJf8a8nb4d/+cFvxqpYGXG0
npbugqTnwHUW0YNFl7rwic9FJkC8YiVFyF87MLLKpdlcaMz0q8XaZ74kBUxNd6pM
S9Np4wcPSgv2Vw7Gq6fUq565jTVAHi6RA3UGm1qgJ/96lHh7NMIm1v8BhLWK0h1j
PRCsrPo8aRCnlKuHvWPQIbPXqBYDfep/cMZLabrcj9s0Jgz7ut+/ifErtSj+H5c+
lUlBKOJ8EelbxQGSDsX7ZYoX3tS5LN8FWm5xrysXaMTlm/Q9HsRyQHj1nx8i36FN
jX8HXZvr6+wRR2X2Bmn7xNdsLdXUQ5lCQY1wrnwdZc+v+BB25qgDePYlHyfvNc11
AUy7k55aSsYXw82HUFOkOHkUdNxRYNIXCxKcf+qZUfboeAHota+uZZe0+D835eB/
cDW1vwse9oQmTRoavgoU6nGSP5YRoHexDD3Tj+Ci2q4Yj4aVfysAtFudJN69sC73
9B23KFG1Zld0OZPTcP43o1glzZ0ucnhJ/0Hb0+tGHqNZqvqlHA++JckRqoX5a6/v
rQ6QWei5olDNrWt3S+mIRrmYirCK0w0wdoOajpdp6S0M/EjxoshAljxHRh/dDk7n
2zFC7P1cdTxplWQ6zcX8GDMq4h2ZKtl/5lUcspn+PiXmkHb1gJ9hbKYkQzZwZZcX
zopWqBk1b12aBrBNcEAC+yDEYE+FZ/Zv+a9Qub89qgT2I2AM86RA3HVIvc9pmXxq
WBKdIdyvEr16g3i0CiDRbdTm1gLr4DUPKAGW656tpuH0RTyQlUm14NMpzD+CjUbF
v2guPAowPsyWq8c5Mc0A/n2jYeR788BIvIPIT3KzEJ6x3DFuaXIHMm/XmMC3/ryN
fhG1eJlMx+qc4Jl2buzvdzyXw+o7sUW8uaXMp3ji7DKxvhOwZWZqjhkgUgIP7v8F
gJn36VDaOYA4Aa1YuuIxJT0FEo8HiRJF8DpWfP4C8vrjXSpo6lGjnmOLK0Es8zkd
8ifo3ZSfIT2OwARmxQUeqPu6gotFLKM7ICZeWH5cBu025Ag8bCikTZyXb/o6b5lp
e0BNuO0g+P0EvXLEzg6VyO1w0/KPNFHZSAGZvPgGOD6VAzL5vCdSnd12PfYz6qWT
hO8J/jWTJAiwqMmjO42c0CVcMOEbrSFOsIoj88Xr7npQPMoDL3uhgjUR056HahMs
9NTnD2kd8+ccEGsvc+bxaibsjGQpTWesPwjDsc+kvCBKdFYyDlo3Ht1fI1uPkxaV
xX+MojHLcNmrVW6Er0Wy9Nkxk2hDFATEA4u2ymD+ueck2vkY1OPxcKcBysD9GBKU
IzAHlSoX5ddy8eIPZFAiea7uegaaDeX7Px6pvm2wAsfdhgZQhuEivRhiCccgUNWw
jWQ6bBRlENlZchqAcK++i10Mju7WqUSptDZUp4EcyJ1yMK8nBge4rhJ7hL8izaVE
w0T5ODW5cBsJ9SGxxgAfDbD1iPAxhaDN2H2Aq/qFFgo7eXQtu6SXbjXt5tPRvKR1
CtKU521qL7xD5fro7BTQuKWDmxo6Iu3+VsYB7hwxQLJFLNEC/aYR/tm7ZMEk3Ex7
olCFIy+WtNqHKsKHDutR8ozE/Q3X/DweyjnMBtXU8+SaWLArkOEYtmGTXKIiZXP2
SFIcQO66gFbsJUuKOUC8Mos+zbbh3owAsDGQ5OfCgQ3p/DTFdiEV0K92O0RoGn/I
hGMTgGPORdhaU1efWLI//ri4imCdI/R5SOv8O9UxgrsW/Zfn0lTy8Y4YeT6iix8D
XcgN9HyEF9X7ZDWwN8vJ1NRwEEwXGzHoNYAZh3Ri6N+ptLSSzAzHKtbP9wGde+H4
WIDebrxWCtXMc5iVnJX5I0FsBsIKUpsrMZejDK8LdasSuciq/+9oYO8Ig+z7Orwt
AFAptjhwhEO/BZVWZrdeD5CfQOmQJU9pJLM3wLVtRM1Kjh3FVgfPRHSSiW1UOjyN
o7uj361rRU6lwaTgeKGrI0i+QMeL4WWTmQKY7okRphkRfnJmTK7gO9nOo/cMbdSY
Ca506nZqDKZsBJOVtdl56i92UR6pnbW+HWt+Qj2CAA/UTfSUOJiQL1rd+ld4lmr+
T9RkE3IRmo5H3VS4fs1JUfb/jIBBsa3CsP31c3CbNWxu7tBxHNt8fLv4rz0DE/aX
LbBwFrXV2tl2RS6HWlsj2f3IWFgrgJD7g2xOeKCDvNB5SdbDLfheHTjESpVUnnIf
qsRVz2XomcebgsMsFlNC3mCEOrjxBaYiLOEe9QsN0cRTiIrVsMiXfRJtuE7zMPH6
r2350aooKsBYSo59pou4etl6NdC70nz85ldur2Byq8EvoBHIvWt+PoAna19Q9V0W
opnSxoN3vjxzW9dPD9G6AmIZDwrLi4NXj7IrJ/+9FYzDaL+ugW5QdckvLCxdgQtK
sQa9FEbWCORK9xfOUwWmwtK9Kf3uqWPupurDvTkrZIUXyWWdIsmxph7wMMs2o1b9
F4OmHCJmWV6zxKXO9HsbLi3E/C1SjFIYHwpkhF0t4Rpv7m8XCn3uNdP2wvNmbzBA
PJy0288rH0vCSLhnHqCz7akpMuX+leYcPOKjJa+D9nYqR5JcwITJjSphQ86MIiUy
iFeQf1l7awFJ/KQ/Bd35uRh15Z55jSitEQdx+HCvw9ppJY+3t7ClG0lgPLAV/lYF
l4YdGNojfjVuuye+rcsflTG62pxNoDlJpNoWONpNxHA9SjAHE4+pJGnPZxBw9VAc
9hRTVfAvM1w9WbUw20bY8snmiExN4QjlfvTjgFx2H/oqWWoTs8mHjpiXslnvYPHq
rakHJ7TauwQoF3i76n9EIquuBRe45npRKHjhNp5Z9L1F0ThlsMHf/lFSnvOuRoxV
XyRMCYabBvrJLsBfaz2NgSxPANz0cZ+k1A6AdbnPn2IRG53Ryjb3FCE/ZesRwgxu
cdqDVTR69ko6aoi4GfI4TLbxDQnkFCAEDJ1qk+Tl4yDk+zLH8GW1SQjPK2uOO9tR
TlYK7EFmX+9RvFtOXqcbuAY95+YBYbyZWhGZtx9XtxNlv7N8qDFwHU5T2MPJcY1o
Hkc74eJ3IqDqAZU5t3oC5JCyclyccsSHwtYrdeu/vHbfdi8PTN50rSfhYDTHKe/M
b+rY3J1+NcPz3sp18K8ccIAX2frVvsR8ibMr/OUuKmHZ8KcbO2wg0Gz5sGxcuByh
0tPSgU7soDtsY+1qae6Vj6r8u2otJ1hjo0kd5BJFR/MsCwwHf92i/SrPkzON/y4n
q3BTanFY4P55Zeq2yQOZL560aEIyfSttOo7YfVSB+CdBLzbxx8OCFucMcSAmsarl
HJ4/XRzQxRegMLb86WclwdihrnraVZpcuxQpnESq+Q89QxDzlw4jhlqdwNBdHwlL
QMqd1SXlX4/KPh6O9UgQkqJ7ZX+CRpb5xxTDpUsQvYtF0tsHTXGm7dKta0H/oDbB
FBWGgAQNoae5ocG7HKwN6AYRMvQqP68awjLZKi7XwodOkooy9ENE+oH0LBXPhtX9
FMT9vTVPUUDwzpmZrfEjLzSrVmlmuNw1wm1rc2kJ9TDsQA/h7sIG3PR0H5lch2HD
2gIw/3g5EbL9SZR9j9+VMkSU5u2aQDF4uZV3z2TGCbvl0ONRDlM8lyZIbB2mZb/s
GbVB3E46gnG/LCNwC0NyCCv0o8koea7kQjZwvLbQGpAY3BU25+h+O7dXQPGSawVa
WbF/rNGnUt6C761t6XuIbqRZPVhmq8PmsFhAzE591EFRuH+4pPUOxvjNUIj9bZvy
AVaXJuyBKE4kvTzMA21EP0QtSIwqavrhr1Dom4sHVXDjDSoYxWsLCW7RCYWCYuxr
XVKEmhOnRMtMbwPxem6M2vejzRNwOACf3xZUzHEoqol3pi5fyS9pXe6GZ8G0bSZY
kv9IGbX2eKP7IdG5uG6Gkl/rMOJBAorBPGvYiN2t28pUVeTwAR0fSgdUwjyYc+O9
gBa6CXSm55YGnlLIqpBZ8w5q1GzMn8Y52eq6nty7uUfttTUX7x5NUhoozovDcTUp
9fhUKAYakb6/0l0X8OVA6coXInBmfum3CGpjYSkpTPnDftXbqnOiUgnV462FY3I9
g8cBbNXRY2CfD+AsCoftRBD0yTa4MD62yFJ2tb8SC7pEIuloFf0fR2SfGxsrpckx
J0tXb3WvYK31D3qpP4kE5vaB5Qba5vGJKgpCVjhEm1ZJBJWJYgrmIpOc/WODqiP0
Bf4yIE8/wa4/kJegeCTnoCM1WRSG7klK+YDG09wlEuKvR/mj4wa+j3R0Ny2RXmKQ
OAvegg9mpWCYAaFiuywnAlobZuA5zKwOnaxnOaTKOXHMzBpTy5i7wkiShwoJOpIS
iD+POdJU86q+r/3fFko0KROC5TCMMqvxNRHQWxD1iD3Gjt6qyof/lauCrznPO+Ny
guRYDBFhjR7BxiRII0M37mdDEgMYlQxB2/xSsAb8UjpEwDRv4JQM1/eYgTIsgoM8
ad59kttrTN6LFgZF+duCLlsFq5TAw8TxT0QHyx6EuyOsY80L22iBK6ZfjQYi36/K
Un4YqcDPp6FK48NYQ9xIwi+3UkWKIN6bNsynntd45W1k3mg3xgDs4pFiwRtq38OW
t+PoK3YkIwOm23CKtfb0XcRgZhFnbF2T6U3HaYIAToI4UdPpH8j31O0w7Ck0xJgZ
vTOJwxXbS5WqqGhSedHtiHi0iS0vuST3cYeUKSdeovKUixcekDey2uBWbnBeKSrA
ltwotH80HQC1us2m3ThLqwkChZLqPr3EPoObORA/dVsKEnXMt2QpjnLDlnCYEdue
JxBi6J6pQyuVCqz3qE/iclZ/87gWHhaZk3pKZFUr1Lddgrx+kwH6tlzPBX7ADtbP
qtwCOSXnF9PJrb99JtjGNigWXhbIbo7dDoQDLpC74nBodGpDWnUnlFs5RDQ5KRzB
vo3FQUtoQEQeG4Z4h/k9y2Ab9hlkrKPh1OPX0IPhZplCHq5EfEQgmQkV/VRsFz0R
G93uNTvFCOL5ByAk7PK+shh3oE7NEyGd/VbggwtBceQH/lGQJ4pV2AjtaHVjelpV
+MJKieGHDRwHVzCnn9hh8Bqa1AXfgWBDky3kYmohXhwl7fws+K/DIQ2aMWdrBySN
aaUh6bBaGx3OBuFAdY4kE8qkiORQ5YD0/1wPYWONo5x4nWTep5iibylmh7IzGhKT
HdBKUpew9Q0ULdnSe9UV3LqzFmCqJ4Zz0FJCHRQ7kaI0GL6YnczSDYt3xLuXA56L
uLPBcBOMsthCa39GpjnMIoAa9L0bo7yplIvHgEKfrJi92DGqH7wWpzKiytGa5+eR
wXUy15EUb4VAAcdR/8dLn7Ds2o6FsPDED9tFghh3Sm5MKooJ1ADLQiZFwboFZv/H
VKhR9NNkOmfGG1nz9b+ckhEcbxrHUaCix/59ORBATGoE0gLaGHHvLKel2NxBMHyD
LLw5T1E+Ly1SXn89mf/8UN3zPu/AOXIaJWU1RSyEQJfGLcHE4cr6CTTucK4GS+Xm
K/OtcNoVt1Rh+uwSSTcqgEorCuJxzV0X0mBy/k/2gNf4VSGgq/7r4hoEehR4T60h
1EQtKqlHPn2+s910Ys+Trd7+UVenQXLDDbrQyHo8WgnWpycqu2KxNczC5IUm5RJX
uQIo5zxX1OlDOMbA22zsfRIp17ceZ4+Gi/o9QGjBMcwVw3AuLN36ByUBCdTd/ftl
+PZ7fAFQww/3UkDTScqmN4UZUhkIQ4vOAhR1lEax38DdSjTB/Cv5rm+/RdaWrRpq
DYeNefKnFlEi0ocSGvTDYSsu9i0v4iHLKCYUB5MykblvQW5K84RviEN22rtk5iOi
05dAJGZG+8Pbp9VsBhrY9zVR37t8qVPB+MKpDyxI6MnJ2mFYof+9mrqvkCi2mdU6
XKGsu2IbS4PFm1lC3H6rHKoICV//IG0UWJJlKTgwprSfjbtG5CsQfHDEvlx2LnVI
FwlAnEJqID2NLZYDLiDGgVUU3WGOrb16mOFzgiRBzLqG5u/bv1WHHEOTYqNt7edb
PQNTFxLZYlg0rahKVaAEs2jL+FuZlgHHQ+h9KMZJRGw5S2pxh5YcttxtBar8l7oy
u7lgKNk65lhfMWjSGGD5usgCVg/DcGyZ8zkiHiW8zeHkE4Up7vq43HZ885nd0e/+
5QwGOv5dLKVqHQU/me1/E25u5gX3XzAq1dVNXnl70zjeZotqrwjQvapNrKG3D+jB
j3B3XGPjC9gLQ91VyYox1iN8oZcuHBcU/GJQAjOVcdxSZYsraYZxlmpM1LssA6jD
XfpBKFoyv7rn+a/42Ks4u5nOkTfidfyqKt/trv47i3qVcKQtZvYTHJ3iVeNvuJJE
A9I1oMdGV/gtsKP7g1HrlN6GtT5hcn9G+bIvoms3JGvZBy7zabGavobNJfIGkd2G
85jfzlzMAlfw1HE6sP5w/MENva9y+x0v1fXJH3Xtv246a7KLtMhKqJ4xbotNNDZw
0TuCvtf6ao+a2EszmuUiE1y94JJsFYngl2HLE7YjBmwxuUNDJMUDuovAOGsRYFJs
sxx3OVKvAg+3EyekuZ4U03pZ6SHkQZl4a+C7cNG3wtbHD0siaBX0NCzaMGOOVr40
tRJbs1ikiOrC4J+nK78AGPdjsAeczhfXwaxPcHYLBKlqhuB1fpIOCPk44Gcs/f/o
iuyB4BsbW9KelPDnFa34QV8hfjBRk2ES5ljwsdlNM9BczTYGOqTquKetNJo7lPsZ
fMfdo3hj9YD6cuwMMJnhSl8Fv8e+U1YewRKQ7KgkBZuXzz2PMJMFmN00BeYdeVoK
rOT+WBbvYw1kzCxC22kbqWeAgiYfI1ULnQoztk4Xxe9foQ8eY3psd/Rc741a+GPi
X8MkNZQitKQulLvBvfsGdgRaNer5Fk7wV0O4vGUOuXewdxWaac+K6cK7Gfpg726b
qd9mPHG7tAQbf51f8ZfoGxv5zexLFmwxCU7H3izEhMKb3+dhqZ6AG7FhMV9CNtET
C4neL++iq2CIROpX0HQZEUpc1STQhsboQsmUhWzs56Une0vSmArHruh+UCP7xfrN
SugjgHrBPLUGTzDmob8NiZ7FDvK2f9h2cy36U10HQ9SV/ckIlfw+Ez9UWMMDHjdr
S/MX9AwET9ch/ygKD460z/BGs1yGA2rMOJR71rpd+R4KVyOPAUrcWZpWj826SjA6
2/ISLCyf3JB8+rXtfYIHpOlDNruSs6ufNeUXuyApcUCCYOztRgOpSGUhITspIoHU
LyQSPi+anXCXLsQQrZwON7ID65ERf7YBcMk+dSOfeYYpi57iUMC8VfAmwvlCzxNn
wDaBuP8Xgm4Zx8zZc13FMIry0fbJ0PLxunHd8pM+N7dHEqr7wfJWdUKhEasx0Psu
p9pndgRMk3vUN3cPwgRg3cBcEO9Yc8AF6R9XmSQLRcRvYYi1zCd6hWPwj+PL1kqv
6L5bIIzqFC62M2lyQP27v6y96WqHmbDLpVmLCtPFr70dB5aghcPQgv9k8LW07BIg
LeVhSj5nDoEgT6qX2JfAnYdjBxY/DWa8pPEeX4naNJE79v0Eu23KJFhd/66W0HN1
v561knipY+4Z4pn3AGumj3KwIv3zrPfR2SxUf9xs9aYeOxYOCZekT6NRR7guNMTR
OdxvalNmRNdiRk4rRsHo11QcvfSFcHyhDLBTANihAl05jCFW9ioDlDtAM08Dt5J/
QJunOyIKRWWqoNta6NoCkssJyHOFlOrzNfZEMgBDMEDh8vKvuynaXBc7Ul+bCdlP
NohSJplVU4bqqB+CDx7V90Pq7FEQsVi0Zqq3gwYo333yAY3OOET657G9cW5pWHir
5r/xIhSnwRK/IC3BK0J2r7AEiRm0reYoyfqHib0QIUcKTN/lfIcXnoXIc70UOtL1
bpjYNG/M4aNilMWH71cL53TbEapM9fl/0rSVmOI/QtN+UAIPgWmjn1RM+Venwa4C
fjTa2ZnfVHI2Ou9/vf3RoH3kX1Mqb7mcJYLCvshPy/OydIpFZADxaxGzGXlh7z1d
/PX4WhVm8KhI9wR9HnbUJHNmbOUKIysOAWzM/BgZ3/xO4T9aNR99MGJbY0ksFXE3
ZF7IHPAvBiPjGlg7Z3FFrxbejfJbIZ3d3c3SEZAT7X+E6Q7scKXiwnbXJqk9R5M1
BDy3y10/0iVQKnTCVn+68fNZ7Azax/pbHbsUCr+tc6jgOqAdCos6ggaBzYE5j/pQ
G9x2JdVtKnbsIATN3uEmaHlx9fIJykjTE7zmV/ZLPulek5e8laNgfOCF8SN312Wf
ygMtZStwdhI0cNz17e4fmKjdXrw3BjQ5IaKFEJF09Tu/rp0Zehxf+Wmj80OM1peF
CFWeb7qPmpdjx+m5MwxH9Gbzp2ufv9eQTmLYkyYvENAUWmNt+l5TLN2X2LxmSUrY
JF9eIV3xMfdVIASqQ0PvPJN1tYQHyAlIsWFHKJNDDjHDeyymJtUyvSsbE3mcwin9
h0AwwEgXCmMbqehe4YGF9BrGWdib1/4cHkLJ7aWmBb3DzIcNIiQWnbUURlE/D0qi
mvwRNy4TT1AlPScsg/Oozg9cNwM2YgKp52rzs6dSzPUt75xmU+6Ud0s/3fqBFKbr
OSlp0SK/7PObNrI7Gx8AbSpvdgaw8IoP1pup3IRGn/Z4qXO6LcL2JC1CuuH0LxzM
UbdJ0RJn+C/YLKH4r9VP8AvPqNGXfED6sZzZppRiYDsE+SpRRXwZLXW2iBZ1GuhY
QZ8tYj77bsfMtgX7vOpKdsazur1TSnPtOuY5I2d8BYSKqLso+c2I2zUfSR/96vfE
jQMTlIcESZTzuMAN+4+AJRkW/0rdLI0rmg3f1tnixO+QoZRR2l3e87Fyu7Zz25MU
5PIqIe4V25PTtVPrPxc7u3RKzPJ1i/DrirUzhC3m0GwvDzUja4R0Fbv1SFTWQwSw
1Q+Yc+RAaT2jwfHao4ocjA879AXFka/3Nt98puUNd38XNkmA76wszaT9OLOiUXBh
m02jE4NKj8oqIDpuHIqjhK13U7Pt55Sp1/1bwXVNBpLvrnz5qv5xyMRKbculBp5t
qgfKfwrvix3RtXo6eZtT6dBKjU8wrK83XIlSF+HHBlRbWSubAfBnmV+jTE/dZKG/
UiVr5ajnGoi/KFZkZ6hTOgIHLDjknJG2njIggl9oyCqkStOxXWDzsTIfIXf3OmNj
rlahSLFuGgMPIC2tSwYUL+wpdcMrwyqvIZFNlNRr9vnbiZtFF/hm39erbed1orPD
CBbz8ca18C/vGLOPUGI4gqvz9Spdg46lfVz133LwO3m/BW9cj7R5S6mbP+gVBTPm
manpJzbJGizt5dj694NTfGoNlW6GkEBmVmBCkcUO5o7l/vTYOVDPKP8aCARBmaa+
eqZXijJRkzcOtrPSStXHgdqM5CVeXDKeoH+5FVxkRh4DaGAUegCdpkgVdpoGD+9D
AUuWLXaVhfeOzI3XP1zr8drscYseIhDy4FKO833MT4nSNd8QZa+n1S3OI4LPgHJI
u9bj7DFdBN5ZqBUJ5voKYnB4HXYiguYZj0q3SqF0yH93iFPLcb9khE8+B/rgv91J
BX72QOI10+K8zTwB27+lEgD5dD1PcjgqXDO20R14DDjEvjgSzB3deHrK10ao7THE
ozEDPM0Jk+zFh0rS/H9K44hNLzxbfJ/39SIYWEJ5feGlB437n3neDWqomfa+LYkp
9Q+YWo9kzVnjfhHOfQ353ys6a9JEjTzs7DyifaoTAMNkM0xvjpMPPoWNxyRx7XiW
bG0swv2Nd+fw9tMfo3LpDByFnowZOVPl7m/wCDr9XDLTOg/YemQWc8iRokEiQix4
mAC356W00Mr4kRpsLiRU/jRcDRkNWcV7cTVu0nj1Wu06YmuYVVNBnPTE6HdyfYFf
x6OWistlKoRRmt6zakAPhGnsW3hn8MNheXeUNMpQCXuOja3giZP/L6rmt7YYJ1yZ
joZVBXbGsRXGsBH6nnzfMP0qwL0D0j+yIf1/z8TIgXvCCBCuMB/18rQJhbBP0UAL
ERsBREOzUZUetr6NreJdSw2Y/iP96SNBfulrawUlAtkxSIm3PYuyFd0v1TsSDsxQ
uMihclGKfpbtBCCwQ5+3ScoR2a/Fowj47op1Wn1rShopg40FV9bRmjnrHrGJOdhG
o6IfHQH2084afiNi7Tq+Zf3aHcuBY3VrBjJIVa4PkpB9O315e4mWRVfmcvIXUHD1
PCwiEbKxeVUo91lMbw6f0Ua45XnTMVjBccUlUwpDo3fwaeIkjy+QgKvsTqPtiNdz
v7b3L3BixL/SiVI7YXcJ60nULpo19WcEzoruezrr0qtOSPw38PmmxxGq7FxRDKe+
xUd0W8YKuA7sfjSo59Jc9G4TA0XrwomsS67VhkxeKp+qHlwDT7AFRXt/1mnio9aK
hpBVoTjd1cnyknvST6gj39wZsyg2SUZvuU6eA20iROO54nc3Rhj93tBwqyCfiLfk
WtcLtENl0zqGv0m/jyvzj/ooj68pfzKodYjpW0NBmqLz6qw2JFXh6ZNk9nXiYmhG
p8wGsEr5aUVbhjxiyVZxyNJelrFeFe4ydrLzoxkN6BpyAYUWuGkSp0mOVTJiomZy
n0Ka6W5zurDE0Awlh6y+l9eDwENqnvQshUOJEo2WCX8AFVfiopI2zAsI3iucUnfK
DgFtEZ74T43ybpiVxBcp7Ffp1iXo2RYXCnMJho3dvKdH3NBLRW7YjFXe12aaEaPN
6Nw/JZM5rC8Ffu65BNzmU0OMLnNlzRo64BaijE2GUP6xVWf0aTt2O6ALz5fZpx6p
TZRd2smAUio4Dad+okEYHg3Rv4qYPyPs4tmA6HW3pO4Qxx1ikvYTb12SVirv0fDm
gS2hv1jC41w+968xU9cavvjB1MKY/Uq2RUdd5n8nyjWiL232vduo/gig/vv+QFOb
z08E+NsfOXWLqton3vQ1sZ0aWcouY0VvDoRNxFGmpeKtmfZRTEqcSCRD0XzM2j3C
2vtLUzZClfIcBQ7rceCpVXeyJ/0k3fPqvZd+5MnemPkgu1CcxRBAFNqkGrwXOMoG
h51BZ4E0cKo5QK/6vrIKkQU1sEZZtJzzfaFtqeukgCxHKv9peCfJbkpkjVz4Z/bE
QNEvu4Z2cd89ioN9ao2Do5HtB0+ydiFqfXkSSm4PLgWyDFm8JG1abp/1Bf+u5JTg
woNseqkIvxiFbvwYxZ3bPcPPhm40y7ZFv6OnA/IUO2zRraNG0Yuxw3GhVYWsL3+l
QEnKhD24m3rq1QgcOd/cn047+WbffARYMfuF17X0JY2aOOhsqUb+RFqBConZ/1fA
AUj7Oh4heBFcCy72aRsxY1t95NUlsd8ENU1+WnO1xDDfJ4H9tSx0hKjCeZZUZUwd
mOb5xJa3zdWsJSLFjkwmPgzYw3KxmZ8mIhyWvX0HF6VEwdpzKQsDobvo6Iouq2yj
1PrlPQk/1JngkxTL+FVHXscpTEHfbHPVKvCPCQo2fXJlHIlWmIuHsO72/H/V8nba
V8T35SjzuAWfD0sZ/nLS7tStkK+ABQYhm8bDoYMf1UCjaTI9q7/mdGNBvp66Ad79
8CsPdQ+yQywg5PWjZR+z5F6luD002Quctc8x6nZ88WqIaii4rCOSv0vt8ncveUwq
Lnws2E0o25OuDW1j/kxugTjA6xM044pp/0WHqU1r4cH/8gaeM50bVvuseFBJA4fv
g0RaJNAuwgiZS7rxt4twj9Sgoxq2TqMxda1UykKex5Ln6lqhvWsiYIpv24mODWkb
9tHGaYugo2dMK668YNPpGRpUzYQVB+3448sL0jyg07PEVfeD8RMStczulTWs3msJ
6SSBrButFzjMA2mmTGYYYRBd+DABPs/+Vwo1LmYyVJSmxzbb23XFBo+ngZNRFfeZ
5vrhfS6Vyo+EiYoqiAiFA3PurGANyvQ/e1UgNDPtTCFNm206NiKzdnQeLXRDlugL
M1/2lUDOasIecW1DITrzIvv/iMfoNUv+Z99Ziit3wIXNk2mo2tqIuHhMLS3X+p5E
Q607m7SuQOU4P2LnIfBA3m0TDeLZ761LPphLuqKSeSdIwxqVr1Xn9zS6DGqMh1wA
bRnDVI6ZLkFbsJG8b5VC1CPVyvpACOuXQ7EOTKBEorrjnIQ/k3XGxPsi+7QK6myH
x5+3xA2r3FnUF1ybKusKiblYfPTENRNAJ81yDk0AmICodsjAbd8JPk5L3xTNVpyj
Q5IPknj/iJB9kZb2Hjp+iu4CNFfQjkulqvwjgt3k+7jhCRnMkyg8R67Ay4WxsJqD
1sud4dEC1M2KyoNMVYWyit7IafsGXHFPqHIcRqtSG9Yq3gUKH1KZpCye9VsGD4+c
gxQtR5bCyCsb0gCBCigj4JG5eOE1ojvKlM5swmqsQppwQ7Wv7daLFZdPAvujPF+w
GzmIDfuMxrG0gYuB0xneW+PVE/72uaXkEojE3m0QFdsWuLz/4YhZlfHQGBdqRJ+5
YZcPjMk2WKQQ1wP34ULA8KdM/OpAEM2PGvdGuqDZj4Y/0kpNGiFWDQ+12zu0pUNF
hBZ/9iIzP6A9g5BN8JzUUCJeTif3Nce5hbvg3R5H4ROcWa7ruhOwZlY1LS5dQ62G
PGSpsqM9iUpzg6kI1NBdImo/yifGEnzdMdQzlorJN5Blw3zZmXz/eD7RaJMeITQs
Qpb24z8ewRUZAaWWvZfoBesxvT5sGeGCUeNzUJhRY5j8B+bKTwQhMjeA2oBKO05r
vUc0shW4HMBmhmC+yMPQ2eZjcil2etKTfDJUPMQ/4N/J1/9I8HQarZ6b0n+AdIdH
tlD43lDN6wmDAvy9WTqgUM9XcFp/FUQploV91AfgwZdneXYZx8ths83SbkdqSbgK
MpEO6vD+WTUkba9Uz7NfUGzdc8U/zX2Zm1JlSxnS8NVHhSqUVjqVgvvOzxoLhrIa
2cSe5XJWmC3cjixH+bWZG5S6aosmOAvvu6VKM8bgoxXphpQkHZ+VtiDepIb55+UI
0UevaK/ouCBFmiyCJw0UMy2Iacjr1PPg3m/MDSqj+GCGr1ke+rYTFXwhN9+CaA7p
3Fo+ZtuFNEx6yp14cEiB8qR/0FpZ3LhnE0WGJlgFp2f7CTVXQsfjF42ngYI/AKWz
GRI++wPVey1BBR7jAiDtkocEG2lqMGTWEd7T0XjUwGuGQVs75TW2E5A8PwmPqQ3I
q1QR/zz2YKdjzXXSxvA20i6XBF+AAfA8KqWLeRqnmA+pGzb6Dnx/U1iuFsE0TJCE
zF9oOqGhR+4gE800awzCfnWkRl9Aj6e79jJz/I4bNAso8WizAXBQEiAFIEaCC5R1
zmwLlrrJF75lFQ9UdtAgeRydpHJNTEHXmHj8svOHKptKdEdX/otCmkDWTXfxvXmu
3itl7iv8TWIeuKc9wlsItyQBJDkOBzK3f88g2BNTk++e7DjETN/QLXdLVQyGUI9v
CC1KJHtY5ygvw7+AE9LbsSYRciMheaHnzpUi/E5T+lCO1t0aj2ia3q0XvfwslfUG
RwIF+LwPP5o+9x0WAV6Q+RxNulcaLgwtG5HstZ25f5Aa/tSq/BEeJRg8TkjiZQDg
C51yOVxGI8qCW868keKYYlo7ZdETbSheKZhnItGc7dkRTrnkfar6vipyXYRc6jb2
dNJRtDolgXP+NjlsWmoMDb4060OVqd3izq8l3Xqt30WhGeWlMIwGr5KDfu5aScDR
sqK1tJj9LU/puhrwohZFJiRb2+zH3YIV99PL3qZNTBMFWvYsb3QSy8tkGeN8rEsn
HGbynhRAgeVWiFIHxHf5egvbpPK/THV1woZ8Z4NAWglDLjFWeXWYobl8hoIp8sfU
CoqCy3reUOGc6+2SHFKR010v9Wkc5bJU+C26P+R7i8kC9nJ1lo31nPAISgVu8eUi
/1aVoywcxelevsszKmvjsubN8mVwU81hJrvmrS5bC2FcfrqNyhAm9OyVRxSAj4lP
kdj3jf8G+3Ry4VRxv+eUs8VsYTsrRAhOTjxvG0pq9BRKRzvtOh872TmoRU7g3K6g
mk7JlOAHJkJX+TrPKZFT0+HndCuHH4eKGxCVj9REWOdvLq8llF9ls6FHv1aBqs15
QxubYPrV+hGF3OqTRj+gZXm9e3TmOLHRqRZ7qoQ5LLi6dEteDad3FOLY/g47PheI
lxaY4loznSbZUmTk83d7/wuoeZORnOzqQTSgSbz/WRKLP5dah7ORC553F4pjuEAc
Kw/Pt7dUl/SXwBXI1uelY2YQml6dwjYm7Oxw85xkccPvlgtmAL6FqG+nNK9XO4Xg
hSvtaaWSluAk+7++CBD1ypibk6mgEG3kc0Ip76IjlAslj9Z1rVOP+q4chVVZ8Z8+
Czpl+HyZ2IG1zyAzJi0Hiu6s+YQXR5JU3+tNMc7K0g+/U5X+2cwRIih6a22s7l65
0BKVBxOtGJJR3lLkJZG+57mWeNR0w8i20Eb+2KqKzoafuZXv4CB9qnZEASFu6Wne
AuptFnJoalzssOfXTCQioxwY977U9tBzTxoPPf2ZDOqOTeU+VVN2B9tUVcnCkXM3
s435eIeja+Ie8Zldha93VEkboi/iatZeXtO/V7x4U14BFxDvz4cgYUBhlKz/Q5ug
pDZu+0cRAAwdQ2WtwoXJWToyPpTLj4ses7cGgYd/FLcKIfSYWTKBOkhMo6rQWS8T
uMwPP6TxgFWLex3etG7yKIoN051mNk9Yc94Jad2L3/V40b/hMEKBIlmCmzEsk3nu
yLnyhsuSm5LdZL+u6pFv7MkdIdzTG16ojb5BhzGFIaXuD9lAsuQYgJrzogbcTwJg
V4SsvxSjiQqo9K7VrWmlyzURebspfE3lA5qFzBN1VqKvV0oPCaPh6QsG3njLDovg
AmAsLexH4GhO/XFcZnYUTdD7COvKZHM29ZKljL95vb2ykd+XaS2PLcx1sCFaCENM
9sMFdJuBk6pXgDn3U2VA9a7BH+VbGf3XFUal+IqShULHvsH+54bnnqpK6rIyy9za
5E2ExiiAa60ReJEfuhR/O+sF6f1kzfiaM+baX8iktm2uz52jDuzBGYfkjOgx7JGD
5m3AwErxPDVeQ/zjvV1JsilBJ2EOj5jMU9R6mduPglpOuVy/5IQGsCT1ZiRS4tlU
sLSMxzzlA+FyAlK99Ry9KXhEhgdCuKlX7MbZ+3ut3C7yHhM4F4iRhcoqKSOeB2aQ
2YLaxqrwTOPbfaoKlQxYRkog1/HCXyJdFaKN5M+bIKRCFj2iHw7qwIi0at/GyM3t
8SXdaBDCKHxQUMydQGluB0Cfe54xHoZ1X2y0auLGgaf+TNAOenQcsCgYols46/gF
QP5fh1YoXw2Z/klHoYLdFLwgmir0kYXtGi+ajgNm6C5XoPsw7U70Numz83dMMhNB
q5MwmL/1htxP/Uu0N3Iw35HjszoM4Re4/UeDpCucfzTMqha2jJR12ty8pueI97Pd
O9W/ahEJyEKo1TCHEOE5MHBn/AXEkoKOPwqzpsvaZgxcUYAmkRvKECc0xq9Kf6w4
6PxWXtX5ThUXdjT2h+e8VXaUnISIE2IFE2vbcipzPX2oq8GYo6k9UFgSN1jhHkYg
ErCJlR5nFsSxOGO9euCSKZJRVm7l13NxZGLgREHctdkk5Irmg+a9CseTXZT7nbpJ
rhYfZORoARl4L5P5C3yEXX2OzUemS7gObFJTnf6an7bvChlgnPyxfRtYdF0c2URJ
p5BZ8n7cnlOy66uFjzBGKaDaL/QoTVRabIv7M80Pf/hiOlPjCfSldOCTZfJaBuQK
Kvb091zgi7ybBVx5Iu8vvlE/Q7yvHnn1zoaqXO+3KdHPND3xOY5cKPBgkmDfY5Nh
/fo/PZ4S4zrsvm+yCg7ohGbO0tAXeK/CJJkFQ9ljbGKTnPN8EwcB1TN/iWRSgBvR
jj2fO8b2Lrtg6rV98D3uyVRbBGObjSh04snbCd7pU+RSPkjrPQe8UWK8PWBF0dwX
h61Nj7FQbteTwew20zJPQx2W4F+p0bCFEnC5gnfMgmI5+BaWuydPbZOFiO3dRrV/
b683rLO0OTGR6395xRvF5pDPltxK0EciCgAk9QEenT/eC4PxT01NcnrTCi9beW9z
BaBu5cHGtAnvqRUN1iElT6kUih2xm2calrfZyxdyiRNvBJL8nWWjhQ3jsw9oVBIw
gGoK8RgQlEgGawQCgPr7ghRdx1G28xFp4khLX4wMLwFd0vH6cGXYkflWpXVX5GXS
vfUw6+KHzYrWdwHAjGJkJfczAIHugs9Z+ObIktT0pJgeImYmyUSOvn2l4bEfO/0S
F3796uHEjW47vz6790ji45jenJTN74nW+3lPLjH1Om9jPK1AY42A8flLzdkqOUf+
vwAyRKHqojjQTzRSmr9XIJnY10dcuaMHBg8UjzbDpF9MAzK7tokuK6HKTaihuiuE
c+/Yjef0GQ4eMfilpJfVFw19NJ0GVP/vEXKZi/brkaLs+gKvMGfWZFAYJ5XwYxKT
TYIcMgIrRM6EpKliUNKf5061eUL2SGgzOLpThX9WOxetBHPezV/+9OUC9XNJhxwg
n3NUl+KUZNNReK53Us+RGuPHiCtPISlXynOtxjPGgr3jwmCv22qksF59pDcEgSfT
s+4pLeVoy+6I37ccYr/DeshVmVx9Inf10Dfak+t0hsD6v0t/E6sdeH0hDeSxYkBA
NKuhhugL4GGKz4jlz/oeKsifPUjdUVYIWqnM9sGcATKbU/FNdNWzb/miDcRzDfdp
QLH9j6Kol7Z08EuGUqGc8UYAIqYeEy3Zj6XGob17oJ0uLujTlVyTxD+WB3fUI1PH
rqhixTXEa3JkdWlBp8IQHAouJHzKMnIv8viwsDhVKg3C/p0YCDUUKooLmTEJymhz
nQFoqbj5xLU+AWojO4MsQAfir5fk5C5BaF0hPsmiEV4COsToLhsRfd0z778iErR5
jSt8MIexmZD/ldqRkQnBerg3OcIYcNZ1axqHRL5eft1De7TdUmApnLTniN2z5Zbb
0B46074fztWV4x5cQpCjZwUQcZ9tl5350oHx2luO8RmOqQwQMyotGcDbOI0Jo0tw
/QVt6NWlEyNn+MdVHWuQjNQQbjuyuJXEtnA2OXNtFXbkOg/Q+joH69P1vdRQ2dKi
8n22XKjAzegdI3HmDnF2HsodvTacfJ+0+KciPl4hQI14acz/pdLBHjP7HTWaEDD2
tTlISRK9eWGw23cgxODZmp310H/BgVhZ/2LoJo+bJrWLNe/HZOuM4gYcw8OkqhEE
6Zga3TCdkGmcW+LEWfKz5t9wCjvOJ/Xai599QNKW/OHsSix3C9AwemTLiiOZHXb5
7ecAZo4p8BujJMFEHjirzRIgDoOFsRznQ6cQaFhe+aqbaC2veGSNJbNHrlUMyjws
hi79TrByNw+6Za891cNEnq896/Y/BDfqghJd+q97U2XVni1d3LfkU7lA926kP+3N
8xBZOTy+vrr5SVStGcH5JjbRVP9ICQl8SWO1wlvb4mLfKkBnrp9eRqWCosJT4pgU
f0dC1JeIQnIkW7k8pTtXs1lb52iOuRQRFOcfiGnMd700QJQLvptK7eGFGg/vxhpU
+rc4GBDNounmsMqcHpQ2ShxcT5mNWfQejZiXlhPHTWZBT264EG3tqg3Pg1QHfaTm
QMG0U3/1mQeP7e4mzGicRC/PfI5WVI7LeN8w8iAop1YPn6HM82i8sEwRE9rrh1Jz
CtIm3Ew/FZJno7li6NrEh2Mf9jn6epZyEuWB73uHiiPqizJ3b2Rd/JDQ7DqcLB4j
X239fZWIfoB6IgJCA1JX+QvOhc+30wPhAs2JLnTni61U9jLyxFwyaDwxg1zzkdEk
SXrPyhwd+wXs6fnYDhzq6V02XIJ0/JfdknM4n/YUmzOxHU7a1lxnvTR7D6RM0sht
77CUUEy6lOeWrqalL+gDTcsY7/lXIB2QAgRBDxO6upVV5wQTdJCKgQM5GQpIBWps
YnImCqHW2I+EZW5fbkbz9ccrdABIlk3fef4LqOmupxZkus1D+9Aol1vCIDlWcd3Y
OKNXfEGV7r0V0jyPMCdwPJ5Vb5w6pX13fBUMvQA+lvVtHqSKsAY5TaFnq4C4uiTW
aIxcsvKUBZgUQV7YHMvJzLk+VXN3DGTdRZyEEzFfBoLZ/j1DPvDmub5F60JL9Yar
xpeSXCUorfbDCMA3WsyTKDfyD6df6Jg+mu6AefNPoAmP/HhD/nnjL8qcaKUC4sUh
Aw8cd/rTJzDq7Y8BepGq2s0HyJyPG8ChbZZa//EuC6NY42yg0XiifioQa3pBXrvW
ESMSjkhUWx0utvTDiZW8k4xALvU1bo3JXGk5fCR/vwOESvnqIOHDRSLEO7l5+UrE
xLN3D4H7nxyLp0MMbTPjH/jDNNcPLfseQFk+Gjh0+3BeyVUJqOOxSQswvbk8O1qz
hcAIx8+KqnQ6HzIa/OaSzT5+gUSz+2iYeiEY81zuQCewdJBXCb/VNYA4g7/E/+Lw
F5PEbsPwxPjJAluuS7808tKHXDqZVYkSarZBJGgKH9PB/qNUNIk83UfbR0+GMxpS
tqd7YAskyD5gIL58r/mJ0I6rn6qNweDtS9kGGaZlfQnS++T7VUzx02gdM7CxGXKn
yoW8XOgLDwngCqjUXjR8WCXmJOqLVEJCTiyxhHudewUpx6ix7X/W5DEjbqxvBhq/
6fIuch51G5xq/2L46dHnGg6ymHMb4GYYDpgjrBMxRWqf2GQkfrprFAXDpTMtBFVQ
bU8nwxwOAmpn6njH6U0I4MSy7+W/QKoEJ/Oqncp8EPw2jIisycZFwT1a4o59LQjW
JT83kJTgD3TSxuzJoRbO7LweAJuOgfKlE95ZZ6+ewOZKjjnf+HyfLKvnJ7udId1A
oUiXNjXRn7XXuVi+HqlQYuNsGfi0AH25jA98vbT4eoiZr8aBgPnZKg/5N+yCquCf
x06AiKRNpti8b7QBwdKSpQJp1v5wF8khbyRxrqNZ28LGT/qXg+23glXheWPm7oIG
3gn/PvrawKYl0CL/lmAALY6JfbOh/cciBOuzFgE1jUXh0TTvujYXX+LiN/qDSmnz
rFIh7h72MuqQCgP69QeK66OkswWZnj2eQss0Qt128wmt04Aj9MXOXdiNTXc/r006
Y8sfokVCKnVRi2NLj81pzNAxxMbRc3WXAXrRnvHLeIfatf8fikwYbjOWvk2JRkgD
wupFgBtj7i2bDicV1p9d5zPf46XBBeGad3Yaphjw5vtfyPmvIss4Idtkpk5UV0Se
F+JuYa4EE4lrx4BYE1bc/+L9UpKPXMMAcFV5pddUHd6K5HEvrzTBeaSVKZeSKKHz
obRpikCcpylKQd3gsMB+XWd2zVi+MyVz+Qkf15ksQPU3rLbSqEO4Qq8uAqliWa2P
Oxaqo6LC1KJlteOEAQJOHqb9lmXramHMfThvMrlRW4Afj9GuOJkwtprCOner7ZEl
LzN+avD4rrBtYvQX6Qhh89SD/T/JPoMG2+kGeO/2nT3LM37oP0b6Y24DRl82fXUB
30LhyTz5eS97RWY+1dk8qAptmdC3psDkCkQYB08b16PiReZmw7R0N6+vwbHShiJC
1vPfarA9m+hbnu9neYoLEM7BJ9irlkU54iscH5nGtzQhIpWmqVbZuJEuDyR42crQ
InlkpjiSqO/K/zt/o4ZbpsdnwAFu0r1xXPw3cvMOBB/1uLbNJK8f+N4xD7kbnM/X
oFDNvn5/yGx3pkl6EJJzoS2/PT/2TWOxNwusLN7MJmeTTvSdkxszNq4zE2fErk3o
DJpIAqWMmsieTtkWuA2FePANp0yjUwp4ZMXfLnpOyvEioZOeX/VSBNUBvP3j/yGz
6e1GlIgchVhFqL8mXCDIFjuVQk1Z6J9rBCP0MgsAT6Ohto6v2TfORWp8SHSeadt1
Cdk3zU4QXGXmaEDs5PxZEMpim8sDSk3jjga43NmK1Byrk6KTClHLgE5K0hSXnACS
9fRdF0OSjS9VWfF174Mkp+3i2PAkQ1LXLhUzlYnU2PBqkqPguXsL6sP2jOeWSfp7
B4ip7cZLyDz0zohEp2J7XVSVFVvlfpVeFHYi97kdTQWSvKvsFk8VIQ3oSDMWAj/v
a/SWcdrAxee+ZVPh/w47ZYn2O0Qf4ECT4D160RZC0gUp9apQEmpBo7zfrGb8b9SS
fpd9R8v/SQfI3v+pAhLkbE9BkfiOadZkF1CU9XYuSDLls6MsrA2CMxPgsxriqrn9
m8hyxtJrQiI4viUplAd+Jnh0Ro/G5J7rxZ8p0e5vhf/7CH6kepDAI4lgyR8+hj1X
uq4KsvWELdQUG1F4VttTAt+35PIwn1dDobFpOTrp0QZJZ6SQBqGvibXcpdyt2gyw
WPS6JkJpJ0IR+g8j4gr4sTLx9ChSpeAcndPV3W/MRRSc2VSs36KIeth5TPu95DtA
uqPOK2LL2hGnakc4QGfprUCTxVf13Niai2D5Y1qDfvwiIJiRBbuTo5ZK8sMfjZ8F
66hZWiDF4TbZjXl74ACu2jM6NkejWvgQjBokr1RY+o37uFnBQRk/AHCEk2laSyVS
kfIr6shfVNDiVtqpKB3dDzMA57ljcXS0kUOYoxOpA9QfmGy5TRZ/+nWinATdws8m
sR09kRSjZsL7+MMS7lS5ZXbqxIQ25qzU+51B7E9U9rryA63MLEks2TFYBP5+vxd5
6RCI8O0L61yMoubY6CIQhhkCPw2jSWkA10g1+Cd6HUPqDfmC5glMPByEwGxqSEAv
vMHnwupi8YHfyqz9MPmsZzHf5uIFDZO6tX8F8eUUDLiAeSUFg/zYKssdAiLYFqRS
3n4SDMdnTIzVVZnTKM9c7GK5yFaI/vHHE3wTu372bnUakFm0uzDcaoiAf/g6d7x5
DTEhy1aFDe/c3IAzqap2xwjXvdR1B6TFPqe/GDZcq39mm669gcNvDTdHnJHgOWWk
jQ0e5IWbfeO7IFxJ/sLJDyD1wP7B5mXTlqJgp+CoMd3Wh7hIwvhkzDZPwHmf+Zgb
0LfkFgxTQZlhaurf33RO2C2yipFAssJRgcjkESTwuXu+XyiG7N3RBILdSTUkDLS5
MAOtOCk1k19gQX+u/SPzBjJS9pRy/T7gDU3UIHx1CP10X3aSn4YcSu9rhcoVqg01
Mh9c2PQAA2GQguVDNDrwqHzMFQxkY+4VCZqADqpuEhr9iX/Du/M60o1Sd1bCE4u8
ujFOP33RWB4v14kPM7SbCmJ/cTAdZrHQQbmW9qwevKmw78EaOljSPB6WIwbMD1G0
zpp1ozQIYvpO104e/eOP0JDwdlPQXeh6WA8V04V6CZte/QaSy7luIaGgVmVlkM8B
IEFKcDzb09W5qhUT1Defsd13jMxXvHs+8cbIInoZRGL9jS5tOv4zqPdUpMlnqZT5
HUv8EWETrwcXRdtSHYQxLew+EWSx27N0XZWxxCL/GRzrDqXFyEoEREkLaPTjFF/Y
X1HcWESxufipU/y/f3CgHIBPvPdzJA7Q/cBI5Z6jkj5CSZl+EFGouI5kWdqHz/Dp
gu5mW1O8YS0a+L/unIrBbI2yxkIvzTIYPiVamAywSOGEhXptmuS0HupEMDi2bzG3
Oxs6QgGUSx4afYf/Hvgcs6AGooGkNUTCW/5E8PMH3w1JH/80zmpYMp7RuwAglKgA
oS31psyb/T4i1IjbG1YVSxBMV1N74iucbQ1brmnfCpgiLH4a77feb/CQYRajx1tK
EmLJ8YGd9JrLPiIG0EGdT9sXqaIioerEu2RTewgrnuuXh88crxGVZOinB+9nY0xO
hTL7fk7rYUZad7E6wdrwOpYYCXx2lGPeoZXpQifxfVRtdNSrJHh2EE5jFfiSiyWG
qQ8Xj3v4+QQm4GGEjI6hS3VtQHJY0ulA9ZGpzsFVzWyjI4jeSJgvO+JMiKo6T3dx
yv5+xu4DlOXZOpMv0rloyNoQT5UjrK3EG7QNaseCOukYLTIMZ6lPcVgbLzZzSFV2
hTD+rkUiFkhY1qmcowrCGnuY96PZvMY41eha79nHpk3iZJLqPupeUPBDd+0/C6Pc
GNQyielnq0FiqxICSf2yqflebNaJX0zya+osk6GA8Bd2rxOYh9UyIaztr1VTXtmM
QiRJdZc1Us34EkKlWyEHnAMPdxnkG5LKdANgbedyNHlt2Ld6D/vp2DLhvp5Kj03R
+NcCXCNwFTYuFKGBfk+zKFYBrD9XLUapNx1JjNyRe8jKwWhFLZrI7kOsAnkO787G
BUOubcLO5j9Arp5y6ntGO8zolKSZ3DOajjr+DxDtB32u+X8h/1DE5LbgLCzXIiBW
SuTyCP7Y+RkEtzjS/ENSYRdUH6UP4SwAmDDh+xnqj/NW6lbboZcQtPLHUJgjEt7X
Z1OCLuYuVbswxpLB+TuwNmlAOJvvfmz69coxgCrkngmFXQZ1FTTRId2hUBxjoTau
crXXjjBhyWfcZzQtporW5dZFumzR6YKsJga7QzM8z/K8XPaCpEyH0XpB2wULEaf3
cf3nHwcQ7sEh8DKadnmRv3r3/oCnEIkg9b/QwHdtNomMF3Y5Xa6+g9WJZqYsSk26
G/04l1CezjUppxL2PF+6yR01cYBYXFeXM+SYVLY9su32chxE4foa5oSQhF5lD0RC
ZhPajPkhWvfMEcC/aOZSL2RxMRD12L5jnDcgvxi/GWsYWi0idmuGfMi5d8FeHVxl
IREQJkRG3Y1N/zoi8y6vQY/r5mPwM0nPhe5+zzLxL3g6Fo73xFTBfpnY3fLhsSrY
9cIMiq6kvLekTfqkehjJ7Hg76goLpiAsMPilnCYfKBrI+1/ERjxFtf6nM+LeMqRd
kBDt8+2ze27KHPDU8QSgAsOcnt3qgMNFm2dqUIAopPbXDvlWXYtOO3JgEQvNuIzf
0KqzhVbPra7MJ6RndgTNVymuLa438l9IWgIUYKTicOC9UezdWFwFCZQPVcXMKSi3
KZop5Tluy0L4zO9kRzDo0HAMjl8k4ATtf2sntO3JfhWN8+hD5KrgOtGpnxW801Q5
z4SmOAfLOC7AwZaVrp+ZNZWBmV+NfZPlvyc88BM3M7SaVKAHTHEDRjfNz6PuoaQR
KU3FukiaFW2cNPQ649djV+D2JtGgFzxTCAMzEDmfJOQAoH0Gbd4FMv1IgUSsNqau
+Rxk+bFoK0FiqG59wDAg8zOw/HEMMQI4NPpbXqCMSy0gAeCpNxnhbddSQfnOYspX
v9qRRfaius8r2h5zRgiZNBBcBE9KUdafDvyX49HXtI4Hnf/pYWbnw1cH59klNDNx
xit4NC90/csEHq1xOUfeP4p2x2lEDwdWArCNjn1r+ga/Mg79C84CxRIAClz48jT0
6y/aX/NdqnlstZwEZQ/dk9YbOejFjZCS2U+Q0ke7vHjVF5si2cH14/4DG88Z0XRJ
R/IbNahZhn9mu242qsCx8MED0Q6MtFhKRBrF0mJdr67aYOydMetF1nStfTksja8u
KKiWse6fgBb+c+rURxitG/kGPvK3doiT8w5FEzlfzOXFctImuk39Ip1FCppMQL51
tbr2AUTkOsBbRQMaxjbatAO/qcNfUd/ktLi0qor9VLwInoG7D5pY4XVYg/X0pQRa
BM/aVcOaaAX0AsYVcMRkEnypKQsV71HEp/hVRNuo0Ye7nRWOlB+9h7sADqYSpB5h
erJi6UHCsbd++NR57hLOrSzE1ECDWG1znMrPVuNSWrXjM2mEseDPu7DejHgE/Lsi
+EiUypCu7DQj99JLA88dmm8AZ8K2w7m+sQzccp9KWwVz8Wim50CpM9/Z3uLXI+r3
gZ171++iJlo6crn/F+a/P1BaAO87ZsqR5vZebPADBllRiVeNlAmBm0y3btTrm5Sb
p4YZ6jaWcjjBv+BIPoHXPRKqj5Bel5dG/mm86CNl4QXO4SS403wEkbENHx78++gD
kSEcrBIR07STTlHbCCM6PWiJ2ZKac5cgvKARPJr3Wc/TMDxzrqfWV8YtzT5eIKRr
F+ppf8YMttIgxuWzryCQ2c558QwdmAsFLr9Efr/NX2YM7Ex/HWENxuLgQX4uzCjA
R4X5qzkPZ2qpYh+3gr1wpZ5QM9vw8J7NitpgQyP1i7/n2Lo0qCp0r15jwecfiUsm
eZoUqlJo/TI2Zp5gG6F3xb3EAdXbCkC6AuhRuAOwOg5Z2T0h+CoBlVJjOxb1M+cU
2xurZj63L97Yq3MG4R1WuZ5ZyvfkKRlLCzI0uNjmTdFn/V7/s0rupPRklrVhjmW/
5I/lJiZUTEMXVr+fqyW89vTxYikcqNT/NyqXR9T62eaCzWytDSpG87euXdr1KzQU
BCAu17cDW8OI/8lJrNRNNiDjbxtEzwjY40+/bSI8tyoUAAS5GH7ZwPf3k9htg+pI
O7PMPqFYvuNrvxD7NDAAYwVtuzdRJS3oloi9NqyDy8ZpRQoC3zcE3U4XPWGUT+Nc
V1NV7MUxE8ogPOO9p1COpA2SLpjGMT1EH25VxgPYyUKMNwOKa76P1m3wfDkUh4Xg
R00hG40fUSMtuH1FzxkcsRBjDrasowijADIBgKcBq7plSDjnPiqT4RpRBrUpMW71
KCubMfmq4nfgkV/T/5TfhfjZcBTcFdgUeDFAs4s84JkQLRrrmPhX63iAPdTAwR4F
hUePp9vLBUdKGox5yaHDTJk201pnwxVLAJJo4dV01RZC/bxsTwzaHCmB2pkMq6Th
X9eljz58rOXS+JW0q496B/t3TiBornlCbQr6+Aqth6x52Qf8VgBOJGuKKAr4e9Vh
DXIQoFstIC59ggfrvF/5VEKCkordh2gEhnsDsiEjzW65EAQO3vBHBgebIXhdQUjJ
cNf27AGM92ki4r0Tkm67AbzyavnTD/jOMtFWVQ4Pktvoo8xhe6HRhdGqzV6uCPRt
Y2X0mVIJKAlTxJ3JP9d5qYRGUqYeLVMvkd8fN/HkUdLKQZeFI1lz8E8i6vDZ9SRc
9I5WBpiqRTASPwCXNTyAb5ERkj7nA2efwsgyr/Dxe/lId9/cC/cZE28wc00z1MP4
hfpvSAyrPzO7J6DHc/4n6VCCSPSn+VGC6fNAvI7K4+BjCVl/DyUFxLgjZ45rTLoe
d89OAeOGQeKZbLVlzpJCPW51aAqgQagLAGwPoOpeKB9cvKUZ6vCwxtq9cEU5WiYY
1BMtNBmAnWQ0+T5AX548ormbwONk4x3X46U+rgXfq2ZfdzqZeDkTL4Oqz3Kx0e67
ja1yPT4i+lUr9g6ymuVddGbkNhkCtUMUal7Ohf9O6S/8JPjdvrYuBdEStj24x3h/
sFvEWPR/+M2Vf4J60bTRC58HpKiz9TLic9hzeRWCnxTt+a6rjEPGxXnc++bOJasO
6cyFSLit8cuYi0ICQX14BbkubeVmefX1DxW2Jg76BQcSWWugOJUd2lxCpv9JS/xe
ki5H0Vu+5PBH9k57y/2FYTpJd8xn5yozkfq0qLPjzUShIyxVS3a9AYoPT2jiGpjD
W68CRENbMFXUAd4uz4sDgBGu0HX/Ld19tqx0S59Y8n7/uoIR2BFRGddvYhqn/FyU
nOdNuM4FcP4FpSkFNlNw6m93yrq5u/+oG4Aw3blOR0/FGRqzxuWTpiLUYjMJqNC0
nOXz/HOMoT/UfEO72muze/DDVUZWrh7+mrpz9zTLEuaL99QzRwBEFG2vvKWVnVaM
/N2YrFd//rrV7GW2jPLgqDgkCAp2oT+RYjytZacgVwjf6NgfLX+b4AGHUuQvBXs5
q5KtmM38esUui7JBfIcOVWuvh+jliVG0dA//crGje+EKJ1IssSbJEpA6SKPK44KD
VYXYKXt74BLEd1E+UUlwRxfMF/ehiYnfv45bdPTwYyfqj5+EGwNnymvlgM3up3P3
+1wUy9zw6DgID7YN1djGSzbbv0jsOZtrQfv+Rf8EtKrwDO3e06q4JKcpWROGoQiL
TWWXl5Sdu9G4kCiH4TjHWRlnx1hKQ/dDgKmA+oX0fI7PmBAjh7K0uRYE3k3XXVmM
wS/QDwjiyStQtEhbqc5XCS9HZ/5IbXX6fClj6rYye1OIvbMojMXKl7xafDaJ/s97
Xrsxaxhw8NM230OQ7IkySRthd2RcwR+L3vCEekKm5nuQHS4qXUF1ydHqMOo+FrYL
qPTmhsdeR78oY6TS00TEO51q93SobtHWPfV4fdFgVo8UmLJApERSnfYfD8Dkfaj1
Knriy7bPf/W2paRkJpJqjsixJrvJ6q0N2TPeczrtzAjpFlutVodXzMAvxJ57R91Y
ergcwSWfmZYrkwC0F4C/j350QhOxKf72ehEmpc2H7yuPctpwjwZkuYRc+2AB+fq4
6j1WpfZFi4973QbNTOXtb5Ioiy7GtzoluUDcl/rSWtXfzasyr72BYvRK00HDMjpM
i6b8/qZXxPLobBuSABhgAXRALXoeV9m0dvLWciq4GKDGEQEI/hG15oTrU9FXGbjN
nRgByOwGOxDEvSi2rytruca2MsgsJXsS696fiLBQnNlfz2L74zeqg2Cyc5meXW2L
n6D4WQnjKGTm5w9O0DtvP+eXfds6BDkSE9xhFoJhJDUB4/GmbMPb23hte8Cbq//G
nuYeiu6kRmNopaIb++rwh+P/d2GTnqlK3fTlvZLFhT08LHydqG2nOgDjMNKZza7a
YMnSyal2QI/EjuFdOxhexbTpZb4ZkZ2293HEfkhiTk25xBu3ykpdjQ29oA5cT7Op
59Xnfg/1J73c5JiC+6VAoCs5vnfO7LM1Oes1JUL52ieZI0bzoj2crgYrnSkOWQV0
+ktyr0/7G4jO7vag9PyWrZcGo1fzD2zTvvNDQYhP++YUoCU4SCiQZPlkuf2Y5vbi
WDCvoJVKSmuvUqLXNpL1iHbvupFx9V+y+iOmgZYFwCCXlt8jXCRek08JO1WAHbGM
orHlT/wPbbzr4vSE1VVTseThXAzE8BwPLhFUTe/tCjhoCw0QBDhMVVkR9rm1PCDx
0dL0dwr7BRX7DLDGWgCKYJksGISXlwsi62M12N5b3k9Wqe21S68WtegmUA1Q2gug
cFhJWhwpmJsS/8RgViMoiIZ2N6c0xFuaXfWuDoBw1spU4vQXH1KSWu7TlcfL9Ark
QBNWZoJXzXdamPKANAEbdCuXNOMiMluol+rkOfqEMZmByUZmq+O+J1gpRh3ifR/e
UTvB5lsLW0dSUKar4i4FTp+3HNAWuNX2T4V1vmWtIGEfW2LqT+gYcEgdXBdRjTaf
lmhtd7+Wjb1oJnPJWyCHzd905Dw9B/PMfXBuDUWZ/BLrUMMCgcMZGcbVWO1LmVfx
Nso/Y0rPnvq6RpXEPoB6oettuGkYlOO1p/jl/RP5fBEXIeWl6jT7P9I9XwLKioXw
6zSRncaltrQZiPM7RkWLzW9QhzzDzL40wDmx0Bw8vNLor4bbsAsBVxEmVvE4IjcW
JgLlWnvTH2UOyht24BAJ8d+mqHhcCpu4FS3G+/231vVR7arpZZx6SzZHoTTbXZEC
kpiO19BO0++irGnIawBoP/HdY/f/9/QUqtHA5lEHgPPRd12v1kxwi4EViDFC+1nQ
l12uqPZCee/yxIa+lzFIzPGJeT0g8itdzMOlWqw5ydkxQBRqAq/4yS1DFzigOcN8
+5ncNCmTgKmi8wPNfJfi16XLdbgRjWI3Mn1dBfRxHCGRMq/UYf8FiswsHZRHU3rm
3+xx/PVfqHfdqBYGt+rg8UbZub77MSxZjwg3vOvc20QWDYTnHCxsN60wi4UAxrSg
u7oesTgZpLgQjREBOxbczjPe/gmHzn/DVY91pzpyizP2+3c4Q7PNPNVYUFS+dcE2
fyQm08YpxmffkULYZmk251PjZVPLGoHZVak124qwASiuNnjSulC9ywDQSlvQdNnH
otY3ynnLNPHdS6qAGFZFXD8fsQIigPK4md+iBf+E+NzdR00NX6a17Jc7dSzUDsNO
dMnlkr+R5aBL5BtI96dC8SufrHEUWKdx8drGJ5LnbSajBqHDs9cEJLFM+hC/6nwf
RFMttQtl9tu2UyU9CJ7kuzjMG4DMOcHeKJu+MsF42vrJ0Ac0m0B4r35cJ2p26l76
nGIvCv7lD1WTdoButTSX35DeM/wraQwj4AaL1HK2vHthcjvH/h3dQzfzya+dojaq
oU9M63vUWTEPv3vHDLNGgmulsYBem4ki0jMAc3tJsK5Hlrvxy9joGUtEF7rM1BrY
CYKNRgBonA7Eyxad4haio79bO2HVyB+wzyd22vLAJUyV+AkwzwoDx1ESVDrnbSc1
Z6wE1FMaSHmE6wGJ3VdMa0ARE9fW8muRGTzMnEeNNewY5ti8H9nvCDVvQVeSZmPE
0NYfuobk/zdUw6FDNhiDJlEXnEGzlNMj1YwnS08LjQuRDDDVmuZ1oJbf65NtxbZ8
O/hTI/FdaHBZjAK58MHXY2pEs9zlmaNYe5iuie3bzSjh3gqQGibxHZHV8Fh55dXE
uF0l7SysCztzFc3jGHVe/idXzJLvcNWQpKP0BZf4MJOkFN8+i9Ps0JTlaPkrNHWf
G2e48Zpov+RRe0Kc3kHp8bxL/zt+e7kTpE175ZBu1/rKJasyYejBMjFxLnL2eL2Q
YY6bFMs8jDbpVQxmFb4KsDAWcPytg5ZIwzyWNif4kEHdss20GZsn46u/5ZbHtKOS
4YLPmGccn0ATWLZkM1d+yeSqhcUzmUuy5yLeXFkd+U71iL2yL9M3isbEsuwAiT73
x4GIVRIkBeJfgM1BV0LGLuksD/N2D0Xi9tMr5FKpi5tLWaSJzBNzL7K/tOEO5SGX
5EOxp/NsXEtXLb+CzZ0Mjat+aE2LcI1P4NOiIYI+fz5BA53IDTeUg1jSgw5p586O
PLr5dOFnntsGsUp12FXP4zJ2pIXXWtoS2UCzaaXVCApE9nKpiY+lPsD4O7BufvJK
rbJjz5+a37K8K6cOaoM7/+TLVuGkt5V77tXKP9juyCyedW+drIov38htsiVPP/O8
tircfWNSV78FfmU/4JMWYobSYw7sp4cIka/FJdWb1wUcAPJWeKJ87uqgbemdTsRf
+VHAy5lwUpzF/NbpBvcN1cAx3xX2eQUAhzAinQ9R9nZ1R/j+Ciw5KGYgzYAMO4GU
kIZQ/FyWa1eXQF/ty+V7XgtaHHNfotMJrISY4Bz1YgqXE2pLso5qQ1C+W+JpGnp+
i6WThpwf76IOjo/t4xOn9lV+ve6oBoPAmImh9KuTGZElxM1NEOSJuaW+kcTmJSGv
4015ni/oLvqBJw2KatR1Q4h/VRrKspw8ZA7GQL13h2P7LalZOLbGB4uvYCUXlryV
12hfJ8sYZBJV0JE+3ECnM5WlrHbzqDe33uv+TReILp/o08SJNVv/847vUoNw6+w8
v0k5SUh37o2sPPI7TtC3CnopxPHgBNkVIZl6wG1G3GENSpoYaCmhVQqspS96Dk29
nMxjBd53KxnhAFCso+1TFcmlUstIJpoYL4429brOb4W/WrViQ6Vpb4Kj2SU2l3Kh
PChcsXYIbCXV1l4gK0q0SxuA4WpczT1bzEYkU9tGKgvDiR5jOEl4HuiCsJdSi0Zz
mZfePpz95co6E+UVmQSvyZpK9Z73sJV46QEHFGkzQCNFPlkMUvmc7gYT21Xxlw2B
s0OG6HBGgreh4wWUceltqP5WUSFN22vn2weHtjlFNpmorD7ZvodfY9EMo8uq4+vF
NCs0xO+r932390T0EJwHiIIhF+rQDJZhK9yA9TeDcrDyUmQx21PxAz9gLRG5kyH4
ufKIOIPQO2BnB1R9H6uDxCPw0/t08/Fwzh3nHTakqccx7LJGXwGL+oNc9uh1tiRY
+JYYkqbT0lvd02gwCOXiaZOmjmd08j+rrIVupP5W4VRsorsOnwE0Zo4WMJCINleZ
I6ntLIb+l19Il0FraqOctP5H2OBoymKcl7Tm5m2ymVFKtmYWUMEuHLGwUJ1zoXU3
M3iW+AnxlXF9TrDqxNaxyCoesb3Apx3t8Oejv5E9od0xLwC677sepBRB8j9uCWNO
3G6Pq8u/T9YxoaQdI+GOS83LBdv7MABDoCsBvDuZCAbTMMn39C3/7qmeSIKRkXxG
zHAUxjurnTqrNN/PqJHURKYBLN8ytM24w+LEDrLtWHyJW0RqrKc8FqIChk0IUecM
HsQXgfyl4Z8grnmr+ch00LDdZDSBpN3mlWOd+1I8EH7Cl3zb79LMEhys4FecEkyv
mhbjC9lqgmSA1goj467p2/TTAu0Kja7SJ26S2EZnvYTKpIHO+wbevk80+rhhzeM2
wxKPdSjRroXbahZq90ICJVFx5yeJgfl+waID3+vq6rwgDLvJPl1XrPBGLXNiY74Z
zF6IKu4FXWqFegWdQtAdhh28GHmr1pyAki78NfyXqXGKjGfApZTs5Y/0fuAhqnfa
HCJ5p90tgpMOKtp6+YnXAIOkt5MGDOiUBWwZfgFCd5pN39MxJuQiJBWfFN8G8r7y
LRi/Nf03zyLjGd9jgBVj0TQmpo4xjOeeuzlrxP+mVGXJxv6ZFEt51nTvzhTN6RPn
r6PDkjbHxs6+y/tkUY1dvAv2Io2CVBHL7a5GzPt3wkG9yuk1PXNK1OKWSihQ1hWn
2nQXBnqKAJoVr2JCgiqoMhbJlLH6fd33xJqnXg9S351eX9rSkUaSxubcvnOo0Xu+
qB6Pma2EDsMVkhxjVsqYd8mIOD5uY2z8tVQWYLmWOLrmGllcLZVgj4o2tdlt7XcI
hhv0PI0P2J5SzW9Zb2Uz2X1t1c8ZMLNlh7OnsMusoBsDY1eJVLi1ofBZfyrL4Daf
zeBAoWy5c7VdeZScVvIWP3xyuPbAviJB5PV/g3dSZEPvTdF2HVD+/1JnCnI0Ng1r
3aHXWEs3+mmFzF0bZFjykXF3qFZnHeWfnkrRyJymWqvWFAfLP3w/Gxeau23sgiGa
DxtZyNsnwArpnvG4icmL86S5J8ZBdtrbbhN9zCNMX8qT5+IY+Wi0XSnJetzMI+q2
hu/FiEqstRojTHyjfp/a4/LSbV9RQS61PyOg6c4zQNBwzgMo7iSo3zbTvLlctvuN
8a0rMVYr+GBEO2b1wlvDKcMluWJjZAyH9ry1cfUhz8VEQ+F5kVBjKZFODTzOUXmH
v66vz+2AL4GNliTcU+P+6E3p2Mr0YEpfVSfPCIeNVlNYfbjg5BcuzwSQOFtqkdpx
jftVLDAa+N9EJjgnZI36yd8EXmUm7WvqsT/k4EgfS3GDr95o4AICacH9RlAyXm5n
PXh9QrARTLk2o+Raf/PRLaeosSJI+jkw+R/TYxFxjnh4w0mRNFpNURyHi4xXRTt7
cKYt94xBZFGniT8dRIaRMOFi0CZS98ZLiIVa4kbRmVR7bbwPDZn6RW6lUIspijkN
U/LAuICb2Jq/dXZVU5bGiArx3X7ywJ5GyoFbqMHMLUxcdP3uvqqIlU+7dPi9Rn7m
bMxwAtSGRtVcEmsIsbho2JycwzlKQLPaq4LZ5GE7S/FrFcm/3ED0FiaNmI1nfob+
gd50h4uD/DC8VpB0MYdBm+Mll3AFQjSeRp1NSMgWjQINkt1Nw2x77DPaa6lkQBe2
/CFK1TbwZVaFGiThhAITf53bNdBgvbQcHHI+R6VOYKWYWiolArAhuyR1aWUQp+NQ
cGDkgvxkp4oIuyUVnihXQAH3VZjhbnypjGkMEwLHTj7WnSDoscljLMEXRnxmD1x4
lrX4LiSsrdPr4fxJPxKFWBK2Bp8D1zKyxt30CGtseIzojqrAppVB005rZ6pLAxXw
uhufsl5lR9bJjbReB73VRT2Ug/xdGV42frsKd9yabOlQNUnaJugd0/xLSB4PwqUu
SmiVnvA01flqEwPgHXheiPoTZcgzIR7/UgZOC7HvDtiIBvO3c2HnjUlSbKM3y446
l1aK4Gz5A/eCMbQaWkqtlk3nWeOo5CgJCrKAM0LHAQQjOTmwHwo2CPmPfg26lqWg
vqc30FP3mF0ynsSYGZXq1WUDMi3eUrUN9qy0RUMxEl795adROKxpa3f0UHAJvHrl
D1ZEp+mRwWg7pZSBqCD5BnD5u5Qxbi3YF1PFFAuKnQEy6AAkRqAK1V7AwA2XC6OD
9GEc/iJCujCn5gsxHgTxL5fgQJLF2Xhc1jAVfRTOqFt7G4Bv2w5HlPDLxAzvF2SY
F2T4HSt5MarMOHmO3HK6eF7jibtAsW4ZW0EZnEujd4Kp+AqxexsZlgAWXOAiRvgx
1YvIcnl2KaBM1pUCVH9gN6tCM5rrnK5IZDElOBpQJttcB0JlpsgIDAoaP8J5M/CM
KzYqtXq4t1vO8+nrVi2cuOcgQNvH7beEBM+0xmRiVIwZxmV9qFq6cmsNg3ceo2kF
LEEPih0v5mosnf1wzQBgAhx4fnActdMzMLp/vYl2JeGC5eoMEC4t7zcNYq5M6MdJ
S8vZW9Yzy2sQjgVQrkwXX2ckgBbyRLtDEJiChaJi7FdzOcTOtlerwW+FH9Qihbk0
aJTamN2+IXHAeDqZzyZEAhlJnQMD8W+9BRq+ZjITRMDwkmYlVNEriBN+W3Av/juu
xc85GM+SRtd4rAa88yHl2NKPoF2I822yuGuililkQ4ifp4iw0LZGYBRil3ZR1p93
uyrzRxRNgNiuWZmlkY7oxZ6ult3Bstc2orD7/8wiOdL3LiOjZNyEPgiGF0sCWOTq
+yP4iZEK4rcY7hr02dqnH6AXtsVs57er5t/7+CGLXb1Vqef5MDsY0l6Hoedk2pHF
CNxhv1INfIiadSDV8H/zW8/rDouhtDzlKVfYWspvN38MS0CCwSByg+DO0Sejfcwb
MpZA+ntQYuA/n1Y5kSjaeNwtQDaX98/u0FM0kJS6s0uQQWVIblPowykogKvLJ4BT
Y0PQpnpxlzjp8dtAyw5lQ2+/yanjhftbwKDf/8bZSARuTWSoO1kZxA3DJEyDjPwD
+7WqtLM1stMqxdAfs4OSGmEug0gTdPLl0a4TbJ8Xox+9I8Ltw5WvDe0i4difgABj
9Dix/NcVujrjMI/F/9eyvwx5kbwspm+JqmDaC+ijlQstnhHIYEk0IVa5U/AV5r0j
jI8ElXkNIbHlCIJd+y7jHl1udbCf4wYmKnRJFYRNOCzWQl0XC6O4BtUaEkwWdLAI
5R7dX15WJcxFDt3VIeXIjNyn/cZiZSprPUPXeJvFle2wiWDnOagrJJl//MS3XFlP
PRVOlwYgkoG9WS7xH/yPD7lTrh8e0wEKoeeINUkWd6g2NyY7kmqUIfIIA+AJEyCb
xklac2FlxWIW9NSFlIlEInjPUsOV2Z64ikNJKo1g0B7j78iqkX3aekXS9NATL+q7
Rto9bZk89zzBVGScsC91AF8LYaBBOn/ciWvgDGABgL5As/LfldH0BfJvAvNG5d/6
xBfjsamCzDC7+p5TWr6s+TFy+sbGWZAIO5VlV4DWjnnyLkuuS1W5DD6suYgoHwDD
iwWxN9OSFHeDG9WI8uTeXT7MYAl97MbxsY86hRpXUpts5d9IFhhFydvIZf8/fDLU
J1Ci15OVWFvql0T94kXfGSKBb4LLqs3uOFeDyobLpmSiKZqGywIvaD3Wx2/IK+rz
2FAnnvMP93uSdUFR+rfH3uK+h7AQySIIMChIYfuEHBei+Yn5AZPrDX+Aw61Xfmgq
iRK1tSAQoE0a6cTHQ64YusIkIVQvLfRpfDKduPR7ceYrhHUCdysOT1TamYFhcRQf
zdGM65T7ngNv+pVN6/CLkSVNgvzw5/PBdtDreQ886Nm++YAPJT50H7//MEN5VCbY
h+oeFNzZMzdvWAzssUS0ItxiKk8qq533o5DFsws5VLQd2/g8ef0HF4r1GVQWu5Gb
AS10zjzqQAPzg8cZAEECds6i5DdcP96UWY9aSsZ0nDbpVE46ydEm1k5BtR/4x4pZ
7OyHvDK5AnNRh7fQ/T4+wJ9m4EhnngKP7TImEQa0T1aaQIo4oXa31hjCHklvbjY+
K1+6VWa/IpN1g7DXgrr3R/tArugSAXr4GwFgUCOrWA1g04yh5M75AwjRKMPz1b1O
aECpfbDBSc5O9s6DsO73Q1PlHrnOOnVjpmzZPOdfFP2cOd9Tav5R2MnaBYJTa0Bh
CHtqYezcFP0owH/Ennfdk3QhHhofewe/mPlLc05K4xWp09SeC0otDQxnEqqS/xvI
IeYNlUZWEW8R3uBZNEuCyNsv9uKhpnrbbSUUGUZ0oKktzb6XJoCWTVsR9OQhz4CC
16/Fb8CyCHjYO9ZavkNXfYqfrdUcZI5weI2MBqhLqfIg46bGyq8YwmKN/z+95K46
FVexE5+nJiVXzhCWWKG/YT3wjCa3sd2ZAS9gRY5aBMvqrCwWxypZyQ2VCcIXIZgB
pxmXyRcB58Z9MsaSKNILOMXrXwN9IbOIJWVlLeqk7ZAwI74rwOPrwe8NSrymWEcu
Sw3pYXU3VDSEPgebGPrvGWKdxm2b0uwpC+88nNGJvLkVkhzyIY84SLLjF/cBmZZt
k0zAP68GeFPa+O0watW7Fj/NimVhdazkPziUOXaSNhCUTKULRqSntIOIkvefDDgg
7MGRuwsCBQau99WBpbQq33odsML73VxfbXbPMadHoQ1eyVDk5txs44XRuTtOG1Pu
NH6nVThW59WNN+1NnjfpB2nlT7YJBi+dOMDWDQe3EUs4cucZODE6xOv/SdYsFRLO
Jo3C/Q8Xc29lTE5SA0Tf6b6Lpbm/JucdwB3w23EizAYzON0j7VuUfkpv7O/0U9Kv
Rf5NOXQFseH/tiRxCpPahY4cuu+za6izJfHKHb5P/rlwLRRoZWoXnHkwCq3Z3nFK
y/EjCvai1HyhFIxriXdr0+PfpbOOwLd9d5HJd3Mm+f75pA9f6PfdQ6Wk+DIde/wJ
WncO1s5CJL7R9sELnENTVgKWMo6DP/J+JQ4OiuLX/h+x7gNJqIVgCUoHLytrxX8m
hdQib9YkU9xDkxkc6EmFTZMgkNNyZBTkWN+kcfYPZwS5TaDnzijl2dXFpbEINGAC
RwNtipBnTEb03P9k/Bp5GO/kZT1CF2xkoPRujEvxxLx9hD/L7++ib8ZAKt3kMxkf
WqXwWXj6RWdBcnQHvYouhdp1QJamllMXdOBRXtbOHOhOXL2OP4QdZqGoHbIG5xoi
vFwIix2WNmjXUdsPE4BCLASeruz2zt/qQm4RjW/SXmNSn93c8edu7lUTs7l4wSeV
PtCvlZWktUS1dyGE0PQL25gjInRVWw0H/3W2naJppeGWLbNgTjLiV7Uu5f+z0OFp
rP7upbBR3VMLhixn4sAi773icJwFszrkMOOaA6Tfz3huLkHCX+UfYzpbJmQuWgT1
FjGAnKHmGal1REqvGvudF8xB993rnoMS8by7Fi0w2Y3+xAK15jJzNvyyf4BAFZc+
7YVg0OerbaiNzedi1YAjMHg3/7coFPnqx/EdLg7RxqFJCIfOsst8I0Pzu6xUstvP
0C9Q+lV1SfKQEM+4asTK/JScRwLSacs3CLx5hzbX9ScGz1/noXjym1xrOp/DR8Zm
uxbP0VR+0bhefcfNlHyvtRC5bRIszBvUVGdCB+palIw88UEpqsq1XX7mPuB971Ps
OCYDl0niUaeyb5qzup8LTwZIvkVXc4CZgBt0ipzmbnZ91eR7JBMdn6Mjl2M2Ljxj
3Ry40WzTQlpHpeNutQ8i66AwbLWaNQ/8wTPf4lsD7/lG8e1b1M6Op3M2ne+z9BOL
4rF4oiC/sA5rQf7C/88nQWoY+1u44RyKjYrntg3GJx96JtVUPl1nq/lJ6SCPiqH0
N1utzLkR+h7+NzNNxmrDiRh9quqfTPLAg+tCyr+XVLBVpHFVWni+1zV85AnePBpk
Ncrsi+Q/uJQe07G9MlqTCw2tks24fE/8Ud6J5u/dhT9xg8jzVF/imEYt9ArU/8jg
MqRfx/J8aCojYqfURqR3RkdqjgK/pDRQPBzkma11twfCUQJfNzStbZpFG2CUnZrI
VmSkiUZgcxUZkUSA2cKrRgd2EzJwpXHAnMLipihuGkcC9wPHwJ1TpwRKhZw2VBRn
ZGyuE5MyxknH+FfZuGfnF3dC1Y01kGZtluN/IQjkRhuwKQcaL+dRoyrVIzQ6go00
v2Hf7d+SQmI4SdOtGWsgMq57oRRSdeyvuecEKIRZG7WfyvqSbTjK9O6PA1fGTuKm
hInORi90S5EBg80nBCAVAQ8Kahpf1lPPqoCjM97mjYLxH6RhLp0CXe2iEQv6WElC
PrIiCfpUiGSDia9ads/BHLMQNxs5lXBfspnuNFrbZKlOqK4eWWd3cdAb8NIZXTgM
idD8RQzxvrcAJj2usV/8o40OkXG6oOfiwMEl6IAwD54MSWC4qPQEBaf3SwuZ9N0c
b9FbDQTBhzVs+4JsEqlp2RNuK+VXI1DgblLryGI0bih9WJ5BevYVHaq10Zov2YCJ
NYH+C0A97k4KRqn2pyeQ0QGhMO0fELpILXzycHkY5J3n/vRx8WrdLAWwWYhCiFbS
kt4k5JLKsTH+J9IJlOqpqG4P+eOSny3okj8lP0EgHLvTkqGaeeoSiK+pBYtEMPR+
rx4y3q5V2ErLkv46/4O42BZnqcTWScWyyow5WJSpPNupAZARedXwrT6dhOPKke1j
961jSbG7q9ky7VnfOi6J6o2Np3dLRm3U8rZMuP09/EL+PH/l6HUnypY8KYl7k5bP
SOGVtRzcTo+vZB5npg57vD5isUIoZYlMxexzBp/mVuDLDh6CdlbVj6QNAri1tR60
B92hNjeUb6ExDlRwjD8enKix87GNiBBC0/RYmXaF/Nvm3u1qoc7M9HKaxEAjG7V+
oIA5UuX1Os/U3/HXf+Gxy+RUE3YyrdGXQc38dDCq65+7ebkOr2TWIgfrlbmN5Wvo
Sw4yXO1tYssJBOFdIqP5TNFDmg6zU7R7fXmew7ksAqXJOUSBXPZLtW2nJQN6Ljme
ZXESM2PwjozvbedIsylxDQrf81RYOU3B4CAM3Ix22du6NhQjCmMEx8MbJ3k8UyBm
J2CeF46ciIbqXE542j+69fabSSwDK16B27Vj6y7TcaqhukBJVaEoHK6Jks2A1U/B
dojnvJiGFof/wuprVAQriTAxH5b51RkGMMMmt+cJihg5G7zzh6hBHpQIqSQ5AaOv
xY8R8HVW75h2YalcyzPhcD95pf2ux/c/7/vjf3Ibo+8eR9GrBGjRwKdOx4afO0b/
tCI7xC75OkXTBd8IBCvV4tgB+wnDPr84As/UmZuZqIkBicUxZHJzFL/yy4iSDtDO
m/7Mf6LKhDx3GyGIKB2dkMB8ppgN6+N6WXsQ9CIMgImeeuZjt1cr/FroeP2s+G7Y
PYlX0wKfiH/laJwep7eucvoJdmYJAdNR58tf75roLaIUNZRZdq/bbpRz15wIEmwC
jsr5XZF36pMgaggAC2c9sPg5cLFBf/bo1jsfHVPu9Ngs69V/KbsPbRtmKM4T4DVr
O3n8tvTvGaW6XPuasJJOYyuLkLbecxcfjsqqCapz3EL7cnZbhYn6jElWmCe1xSW8
d/bEoqdgQmqVzwdON2i7Xch46Y/YoqPEQOEFEYqtEELqo2u46KMgyz+lE4qQoD4T
7t/5CD5kOFbA61S+OPF8i7jt/667EUNpND30yngYnbwrolPZ3XDECZAaA0wvRYpV
COgKvsz5H9JrQn4QPTZtdLL4c/5cF8pvJ+HDi3itF74Vg6X6/JhycG01AuNfzKSC
BTLh3JsWEo+pi3zxyXfXUUDS7d6489gurDNocAC0o9uc8cLkrMLCz4vJ0IbwGcd6
Y6MYaBK5l7++B+8d/+yTZNTHMQZKp4hUiNBYp1nd1ZO0/fculNKo28NXqADBa5Xb
EJsKEUGIYrX1StZ9vmsVoB/yHuRcS9H+mGukU0bOBNRsAKXXj6bI2VLmxUU0pRjB
JocRSYN8AyYXydVruiiUSLJkEYhph1y0ML4z0OQ20hWuVYg6y8UXTkNiSVHpMAT9
P+2N4LPxCaH8b9Gahk09aqT2ieLsSZDEniXCnSOfwtXXNncxLBMI0RtXlqFYL4SQ
/WJx3m6klTXQSQplRXqsl9uuqBi3dL56TjFanB0PO38lgTfIiNkdzmWCMVnDmo4q
4K1XFcykttOXdmBWV/8Ml/V6mFm+P7Rh0xp5/k0Ity2Vab+A/CGLCf9Io5kd26pZ
71eMmIhb2NLHzyJx+L7kPYdAiZj1ZykJz8e3FprgCmyGIwFBV5yjiAUPP5hSP+z+
AQd8b8qfLydB/hKLBRTdQ1BNtRC3OtCUCL0/j88/3n+7hM8F56Eay5drKtdzZ7d0
cwbY8e2j2ybtTgMJja76rGMeCWfrIRwNY5bATujPol/PzfztdYgyttoGZYvCV/KA
uBFoFaUFdYV8BThPrivc9ptXBD5xIiZMFEbgQJ9U9OJnKm7aE1AA23g4XZVrGI3D
PJCEda5UZuHnStAq1K7LewJe8Jp+uBSy/WXwMvullH5i0eDuChBsxC6sQ957WqSx
n7yWaB6kZYkz+BNbVBNFN6Sp6sd6gaAA/rYpZpc3UpPfN6EDp85UPAfLMHZ0SwG/
Mt7D80ZsqpOxplKIGYnMr26xY4jSDsDR8P+kaLRLkEsHSWhfx43TlES87Iv86bfo
i6XpwRHl8mf5qMdlcKxQ113S8gxLAP4slGloIt8Coyw8DLy81/TbFtpk5agr1/+N
9LXx0dG7erkWYwub2zSEz77hsVys6f17x+bSLy5ofSbvC624ZDLasYb5WvD29xUw
+vqtyfh5RC/0yJAPUXSsjad71gtHMaXcNS5CHvHywkD12lrqmQb/JjzBMB5h0Bhp
GXrHNLfwAraJ3MSewlzPYDgDbzfzpo8J82yN2PxdVXZhqVa+ayh5GifJy4yk+FAL
kwdx05v2V7y6W+uZrXxS2q473GQcslk/Konv/Vxj+XDMLIV/dbvTomxTIXKPFIZ0
f0lKulleei5yJjE1XjT1OFDzVExeIPLwgEaUDPqzePMM+UsEwW3xzj/148LdwJ8j
Mv7Rqhn4tAH6bHoiZJL8vpCP8/jNsT8swdbDx8JTrVYmk4rCPmlH+hF+W8CbpuKK
g3q1RINi7G5Emb4hxpVo4aKFBPx4J5ZxBZywuniAnU+kETyNc6nv+J5QZ4R8QdTZ
/TYcY2v2guoCkNaemRMxwZvMUw54hHWr0DYLuxBQhf7r1TB+pZEBY90yh0di5d5E
63ggjxnhAHHkhX+QzBie79NPxsRidh6Tzqahq6U+CHKoXswth1Qv2Elx3xEx49Zg
pSU2TeJ9UwwfTO4PHoQE5oq1R8pWrQtHWcLOv93ySlrK/eRKRjr5xR6gAWsazVx6
H2vmDb8HlJPaqD3qUyvBoNLlzVUgqPVv1BUl6dg+67wNt4sfC+twhmGqg5wV7D7y
Jalrq6IlYucvYeSnbYtoyLSsWJfNAlZd06YhkljqBxvPy83Z+3wqBpkG+D5lHblq
I7i6J8nYE4mz8XJGPZ7QMIuyDLeqkTggiTBA1+ls85xtcUfykQN/AFtPeHpWLZvb
DYsv6TKgQRm/Y1WR8AzzNaB+itd+aG3SKd6xyb1G/jax2u26zlLohb71op6tr3Sw
3gVjJssbAwAm73NjcBzyh9oUQrEt4VxA5sUy8/eDHpQdIXCoZnW+5BuveRh71+BW
ZNPN+yEApv0nyh5i5Rp2/NLNomo37ZWDZOAbgATQdtoUHbdlBX+PwYFstalXD30Y
U61loYWKj4gDYhYINGgXoYq/YtRkkFFl6jau9q7kcor1UtLfFLnsPLb8MIfr/mRE
EHwI5SoYISdzN/Q2OwXUmZBHcSwllqyJN0TwmqIeueIfuhk2yxg7DvimsrrIEyLk
f1PLgsSmXVGSm8oKJCrkuwFumcU4CPdbKWzaEOQDwvo4vZc/zCjJXDb1PusabBAv
ubCNU0YRa9IHWpPj5pk+wF2o5zApc/8+e1FLJsgqjixOMSNHUm/ZRd1pGnL0SU0i
Az/5+RJSTMW4kYKHb3zMEEhdMoXkCcvJF9UUPiDyCuyNUEU4BP6DepO129HKPaQs
yeGVxl0obQ2pHejuNY7o5voKiIFSt2VTP++TXnAE16dA5Zvv56pCvYbziyWp2tTG
51oUtZ3VUYjjNx6dRnyIkGY40MH/AVLYQ6nW5IAUEAEdyviV5IZ1Af3+trChKeDd
mvVHrt8W0ZAwo6/jYAUELLVxxSxVmuu9vlllBY5Lnowu2kHJfdpFwEZaWPwO8tnA
ROdckUJp+GSZD8Bd0rgcB0zmCzIsKVz2m22iUobOYjvMZ1leeTDz9IwkKGeiPFUX
83aepepqWIIPQ3nBUsJKhFdcheT5WpirMwqsDTotjSzxkN3FrKrPjgXhtDucYwyH
NItM/9N2yp7tH6l70Jb07ZFtwQbG1mu1sxLA15nPbIlPzwdL8KSnEH8iLhTYDV1p
b27fDYQnYdsXbB1J10OFZ4O2yVFIIrWGzHuetim9M7AYY57X7s+ieHjh6d3r1BHU
1EZoj3llGT1WpAFEO31x5J4kppKomDmBKVGMb+4EEOANe8XSK7byKWXvN7KxfXfW
wn613tyi+2ouZ6Z+Qf59gGI86VLg0zORG9eRomw9YobZz0732BqQNYFEkbvuR4ys
mrvkvtgtl4Alw7PwY/g7mYUdrF7fmO5hbJYIFmto9VPW1glql2kyD6xktQIUodaH
xSTC64yv1w0SrHervaYIFjAtk+AzXPkzJLrFCpdJUw8G8OLlfk8s/ujOStWWw8VZ
qmn+Nt87wNKlLuPv2ReopSLzHxwO8FaHfm4CMX4lTJnhudrU7GtHDnfe8J8J+hOV
SVC4WnV6NbkPJpPyHi5+SmDVTs7yXKDHKUR5zRJK8XiiAMVpNxXO0zEShuDQK8hD
c0olkj0xX64CtvIxD/hc1lv3TYF841VcKlWGO2yh9Q0CG7nybeJs8wERBbgN+7AI
1TWQOe4cShdc3FqFev+tNAfjJxm5PRjiV0TtQJvvEN1FmrKKPkbf+bbZynHgrxmk
8V2rd8osKw6Tz6ZpJPwPzsCUL67Up14ooN/Lkur/wv69KSX2paKvH2SFeoiGZDS9
vVxwBHLOvUKYEPa7GEHFfseTsRnGC/qrmHJ1LxLRYwXCk+arOHvAb24lj3PLD5c2
ZvBCDN4QwB9N4WzJCkcFwabI4/3pBUFDNN19HZF3UnMqYirsLr/pKIqteCK++Zsd
jE+lxX/3E/+tsheEs+VN0g4Rhk16aeIrRF0CEaQ5mOO8Kg1ishhNR7zlYhhXWx/5
9V3tjuIgHUEPF57GiIMdRigTtpbY7aMdh8UID4Zp1NDfutZkfpuNq9YIb8xcsUrz
QtLm2wI3M1a8/iPlVcPX92/l1anqYPvNsGgYZppwQU+SKEfIpBYqipwzf3cHON6/
MepZZPpS8EcKe8yivLwaMHWqa1sXoHdiHDjjsr5ln7zugl7dqRhDdnT35v4/S0xk
GChrAw1iWBSX9V3fbZgD12RSSAvm/wbN2KY740PPVAwr0uIY9o5w6XSJRZ4sktfN
2JyayyNoXCf0da2wxZbGxhBGBi8/1r+yUR2IAQn15x1j11/989nPkGDuYZdNvBhn
NyS9tIzwR0Dii+M1Kim+FNKka4WjFlfLOEXPc7q6Qar9aWw2fCBiHf/61+k11ilK
gm6L1obDo/YcYG01sD6/vR+AqFW8qmk7FY5MBmUDbC2QGtiwRRA8FFPjWUBOVS9M
SmDuIEbbyNZgX+NBWnexcHNZrCjuxXU0HPdfla9zO9CBKUb3cE9eBEwyD45VxE5n
zoM+4cHjWE0xf/yeBTHjje4qJA5jTlzzg7HLpbw5fb2q+vYa9ajKKYiQBX5Ttq8G
VJ74uIGVthmm3BZNkFgKXZKSXY/n7lxTsF09BcgAbKRkLcq7vfXnhWZJ8uXImB7q
XJazOZYbokWnnRBySo3nkfVpcD5qOlGF/9Y34m/2Ewt0PGBslN9nSjLl1jiGZLnu
G0kjB1IIrPikQh3CXnDizbhiRrFa59whHU4xzJYd/SQ8QHTCVO/ZsAWCSByI1DWG
ldKxIP2ax737gyADvbRh+UaTXInFwnrZ5Mk1ey+SPp6MOsOjryWXm/zkzXVv2QC9
TeGx0ze2SYK3/MO1gDVJG3+PKGFxYZFukSbjH9+T6lL0WfcD0k2UV1oeUe7k/r4t
l5KjutKfbiuJa6C8bg5Png3pMk6ki8gCYZ3dsZpVKI+t2Jq4pgGUe+hO32TBNTJI
VqFau/ogSs8QWCrQDVFJwFSLOpnWqsGzwASncTPBe5Z5Xaj2kkpnOvKyBwm00CNl
2k05TYrDyb2lbTkQku4ay6aUI7pUHU7yo+SfUrxh1dqmqMw9HrEGO8Bxb4BnoGcF
M1jfGOlI6DCaa0omYQqpt/Gh57/5YNgpurRj34nlp+gmiS4r0zgnH6J0iEMMiwzz
XK5ttG/OHi+pBaZfIzpB3+UgAi1iPcxNWaOeTugq4gbCPlNwHgoQL7segOBKlET4
O0NDv8b8O2GzjzchDu64ofHeyeDG9bV2gNzQkoe6QMjeoc3N6eMRhD2+VBqlUlb7
J5iUbzIRRD5wHRfHhosvAqTiORqYGgkXmP/AG01q7MvZVQBxm+S4ZO9gAb9gLq5K
dszi0Zl2PZFy4flGk29MePzOb27c/CG2S0nRAsg3soXhN7/yJ1MaRNeOm/2pHHZC
q5BblXrqTSWv2y704v7DUFvSarMdEMwo2ijVJZXg6hvCyxgNM/BAM2wsNYk6Aim/
iDsC2/rJ+oeQ0nEddMJYndpTdqM3s4vKLr2L2GJqGvC/EMG6QcspSXMgocLhAmm1
HNA/1b24+LOpZzx5y0ke2xDoXPxHI99FWZXou5/s51ObJoHQpOLM4HX3t3ug9zO9
k+GN6lukFHMmBWXMXKCCJJ0N4Qe+J8IpDdaz2wvofi9W78qkm/z/7Y99Pr8OMtEJ
VBo1AsWyZOr+r/rzgORFhXngXHCRw0OY6KTq58zkX2SUrqd92KTkpSATXkud7Buw
G6YW4uHaAkQ0Aw2Av9zPK+0xRZeEBRksvLXMYMkgSGH4DGluR8V/UayLX5vaQPXB
0R8eZVv9nD3u95l1yaYp4zIhdkTv3VASoHYecRILZ15lZ2rblYtKBpkWiHUCNMR7
r3IR/1alGWQlVDmT+8VdmoUZUoRXb31ThSwGuwpFaXo0T9F84pqyGhYVcHVKeqd1
1upzYHjK1Tuz3DjF3QvbkQJ8Lndrts8gfUN7QVi0FACQOl2hcyYJznEZ/ay7PWBq
yvV8bDg2FN6wvq63SDN6cXm7/ciSS3+dcFHsLv1rj8jHUnAPk+SmEQo3G7fPRh/7
tg8/S6fuDgSHVl+0XYnWZnrHu6CwZAeTJ1ndnW+jMLu1eWVgm0Sc4Ahd35ddtNe1
ZvlZ6uYYwdZmCcqB8+zNOk2vKievCImi701RHl09RWkLPLq7D1SIY+Hl6SBdgM7/
mMZi6LsSjvE3l+T7pPwtjtwHwvLHzhRjm/p/eSNLw1rCoHek6jNDejm0OKhXsnSl
549JunTjmVesR3PpYhw6tEM46Pz6atr3YLnXbEe/P/FfE61Vi+jYzk9CWeHZtOSA
feqYrLUGwhE2c7xrmX13EMY3J/iPNVIw3YHVZi7A460t+tCBALElbmvrM0WWNM+S
F0nsUpeu7F74ZSTEdz59+3cNmtCr54U2QEYi/iFawBte8U99QiFjzFrSEmRm73HA
pPehCgPGqj3mM/ih1b8vJ4d9j+7y7Xy7Jul8VnAqi+FTKaA46JUl1d0QcYlRLipU
Iq5NsILDO5Zw7fBMDZThfSTBp+lotXkjKpYl55GjclH5YMZ8kLchmgAMw3ZANVNd
PsFYcSWlOXnl0ZyhQiB8M0ohKPCEqK7qyqrUbBH4MFb3JXVJ3bdlIzmtjm/fszqR
pwxueUtJ215Tt/thwnkzOFoFP44hh3b6TXgRSSR5sjKbVdBQfoSTCUQIzgijwxwe
j/i4UxbYspiw/3nRWTQQi4g38n/Sh+dwER09z/VsWilcenYNxrWpMJ2q2cMsmubg
9KWHxy7NkM8h0FWmSEP4RUkvDJBI+TPaOqJr4fBmKk2qVWLKCaGQUfHhdUbniHI2
W0vVkjv7CaxjaLAMHi57+7Aki3YN83dm6xLCl3DLWxXEnR2v9hOEeAyI7zHS1LRj
Gj0FzpUDck9ib4MYSqpFMmvEwtg52LZCIyt5ruVgyPyFfkX1A103jh7OH6hETlDG
gTGaaxlEQlonbIszO3Z3UOq+gRsoDM0ldOi7rwHPN17i9JwmDd18zRBj/D67QAYE
WTGvWhth3eL5z9TSRsSfgoSSE/D9uTcFllXonFk/lnkoAMmA7O2vvAf+Mk7sMDDT
IJoMvvx+J2HnE8mxMzdmnHsnbErtTfuDSo0hGMrq8N8mgemPT82HqF15sPy/y6YW
M4uvTwm/HwHQCT9jl1yRgRUbBhEk1lB2W/Ewmpq5CKL376QeXWRy6hbsfyiNaY4V
Os9G38KGwWMvkeFuN1ePoPHF+nMFos18obkXgZPObbyf4BLC1sC8daFbQ/MI8lBb
RNK8KFbcCDidzsRNmESP6pIgt/c89m3bXYPIeMcxmYjhZ9N1ryQGYg1wGKm7R2wJ
O0VTZxSllPL4jcKa98GMdIV1ADNdQ3IWIfUE+rF4rypi03FHpZIDQXQXP+ongJ7s
Z2z0/mTSY9/pmdK0WPtYOLLg+EyJJEBP1XFO9UDWZ4INaY7ICyQyjJ877X4yYVfQ
8/z/vYyyNr24Bfi/el6QBAWI8I/sRuWK0kLcU9Ixu9X+60GgMb8NvJ49skJhq21H
AEc7aQVPMXdeVmXMLwMjFTKWD84qOlh96X9Xyi9QHPxahmqbAxnSgK0OawZNTenV
GqpjJorL1e7WLZiOvbABjk16DSHTZzmzw30EtWgCkEny5LegBBRrhzhWTT/twbxz
t1V528N2Kg6oTVqlpD+DG8oE+8yaMwoSReyCmuOAjMsDJl7NgCwhZ16ZSNoSFIeY
n2zdXt/WmSbwgiBMdHFht1yaoyAEsDgqoHxTyS7x9HUpXVgymIMU4TCprBVGoHBm
bZngtwgsr1QPo2XAwjrVpBywnvXpK2BHUGdSqZgOjRNpFX8VWdSyNPb0zX2JJ4Lz
cOAT/B6aoKasOLnaNPSdXRNKP68QkrXPjlLRMk2JoBO/KrVKaDKESzNdYD4sbKJ4
kAu4H0BWrWluVbzIPhPYtoQSIryZmMhSaQRsgVGOSikFZYQOguK16+k5EhVi/dKw
3wRtCl2TmiSRVLH+uFnFm3y/Gp5twZ4Q5Tv4Qc/ly6oDBKHA4lldXkTkz1po6fX1
ObSfLOOWYZ4EdOWJoMNCB5lL/mhWYf49B4wuJlgVxoMpSCyd1o7V6ND2XEUDtv77
KgK1Ha8tOVDxcWf/6UojbR5aKJD7MRKFaPd3MLv+epsM2ANKlx1DD/C68PSi82bE
h+MX+h/LQdfDLyUN6UA/4P7sfKzJNOTizQqFdoqfA9nVbqPdlopM61cR8fpgvTVS
UMgeYq3jonIR8/Rlflij3zHeNoP01pnVGqIL4+ubL83Tn/QgPgCujLljaTlS300h
Zn85TxZch8ktS0Rj5AJoShkmPnkQPRTvq49U52h/jjF6iTBA04eZMcn4yE/jkgm3
/CnnFMbYbtvUTSmxdYIQk4BCbiFrSSr1V0K2LP0kprLy7+Xii9sJn1SF/anmw93E
D6AZtUaIy3i18LtJb0WOf+t18ndx4/DT7PhztZS8vVIf7l8wNEvWpQtyCdkihdKN
AX6udy1DlyS7Sm1XG1+w9rG6CC//+EIr90Y3eFKwOgE/IM87i22JMoRx9HmSAg8G
hbZsXNTvQ0Bau4wGctAyJcm72enOX/4XTNyveKs4MpA8gmo480OIdMm7ABLNAcXD
Bp/1dPQvu7SnlH8VxeC5hWapGF/lM8lPIs7D/qUvf6Gs1M6jyQmQq+/LrkCU17Xq
v6o9SjjmfR2OCEIqZ6Boz1Vc7fJI5ngiQ2RSAcR9ENCJRdaD0xjulepIPYovwdMI
jicMCpfQ+6OE/2teAodw4AOSt/14tAAO48lUJiw4Vikhs+Er4Taxm15xrDQ54oJD
4ocAoGIoIb78SPcayTHeZfgG8FSKzx0ghGRuhUPmsGKuVYh0/xwq8Maf801KuENh
B5JeWubwNxXlyLb58kkaItviGckXqE8uYX86UY8m8kzC7tQAyiTdVIgtSUQp7VGT
wP6FjJMcjzafe8l2IrjdsZUoakpOHC7oW9z7/ivgdJ2csxgX8t8xFafnQ6/IWCO/
9Ldbuh6JwHIWirW52pIE+Lfe5vRS1dK41IuwJz08yjGjkNvpXvcBClVGeIrP6UV+
8Qnme7hcpcCZu4oh9EFOxEtNz4eD7Xb1yizVQyXR2wK3293k2uoFxdFmKJmfjYIs
N2JEgtgRCgyYgMBufzVaQopQd6N5SaBMyptRKv2wJdWgAVcVWsLJECumMutnsJEC
Io+WWnh3B8SaLIVSyA8OICxWMoeEdFJhgVFotSZ4/5FlJGUhq/FxBd2JJiycugmy
eFWaH48dUF/eAj0bJZA8E4c478sv/FnxO03U6xgxecLJBBOPSYR1pe8OyfvMLgqq
ALtTAqZISfCiRUcuP489QjZn209bZRQFRkRAnNsauktm2xh0Y5IKl8sBFohhhglr
1I7GKJdBEs9PQAVwzwGkYk9Ie960+m9yy1fjzg8+uzkmLja0e3NyteBLE54w9AxF
lUBQOmftqDPE7MFavlig61A0eiskfccjhro1+126+JHpVhqxW+s3AVvwfOFDKz5H
C7PKr8tnuD8qEVm58sHqB+CzF3OVXwEjhIX3Q9E66sNZ8duPVNX461j2Y2tca9CV
jogZRoRGEEWoWgrS5PxLkG6Cz82TB4bnL+aCT6TqYg9uVsbXS65gqvCalquek7Jv
cdEUiZ8G2WdliR3n/DkOE0vfWOOkFmhQMr6cDXnRUyaxIiUG7DirR9acosdkhBo0
5/ehWg0t36PSE292xu8Ib30kShskSDkX99D9qgWCKy2cBWGxuQWxZJduKor9n6no
feItt49BgVzGNV3FgVrOOSCk+W1+YOi1KAiFiv/WeBwp/3We2GXgrIM7oX1BKZt+
eJ2SBBCgTaA/2xqKFPhfcoXjedwKt7kwosMLFqcItj8HsXvzgza6gPLZcqPCX9Rh
+qgkoy+UfoZecwrdtJIeR9JiaAEJ3HOzQsWFNALkfJIB5BLnH3DDkw74DIeePBNK
jlTtkP023BRl7KA9o/p3ZIPFJ4aZdUVv5hw3LmQjKObR7NoCey8x+KBkRwbghz0Y
FGgbfmccTLUIvfhtzEbsLNn/e95+ikqWBrx7fQe8oxHdMu0dGgF4xVntJeP4GE0F
Tm0XQKHSJDmUAaWRUNphWebKN1k5JTfCrVS9N+OUZcE/Vw1R7dEnXaf5J+/3wQ5Q
+L3JrY/8EJCyK6G0QA7R3xOVHNDdi1euEVFYAlaR0oL+8b3cLpVZArbNxlJGFOkV
kgQO6tFRKT5MF117NoOxKN6UNgbQ9fXupOwZevY+KmIE1AyebuOB30i7VRI2ahuG
CIlRusNH0S45u/t/1iSqTvBrISY/4sdx368FmzrY1dXpKU/CvvgYON6QO2ykxg7P
TjUoIlUvBYmMyqp5In8v/plGxlLU9+rdnHeMkDUawKK2ZnLO4gC3RQYsyus12bm+
b7z1UmQZaR9mkiIgs4/RY0Jx5qdTtU69KqyHhXB71nGV7BVxVyhAyOvzCXCXXwwE
rEUC7fHl6bSCgbYkiHKanL4n4/AIlqS36M8E5N4kKSNizDCfjnMyl4VSbKRkT62T
vLSnUY58GkgOalYlWRQK9m+qmZqZdLYBmKQPEmq22VjnpyAjKM87XeItego+uO2B
rPMfBUQgecR2lOO1xqgJnqVP5eScztYfFwL2QYVevobrfoEMzObmkbF7arcR7Ku7
+QHRqx6MlyhUytCl5udcBx+eIfQW6hMpdlav5XBSZXuZFvswdOlcPIVvdm7JQalQ
Kz0Mi58Tukup+1OjKW8L+9IQ2FLiTghd1I5atT1KLriOtXdGdDuYzL2Fal+bgJOv
88VDRnGt2EmHTDiYOTC/XqD51zA+73rvF8pxNtBTJcVuLJWJAfp9h/hKvkl5qOLG
+nwZRDR4nJSrr3QWxF+sfN+Rd8FE4Ih6vXdHg9dBnmgan8rQgaSZzKD/YrzpPm51
7HfIDSkhZZPaK3fAH8BM3PRz5YQWjAfyHUXjQub2r/XGdc51Lqc1HoltwSeZl55i
+gv0l3RPfbvR9cxErVM6bIAcOZZzYATof72jNHJ+wC1UEo9cwnKag+YTMFG9w0Nj
0/eMQCqLdpB0h5Qxow5BMY5XojMhBtY7x71dUzExHjEgrQ5xOhsbnsMTp7MNUkf1
HlT/0XsrV+1t8kJ1/2ChhtsNvSxR/IpgYEMoBMp0gRy+FZ8SEjYuqZ0qNuJ3BbjY
tNe4tz9CPwZmBWV9Es6Idb63hsqsgGDKscyH2O0aM0aOQtGzqv6nf4JRbaUWEB2k
R6Rexjluaa/EJ+wn/TR/VhKWVvBPH33NMPi303uM1GBFUeYV7ZhxVW7WiFifvlaZ
E2pzIYeqVad8dacMmhWlOIzHuWQ0FLPcX+DIaKcUbxiUc8Me59D6coSK+T6pAscH
mqpPlKcjx3woYO1lKWTIWRkUPkERY0rUBtqH048GyBGhLmk0m1NXpdO/pmNGTrJ0
4rsjcBo2plNwd0m/WbkuaXJ3tsh3qXLhyl7Fj/BDhcukFuqymN38dmFv4vkqGQMd
aQf/fmmVX99Vwj4GRbdPWJMxbejaV7V1G7AXZiqRG/KvD/fdMcFcWCYR7gyBHise
PolNJK8j7KU67Ud5wBSTgT2rXEeYlIM42X/DBWRd1XYS3Qlxkfi8ABn4ZdwqJsnb
KgwWQKDLKAlm+1qElZKwTnjGbZyol9yrZMjbApv+f7hPtV9OS9AHkIwwDZSPYIxp
xdOrWqihmrpF0TnBmiAc7uTAiYsNcTo5U5gR4DyOrRNZMWqkPW+/s5gx+UuIjfe3
8q50tcRo3L5+KUXB+1HbUpBvJE5HO4uT33hTvURsCMTodcyj5fr0iNhP6HsWWhkT
tPuvcTaP+Knb5un226Nt5tJLSRf0+Yv9+IlYpzJXiFqpmw+rXBrHsEbZQDIO8Psg
GR61UmCeCEVMi5VuoN79eZ+KxzKEr2KeTDE2km+uOaJMDEBOHQzL8aqaHYKF3p6y
gsE37Rve/zpbFEYOIsrfmibCBMVH6ge42KXxljdEan5xcXK6nFYwykZYj09xS2sL
yZlB4uAJvBMemShRoujfz8x54dICoUaxRGDnguK+1oj0k1Lfh30+G8duFcOv/PAi
wJv8Sl4GefNYWz1iKggDgYBo77zWfO96RbmNTrlGwGKDhlCelMGasNoB7wUd+O4z
26F5C9VaVZoyQWfq4+94zEq/xHrWn35QleXQBaioLbWdpC1dR43//aQdIV+tZVkx
Y36gV2t5arg/rWZx+9VmpfipjDRXlCXQ3AGaE8QI8aXaey4KgmHt5dryQYxqcwrA
0Fw9sAziAbwBdHKWmJ8f3Gi5wBWR+R8ySrPsXEBBWJ7dIalNsQCI8jBprRSbKoj3
MSvst/kyx2stWAFUxR+t+A/ifHrSY1tfulOH2m4/T6Mgt0wmXG+WnhOtHTenGai0
iRaEPWvkOwbJZrLtKEXFpiRDeqBdXi9nNS9ntkAzFYdNqR+vwKgC8RD6neYHxkxr
dqjAA8TAJKP0EDUnRxhDfQR2Dd7T8Fq2Gj7E9sev/MYi27gNkF7TkPMpF9NNmWQp
FIGWVKXzXa2oVCBfyD4TCoP9RKCVDV+sjj6/VuCJh1gvnrws6wMob+y5jsiXDI4+
DD95nFQvA+WUWaU5nq8/pRG7P/FJMh/RTVKqYOAueBkGMvtiudLrcrFV84XS74cw
3T0eTSLfvjq7got92iUuaWmOxRF6yMDAX9/k3CRogkhZEPcGjNUmbr4WnIWnLmCL
QKuBg9pHy08hCEdS9b+UHhZxkZG97xQ+1IzWxjpYQg7nwRi20ivg+pEJ4r0ltI1A
0/xYQPaQ9y/2quyLJpoglbZG11YQInYJ0JjPRELD04XvkwOQlBgVZIn45JicG/8N
7zgcOMefFOYBE6EFQJNfXBOND1M79gEopGtFcOANUlXcHsInQ0Tp6gEZoXVfflD2
4sCzQa/WPw/hb0l9p0yGLSvlzqK89KQaXwD52geHwKDtCRBXAdtlGlrO8oxcO6Iy
BRBn6rLBDO2N/N6Q5j6kNpeP1HP559jNKnKSO5BYaeaFGdilkgx4iny2fQ88AEWE
3jKVi1tNvDK1m7OWWLIcoE4gs+Xn9pgp/gq+0RV/O12+Gy6h3yFgrsq/d506UJIj
gnU/X+xXkEjg1BnlHxcBCduGHTKauDK5mxWLIUXxxkvzk51r9SWDf3sroAoaPoMC
/pPWUR/+jZcmxZaobzz7Q9Y7MXc+/zSsIKEOU0DJmkV4/FCl9k+ROWBhQyfw6jih
BCaFIgoSEvA09IVnyjEAd16pZPDWkN1OOz5LyIOT32Is9DbStoNCtLieB2PazVOf
kLNnlCj+etxlTqzdSxsr5AfSzca6pgXs5h2UaONDUBnUas3G0+6Nkjlfu8X8gXqU
lrxzyFUMnlyClWsVAM1ok4eetEA4ua6T6LzB1D8LO39Z3nF0cJAKftwbwiBeqLHx
sQMAgiss/O3UgaToM5oX1Ww7bIavZ4gsDhpJ9k1zjq2hdaBVzyiaErHSReyAvv21
dA6ubc/b/pZpPqv0G/YynOLY6ePNzfNKe58O21YrpVkguVmcGr2y/cfYP6LxqFdn
c9mOImKPGcxYcVD5xPShz2Jl9OkGToBY7p6pjR10vNfmbCQ4ORCG8bYIJU63sgDh
17Lvbq7ZXD2xt0/mZjbl+kEGfEn+v7sanvV6Ayqy2zqGpaC3Rj70eI+KvlL7Htad
JxEvo9EdY4uXHTX8KoX3jv2wZK482ldWgqeNRqS/U8cw1UgtSf/eKQlvxPXlr7KD
ripfBq3Rb07lIft01WgsjeCw2j3pNA0N8v42rIvMfwIbpR3XTpvIox2STpXF7LHI
MaG9kPBmK730S4Lp1hSu/v2+PoWnfL87eCa1R4+UGQLT7UBbMdZjzMyGdpzAQDeP
ekuKdd2FdJCfvUG+9sj/CRaCFg7Tn7cgPJWa8lt5DlbqsFOosi4gSl16rF7nw0Rf
0OKxcNrPX0y78vzinDPp4ZLcYTRjHQBZRQiu7Pp5eCgkXrDr2PM/VevutEdls6lr
lNQz/s+pGXgarZa5qw5ZL6ZGGFC7HnbH9/LWTRPlt1sNmu4eCg47Ta87Cb/M5bDV
sLRvdqdvAeL6cmWYBTlpPK64hXYWv3MnQiNqDrATfc9u+n211q0vfh5fRL1Zj0Qp
ZwZUeh5KVA69pfnHOBIVxR3mQ38hKxPpGtvkDpRpU2y0/ol2rzlNZWAqrmACSK4c
iTCN3DU7shgEaV52bEcrN0U13fsFMVQlCpe5UHhhXEwWDF4QoBP4C0WdxTRkiHg5
xbxKlDDhf9Vx2eHQ5saeaVHeu2tZUK39HvrUTLiG92ajBTzrniZH+URUOuf9Hm+r
7Hagg+zQTXX125C1sro6lCfyxY7nL/7tbpmn2b3yg4C+8jt2/vr13sgQqa32u21V
7hfXRbAXJczqYZjhTIJ7/QwVlVXd3aPemByRJfBi7pwQyZAaK9e2cdk3NI0ag8OP
t8LGnElKP8mLWvA7Z2Ga7t7rhn21smK8EQCAI0NlrFxfzki2XQ33E5foB0ywRTjU
mo30kDivfzVtxe/Ec1rov4SCp2MY5jCzpDmvbEKXMgYRkKwKAKdTaDRiiEDsCblv
ufdsAee0vqBbJ3SXtwcV7zZ/BA0tDKJLl7S15DrIcA1HCU+GjEhnf7UdDDukAVyJ
JWoqaKpGYE1ndSEoz/VIK5oz6mctK8ElC6ViuByCZHJ26TMemDsQAJ/s58j3GTaH
jF4kxqU/UI8fbwGWr87IwfphAT6vsUDUl9wFlP9j8r6Yri3KcdMHLHyQ6LVmCr4/
2psgcM8IMu6aIwE0TWlPeP1qzd/8XwNsqAVhPWqgMMbsUyhFFfK972WT1XxxB0SK
LQ9hkZltcRIkvDVeFE2eEQXF4Vfjs9PWK+Y8Wrjrmms3JFXCcoaxKiBnhvnz++AE
mkelgtGTnc1PxJqEUznpscjZbpbBIf7/eI/tAK3GnVsBor78NdxbbInl69/6WmmO
luC4l6RscfDepxCKIW2u3dhC+HmG1GFwr1tTKNeIbPf5pM87tu/+Jn167xt7vujG
8E4CesmlHDMx5nDDAsFFYLabj6Vmb1mGeT3Ikfm3LFVmOuaWtQWXZAwD3eKKO04q
QY5a1IBj1Xo4bJjc2r76B6whIRHoj16M96xL/B6B9/+rznV6bJDcuBbS5uqG2hkx
cdaGU1QTkCBTwgGY36m62Zc4IsDzwhhfVPn6/JE1HtikVWepzPc+VprFe1sPsbYm
LCfDHi4NkPsPbMl34EC9k/ybnT5XFOeApUyhNGbH/rps4NLTs5L2EyUHoRMw9OSQ
hM+HKEZYWdmeVo5Jc+wfh2RXGnUTjVBTGGv6hbra/SvagmKafC242OohTXNHmt4J
i6h8dq1KrA7hSa1/qAJ0v+FwptG/gP+MvYJLqI+ZWQGcVSf4ziPHxmsWM2cfl48c
UvPoG0yN5qd77AsT4aTlTGl8/lMpIDLfPW60pXc0udbMKmcRKsLs2H1dBSvOda+g
NyDVadv/13YtOb/PTq7oGxQEuUhHoMQRuCPDNwGdt/gTCt691sp71IfV9kKHI99Z
OMIPEY2VgpitPQdvOj6evw/6JlvE/5HkYobWIce09kQLJT7S5NI3axri35bqnXKJ
DieqK9kA0mwT7x5UVcnKGXeIDPyylWdLIK5BddP2K9s+aQejJl33BiEydls8ElKX
RJGkZJUmO23ZF07m+Ruj6pe+3lRm1b+2Whaygv8e4M42rFX882EyW979ggfilF1n
JU+g3cN3owSAyT/PfsE4r4Sky/kV6elDOVhMGPcF1pxy4+jw45rR1DHh/LpgEVB3
FMIkSnt5jtg5aDDtGuv3m8LqUuDH6AyAIBTql7YycyRLdzEd7rAFSkWoEocSSKUk
BvJtYeojxWviYLX3m8ImAK3vIUUSS1o8WMY0yjaDW8D3NCE4mqTuROek3rUQNALj
Q0Tq+9vYHImPkTIibtdUSdWNPg53Q389uXbs8UjGWrVQwi1S9HaBmL3fsgoY9N6t
s+ESmQ/4qYQPbeLTzhz6q91AzMTtVuPyH96rw/x/GTZ4NFeoqgdDWMkJiU1LjL5Q
6EYDd77Jyk4xumWnGqcHSGkUAnBQ+h0DKEmbZVqbg+qNmJMFqqrI80QHikE6gPF8
pP1SVPdWLhC0dCuFkDsZu6Fdgc1BgTIuEqQXCAnN6i2iItpnUda3VGZ0zX8zy3lJ
nPt3trBNU8Bof5Az2+r2P9geZNaGcDRt714q0EKS0vlDjUoHiR2G/mHmSLbr0jjU
vouz5WTux7zqOGQxX287/rCu9cu5YIhdIACqBhaqZBTpXTOZBqiAvH0oQHoKzxpv
jNjWC0ru4JQMtof4aFStSGF9UZCYrj2KypeD7r4tFgbKNNz/5KOlhHQN650dbTnO
vXEduv/BSFiJusTl7X/krdizDKxAgRx0yiTQZsDA+0UY8SgjnGrURTzSKzgBR7Dh
CTOMz8cqKDSxo01iaxf5aWAhEja5Uny1ehSiZ1MUChiJOFg8/01AITUlI1ssqRC7
MG5/8Xchbc3l2qIa04x43QNGTj+P64eE0oAICZ8HS1IGnfK9lCD0zKOT8edGDAeu
teY4FvwxU/rsYynwo9VMkBaZ1pL2wjKZ1HrDOdADCHHKqv/RPR/V8eoCZNOl79Pt
L2Wc+l5ot8qwXt4sHyRurSqxtLCnkcDytnph4kz12z2o4DzdzisYb8k6Y1QH969Q
8Yw6iDbCopKHlSVV04SyLXz+RC7mDQvgjiSIexreOSZysyTuM5jYDK47UWngaxfB
L61QlW1osOStVRslyseo4ySA+CFyVmvU4SVyiIR00/yB6lbmyy2hq4MOQ5hP9etc
BV1oBU/qcKOzML92qOCwHvCQ0mTxRgcP4eAER1qBR5nvY/3AmqYq4GkZAxj++FXG
9cbWfhq5IJuwk7eS3rV1dDsUcBkdaPlvmcz7BWsFZ0+9/Ap/pNzSgZxhBkqBO+EI
dcjRbV2Gg+XlfT9CAxX7uc7qO5RqjhlEbWmb4J7jS5vmFHBdC5cTFWQoZI7MYyoL
J6BRfCrNi0suOOPAOOHK/TWjqZGn46m18RzkXGT9Oh/3AZZCRuxx3IYVf1f9FXT+
ULYff/XwMQES8bjF7k1r4ALx14dgv+KGdRIUNTQ3SOvpYG/xsL/+tOEz5hdpFRzE
QOy/Opospoy8r2g45TK+RRGDEkinb5QYfDJSCnRRmtdqFVAhlJEEfshs5fIf2RyM
CxBaiNkAnUdsODYKhCUAv29sDPwlSIxgIp3Z6kKQ9YuwTsJ40G0/hSjdtCE7wgZO
/BaqS/E6YDNRXC8fYpqsHAsEeIn/9FzCGmY/1opOhPdBVsBChKht05f2DBh9qRYe
M0kn0dK9XGN4awcvvkdLWiVVEmAPRL27ml509VDXwFWOec9WSeJVf/PGGitYjolG
gU4U9p1bmY7MwMNCcZcHf7eDjOGkKKFBvCHesLJMItbqrXYPqPK9ytTECapBGZmi
sGeUWA3G0nbg2tOiea3ytOGtAzCRVMb+Osx++TfcLk0m43yYxV4esKlciwQUOK24
l9+cZHqZRsPluD8nJj7M9LoM0znfl8ZqLlclWU04nQFe5AKfyW8s6uw9iZxtyZ4r
R5O3gGTDn0TgmwTviAvQwhXSSpD4/6LZqpr3MelZT+9jE8vxbsbStTdLmFiA1s8m
vLWEBs30yauwxSC/1L/mNGKqnpLdFqSbV72Fb0Qu9BmPhnn2ULdFWrhZrVU2RQ4f
DJO+OwbzGM/sFLiao+kU9v88jC8GTVPmMY8JYK+XuaaQMmiBNKqK+CWfC2ThB4tT
RFOmfng7oUFRy6KcZwbOH/pOns/xihz3/20KWv8iON6a0hhjEGFbj20wvpNh82fb
SC9R8yOsGS17qd+80QhiUOAxyJ5x0WsdveLg+WnuH0+JXX0zGlJ3Kzmziiu//5eC
1zx6YiIPeCMqYg4G+p/k4oBzgBnWQCm2mOvHxeuqeyCJAcK8aLsfaEGcB6vUijkP
jyPFqVO+cpm47jrNBKodYVLFSvD7RmuIR9ife6/6S10s28d7Tc+xZEX7I258SnEs
ZoUIcZ3FrcLEQ1KRBRKCzpwNWV87w8ML9tKjsF91ngwi7/DveMWYTERYX1V/y6Sm
tI3PnwDuj6bJSRzxxl7uGnXAvWOpE/Apiksu1HWCuTnsjCB4ETh4XrVNRc63oWF3
bdBhVp2Oc5u8NJV7l/XHKcinoDNgRRG+Nn9pHba8GH5woaUtHIhK7BvLAazWCpPP
cb10WUXaHGnXDs2NX28kRuuuNpp0CnOESEr2yx3V5S8I+WwGCJudJFWcYbKtyUtb
mxC44pDbve50ns4DHQG+Msw9/495FqfWrkG47cYqJukrggLcC6juCAH8UseMQUdA
lzZclJ/RqGvmyu2nmuQB78YF/MiFPAlky2u8Q5hVaW8exwQIi/Z9hA9oVMkkGPhM
8bqiFnOx7O51cdVFM7Y2wc89f7EnrraBxExyvql9VISqMFqPLBQcWvsuCkbOtZ/C
gJ74ACtd8QafsjZXNm8i0B+FF2yz+jBecLvSZ+sRs51yCAnxc36UzMsifsotXC2I
/gta8I1TzZ/NcEyE5Y5jsL1WgH2wnIRD76nJGoI6yZrnyRRMhQdvyn0ik5qpJZt2
v+Rv5zNN/wLtj1EiQ3RBefMjtFFlj3CEUKdnrpMoO1ko3/i8eCyvxUDLstcXE+Lg
9WjqYkgGVjOv9sklWx8Mh4lCu2/BIXVyiTAiKSGwe1YgMrl2chbDC8LxyuSYYuWI
AJt3b9ArFI7rWoaZYL32fMwm/ezvfAgrTPHyixBglc3qZLf/WHvQb/tqh0SFKIcS
DWLeujLSBErx+jZLdu2uMMA99DjHMdtBOpIQ4b6i25QYhpsc8AOFh+7SxAvns656
k1i6E5lQ7O/Sq3FXXmgt7rQIEa3MVvjSfKEvjw9NwT8C55chlq4ECfADtnUc+yTB
dzdG/scazbvfGwPic+MQeFtY5kOa61J7DVVZRXowNjYqNiDlVAxecSbBxtAKX6sk
x9DGvkN/krDQIsoCDfjZC8RWFK4J67UahD9B+XVBtQgOL5IDuKl8gHEjeqRrI64u
VYjA+uAifxsFwdgSnj42Dq732iXC1hXD6gXGJHppF+I90w5cEtJW9mnVAR2eHs6U
GjNrhOoYUeTaMeQ1sd7P5U5gDYWBbuznBl6xQ77TuGL7EgZIoaEhd9A3P66SEjpt
PkefIxQM+CDWAGYadZRbYOzSRmMgov5UgYzf1U6HCI/4gQ4FpNKwOUQFmkddqTXi
exjBeUmMOyGqMvDS5SJuxeWLXZpaK1x/IDbmmD4NPdcN996h3y8AH+k5QeuKRVii
qq2HEFuCiTsERDbg0OHXccjmrYY9tVFALYYOXt4beJyZru+7SFTAUT7ZjhH2gAKR
WEjQI7ur+a9vlUnQJgZOlcmuzOI6euiH7bYJTYp4IUbrudNDw35ZEWvcudVq+U4d
waf0I4RoVW/HVaNga2uaGdO3CDUXjSPUt/MJ8IZXSfa/8pB05Yvf4YZ15OKS3qCE
DxEnn9aUykvrSXT3ecA2KUOnFZhrqCr7c2auGtrJnFVVQXUn6a2toNPa9eSmz51j
DdHJdHoRffioNuO75wJkPrBaAcuZQSF+uzlUTQ9+zxgbWMVoDlXDCEzE0zAydVpO
RnZZS7F6t9FFr51zRQvtok5KIOVxrsQa2oI+1oo8ztkh/1aHKP8ZoQxoabhBE+7/
c/r/86CB2IScyEYk0NJ9I04jb+C/GOtGz+f1/rzYzd7QMGtI2SB7YJn9NuJwWgwa
fNIMVF0IYv9HWDCzFi0SoYre/fyOASWWI2j4bbDgYfEvsEhDkMknOK3TQDLbIfwG
IX198yx/d+fXZr2XfYgrNfGaNwCQibtsGaXlNMtRwPGuSjZ9JA5X6Calp4+Mq/nA
RN+rk0Os4ncqwCIQzTHUOPIeolqUYQDagcjxwx2ljQGcyv8brdCdXc6EkXG6Ulh+
8BRbx4y7L6UrtmHBy6w9HMxYdRDaAjD8G0qMQejFM7z3b+HdPIpl89BOid6aDq0G
jOOjM7vr/dtGmj0d4AY78bwEIpinLC/pf93hs+SyW67g26p1i7BveiQ8UoSjNxPG
ZA2tzsxdS2U+t0QdrbMb/K+fYgROTqyyncbMWrkNNDYesIChq7a0XiO62Rdp5sXp
sEyzcZW2NM1UwwROKA2bThwSOj94RMJGTIan2icVJ3G1ObEdx6XTlaT2b3eo6avf
ky1oXVPZitPnEWvNj4wroXIDfzG00u4I8zWWzXMFl77Naq+jWuir2qHGKlkveFcC
aCCE8U4JS0EC7voWQ7BqjYxd8s1ZvA1TC33Vi9Rfb/iZEG5uUpRmz2WbbdOMqUGl
8w8vJw4wjwWZolrYE28jTljAj+pP8EBsw4/DoA2zzFqwLib4I1f9mhiKj7u9seU/
NJqaDPrSSXsijt0bGOMORd9wozEqvQ+jvjp5KlOlEGhd8YDFgqQjrxiP/DgnzGlN
PM0Yhz00p2uP77AhYWtOesbU+DXK2ViesJs0nPhbKST4PdFxIg9GeGR1SL2zla51
/ZLE3FwXcCmypX6KRmzEClnUOoPAkXetCIjqlBx3w7tVzcaXGj4y/hkwyIhrGcGY
kDFK5kdzi+nt6/16gtHTBkWE8AgOvYXw+ETB79rEYRnq3VQyEsZZCirvE7aEGrn8
aD0Chf9PzTb0WQyhgyFn72STfIzHoXTMakyJFAMVyxR46ubisbUmfTdYxxFuWaE9
dtR0oUdUJ8tSsIokC8fPyT4Unq5hTam1KqxUS9hyIokR3gsy2tcN71FjuVDOUfFZ
ykPmR5uE8TD4HMgWJMn5Z9zJqDA/FXBRZ+C2qepP4MqEkbrLAd2kWl6td0fSdYhp
kLCJjMlUYFDnfGblZbECCg/4bt7Pa2w1DufBDe+5zRmRyRxPD2mXdZuEDQWhXwg4
3+qRx0Sesn3yww42+Ew0KeNvJV3DltjThoD0BKj+kxMpE/6CY7kKLAtE6u4E3QAD
alvzIE93HHEMubH6vOe3eTfzWTNfnF4HYv+hE+IF3v9EdqAzBUDWVxjLneH3JGXQ
39FNXr/VoV5YjNvBHnzMU7sWQW38UVxS7ZwGmf9VJXhXyh6BKLgToJO7D+YkRdMV
xPv66ArMbPtR1RIpLBWQ2QTp+eD4m37+YklVlbRQlkMo25CW2q6jN6Dp8EzgHZAu
9K1STWHO//9H8Ys7/oVAnI/MHRfYdfwAOIBTdpuyxwMV5RXRPsBqIFEkOntBlKL4
KGEtcQRYu/6SFSZempCReGyb4AmCb8Xf/Hub6PjsDx3EYsml7jHB2ZPXfKv7ybP2
qTaohU7UQE6NuLEIlyTm9WzRdqJf60rRvoo6Q4H6K2pzBnOEoxEl9gXfPC++GeJ6
wNeISXhm+txXfcm/oFg93kpFIssI6t53+63gvFtze6SQ7M5sP/6yUHkC19apAQNQ
juvyNT6dp7Nx193loxYnBTozN090Y9TTU0Ws8D12aC4AwcJhVh3vrKTP15x1cg2O
QvG0D9WWlHmZ3y1FOEEovRw2/XPmpSO9N43gEdzRf7np+4/lqAJM8JtaYxduFU2Q
WAGQWdseD/aj8U4Vl0M68+P5E4exPh04aNyRuUb+mdyXuogKc70Ot4ofOQ0q6yQI
59IjUUp2y86SdIbc84gWPER1fBR0cvZWC7IqllN7a7ty8sNUNTepjVDnIgJI98eL
IXA6TGsSIddfOWe3zFSxR7TkYtrHvPEUn8/kaaUnZYF91+M/cW9S/0TD5cA1QvXI
LFn408oz5KEBI0znv3rcimypPQJYJshhOEbw8DAUtWRD5jzemddk43xhWI2qx33s
UveG9vLirT43bXSJNyOK4xjiMINvxbnViBjCgIWSB2aQAX4oahV7pNNWEdYrx5I6
qSe47mDri8f49KntCV22DGPHPK3DaRp2h0+4GJybWk4GLLuo3btAgQNlg8uf4Aq1
foMZgsls1qPFbfEigxL9vDNSTbcpRtnjXP47HZnBzkzdqIZCuXKd2qaZxXLfejeq
Hd0fDDcuEEVgsd0UlFODF+9TUz1nb6QNPWq8hD2FEpwZShy/rFIjShu2fYYrlPHb
2Ylt/ep1HTDAbb/p2oJ4wMN9voKiW476bZe/Ww9EepWDOymQNShcSVXqoKW67EGG
p80jdbW6O7FY04pz8UKCZZ+PUhf7jaKklkiN6zHs7Aa3NkiIJnc34O6lRzvlUDsn
uncljmaFP+9QetgE1xVR0Y6CrtCoKKLwd6VSksT3p6ziGfQw/3JbJzME5viERUkz
O7JE04xtwcUvGFhAw4Pvl7L5UdLYot/jbn9uSH6Nt4YEMkxZj6TsAqCb8az+MmF6
oVIysp3q2WM0VKmze4tdDtXf5qXzi4Apb7McrO3lKpiUatxy4yKT1rjbBX/vx3ZH
NqqbkpTraHmX0ibfUoTYdUyv+0MmUOXrahAf4M3E7bW3V+CFybSwmTly/pb9FChh
srfsbGMa8nFoj5kcHhPacZBVB7cCPKAPovTi9NJUsRNnReNwsTN+qTSuj65LOEyD
UD87sSMWSxlsp270Ea3I937RZ18e/V2nlV2XI5appkPUldgPvXOd22culigaeUPr
CccxUdYdmarNawSFs47oxZQyCohLsRxdO6XnYHPUc1laRPheLAIA3sDL5yBIYboP
427LQ4T+0fnWxKfLganuUPnLVQrPDcqfi/dphOIceo+nP25Na9APeQwRa7xm72+k
WeGMm1Awv+1Daly8Bhg5qujKrpvHHcSurEAEqKwHTclT7WNkaxjidWLsCDwPABUJ
Hp5eoF6zMfUGzlF4Ld0JUGr4prRLzsMQxOemtyrg/VKpO+T4KF/brROLeqwNe7O5
5XCkCCIFt3COZrc1iQi5X3QaxbHrI7mTLqM9+FnDqBArEa/nymrIDoIfoUDLeUW0
KGseJToCurZmWo4FNYF2lPPxgH63egAeD7+V/qQwJnvWDQBrJU0o49NjSJBGfWpt
xOprEuSuIsA7L0U5w8BSKHUjZPTh+PeI1HyY1wEMumOWu7rvpIYltOf8g/i49MPJ
Mm9ZLgmC16hzPFPerkVFUZwnyK7Dk9O7H4ZEi2BCVbtsaF81VXGDpDPAW3EG49sN
Bnx+bLXbYoVVfFqcyT3fRuc1DL89Wftn9OzPDnBTNogjGXX7cxskedzeuV641rbH
TCWZ8S0I8Et114xDPWc7jArwfNdlmxVVj90vEQ6wvsibl1RFIMI6P7O52qV9seK5
Zi70h3LviQ0lGX01ieaYIln4QyYAqpf6IxKGcTi4Z1quEkzSHdPRK0sxipguUJ/A
eTk8N7zgtFPrsQE85JxqemjvH0ulLqxIf4Dxfvx9mtE3iOr59TirfRfApXGWZWd4
MjWAf5FSrDSrLjBqOEk/x1RmdoLPYise3ru3HDyQMWPRvQSk7ssf+ClxA9ECD1LU
f64MAUlJn0/unQ1eATi8YorLWZ9WXYHL76rSnsjpn/VGN3bUqaCwgqzenSj8Vhx1
6MiOndp0D4FlIZxalIJ6DGJS3h3M9DlUMmM+FeQFzubf/cPa2qFovHJRS+xggApK
ZpKZEb+BP3hBC/s9PHJ+7vh++hFkSnJaaiC58GvfDoq4nQL9+8Oc3OjcNi3+5Cw9
2BFdfuLP9igpOK+tFdiVNTfy/SFin+kjux1rxBJrjZMqB21ZVLRKmB0vKIDN0Ta6
7mtPcdfRJtsia2wWgCBqL1anXFqOFOWrr1Y5LrurPmd2mPSzDfSLcBmKCIh8H0zj
1bVMiIJFK38d29/edNy3+eh2UPhv6qQf8I2dHh/K6xI6nVOLRcNiMe+hFVuOMI6E
qfqoBAnKyS9EFbN+GvA9g8N3ExBZUq89w7wixsRVI8yMg/zRjpPOlgTL280k3MKd
h7N+kgDQFgmhSNSM6CMmN9bJ1jaDGIzInZL70bU+U2GGq+1NFyc/noCv3tnp911x
u6wYRYThA1P11dJr2rrV+96sH0UMW2vXa5hr8+iKlucFr5Mdplttt3/XffFJ/KH8
TLR9hbbLzshMf39ZVHfL++L+yBBGMumCM84aYcAf15KdUmzY6FEGvJUpctZ6FWyH
Ryhu2rgh+Orfn8CWgqiSI0b4uBZIFCk3PottQ6gi7FMMjyqpP9yNEB9k7477S78Q
m4y9/0RHd0QIyMYh1znBxI++hATEnTfXrayVjNoJGQUCrxWV30NOadYpwMIHJOm/
r3FDvLME7YNqAA16i9FCuh69Id2vdKyNk6Yq9jhdN64wiincB9FOp9GmXTq2cJdz
HpU6SOx6Pq1AtgrjqFpQMHl7ALBlMZCm1YCvH6AiMptGjurIIyxAIxI1D0LuuoI6
rU1P1HomiN2q39Bf3BILhnhw5nO4VMhpP3quatPGS/LYpH6U8A0AZ9WvnYNgb4AI
raQwmbt5FqHsJBvhohiROHngWJ3dSqBsjBLehUrVpKPNldpI4vbwVePKMCnlw+Uk
P4c/g2wlAPRZ6vZ52OpaTYFZ+ohVzb/VWvxnKyDkl73VEpckYWs1fzAGH8PMj4uf
Y7aJghbZcqT8vm5O2iFYXWeNNujBFZ7IKjb9/l64xsMOg2geROIqr/i250nOsv0d
JmGHZjiotmnFPILv4LsVR4PXg3XUK8gF7kYe1s2XjmMygZX3yOEeQC4mjO4bYDCu
w9pRZ/btM15gTXs6lmSYCxb31F7OAEeqOoqhGb3lyVuMo3dERFtVRcctkV5XNe7y
3/HCwhM0LKdcpR5hVQHRPKzbA9HxDFOHwESozfGNRTjAnLd1qfLpweOCNTZH3z4O
z69TWCKpOmaP+5jKo1mtBzNtYCOv1Nx3Cw+Cdau/jH9EuqG/81hFNym4ytIMBCAt
N+1XtzjC/yErUQsn0qpeYhJ+LvVzGFhBfmeohV9+2HCZixvbZ2LVDslEcELfB7Iu
IjOKSUQ0rTw/8rzZ/oRVbLyfR+ib2ULgSAAjA8qZhkw30PcrLtKu/Pao+jxJSwsh
KJ9uZ7xXtsij73aMuQKWdBRhtaBk+Kjqx7yun9jnrlKC8Ww5TIKXVkmWofTxFqKm
3XhSvAQsg/rFOKm5zDSPcAyWkUhTMDipoekqA+0aj4bMUS+PFFR6Jiu8oQmc8lCk
gT531SFB4NIHiW2DlqcPXZPMIcKl/tz8VRDMah7XY8ZkH/PuA6q+/TYTJVnjZNZM
An20G2Hg819pUbOc5s+d3PhBDbtvNYjR7rrm2HSrsyxfcvcyjiKGzwEDpAZMqUmm
TL6yd1w09YrdZazs3/kT0BNzvNE+ggPfzVxNyzOLGpKnYIdh7gqle6wVK0wiQxC5
tvxOPiPjqwE1+lYENoXZ787mxTtMOQIZpKE6ZLeS1NGMqvxBhyqP9ie986otvGOC
8i45e+lk+9vWIIZFp9+v6/6Iw+6mnBqu8qemSLnnRfbU+JSCta8Cr/iDGNa1iZ9t
6DKiWTpvSMVWMSPgpg3sZ5geZtZMafGemNGJ1ocnh5QKw5EbNc3F4thPOmDtM8RV
m7khaA0ow+GjKqtGJ5XWCYBIbs2WOnzEY67TI6FdUa9yzjO0DCpyUcUKI1tTYaqG
i3QyppBg7M3grGkliRNIeLaTqpz0N5/SMXVCuFpQ7Be7i2XX9zPwG4AyuevvLF19
xn/GGKQjprj7z4KNY7DtYFy/5hmCgFD7l6s8GhTDcMDBcw5sth68DxAaMCy5ip8v
uxLBEFx/Ifpkdgnkshu7yDsqw0WOuupMyPVAMxWUEixBm8XcAt5nx7nBtuCFGfnV
w4P5xEQkonpoqmRvl3sLvmZc3+WU6FE/ul07PKN52/EBU1baBgWZjXbxgb/58D6C
mpddoHBDuZaPvtbnE/tKZbTUlifQEfrrgJN7/VsuCdPnwI2T1Y36192mTID2AE7R
99HSXy2yANJLwgePE9PUZz/PSo1KFNUTvQ3/aGQksh+gEbTxhS5nGMm8Y8IKghqQ
y9+UtrluOK+HnLFS+TxGKRLUJGZEhdtXv7pVdAUXNEbDdyaeD/eDpLRP9ax9gRd9
vy0LxYgRgDZl6gr7oNuxLyP7fGeL94G5VYEdiZego6bHgfJccf14jPwOshDAaheU
50/WE7msTx1OZ58xmVJgsle9hYFUmPihanF/S62a7LtHrvEMsHSBoKeKcsNqz8EP
BV1eQmF5Oc2DY5r3wzt97Z1WPgBULv987OWbFCsDF32fFgXaJoEN7USK87wdGbH1
Jx6BBw9aVn3iUC7MAy26HqekscGoVyCeI0/1Lp99O7hq53dYFU/cm+DLrIiu8LbB
idZsf15BvmA7vA0HqD6FjiDJhGLjy9Z8A6InzXQjB3c8Xevx79Qik5+0/lfGzx1b
fSmSNnTwq9/yIz98p9wnX8dxtB91n7AMnzje/ewOxnRFXVomw4kNv6Ei9fasrhgZ
v8CoghEi21J9kU2bne1uG3b7r+4Y0PIy7Ma6ZQoxVeqslKDPPFHJHHycNKSZlyWJ
oiqEMP8FHSVFhJazOUM+LrdRXzpBtas+VHKd4Oyx4B6+paOlMD0WI00YbqLhAZmd
dIQCrX9latWoQU3E5abMTE9jImS+sS8Oco5EIhjXF3EgAlnqEUCJ378DWB/JthL/
BZk8zwVS59IKQ+GmcfevIptW7DlmapCUURKxra715Drvs9nag9TzhVgRhlh9wmzB
9760DGfmpGCB6kTpFewZiBEV3YJX5zAi8QJNwA/BaVOmg71b+qMfWPvMe1WuFW6c
G++9RI4DqlLW14tl0Syqe8qOgRMJk00NO/+irVoQGauohCwNFEJX97ufnlozQj9b
8q00Sf3aNjMT5jGgGUspM/kRulMZ0UAreUwaRmgPzmbDOi9cSsAVq2nd3TRRWisq
kIbmF5VaNEkzBxFY/6USkohDHezzcXiSwXqkzNh4XLxIBmGAQcgqw1Q35uqUzKlI
oJvluTDzA7+7fSQltNZrVHWYg9+SoZ9LXjVKt/69xhRGDy7COX2FMIhGTJR2K7p5
Ovs/Bt07UnE/YTZ7wCMYeK93QltznnuUcJUfQbQsQoxihic4Q7jlCScI5V0jdYdl
vWHBvvXW50NVASpYDIC4ZOgp+neE947KbK80fqcfMr0Jxm/GvMiaXbFK3y3IztED
Bl3LsP78LE7DVqfS1di8CvsaDRrq2uwNkHkcBHRPWmEa752PIlzUJqVMU/7ahAzg
T3YnPwmYxjDRBjE1LUHhpLAMJ5hxf7A0SPKFo841KskNCPHVb0NlKoUeYqP8bVjT
GkbeSrL+eGM3/7GVo67ulqzbUGJdBeG1uZvZKxT2W33qiB486O0cIBNUJwJqYQqt
ToUfKi0XlXMGI4+i5JL5PbW6NHGSYN00xN0ADzR5WXfnlb0yJgxxwTQBLmF39gdj
3ac2oFZJogh823m1gB+1+4rIbX/KMsgfbVSEfKNOtVhYmYrNBO5xAmFUO+RshMRf
WVlUwnl9gUNqKC6qVLF0xDjkGHmyzzfye4JRPuXfXx8dTjHKEJ7aHs3gia7parNq
hXI4kvMnX/EZblZME0YWdZ/81y8EZIBO6vnJ8ImPyMD8I10kpjWqWsONU5bX61Zv
mtBFYGHEjrCIyPQIRjKIL78WTs8iWUCXHJ1dzQgVCEhE9FwheDQa4UmPkrBSJoqq
JjhZlLLq0DDrSbFmm3lYqHNOMyvvUO6/O2WA1reMNWjYFSCvNPoBRLXx4Jy6Ril1
Y+ESETSpmOKfuAn8KvqFNp5hUnjSoFqr6x7B730jMKkGVutM+Ei22po2ieJk73zU
FQCk5PXBY0EiEhNcun0Afu5ay/rOasE9PmR0azXUTepw0wXsxJUeq1eAdqbGOrZT
PdxkWWBHMWzzTEh7yiHImVX1Ffphwdvnqr5hLyBwbl0WqQ7bk5rdoUjRm4oEgDdK
CpVt7TdV/lt3TkvoBKREr/aqB+7ACRm51GvXef4zw2xMIaIUbGiTflmWbrW7Kh79
JBiPUY/d7VayEYNETaoqvMqQhXcT2Q3aC/qTfRLp/lnL/21yus10RkHjSb3sJLXZ
NAmBye4q5v/YPrUkOXOue4a3ictGG4YKoH4urZtbTLCQ4KGD9FctEZS4fijjwyCh
gz9Cn//swaC5GIghdO+nkF9lFo6VG7xRC7ujmchOsKNajwNebvbzxWdM5yzgWWP0
RQmA/3LPuLVUVxZPMKROmP3YPK/zS4FkLxuf+at6OnRk2jBB8EeL6S3jtPRY/bqD
zDI4thHX0aREB7+a1b5Kb5pDbNbjyFrqln0mZzXGREPVSOWRfOF5/F1e07wKBI2t
0TPGggF6o3BFeXILQAUHLBBeTHkfAnqHldnvgwWSaw625tmsA29mIuLeAiD5FkFc
pn2RzYb3HlZjK8kahlxGY77tP2VNoZOttxGYPCmA+GQWZ15Z4QpsuJ0IjmqEZ9N0
mD/nX/Oy3CQF9n58T6jRDT050vqtr7rOC0tEBuRS5h4dQoylMCcX9BciLZ5SrOC+
xNzqKhQIn3lLNHSaCUoxtTF5uVAEZzWlvlUSHLrw//AXp83Wvp0pmBvdvq78agHV
l7Y9sQStlLLK1x+Q36GjG5jj9QFDyL7jEURiFY/4YVlhlkanAZjEnzUX/yIqrNDJ
RwhytMmWy2f5+o9/GpU3zPihZCKum97e1PUJMyYMLrGsgTqiM+wJACsHJtEFSFKM
FuNyADhHGEmdeIehqaxmNCFZGeEg8Zt2XxMIVH8nFWNVtvxNh8tlOAlXL4U4cVuj
o5u9CtwoMuPhXCW3sYdgBi8r4zZ+JUJh4fPk0fW9mc3V/67gCvADOb+2SId88cEa
NfanFO1Z62j1RxMvJW1kX70G0WzD0clgQeUtdA8MP9nhVtcyOVA5Pbsn1pfVSaNO
c+MApkiHMs9l+2gBnNal/9/DN+KHuzhAH6YC1I7K+zz3v4wV2i84jOaS0+1MhXNs
4TZZPJDuVPxHp/sBdTDq3PkGKYScLh+QJtUGnvLV66v5CIaZ8gSjYA/FlatltQou
DAjX7Q4uHfC2pxjpPXHucSL1gjrBf5pqMy/WWJ7XMew9Ftjq02mWmx04+gKvy9L5
NF+bCtaCThlslZdnejBpgYuNp2xVHrh2aoF7yJkGFzjEbfCUHMAUO2cwKVdvdfoB
z8Hd1lVchg8DUbgmWUb0mtovm9a8KeycT7om4pIT0InFQZSL9yrhzwe1caSMuH67
PMMC6Nx6YGLcEaYRyutry9jhMkaPYY4RhgxbsjjRwP4RTm0BROpMNRiT13rRQr7B
ePJLJyALb/YOxMv73FCY8QG47n0dtQ1a8u7QNq7SRGAbCXJgUuVco0ucn4K1R/6/
jH0GbFEbXoSwORZ/2u5vu3h0xfN1J5BEVTKWMqxPYjNXcwQKA9THeTGGW/LMUYQo
tEoiGKKuXqJBeXvyTCYW2PyQhyx69+/IulsL/wNR46UhYOHT/k1zWf1B2Y2U7g8m
1czx4Yt8PrNtOZ7VmG9LMkTyzCA1+B19WzkTZ5JuGkLVLNQD5ZDpZWc5gZ4ww+9Q
NcbNEu9gOj3uMoZ3jK3OkKWevC1tQp4dlXOcoZScq4x7iI6ak4pGucPQ3AcWHj7F
pMBxY+ziShJSbNBkwVSt3iPkpkVesMkalBif1qbmUOKmGqYGd5eK6+UjbvIHwRTH
Eew9Wv+Drlqi9BaQnHTN8ina4kLdckZpTBM1iICLQ2d3HGJCxBnaLTYh+gSSrywT
9Ly/ouTlbzKV7XlP2cRRQ/eMNNpYLlFphcGNtbQMt0np/HwGkSIgf1xvn5QUDhaT
ss6iFj3027/GxsI9ij5oA3r/LcKQi6zA8qmr/bIijW96FWY6weQ0nnJJmZHPEwBE
NrvCHAwOmwwALl+L89tBsmX4YzJkEflf1kfq4Stz/kA5v38vsXkLzuqO32o9e3oO
cg4qdXzS4hWsvNV7DJUy5tONJwgJj5sKdMbn/wYSnEklyvPOTH6aYl4HAuCQyz/G
RHj5VfyWcxgjiAejN0Jn2/IHKL5v0tEGpATMnSULsKFa73YWo//REM3KoV2W/+Qt
kh8KFs/+xWWBe12MCbuPDEZC592WlnvDDVCjzzVxT2ZNpCoW9DVDV1jNasEp0Qw4
r5eO95miz8bbZ13nc0P0KKOJSs2+xmxVo1L/wnmMZd588T0VnN9HOfY3jPJS1/2/
FXUfx/kiG64SsV5s6+iwGy5/QuaWnhiCIpt4kWp3mL46LIHS0sSjyZVVUWNWGqLC
rzagsygyg7G4aK/KnmlXoBJq/C6yLJH9/ILZY2WioU36pu9Zhci5z3tKP5TFKCjt
ufpf1N8+/LPLsDQoavlUzfA2j1Z9xqdsmvdR4Ng+sMdiijYiybU75L47QsttKQ3D
0xkHT7BE8YjwyK7LmRW1e917KAw7dSsgr9K7/6kCDdT4Iz6DiGX9nvsHpJ4RrtTY
yQoPx9NBIKE86VASlLkTtZJcFgBGPyFm/XgEMedqv03EKq22hyMB5WyF1JGWo7vC
9PeSsIDLKg07NkUcYC8ZmSjAbAkXol/9xWApztR6lEzIWPedbVuVa+nNv4e+hKrG
3OOYF8WgM3Lzq94m3O3DQWZEbcfrkusaNwxrjcAJU8qK6Ym/s6C7FYnBg0uwhHd0
b/7Gzg+euh9tz5naN7uYDdByHrk38qetqMPKNKeaAmjVhROOVk8KHNvDRD5ogRnj
i+5jhWsLJtHoWTMON4AazG81y9ZxZZWVQpj/7isIh8lDbKtfZcgdy+DdPe1aVGwx
2Eq26FhVYgQDYx+3EfhVLzrXjK/8wa4RW26hfIfapd52zSlAyA0x+D3JQHm7iuix
Z6x9KCraHGjEOoSEZ3xIDi5WJpmeqbCLFe949Z//gGl90mgaJm8bNWRmvESee+jp
CpSKsJy+wdjX2nDV/zQkaCvgjhDULAYzEr2fBNZAy7S81/HINGMiFmzdVYv5QJMH
/SUj8Edw5tq6p5aRMEQq32u47gCiP541gsaF2GzAOQzuymt8uGDbluS0KH9fecL9
TSlAN08Q6PhimI4OGQCOeHYNvrN7PLjEURYWTtN6LwRjFGtdvZzjyvtxBxVNoFTf
txtD9GL2bhNxqnah4fjLwUowoj283FxQxx5mk03urgYDml+9a0QVXLaMcFpqW4p5
Hs1gKEM+DFI6FE1URM3x64sc6XA2jQrQnCd1lFHnlTsAmED48QaxZSLYIRSPBLDX
IFw5uStLm82buUUYAa0o1sjB2cjxpMV1lM8uv6PpDTElVP3z59+F+FifhdRvuq5i
ndR8iT6qMR3Sjn/Mq4kBGdXJ+MtNX9jQT9PHR+q02xhi581qukEfas93J7Kogh+/
x4ihmWMCARPyU60/I8M8x8yIBA1NA4/mCDRE+o7m3iaM+Z4V0ZCxkg6mE9k/qSEF
hjCgU+ZlZuJ4T6gi34dD8exuVUsDYBlldETFAusJXxVwkG0SxTAOEJi6HQAz7HvU
V89Sp0n6xUcdINl5hMllYYvx0Mm17dZzKJL7RtdvTxXF0NQA1kvA9qktnuflUicR
w57vKSLSXDwFbYEOOo9GAYB4hp76sgvfy/alyIbjfwb/s1lubgndMJ0jUKA7yeva
AhfjZN59saYrhruTzvO2bzXlM8cyoaIgBxZyy6vAM5r27TT82Hw9igR0MGJnV1tO
gTXfg1GrJLpq+RMayCXZELjhwduxitXI6Thp9DCgDDCW68OZbeAiAwhlAOAV+7rO
zuxRsDvK63a8m0zQny7UkzQJnLXyjeB5X/F0akBjLOFXfSaIfXlBxZiBX5YAyVTV
uKfT2biIRVbMGAvS6Qmj0Mmmn1osjjuWOsHLaiGTGFHyZDRR2D2+rtT45B0MsikN
+4a9DLjFAd9AgZj+bvLp4PHvEDCkpKxyOUL9qS1DvowwglcUzlksG0onQX5D+864
DsW7G/U6wbIb0c9/m9auF3AnIm9U2/47BgyNNESCfJ8kkueTYqwKOheGxR9F3/fy
+L9D+Xy5eYrogG+CaO2hJpIZ0rrUsxalVFajt/zFF0/GafHv968AcxKTEDLy4xzT
EesmGiACnu+ecvQd3PmCagnaGzvEOIsi8zLK9TkgK8Gl4jUXBl93FlmFzdzzXMwc
J6C7p53MeBbQCQ9icVHRFiDxqcOinAP3a2h/4mihyKwNYn4qpSLZtuDtXQUHDsnB
42mGCbsg+uuKBhBwjLd9fKmH2B8Mfx7BswU+BpoIOLHa9iq9VxXyRJdnjYCWpk4o
EyO/I2r/JuSc5Q3WC7sU6bdMVFMD1cizizj/j5z0l2WSEuiLze+4wmpdcXd9SwpK
VIC3bxVCypL9erFkqUI7fs53U69DkQphfgM9AXlTTxdWAxvNjKmoy8EQLr1Tbxt/
ja+8070axgzwbrPwrsH/iSqAYfM0Arh/OXYucUlnaG5nnZdf6IDhoKZzYSGjvYI5
hc6lf3L60EJuXEjfRMJFtnuIh//1712VWX33qPGZOkJG7YFlUwWlnnoW0ZdXI4y1
eedrlTG6FRHlF5ZTubofxQM+Y/z1/jmBy/dxaj88P7ycTo3kiAL9Ziu7P/4MMqKB
IxD5L9NgSJoe5+L+Sxoa056FK6tlX+2EekTpWTbn5Da1pdr8vLFGe21Aecs0P9d7
rFCVLafGgnvTvgnyUi6+LQZXY3hHwHvBQ8jn6cIketKWcyppTMOgr6hd4sbndpSH
Upv4ze5J8Gft78LXYDaztdq6zRQF3K7vX0FYp0ztVu58V+8V6BjZjj30S29edu+V
k4gOloC9J3ISYPB/47C1HOhr/fG6IHnKyUqrBrOU9xquNUz6/Ci2iAgImjGgX7Ov
qxfirVdF1L6dkYToBjhLewDow3cZSaCw36u+qBtUEcJszJ3ew9R2+BGtylZ6UZIc
1Z1sSJe/15wGgpjHheddSEUwY65HIP4dhutAtLDm9GKWbFUapYOxTAdpDp2uJ457
rU1oLVwHEVLM2OFAOF+XY5gF7T+WG86Rk8v/rvy4N0DFuTpaBDyFYs5wppQD/fJd
laDLOPOAfNUVkUgjFSOiyHuogg4IxelNeLM8ZmdiRFxOXsJlWo1geG1ZMXOPOKEz
iqMpa9QDy/qCQWFuNNbq/J4auB3jdQnQr4v+Te4H8/LtmlGhu1rzBcIxvvTQwxie
4JnIuMv2+B6tVKXaVplt128b8tTNE4NkEL+JHyYCzHZe9soj554WG0n74ir4zlSe
wjexwvc0nDeZTy0636pWcHfL0wUGsPoB8p7qN2s6hIDnufjKfdx0vrmEn2KInK5x
lP+1G/haWO71eVNN+jr7w+7F8x8WobhVqf39YBgtj5K9L5ToADxHA6RA09rpYCXb
P6pADEvEj91xtUED9Kokq13C0INBWGNeibBG844Cm7iYMwFhCzPYyH9rLmwYxR8C
ij7MVBnZGuY354QRfoe/bjks1W0488rgT5quw/r+xgCnrRbzBnJi23++OdCvcl3Z
D4mrDGVR4c8qhUw4CD/kxUcoH1nbvUTqujfk/hz+6L7DsmINFhnzTsnwCk1BeDah
p66nkhmf7PFYGHu9xSBZEtjLRLwKv6r8ogPD2XLNBz2kcoCxiieoWV9YtzYLNOzx
QtTKZL7r6CxtNLjxwv9eFQz1tVCCoKxtbjnByQDHVFZdtLWtnRsMPIkCnJwUzeve
U7ro6tVAbyV6i4bGowRlGnQ5pA/GDa3G/1e3BAsmQHQHdnvZbo2oTrHHr594dNTF
SAmfFTaLn4KTCZzKAqvOjS6evgRG5XH7dWiR1vn/CpfHHMQsetA9ZrnBW+fpPzva
QiYaDxBGKHvrO1ZuWHwFx5a12YNj6WuVHaOMPWOA2wC4xWnzvwSblMNsHS4+JSxQ
8j+2lb0YeGRFhlZ0zI4BvNAmBEtHWDG2y4nAiiMlutBpsL/14dVr3BFd2VyEdrRq
xKvXZ1XHIbuMPu/d2GTpYxShwUitv3K7FcLZZ1vSj0+rqQz0tahqqWeJX6TgQ3Gx
+IT0yman8N34SrxDZ0oC+p3+Z4MRgAIBrLTaNFtishAXm+olfvCD6qPD26Aj0H2F
R3k2IPFvyFBoK8lR1csQW9eQIKRGfHdMr4/GoDDBdQSlXecTjAOzTbkzLFk3ZllA
xM8tUP/6o1y6EENSl89I5FKwlbRPiGvel1Ky3/xIT9AAbWAHyNqxQItvrAFluDim
2sVhNByJcKWHxbblmxxVozkVdH60Qupw/zQdPWxPVDdntqdFFGJq4tch6d+FKXIn
7W1MAAG5Pzq/YuTTv1SHVYzVs8XARGigsRiWIK/iJXEU6he9rYnjvtZvrc1muONR
1KwvHskgGL8UeUBNnC1EXwxAvmBqEPeULRNTs5X+Jjo+9BRtteyYcxT3sj4xhOIE
rDq+X6DNSlodrcIb43XAIeX0OCOCY0T8U+q0d9tMKf9UAv7h16YI3GED0Y4jdvGb
YKxH4JN4Pqk54UP7qKtfcDMkLz71UKzqhIy15P+4egcCPidkefDQQ3doEWTefYr3
aH8ePdlWWNDS8PX14JJL2DWSuPe4r8zBsUh3FXJfvLuUUkVIHO7UeVCCL4NSm9oT
EN7AvpTrpHpbY2PzqOXhhoxo3ctSywNjPsZNQjCKNQLKQPGMFPEMFXkH3kJgEK1K
shduMvCmXCh/2TlQRqc8ikjvUHTdWXUFbA6Tzb56ZWyDTi7zxoMwtbDoFv6KlXpX
1t+1ecfNgp0Xo6szdjqUz5WhI/erdh6C9jNFlXB5bYZtxT9b57kd6xpN694p5oUl
Ryukosx2yv2qfX5PueAcOsUWtI0NClox1d7/rKJGev9JJh2/9/4FrgWf5MEEamJj
dtzF+mc+dXUi7IlLQK5tnPXzhumgGEgWCvfKndIi8fm57RQeXZXPmvq4LFkwb+Gy
SLeDCrE21gpOzNdVh48vE2FCuHxZTBCODnWJugdnRZz9RHXoolF4Akgm/SglBFYQ
V7VskwKWAPeoRgDORtFD9oPk9QWvVIkhQDzHgbVFMJoXmvEUaGj3UKKXBlU1TDCd
2bnD0Jzl8L93XgiPLjQ0CP/Oo33hSofwf0ECdo3erR559sgekUV8roP/Y8yXGxeI
Nae5FZr5N62t10otoGr5BuCZkhvUA2TJiuf6WnaS689GnwPWUqh8kJKEOR2zXk70
j8rRBlFw/9fiRHATUUELprjL+N9aiwIRcUKoMejTiE47B0nQUL15jsuMdZvJzpgT
zr0P8v/mxJ+TWxDJL86DLdfj8QZIzvF9SECs311lBDgip1Jcp4YFcnZfCP6PWYyr
qeG2dz9PiSWEXOKoOfYixjYiPZjnFIDsle6FnKunJ2JaQXJuba6uVWYU1afGKp/w
rc1vUooYSnpWQJX8XdTZwvSXTId+QJG9xXB52WQihRveXGUEcmp2ypaWJKpGkmQS
PTeL3VOA57HZ3/clUMrwuDZTRBJTGS6gY4djdqDJv6sI5msWFaReGF/p5Dk3qVvL
GJ0YiQi+cDRKeCUNrsGUoBqDAc2TDeELhwuJ52VxvEca310YZK4ot6UhfUa+cRoH
8+1c0Ms0xSY9+DPSCYQfgOmQxGMchnWQUkSSKSKuG340KrafFMnTROpMpfbaFi0/
T5Jk5JBjIh1KaLnT72c3s9hZZEQdHvubHSOHR1jjN8/E29PKrsPDeh0g2zyMeXXn
YjD5HonbZfYPrOBTnTmGPQLHrMToB7PUlq0Oo4785BbUkIH7RJGMJWDb2aZUuJK4
1kdJr9Xn+Q3IBz/ik1R2EHkFW7HwhmGDUMGDNMMomdVve/Jcu16UYsNQdKa1R1xP
AkSPwv2siRZxcVpgLqfGFqStAnoImJz8twHx3T6UGy4cURKD2u3ktfeSywoebXoC
vu3uHETipf5Y6gzBunWVhx4O1fA3JmiMSwFFjvfoOkya1Wr/m9w/Jl3jxayEK2ot
gFq+NKxm1AIOfbRHgYVAC+j0+s/ZkqFEf/R3yw7nNorvLDiNqnHlQ8i0k/Jy0Ba2
abZ8NrC3gN1hjC6c4g9DRYTWhIHcj9vbFx/zOuanvnw8QvJR/i47hcUjCxQmauVY
8caOJblb/4AElYOLGjoAqi8j7KJEOKW7kHHpSAGnqFDExeJHopEFmOrJzWqgAhC4
AoYxO3Yudjp+ygshTQDMI0867hC3l9SXwe6YpSVDuoQ+PmQX7TeSY9H9uH1gAk86
F9SnqkfZGAIToktPbhq1Spl1xm45ui81UhrscUL4kioXAPpTPYD3zREfTFkgNnfI
R89wHeJddkPC0NUyFGuE0HLU5AsnBrM0soO8OStSOiGqwn/sO7R1nXwJwOj6Gmv4
ZF0lQIO/eWox0UPQzhat/lYULwN3pD+xP+MF9I2/tvgEeDUdcLpJObBhl90Y4Esl
XfgBK+ZlwjaDJm8k4PbJFLOoYFK60Wrh+lb1waIM40ovxw5lqORIoKEMigb0dJ22
B3C+EhjkHxwonFtUrW8uLmdnH2VrD6v7G/QXoqQ/FWwImLczmZwDqkmgoodR+zWr
iqiGpPWTKBej1PQSbo4ca8LNQ4+K3FKaum6Y3dXDD3cYamoszryAomJ9o27Mh/xn
M+YrZxfioTwSLo+rOz4TawJYPvHjJ2nyM9Ks8XtoA1O4eO7hmm9VEbzJpeCHZ4Ju
5FSEJPglotEaK3EQ4+M/MqtDTkXNXWqjwOUM042CeDau+K+AOyLHoIBkkLjt8OfZ
J+I7HV+A/JVArsXz93tuaJjZU1m/VWOfbOhq/rpRxd1s7H+kOdVh0AJCsEsPVjq0
u309lcPRwYtqFbZlWbz2cRDs3Cks75MHKe2flxgN3zQjbE7WXmEnn8BBpTalnYBL
+JI91PJEUHi/NoYQ8F7nMCGkQ0grazOkySGNoJLGmxpf7XeUHxOzsRkpjPz9AKzd
ZyeJiH02654VCv8Bgty15/adMHrJjC2ClQQPdtCmHobjE5wAGxMDeBRqr4FKJFi9
uowmhLT6GAaQhSZ10fMrdN6FTq+cwW1fKZJYAnQhH+Fb64ZO1NzFKPjb3YkyyQ2o
NsLDYx9ILWf4JnVp+dE+esbYsiLuFwjEwQ/F+LkXekGvRadGyJnmPK57zXRUJLGA
R5/D8zUSw3Oz6MV75ZNj6WLsOggZBmi9AUvZ5kPFrCcwUoXeBHfHUY1PhUaPjpYE
AqAa0kH/FhaNWQP9KIGQ+NrIiL2uZlGpo2LBIG35vC8ED4wgJkiOns0yxcJMXURD
Y9GMYqD6DOI7/P3u650Y3kGRueM7WK9VCR6y04Fgrxm16dqp1CVktgIQt05XTqpu
wCDnBDlO6QfAMYrzGGeEfjG/Okz+ozSD/ndYfvn1iq2+cjzcnmXYDRxxupIp6Wxv
VIO9lWC3VgUVcnaUmQY0ICsLekwQS8HpBmDmIGGv91ce58xFihf1e1jEvpOLil3S
JShXSQxusmLcLNKu04dtbY0dvn+za5Aw1Uwl+rtKu+wUr0hrOxUmjj+y5f2Hy1qV
CT5ATjDrtuPfyKqafsCLhfIFpWksmCURaan7mvNdlPEcLi9tKpedjN8tI1R/Xm9k
2cYvfCa3W7uvZucOrH2i/1IrGRVbZ9JBorsNFJ4ypOkG1QvC/anx/rYtjGHsBUH2
NBeBNtyzcQfrFwI12XEgtvyT4biIjVASBBhzLNKZwqaL91kSO/GzqJ0DP7tfT4mk
irfIfI459yqGaFUhxwX3KylGX6V97YPWr7SDsE1S9jszgC3bOU/xmLj6SUv7Tiad
DwNZjy1HzwGMRa+dtBVpt3EnxY/E1f/N6RkGTFrsv1UMMqbnluWClOenqTdWffPz
Qt1+WsbM1KQlffwbXnAYnBPYTfIUXnh7zZEHrlADSPnuadtsRAHt3hqQ85EGREeh
+Tgfy31HB3a70+uZM8oRpnucy/MIJkfHxlgmFVRdM1yIocTRNY7vRzS0/MqEWnAI
grZE6X0KfvvVzM6TWw3E3hlAznck1YjI+iZhRhtZ8nsEnLZ90RGYUt2evrhhO8ZI
HjczLVTqJK5GWMBX30x1fTHF0ToZd+kd++RkMHrkHj/OBpcbba38lBTWVlhrXUup
gVKrRwN6nKYf64WFJO9Fm1LHsOJN+UoxdqpbV2k7G96jSQSg3YHpm3dB2QUnIh66
/DVqO3zXXjcQfVOKYDVj5JgCyB1woavnQmXK/lKF3Crtnc/9Rp0x39rilJchkmGh
C8wDMoO+S9wAtGYpg024XDohldBs9ACAseNgTROmKz35YGW+IZJuE9nhva4yAnmv
qVJ5Tpk6ljHzHMGVkZDTSg5sYGTxBdjBXqE7Hh7G2HErBPWlEjGkHrEtoIml+R2X
x2ZjnTA+R7QH35wTwxQ2HXzmTWPSuStQI2/ecjpKGKr9aV8jUyLPd/diOHfGo4au
RfBSLYZ5IQRhiWO3b8roJQonuS0D2dktjrmN5SER9zNmqJa9Z2qeuULZ/QklhGkm
ykPHXPPkqWNfToq7LCjPdkcJVbInwEeAK3lHuWZ8ARNJIPchmSJYj7hsHb2GP9+9
dSouZl3hBWIoVR6o7zQN78mCPdGfhzhzBNyfSptaxQ1JxczXA3nPh0Tg7b9qZAkT
hTiYaAvYeblnIztY6epjq3CWUaG6IoiD7G9ZhAoAr09HSqTG6fecNv1s53Cih/U/
fyR75AaxJY6YMfMS/Km356v/OoZUuzmJiD607E3OnyLkfTA3Qr2vphaKZFPGQ22v
WQgyE+7XMYesVr1AywxSuqrqbm03urhq21Q4jSvNZhIwJ0STdZtJiTw3mS+qZMTI
3OtefuAQh1HC5D8gC0mR7z6yElDcQQPDDHjlr7eQYOJCTMmhXvODhOajnlnlSZbQ
gqLBlMLMQmmySRWUoA3LLjOBx4HiLmvChwKil4OOrGv1pUCUsXH5vVXdbJbY5KS2
lf3syxCz04ogZPlKnri4mu9HShaPcaaa7ZTDb5r4PchVDnwuQeqLxlou9U6BSSOQ
+E6/cfYIW5i0tufG2cW/53KpR4rck9KWhwR5Z6ZwFOkgupeqtH4tYauDuEwIy60e
wS1hiEzjYbQ549YU/riPcC9jnY94/O2Beps+OyCweiiXGm40GJ9vCL4Dh7MuOnj9
CUvq1iMfNICx0Elo5puAi0lvzdSRE/XIFXNg/YvX4BH0ZqcGmCEw+pLwqAvyKSg9
4ca0Yil7kAkOnJ1I4HHcn4J+RE17P7AvrA0g40KvZF1X20zun3YThUmQvnP5KXrv
UxliJKzkKBfdwH++HPRT96k23kzg1ossN4p+n5A8XTENcglYn0bI45Jz2KQnlq9M
Drs1GxpKg0aMQxMH5/k0Oa8OuR2Dd0VpSupaLgk8Bx1mLk2XXp96W1XmdDzMhaj9
I461S6AUOmA0RHEj51XrRX/Ov3iYLi0A5iNj8gqBqwSQ7CoWq648G5PCJzYww2vV
S8vWdADyYSahfjAUYjlgTgxa15pJ72iK0bQ6num2wl7t20kiDAdaN+3kViM22sDn
vO9RNyR94uMyi+/UsyVNQU+oDwhXlYcPKTLg9vHWtkZOvvRIlIFcDcXBK+mf2lme
Co6aKeiWht9sAv3qG+6bHeUOVJ9LsczV9HyIA3xXqurKq1pFMaRFhJswKTByJyvT
QaCVSjvb/Ta8PslbYHvShktcO2zb2pgfK16Nuo6rzrCIvcmKGgDituJ0dQmGwah4
a4mjnPD6nIKpijtlBSfGZFte0haqNiTmic0mJRjLybbv5u1YFXHCMZ1a3LVjwA7e
uf01fDtRagSZcRGHNhLq163idggsSdSBdqmHV5L+fcsqul83f47iI/6NQRvyzw7w
mG0dXnBDsltLC+9he1G7NdTMnRlYQwtlO5TmU67CuZ45K6rgVagZVW16SxcS6mKk
7I+L4sZpfhdKd1wAoWQXo8xeVX5NmAVvq6S+2AujNtchflizgYqMfB+pnZaIAm9L
tkhhw6HyLXLWq31x7lTcz6pZhcNkwYvruHIcQ49v+/lMD+4IZ6+aHF4VfVVlj2+F
0CwGqq11TlmDAKspu+LbYjKDc17GsAJKNhMWK6UDHvWFaKOdzQIPeP6PhGRgr72p
kLW0f3JL+70OKW26TeftL4B8DGf4KT+pa0og9yogZuNdDxxtRDHndl5KR11ehcm5
sEOYk1MMS5qd3SZwDV5o8uePzywbWc2qlMY24hJ5G0/H0L2MeXZy55XbUhiu+AIH
aPOoMeQ/wjR5UFwM7uNnjxNxOhxXhei3OfndKI1B5onBa8dwoKrBEHKyJrAC/bui
R9v58lYFt0JjYjRDNnStPh5cydi0I2oEV1h9Iu1i7Mo0QiLplbpdgi+RJ8RMXQgo
9BehARV/jimDYJ7Iu5I4diHP8LLBHRjJC00xouIjWq6dk7zpI3MPqJci+CJurudE
LgCDQVVKmWkNwzSHOb1fycIxoqAwaM21Yeh+k0cCb7Q1iesRoIQ3G+j8+qIlOaZA
/AG/OOfj1k38yRfLTwFY7gimrNsZHL9AvX5OCcZrn4H86TFWbF786RHorLy3KdgQ
koSSRVHyHGe9cEK4kRIFZmWjItquTfnYuLJ9udXVTVH2qvx5X9IhHV5VQOW7QsOb
ETGaEAmBb7yIZNm9wJ8Kgg/xIAG7jqNJebeN1VfKiFRM00aIB1sQCbnB5arAHq7U
HGZl22lpt/eNz64tn6+pX5w/Kq47eD87qPhcPxnERutg9oATF6lAkVWe/eSVsxrM
CuqisjVZYp3+0gBs5meBBrUdHaasbKKFpL6tGConVE9gDjffaoUtRzNdPlX4Vk58
gFTKMmDmFQPgokUMbGLaEH2q7iP8cy/lY03kYtXc70NIFzyQ6IoT6Ff60jYTnyr+
VEj8TlXhnaROzEU+7J1tmiKe6pWVPL/+eCPAGA+XmTQIpaAjtFK+RPXUtwT4G0/a
g8J+7nCX3nVQCHl3sqT3tpay8TkbiK0FUxCF4nCOd6pTo8ioO+XiL8ZzEn+azZ72
2hTJOrs33X2DARQOo8/zspkepswWb6qy6hVYQ2cnPWLrxltSvxgbYKfBanxegpuU
ScWUv7P4f6U0o8HOd9qHEpsKC/M0KAvRPanJgE+PskIP5UcD1NfhhSIpk2wMeExu
4bA8hLWUFyuOIpXLwwFFTvLK8Ti80g/TWBoe1O1vHQDiYzunVvbKtD1x5cJatG9L
1RE4F4Iqilqk+FbW3H/L7VHrv2gjgCYPEsOOPexBLx5h5Pho+dO4GKInIsa+jmCF
vsZYYhkc85YO5/T1nybXmc8VTemMoFL5URasFql/zPzPZUrLCcK/gdJjW3U0MG4e
vcE6TkcyYkVs1iIJg/v3v9BQDHY1I2IQAI8912jEqPXB7gtzZaarJtSxeEVY3ZhB
1FsW+0ylW37WExGKBx6783knaza+Op0AneeXt3Wyn3+E1oG5kG49W8hEYox2ut+O
nGu2pF2MWMHXyE90KVPrP69F5+BI6wuwEU8n0w5rFrQMcfqhFunvDxykTC/TH+eK
R1K+9EMghT7U/QQ6BwrQOUBurHFF/+QPaJ3QJumQpi/cSjcnPIz6mZwkB1l34PSN
cYHQZO5uMybTcRKJBDEd/U9gSpC9qc4Ei/KW8WlMpYwNvLeXI6qSDnFMKlfCuOyv
7aikKCV1YjsuLCoWNGZC9k89kY+tjCfkMdH5MkO1V4Zpo/MFD4BL0RPrKwUpNO1A
90O5PpPGQ18JChrFxYSbQU/e55qZA7XgxCb1j9H4jZnR1AjKLmv3M5DwlM56AYzm
ZDRtIOCPDm2rgpErbjl3daDFQhh2ROm0CiMpLOZxtgRr58ITk1MlnFxpFftcdTwf
I4MweA6L2Ep1JZEhEcwrd6FoA3Ll7m7Z/NAe0IyuBaguvD79msiLI+uKen/dc4UC
ZH9/T25sm6y9lDkKBqCVELWV3TGWHLMGvkP705S2+/Pkv4NRrO8uLEyeTKyTZXER
GH1SK7KCag8ZopENcX51SuYgvm7Pnpd/eFji1e7ebhiCN1Gnwhpd3sFfIsjmBf5C
D60qNK5E6cV4Q96DIs8zT1l/iihgZ28X20FFJACnEB1LLIBrmJzgubOjBuZLsl44
lZqAjq2agfm4yo4FhzRv2JBh2KAEvp99bmkabszUb80fvB5/961kp5VaJROhiuDB
4mhwFwsw3wRFrN4MboXJ7f0J/coN0m6PeFf+kMGpb6gtMbCFLD5uCqIfcsdrAGZt
Um6I4XMlKWOqBeCk7pvmL4Y8+N4/au3zsSe0aM5CWmJohYCAhRMi38zKRw3GPp+J
DjFRh+Sf0yui2J3Yf/MBymqjJeMGUhG36KOPnwNyRgVQxBk0bcr9WOeJvMJDOPh2
pn+Hq1XX+QZa6pZKDnbiR8LftwY/zDTUmq7Xtz1hHjc3epY3h7mtK/0YBr+5mD9r
JIUFavGvDJKVt6pb+nuaQbky63fXrz4kYcQEVzoAEUuGlb8for8yy0cXA7aWxAg5
vqdSqTPZ5EG/xm0NAO+PSS0Ib2G/GSaU+3Rdw20vTg5lVvrUmkuW9pkp+qhUAHdb
K4/nafAxp8o9BHBIMxrNXhLIUs4u6LSiOtTdMuzEQij6VIm7Er1xsse1UeybNd+r
SaGhYhjthsLAuekQo/V81RIBDEK/XOzBQDrG9yacJaMkQK392izw33VknFd8DQ7+
boyNacj7rXI3adOHm20CTd+2lotbLAAgubNE5CqKYyUks7i8J/5GcOc0vqaf4D8B
Ooz87i4dtOGPhPJZFoy0d82XemH8cZsRSo5pZjntPBmkzZkrIvnMxEvebEFfIj3R
465yIjhWDri5A5rwAMj6yRrTSmznFpe0ZrZTXpwMkDvi95IT18pl4pxLKxttcvYn
Evb0aqXUfJkwUq8CzHgUI8sPXdO53N5ofbG6LzcSbqbk8oyhKn6IFyJV5wOGY/pm
uuUiade9ZlXkT3dmvcQBgPd7UUXt7B+pd4XTb6M7JDd5WPVGC5XZXjTB6wFQ3b5r
U/IqYZjpKLq+uDgf2F7h//cwoWhY+hXS3B9qvZyAn1FaeJxkdQdR3SmqkO++8YDU
TtFlnCwy17mfRQKpdnSupKNpxRC/6Z8x04lA9VfjRRF4xhWVuav+HCnY5UWvrAf/
IwnkKjfnmZidwJOqFYVuvGKT3fj0Q0sYv31yVa9RTdBcqNUF/fGEjwTvo40Q5UlH
EXQLjPcK/kFQmNiaEGyl4yOdbmZF5EFLnPvzibJVdN+MaFxFRO7YYjbawV182Y6v
cZDzBlQcXJg8hsH5uyU9soouZWlelHU9f49pj9C0dz7Ixc66AOwRZnVkQn9ghADJ
LczWdzcghKl0sMNJa504aos7nqQu8MJb+68PtAx22PuT8mtzyXM7z7Y3RsJZf6V9
DTT9+XSv1T7lnUKRXOBPGh+n/1i524KeBKns4VKzX+O0RyR2Y7Y8b3s2ccKpRzWH
GdKdZrbtUUVZ+5gaDwTUW44I7LsuQJlnYWFL8eToERH9UZ9PzY1+Z3yfnRzzpDxD
WBQ64aE4c4FFYqwczIRg6Y8/WxfJwi0x1SYWPl/lOximiTfpV8j7tFRlcGMwUw8X
kTFyn6qpxI4WP9cYO9HEvdDC/tsTeIbv25hjLnopcfq8QMuqZn3RFnQK+X+nLVFy
UwExNWhE9z/38Gf5c74N/6yaTtm2oMaIP56CQl0ZU5ZMMGWS8BBv34XjD9GnLeCQ
McpI7rwoPU8JQH27BYv+t2utHi49eAC0s/xRuwSzwTzBD7dikgo/1MguM2hdz4CA
TkE2Yneh1WqurIWRcsc1s1+6yO4QouomXtNriU+C6+lvwX3xDD5A/hiBiePib3QH
AztS9IKxnnFQOuVxbDACnhh5NxiTA0Y1l8QrrIeqS0tKWUGNXe70jhE3dNxkEq1t
C+UqQOY28VSBucgE1f84Siq72vzdB5mMNSHz7r+oOWmUcd10ANFuYAYO6CbYLHAk
rtMRxXpto/GzA/bW+7Y7/nCCg9EnwcR70ZqAszkdUe+mRz+9hKfHTYoJ2Lr269qm
Vm3rlxEK6WLM3K9wsd5wj3LQWOWGmywZk6C0W8xL5etE5pcW0zbYfo+UDBINlM0V
bgBM5+LLagqc8GTeppIe+wDkyfOgiz/xsCdK4v66DOkmNt0KsU48g4aX61HFNmB6
jxoj4kdNj7XMnCaey7rtWBNUetRNKYoH5VDieFSy7SjZwoTbsVxgbbHHFNp82z+2
9uwk8nebzaJL5EAul7QSxI5ZLwztw8tryHKsPsatoYYceASWZQocdzViaz0WzHcQ
79a5hk0F6aCL7PItaXmq33b7AMKXLWoFX4IULcaaGWxNhZNee86AMoAgI8ZD6X4w
UuMuLchP/IPpdUMAOOfjrFWF+yEf/kununuCfe4HXKzgEiAk/p9o+L9Qh0jmjD5P
Fjzu7pQs3zp/uU31bfQq4LgvVzmq7MCIBMmNjbL6s4hbE9qC0oH7VshZr57JhrST
51MZkwM96Z/N78MtYPCofIeDtZ35jcJj81+3GP6uYKQObsmpjO37wX3IFGLSWpuS
ZvLRjNHd0eGTHk+w606SpdoldCMTaOR8eBDSxOZRPa3Z7ZXATxf7RUnrxKNXp6HY
r9mImjKeev09dNoK6DALpDS45TTJozEhWYoc108Fc5u7hrw/v8nHDW6TgK9BEA5v
9qchYJ2qEMRsWHfeC3cwa1qzlFyWoyqu3Tnv9rrKWhFBwLw/cxHyRMWHI+pBJeDk
ZNpSx/waMJ5JPPO/dGuHzbO2I5X1472lemJnhhs9UUb2ACmy1SANK7nwUmLYqT+d
0SetQE6mrVVCUDlb5wigQf6LCngTBYYRhLo88/Ry9hLnsadEbp6g9u1yWzD8Ct3F
mfO8Vy8gjUBRCcZAiW+U/2kCaquRAIZB7CPRPIEarDxT84GzXSK826HKciEcHz3Y
KEGgYtbZgl1zkbG/DhfoRwdrah6Rju0TmMlOZ7J4v3V9i0KkxsdcWK+cBiezDGZe
xpcuB1ULSZ08T55x96TgPb2d869kv/1EjbIbfEAezGI4wb9yJC6oDs1Q4e4+djyM
Im+squ+8dlSs/UHt73cJ0+m0hfjtq9OC9wel7mc79JHfhe/vyX7Is0NZglzXpyYi
tmrVm+wOqqgIpNDnzEfoGaCzA7d/ARaDpC/UJLWo2RPBW9dU6aPYH2FF66v9mm0o
2sYfuKeKbij49SZC6npgz5u3idf4c0xMHjFO486LJ4/MEOLBEFconuPe7EdNPrKJ
Rv+Gf69aMv/xo/j7B0qlZkrw6w0Jvf7qVyIaxcR/KLEqfo21R7d3cILN7zXfs0Fb
eUelsuCHEZbPmDNvJ9ktASea1ve33hzzeoeqHrqauPDEh7/NYaWjcxlwoa4G5Dvj
g4SA/JDTTJoDpNeGhaz6fRn3aIezddAoxe1qUtAsWLsTijb2b+FUW+8fgONbPSm5
oDCwAXAwjx9+3Kiv8TFgESsEdr6h59/jy8rAL8ca2Go79qccHNAfzfiR+vZZeGF5
KwL/C3GWUY2Jvu3W1MEBdCb/MKu3EKm0NLYXZW/jHxb9yrtYI9e4Ah2v61DEhKe+
Dn5UPEGbgeZOgSNCv9c1fu80LEoJuBLaqkgOml3kqYwWcpzFWn3DK7piNfa2bcRI
Ui31e/ul5RtkwPYjNOzuwm5/Xtri6+DJsOwv+0H7d07CCF4FXeZFfBKz594WzRmv
7dMUYhGUxviBuiibVen8VVRfPHlg/lwZoHuh7H9NDAAjRtcNjYBK45qmA5AGCDvN
WjphGhZphTdpfVQ5aQIdyfDhhYqFjexIlc6EOvmLcRgAIDXT/cCL8gRnkcO/1i4w
XoYjnX7x9tD58bbloqozFoFQmzW3a/tjTYeXKiAg4/teYRlESzpSewJ1D5yt2WMi
Qo6UVFvMTNUS/hUa9W+Fl4O2OetIndbbuKeuBSHltfghfDWAJVVLO/qJnPy8s/0s
ise+b7v/ZMaz1GfBnmK0Iz0bM3Xoil1miRJCVZGPt2rCmul5/WWUii7CLgg/qrYd
U7xPYkBUJURSY6uTkURYQ8E7ONd175rAp45SdrxIF56Mm078dpsiG+hf3TkPjSEW
TZx4Tj+z49f43i7sWFKEZu7xH/rkQfKZ15LKAV0YhS5tHpeWc5nGIezV9T2zRprx
x6z9xmx/npq9zpj3R/ssRBsEsgR6h3wo0P2MbfoI+rpfT5qxvsCH9wTniCPrvrUX
Lv0z9NblNhjD9lmIEe9lmiRarvR89aoqStbHhdFj0zk5lWf6qT1fGlco2MsCiUf/
n6YiaMSry1mRDq8n7IBafd4VuC8EYwdInL2oqRgLvQJhF91E9QjTyzzXvprwbfUu
f9SGoulVRpsfgJQdpXe0w++sj5uNPJAY9uF14lBesyEmxIC/HVBgVCwrtPLctL9j
aQcLba+J8XzNiZnBCSq6DSq1/0be5LT30svdCmjKr/7ZyL2hOWhUYOzk9He2YBPK
YB2lL7HQIWgvNPPPZY0hZba1G8we0JqiFxyII49IF3AAVyF2DbP+DvvDazfN/QGv
wyx90EBtnoGKLKL5IhV29jS2hx0nzM7KFyYDZjmfXw8NyAQqPjMaAyhoan/hzRFK
1Dbbn1a5OZdkz/xgLS1BKOmqIfxvQjEuI8EgHDaiiO67+ln+Jcv3TybmT7DcrMUV
SV1egr94MRdDYuEk8KKXd3mmDS0SSGy3yBCN5ht9yZxTlbWZB6JhuANwuNJFMTW4
PtlJpLxpT7B1gzJy2ZoC3uJdcOugOcmwo/qIi68XtoKBPZNc0yefmTbQKJcaXlYJ
oyhKFtwM4idxcp90QTZzwR0m/6fvaeXLxEXWeUdcrSwa9XIxvdOVePsUIpD5bTEk
pufQQCcUdF/FegmhwhTXVpmvono8OGIl2Jb+TdhBXrIwwi827HewJs8wS7aqQAPU
NSKsicKfd5xZbbmfwKkY3Fg5UsIp7m37bnn5BHB0ChJQNT8U7UQutJaSa7t1RlWj
nPrYCpnk3S538wLbR1eFtHah47kW6fkSzGmv2/qVAi33foPVDh89jMqDUzSvcHl/
LeRXu20pO/k3Rycuse4SUVnw//k1+679gCDy2XLqOS6CetMa1WTen+JODCFLTjxO
vkyXAi26QmiG9PK/6mE+YxZmRSiIqMSWPgsxCiTkNH8kdKhmZ9Aai36/AGRZ8glk
ep+u0PEamHD5S8Ln5s6gWYWOHDWyAQG4IynlgpiT1MbbObZwv+d7G8nJxwWOTtVX
a8V6RfAgJKoRmwJss4L/6Y3fTF0bE5QvSqvjMwEzYo4ZolqxOdSaWAKZHcGqx+/Z
+TO+v9FbkUFtFIm6nGVezTbDoNnosYomkNS4AsXaPgWLf4YJXdZ9t6ooeoeV+mms
AQgYQIB9fqkOnk0z0n30fYtGlWRrFpbS6LcfwfQp95loMKvmyraWlQOdiwSTQV0V
hssERKrn0ApyYLAygCcdxJrgkQERvLp6eX8eKsPfJ8dJ9VBjNFCpEJWtOdzm8YZm
4AQDJjvAfvJlu/HW0dZ1IROLv7n+Mds1SimrSP8xd3XlOFeFiSYn8eE3DU1rNztd
zPNE1tBtCW06DDgZ2dDifU+c+hkfMtU8pj5mJZ3j4TVuawoEaTtApJ2fjcH+A/Tg
w88d7wcI7M/Dtfgp4hlAO0wmxfWKGdAaoCWOK0J3PTsgjwWYkZsaPvCGehxBphvt
RW0xGnf2KVMaEAKrY9yjBHp0vGqULLlU601PH0HAlyxh0uneHKDGBNx++/rqhpaI
bnYBRcxNjamV0k4CCyyXAdWiv1pfIePvjyaHDyBTHQw1/+BA8qd5UHdSeNFQLG4Y
mtmmBmyLNjVxgGrvX66lWF4a1UgT2spDKZYtPi+S1Odgcjzh5EuxUGzdQy8t+zxC
gdsGUCPNpizI+zba1ffc7tXBUlQygVzfDlLNgDp1Re0GbCnPBsnZegY0VevL2/Zb
BVxPVhTUy698SxZxbGVOCGIl7sVNyoOXpwGNURjFDt0ulfB2LPa4xgsPbXSfvh1z
AzVjGV96ibi9HgHMsxExOEaKft6DIEG5NEzX1UJxb6Sy71eU6hyZXIRoFMu0BNEd
GHLxD9Gb94h4WxtvPZnM5Xpu0o4i05/evlY4LmA/i+Oq6kVSi994jNVtNXp989+2
T2KYsmKjsokrr1Zfk+OCMuydUjO9UuuGAsvuIJCGuzae9BG9Mf+ddYdaKfwH+nKw
+jOd428zV/yUZ804d5Pt0bYALpnvWSKuatlEGzmMhnmKyQNlMeSjP8RLbdzd9BwN
XRlz0cBc99R5UJQYZiSOtSb/Fs4UKiz7/TnjEd7hRqqn5ymJ08U4CXRKtHYsCFyP
v0HgV+MEHYFHqGD2zhyUgqZFpi4OmEpojAgK0eFf2bjNl3Zllrhv9v4ibYbe5teb
B4WUkeGA2b5OKDM5/ohcsMYJn5rGGSEg7VyTeAhQmGTkc8/fLXUaZMtY26Yu0fpv
f3ecZ5NA5QvrZLdfnFitw6oVGzJayijSkrkBF2OXHMQ+mBOxQsFUXhn25TF6UdUL
1SSM0tVoyXp2fq8z0Uu4nxdU/gWFxaRaS76i+B8lwNesxC5KRJ409rv5YU1n/RHi
cr0/Wf+LqgiNbGTK0zPI2p2+mO38FOeVOJL4JK3hy74S0cgFajX/N8z5BTROXoeq
26m1M8Z5nm2pNr+VzwzcMpp/jGaNVFeSgwzdEV74MtwF2QdooPk4L93mr5sN0UIp
yPrXsr4AZU2gxqW06cNUeL0ALzJ+Zhn+9vwzK9GIp6dXtzGBkyA5pyCom3zvIa5t
KmzRXqvvMosbVxGrmVkxax01Z3oRAF5hiL18gom5sTBKkmEKgyB7la8FcWTqOkiO
qnbsLWSg8ofyG1GuoSzim9UREFYEg843xYZHXBufVY2/CPxPQbPMyF8GN6zS7wBp
FelegNegUYubRGHj3E9ftKJ7Kwq396ARGyz+i3slW/bCvIShAeCUDpKS0fs377Ps
ZVSzl2r+RJL4/K0Xt8shya3MR1sMCNUdOFAjjjIC1F8h9hwX6IP6knk9QE06Av63
ox5+A05tkpVG2+FXKgTfGEfxpwR+WI2yO4SPb3pWJ8Mymy0qRnQPJYcVMGoBmmJn
s4cLFDeZAgccJtDp7hJfCZMOXChKnca3IaFuhTFCWuB1UZkNzJqCKob89y26Iudz
5NRtHoYknIS1V4cXwzl+vp7Fnv2VY/pUyQCh9yEsrI5MWKiMphdYtP+1UpdWJ1qM
RpHbjKdlh9ATh+N+iosebumjY472FB1PTW3h8+yrcwOILcOXMnJWEMMISYpnSIOo
fTJm1BUQH1F4jPaPsvvKk+URLlINVYCTr48LWyBdnPVWUK8E5MpNw63o90vhRr7b
8rHwk9g3t2nnZ5Az6b8e38r+rzdPwEtEkU3phnh1nzPff8/vR9Uxx1aU/vw2tA0P
SpVRA1M4u6I7//zOK2KYaHTwVVZ6hu9t4FHWch1NfwsksoT2MABSFhZbb8gzhqhV
u46hqx4spl/OMhPEuqU4ErVek4/i52iQhJlz/U3RyMFFf+CbYzPX3YahXGNFi53D
javNuv1ZEmdp9HcRZUK+XRdiZMCTiANO+8larWOM9dJuyifrx+hoX5EVCGPxalXy
83sT6crjGAR7Am/RMTjVbUPLcdqmBBD/6MnqHItPecU+eFWxYQ41u6m+dnbLCpL7
mOSK9KvaqK0urFU9ud0Pmv78+GB1mkTw7dE4s5sezOvwM1hsNrPW1OrmMZvAcAqw
kBRqvay/okbXaRN10jtJEhSXNA9YgXfgQUYncte9cWsnD1QjBkpjcO1kHVBqmcT9
iGadcwpZyPllzhnpTfOWltmt48D2fGEE11BHT9S3rEWDBnBsBDC/8I9bU1KMQhHH
Rmo7kCqOrDAxCSn3RUSJmv4kLgtbYSC5EYmCjlBu5XhH5RtG2Fcm7wprHLGJOdkl
reGKFCu1tLGOFAa6enjvBG21MHOhI5U5lerJsACIonUAsdrCQKrzb8iOnmMvs8+r
csYnicAoFDmrYxIt/uqCUbIPYeraqctvXtkQIvUGyGhcjh9BQgutRU3w/lNVsJRJ
ZLiV7KDPnGmj1enXvUc9YJ4nySaX1yWedZ31ucXv3IGoH5dTZ0fc0i1Q6vfTF7XX
dX3VtkDjmHxHrUzOuI/bBYuHMAO8DtLDITXVkwS9qR8gixTKd8qTIsyh98BAHFUj
uLNf2AzM8a6rzLAg5ZxGRq7DVLWlxuo05XVUxtoReQhiMURUjUSzUB/hqbEe9YEz
Qee7GT5ywQ/CmkgI7HSgCJdPhcFifQtSV+LpW/x1EvDrp3NJvHt3kL6wXDR7+DgS
pCwoR/kfD18uVCjnJyytiOaPPtes4I1RVuwNV/01rcUHLGMOaTaKUhnZwplCyBDz
O1acPoA4YGtG5rOhjAxr86k3sxj1T6q52HvD16F7NEe0D8Ma2owIWEOwlN2BhBX6
bXv5MOYwFvEOcUVSEmOjEsjkaZ6tW7fRNd+HqxftfMGD+hNg1LrU9vO7RTuTeus2
UxoAL3N5n7+LYyqNjgfbPNvl0v3XENAnLKPo/C2b0t8r+8itK+GHWUp/yUusKPHt
trK1ZksbhQ6eIlPUTA0Auq10ZaW2iPsMhxP9NGxpKoHpoDFLVSJGJ7BCPIooOdLa
1ttjbj7hqYV5bLtx+1lm2P/gtpmXNarzBncnGRLBRxaCKMsScoZ8JN0D2sHHLWe9
eQenJuFy8bfAHgHGeL0PKtQPkTPzGJb6r5VatLPhhQ5usO411IJZ6VgvP/SulDEp
Itd9bU5ouHLnrELyqFHT2fH4Wf+ejH9U6HN/kYkg4WPl/U4JGW7FP5zaOzh/K63c
WMygBas+n7YOvG0CTZdENThKgGQtzHdHongNXenGrcAUWSByLsrQvOK6rh3lqOHh
+pCOB510bXE9WEGcQnG+uvm78PulS++d5PtSklRGLh6gVWS57JKlkbnthoChwE74
s88KFVMLXh3E7dWr6MSzytftSWdumSErZ9QeO9Rz5OeSpcP3z4QafutSdB9uMs5i
l6wNEUCmB1b2w8jz+ZzDSkjlkEFORsi3Lz5YJmTo4gI92e7YAf/a5eg380ZpgmbE
/ApSKTyujIYHDGk1CyjND2tA0ksgF3WYWowpriAueEo5INSWM2dhFViC//HeXmVU
qv5PzYGe479cFEunvLOuEUwrulsv0hcMgYKDDLM8kq7xMhqe6tdZnk/S+h9v1vpB
pziKoA1tt1LsijNPcC0XvEHDHAyn0RZaO9JaPT274wt63NsGgpFy2lny9NqVCdO0
if8pM6kDo7cWRA767UDgGS86aSdnzg6ZnU/N2qHVs9hod1VxCtPZRVIuaUkaqrGW
d6AqBFmfSvsWXG6PYr0ILqvQcfJRDrnU+F1BDvoSa8ACeBXU8E6i57pSChveNE78
9KqIV6fCWkkbM5UiSGguEuiIDNPgRy0IRpcHJDuv/t6Ouy2TZ8oFqpe40EPxABP5
lL2hQfYv/oV0yXZ6Rm4pGegbUHHTXMt9qhhBlICbA7MDqVKuTCJX51rQAp12/v2S
OCw/dtJLLgq6purfHB4j201rI1o1tMxhbZc/wjfDoC8rWI8WIMRSIVxeqBJThO0q
eA2Z7hrjCxTGrRMZSBb9G4CZSX8JFgduwln6bZLL4FT5kq/bU3Gr5n1LGVEs03Im
Dou9Qr1e76P9mhWg/e9FuS1SQaZKnwIf9fV/ek9frAKjWL/r0rcJ11Vuub9qumOg
R2dz1Em5CqPM9zb7E/4DT93rHJvjcBV+QscfQMr3LJ0cyBtY0igzFlLjcDmpd/qb
USxana929QJNjw0loW58V+Feoi7WiKGtR82wu3TNYzCPRmgjHY2FzRQjeEp+ciAc
RMk5L0lTmV5JeNgor4tw3kdGHRiWG7ij3t+C+DwDA3Uq/WJHnj6CLEj+i1c0hqrC
1joCroVyMdiCiaChl0qmQGMDUUVD4bZK7ptR2iNwf+IaLJfN/OSel1SL/uFPfQqt
5nzx01k9/8/7kIO6Fh6mPzJXeBnv6KER6zGbunc9iRAWXhOyrpqBqyeg/y/PjjAe
ygL6wlL3IDGKaYxqo6mS/NgUrH5fKqsQMxmvJ85HS/47aNaMI01pi5MwrGLos3k3
ZieJg1aGECXHqikfNAdLLTSAR3bZ9K4WXZQ0hZmnFW49dvZbWGOUBA0O7lcgZXkL
1bionuFW5LZHf/hha+bdQgSljdTRz4ON2Q4MaGGKBl1mf6LD43Zt7lf/IohrjfXP
nsY2PPa3CwDN9Vegd2QA3tl8OdsTxtVB+502s5GjAOanvNnkDBEVaJ9lMA2OrxjZ
zfSeoGU6z+TBksbrzoMHGy0D4KroJi3v304AAwQuGbL+C2UGrJ8VV9LwyavJChmu
miiazmL17adEpZilNFXeqs1KUrp4X0jOJVaVHDSOhO5Ql96uwk4RaCA6eNkVlPDJ
O/3O6KoCwtq69gB4vwXgwgWsNfgVoTMCOP4Wn47CMJKouC4xnqOPbnlZqa9wwSZr
QoSBD885ZCUA+gQh1GBqZBnuSF4clni2PmTiiLs/WGmKbAo1CzVvRj+xJSo1m0t0
e8wkYD+eqk+56vz8s7fw9LvrpxIkJK8ThUGSZ6o4TOdEgXTavzt8QMDMqSIJ4prn
LhCzd7aCG+FaODJvQq1hkk5LLvF8MeeXO6DaYvo+jaQd3ElI8sn8Dtc4MjuNAWsV
qndmOXexFaDkXMAuNfwpv5bwL/lOlvCbzy/qIAezSp4A6jWnKefD0jjPc3FqVNVb
VgV9ttlYz26I6kd7CE2v9RQKkKHK0E4TwuvVODzmfwc63SUi9h5UY9IbRc3/Q3ZC
yWFSHHH2hL+fVkT4BiHPNDnf2i9dyUnordF/iCOjZdwZFVSNrgsrpm9QLRaeHxRx
CII7phVxdSm3Oublk6KBI0JlgRb4C9m5jrgBpqDEFRKhZ4G2CgGG2S2HAyoOdWON
tR3OWMLVapyzoj/DKsT42bbXQ4fRRpuqC9JzvKCohoBGyyqdHRypdzXILyYLR8ub
ICmz4sGwFR/8uJv62C6xKdg69gDe0NegIcvf7aebmwcpwxPnACiyQ50pvbjnWMt/
jSTkdpfMDYZiHAvwrTi5LicEPMjwrqBsg9QMZqO9FVs24qItBdfVPvsVgOHMw8Dc
Dmus7gQ2rpnRiX+XjgnpUM5jCNhNP7LVTNuclKvWSPOLxo4Lg2OHjzb8INo82sr4
bsydxR7XoYtbgtBQuXwRkZWynIkV3i/kBaLXN8erg6/+AtPbXzp5mZlwZ+D5cKYg
r7mf5vT2bfOMj+XmHrMJ+xETz+mpEdZb3DOcsrPTzwjaw0/aF1ahPKDwYXrm96Fh
vid02FEtt6bH+8d4WREeTT3FR0cJGEXlSV90YgWzUsWtkWg5e1G+Q+ezzZwRTKW8
xnNhkhP8YD7ikZLU/VpE9F4JkBa8iT5aHPgytzmH20650kmQhVLv16yfxLDypOCv
UuTBEgK7MqLFmIoDj5A6lkvD2pZrBHHsKZHrB8qge+igtDJJYOIdOqfe2kmFNzM5
dkNGTqpJVAE2NT3ZR9cWxWF3N6Iw2IHsBoRNN1adZebL0XOEz20X2ro9uAGXNprO
2ZFHn7rSZ29ApxeH6WTs6YysouEuh553eQdF7xAvddqTJS5SFTARakquBXVYdYwh
2SnFpSHxPfIFQ7CHpjNBNJIdgUKpHEgcRUAhIwGL38J0ZpyBEXPMbQFSXFINBPx3
uTns/+It7x8T8YvQDnfukJWwGBQk7A2I1Tet7StFIZ5U9a3vKAcf7hNZ46LlcOt0
K5ek+GxSpSMqEZNnCGTbstXw16tVTPaF0ZvvY7KhUiM/6FZJTnJ6nGtgfpy8Z6fR
9z8sFvv6hM1HBte5rQJyid8OS5ZSfskqaTT8GbvD3NWJDF2ZnF/6AQOvl/IYxrU3
VfklIQkKA9qWJVA4tA6R13jnZnEWJd5TcesoM1boKl9F6Ag0ee9l+vUKdWWNLbcV
AtTtnsqSH4XM5SJl+DTL+7zzUzu4WV3ps1SOC8XbUme1WmC++KxOPw6K+SG8W6Uk
07RNkQFexHOBhvADj3QsNoNNyZC1s34g6u0xSSM0iJjX6n7uENLtF+tDfpJ05xAY
iFE4SVDM8oWaHcenK9Hm6IbaNLI2QDW49dOfw38RZBjFkeaoRHSw2aWJI/2mrCw0
Qs6J39igQDhFWNVnEX5YM1/n1FXm7Zs6eLgv6ZVR0A3rI8CDSwSR8KFBfcjN0Kvt
BL7SJ7r/wf4elauZx0+cGxaLQzJW4Yq6t9jaLS7ljxhdq1gB8ELM1tXx7sfHuohe
v/+ESf4udL+110qXDVlcPaMFJCIJmFQryvMy3K2eO+p9tXuWg29QVCwEmjTBYW4Z
dwTIUm0a51xALI+Bj73soIpTEEmqZvStU+ZJ9ETC2YV9kpE3QGr9vmw6fMhw7fBB
k51D2AMMgk05ZzA/FZyogjKvxgCh000Qdw1/QbfvWFu7qndN/xbMtMk/g6ACwG61
LrmKodl7+Z8+7rhY5BL2YxvIbhc6lqpUodu4hpRuPVxWqjACZOPc8KKNKbdUzPqt
+CjYhralV8BMWDBqEMePF0jq8KnkLsAhZcO+X+XsaXvShpIvB5Yl0aiv7XY6J3y2
OieVLkvJKotm2SN2llpwTp7oxC62D3tqJMMxGhIUnuc0A9ROsoig2WGsng4ZIsRI
igo/bt3e5gTCSrHp9wFiWKtllir3DKI2oZ7K7zp2nk5h+S04anlzFtYonWgsI2Jc
OkUzC2wCKeZtg3HYvJ08K8ocJFzeUi9odMUVA/Qipf/39akHQkc5tZfSTsaEcsqE
VCQrmLwYsQXCTwo2ucMb5bjzlcXf+HQj03WDrKZkhfZ2tMbM33gSaDPI6O2h2qK2
kQXfog28FTZKdarBT97plytlAUiBb9q0K48+k3se1R/D6ExjaZS7JaRDSiYzHOBH
8pO5iEeYBdUgA5onYLNAWOPez+y3vPLFxsaymyGtEgOlMdvL0w5kD8swAErELznY
XuzXFInCLAlA2xvGtIWl3djQ3ol66ZfshvJy5jeNsk/X/4U4hXd93al8+rH5O7yE
WWThZD+L9y30DLzwPxkxOBgsJnQLqg0m3DWAvK88gKGJYpYT0QHlD2INNqcEx8du
HXTRcbAfqzyhNjDr5617C8xin+K5YbZg2GME4gG6CC5/Bt5T6CVxP2NwOpwyXsyl
NpDd2awdoLwadcWleLrV1G/Nqq4XZP3KiEIRvTFGg2PN+pjO19tW+M/9tm8zIi4u
CUsr1Cs6rnLRWxWMbLsvdfftjEjxR8+JvcptiwACzdVOzNfzUUpwNpiET0NPlqIQ
pEyBhPRgzGXiOyZWZUHATkwFDSntNI0xXx/UbVQtXIdBYFHQDf8gbEGs4D9ZK57C
v8oNZftfO07+FVER6Ifl5scUNJkVd1fZnKD6U6OkfKHcpFV77iq0YvxmQpBpaV32
7lIjZUnlQgn/38wvA62wxQsoY4D36M/Er1MBEt7Nnmun3MVCGMB78KVLXj6rHl3v
WikM62KwgSIj1tgEtimYc9VwEKrmrNyyGfTHpoC3uVz+EV+PRN3cqcS1+xBkfQmf
yHA6LAd6m4Ngszh5+h9ZdejfnsBqlE4c5sY06JUnbDmQ207jz3ycnii3WUacHxp0
jtwqeOcA477EnPIeEa5I6qWn/PitJucilNX8AAapbY6dux7lq1TjJ0BkjLzqzzeJ
7VXAzwFm3KqZqvxbbhY7ZU2Fo/DVRPJ3aqW6HQ8m7HfkkW9Mff0Tv5/JowCK/EEc
RukPoTnM60pOBBKDKa+SkvhEoQftfy7jAK0mOyPhNwuC9/8+0xHaUzlimdfBWDTI
mdZSiLfIi2CD26SDx9y62sJ+h1kjBhZxBetwuD9kBJpUzmqgpSBo3MB0ggPqv4Xi
vm0a5NtRA9E9G5oqZzMcJlCIGss8zyZ9y/KVAzY2QboymQ2rDtMLoHXceU1m3i8V
KB/LiobMSKZ30VqxUj34t/qHKzcj2Rs31zdcA7EY06OLsRr9y51Y/XC5kJrmc+2f
vH1kdOcj724Mv98VOq5qanqk6Zoe32O3cLDOFLOHw5rPsnS5tMa17vedgNurTPMY
I7oI6Ah2HxrVQ4ZDS8/HwgE5+hjwBb7euO/Jl4FGtO+BWdqPP3gRItdfS1zEf5TN
qs5GV4W37OIK2Y2J1iunx1kPlGUnEUJzSdjFAn+znImq1lb8jHDKVF9HI9bEudlO
OQklLCmwld3OEmz2cc+U3Haxag0E7UsSv7ROwUzzdNGle0POkeotkObwWWQazpIl
g7+5dtgpHEmVdWySKQcw7kLU7cPqKbBhF1iluZl3RMnWC6ZmxJSYyPhpcBUrbscJ
Z3UMPgg+Ac1wgUZltUiHT8BjKWlzYoXf6Nvyq5WxDScerHvL/NtcoALvgJ9zQm0k
KXPtRfe9zJmxCc6GsGPAW+S6a/ymSzNNN2cC4Y05+Fmh9V9/e10bx6sdTLxliCzC
kzYuRd83wXQGiKXpFe8QP49jN9ZfuuIqjjmkb8eV79ePeW6bdsfAWZNApqZTl+pA
33UKuqGT7+5X/wKqJDyPZ/8aknsU60UgJigGEEotetMs335rnmvsru54Xe//dK7O
4ZxVa8jetI/pMq0bCEi2cnoQN5phP7xiyBkaXK80j03ZltlVC6zBcT/VDQ5KqXxO
YeBAyY7SwVTZdLzZDzLAq6FjesV26JROGb+7ctdvJrlLbV+lX62dspJtywCeIl4g
/uF9R4Up3el+iuVf5xm0jNPF6OJCamY/nFUlpmrJRza3Lv6WiWULmKrReZx8NZ9I
gxioT1AuIKdAbK0ac2ppByvI1kbx7Oay3k68cymXBUkKPF2T8Om+npTnxBI54eI5
V6EGPD8b6Ke6uAmkpziPrZWdx+QJUC6M2nNXn4+7UGz8gAYoXorOB9fS6MhTMCcF
oQDXz8mbEj+JS4F/zOOkZ8ttSranTv/YCMXQuEFtpd7VU/C//gglFFtjdAVNqqcU
M5i6f2/pimyH4z00CFNKtkk1scNWB2iC3XrvhV3xRaSr4+zrFe6tBIkhqUgVFDHP
n234Vg6PeOursmy1m+I3kwCgy3OfZE5m+9OHFH+TR21jUnTUnrcYTnJ8MCeQFKZi
CUy8m9qMgEaSXIql1QbPaEE9RoQhCLwCYqGvJIZ1pK75ni9CtsnMZSfYwM1L2X6E
UHSWRznVbE8T0RScmMg+5mop/2fQPP74j31I3oX8b+bxdX2AFmDrecr+GJJ01QQu
sncwGkas6w53ZE8rVL9SBpFH5UUyEkKnwCVaTNmvdSchHQrYAAGMs7ILMJ7aCRl9
BAlbvgqQX220mTbZloNbjM0UJqHEPt1d0AKFN21FnVYrDZiJBOPeN22rgnadhOEb
FeREX7xU55+HSGhi2ilvjnsXMUu6cg3vF3W8NokAtAiISWGNJMWyDfUWNcypqDkN
mad44xSYegltvN5kgUgWmvs2BEW6n7U7RUV9Jjr7ivH21bFAdYA9kJSsb9O9eX6H
oeSsH6DsCZYKbdthJzguh8UCHZOM+czLCTqr4ffUxGIRzbYGyiz4so+HjiPjiq9P
yG+sNK5ZJCZkWn4bmxYOaqaOvq3t4Kr8Ay9XteWuVHwE4QPY84gCBjA7ifqAVr9Y
LPXnpNwvj9JkOuTrZuZe+v7elrPG4yB6TxyEt1RH9iYMaWpkjIy7V1/k4B4XB/J2
dKl1WfPKOCe/phZexCWgf6LrtZaZS65fFHha7l0dkUXVF73d3Fx5WgrPJH+svpeX
WUSYn6uGiM1rNix8AhnaF9TyPdYw/yKh3L5jTPYVW6tczNbJUR5Wr2mKWVk8uv+0
gkMYswneXU1Euzgl04vUxQ+v4xfIvu//MD6Q2t0cxUuxRhJEHEFs7tnKAktD3+6D
xRXU1Sa4EZv8ioLeEsLdPt26sIihuZ97h4+jriM7Ny81jYVKuwdWbrwQyQtKoYQA
L/rnDDaoyKmd6j/iDZmMTYpNmF8DoD2a2bEzlpsP2DhFK34HX8k9K79WKl/nkxNJ
gtR54XrbIOPzabafcw7JeqTYVXQJiUG2hEzqkqq6PJQk1QLhKrjWyC9ewqg07QvH
N/iGr6lR0sts5GCi4S1mztJj14owjqkhuI64Ku3ACXpvxa/2DBZNxtDiy4+cQ8w9
0gDBgqKAih8oy98Vb5DCf/PcPlLYh1Z90eb81cAB1bvyv5DseumjGzsRS4n0MF+Z
K9nWZ5wvdsWG+vCNeBsrbwlEgmAK0vyNd7bX7bS9q5KTBQug+xTKnPVU9eLVQ8xh
ppstGD0rQyXocn+6roNO4E3coSn41K+4Q/NVynfU3Uy0xtAm/6l1FwatBBU/9bmC
G+NHxGZJ3RipvuF0v3ATIjNYvJtbBna/RfFH4KscxTYQg6ScdCFQBTpImsirRVXy
X5tVryTQrQjgKPQQtMM1l7XdJDujJmIenqBwy8jrxsniJHggYvYwBL5oVil2FFzD
JErMOmjsu69RXph7SGZ18rkd7Axud3UPnWsE0EhLeuApRuCSBuT/s9RqMrJP5fqd
3DG4H7nk6TzcKn3kc1cDo1fSOzpBMo/aaGhSVMUs5fH4GFjmR/9ptdZpmAiUYTYm
vuxKPVAJ1gvJanXZnpTKeGfv0VFkzA150h2ciNXwcSCxWmHZYa5cADTP3OFnfwtp
f507edj1cTxUcg0gWO/As9GM3mbHzFroUhR5UWM807k+9nYX1TaLmIDOO4yt9qdw
BSqSLqi63zKGRSsbkS1t6j085WqEGNfIDSbSJEbhrvCnILAx+FlQV/8ICc+gdqOJ
EIvxF0WsmykcqXoFYKp3RIlGx7SaBer4gmNBG4GdsN//BMxBK2r9DGk+qGzjEAq4
mTOsXINy4AnQz4AkD/d6jLmwhaASRFvZjvjcHDjkkuzv2lnlXoWteMlsZeJDYfZB
f21dhLv6Qz2dszEaXniYWfvo4QnQriIdB/asrF5VKPW52tz5xG8fe7CyyRx91V5X
Xg4hzD9doddOU3PRJ8nZCSqDcy54HPmwgEqOfj69/NqVccEMYIaH18XSoS0hEJl4
u5VMhMh6wDv9fznK4g2i2LkwhJTHRwoiSEX6H3r1/6uFqK+Sph8kisrP3vHJN0Mi
rgZvC1lqlaUO/QX/DTuCPAI5mkWN0eFdJn9MphkgjujPdh9sZBVZMYFhrUmvmmWL
lWNkNVriePre5DnDLfj0sSt6doh+fcHt7wMnisD7WBCL6vhO52vSZzbhBLrbBo2d
DR/Gux4tnHMlilZPAacdEpgBHBvHlVtCTEMRctoGix2AZ2290QQnmRHDyjYd4CRr
sKOw1FIM3dXnS9uXTT4ay24M50j85H1kfHfUqHVlzClb9jhsFBzE5lBy1K8msEAn
oVTvQQVucwt5+x4PkLim9o80TAGE1Jw066OzKwdEc3s48ZaNN95EwI0jJuK+2tEp
26yS72JTsMSZOUx9AsSESCa80aO5Jt7GXEmRDY7UA9AwFPppzZOP8mzNbfqyfN4o
DVx/a4v4nRgfsfC+rXglSHEjNIQD01NWsZ3faX08OtehlN+KAVCp8rOpZORSLs3h
jJjHAS55FR7DoOd3mJ4D6eVBIZDI9J3JOBSgTfQyqlvYgpXwecMPunupW5oJTbKt
kjTFLEIxpIJQuAf/Gw1AN1LgtFgMk4hauA3CMjF7Gp+PD80BIK5qZ7ylLSX6A9L3
oeAI98/sM5AiA3Dl3k4u8DgpUu8dc4Vx4oX/4IFDGJoGJSBNjDUKPBksuoDSfIwO
QTuFmHT7Ye+OBTwxrDEc3dtcbRjSWRp8dwrtODiNjyi7KH2PZ2lhixx1xq7h89GO
z7OiHEk+Kp1Nhy01VIs0UDy+461ZPT/doGn1OA14iLt3BGVDzJgWBix4sWfaatyZ
ZAItuRDdcqCqpyxzK1gFYz4hhuZyqpbq+YJ5ENw0cynygQdGUQaha7z3uk10ZX1F
XU7Y+q4r1CbG2mkuKKVYVsByryfmmbZi2DJIcdv+b/GbfOS9+Ik1z0oJ5a6ngfjh
BTYaDU19WflwXkTqQBALqsluM8ayg6151CzqKYJWM1qxzTmvd9W1lq12rY4FAlPN
UBihjOA8PZzYmmAu0CNFWx0TS7fyO8EtGwuH7SdNPP3UhpJIiCRKeIt9My+1UrJK
A6E+rf7xqIll7cKwzIucX/e+aml0UUuUG79I/GokAdMd9WfH/bS6GR1knBzIcGWZ
34dB4PILtJjfJBlb/Z2pbSLLYQoTosOTimYWWTcmrd2gLgxenPoMQkiG0hhrs9Fm
yiApOUu17c7VrR8vpy6ciuItV8z03GPQqls1+hvBsHSClqXGKkLmJnTBjehF1NU2
N59VbXVgt11FP031MykLqlb6MaLu3EJ9E0VKjEHOt1ST41OyGaQTlpy8Q7YUAp8A
G6bxWGw8j9MPZjiAuBbmkvfpwo8YPlU7Pjqs7kz2TwNtwYahUfpfgC11YNs84HNE
bdeI4sXcao413lsPW93M5lj/25inCCQI68vozG3BtH8TCrl7ArcAN7TnUAECA/mA
X1E6yUFR1RXqVeZGUwygqU3tAgg2lGN2nCR4NNvj7kjuKZD7vH058NOGiMoowzmj
+AEOBVFOBbraI+5CCc3El0Jv17RDd8zW/g4yH3+jPFOqH0PMBrp6/SjXSBBPg4pD
RPZ3fZpCk/hHjmNflxiWgbYr8sZo8WYx/YUjcMxqd1lao64SdVbNCISGzNNntYDM
SYljxuo0xR60G+5qrhUHbogh2AlrpkjrSVAweCLtsB0aIn+g8SPXZDT3xMLoW8e8
L2WKo6Oqf1KUyfyZvNLeDJhIIf9WGDawKQ8aGf0xDegXKfUH8MTdU70FgnB9LrLl
0qbHQ9AOY1YrcDQGCZYRhYELLMa28pB1bhVmSsYg9t8xFY/rN9Ldrk8iImJaHFzd
P4bk59EAavwkPu0QzU8r5nV7n7ADK0Q668RjPWeGb7CdNDu/y62p4JyR77O0/BL8
wlcPE4ZAPpicps63evftokF7J4bOHdq8wsHd/mRWvjG6n7vlBcXO5zN6LHBs5l+L
tsJfBTJ86o1REQSVShMxM9YibN55z4R4M/rGR84qSCP4UunMqJJvloGdwdSQBcSV
ne3I6GNehgcZIj1g9jtlzFlrb3IHvPlmGYgeAcW4telK2Ufc74mGcOdqJpwhBE6l
KnvlJHWGR2qmGwrh5YmLqrmDCDfpGMx6iVJfu4mXzLWfph0P9YZCregv/xGSjSU0
vMi9H5i1iOqMgbxNeYmRajHWEX75wNVBHIzpnAaoGBDu4K5Lma33OWyAzyHnOhS6
iRFn7cLj/Q29YwfiClrzGL5dAPlhXCyag49/y4AVORjatPuv16S17/8F13x0Rpl4
hc+h5CFbRlnIOGSb3YGcOgqA+uaaFwckqQQ7Br1NAij+2B1MV+/NQym/b+FEkWAK
uJJeynNEV/AEyxsGYpozWZX9R011pnGhnQ0N8n2q593JkAlHPFujAYRrF+sXxfBd
bXI/jsC4YS52bMgR1sU8t2rvKzcVBs/nqGHYm+bOLzPShvBppoZyV+xO737/lpfD
FPxJBeeXpsvUhq5jAAdeARiiE1/CkJi4Hbvdm7ZqJhTX8Fhrcm9T3FHm0kRiSLXk
bfZmwRncz9ykGoZHoTh5pyrRkC/xIVvezJUuMVoNABSMwbB0Yz69tYhl70g96fbm
jl0lpHEuzASq+dasqkMMQeSYhIvABmOKXTh6fpytAdWcsDi4IIl8O7bndlW4Bij7
5mvD9cQ+Yh5HSpAguQ7xQSacaBX7rLZ4NIhNHTkv7UaP8bzcpR16HrSHa8xM7bR4
KdtYQW7HoCMYxnF9TWoD7Ok4EvEiTnSa9JQXAJravv2vTCE6Rv8gEt6TatlwbyBZ
FFJSNUhFQkBmbf8zER6/DlYl3MhcnLJ0Q8pXowAnqiJAIPStHVZDnRM3eRZj345V
NftK3adkZwgiBCd2Y179pb0v7nWeQbfb7JTKw0RbN0qOYVYVb+yFQJi9CDj48H1N
TnIKv/TJamWesXBR0Am80BI84HSZS95GKlmCFCyiR0Rk4PPSOy7DApA/byabuq+L
YsMMYcMYn6X60wumKzIQkJKhIdMQkp70h0X6Tro6MT1PJQY9VK7l+dOBFC9VlNFQ
QQ1i4xtXBQm9W1i86+dtbYKsSsvpuwu8E4Y/a5GOdPc95VXuGb7iYdm1ldbpJCst
kgttGDvaJ0mQyz4VUCrQK8azrukrRu2spVmcfjJAkbmkNth+dxx+XHztTb+vgGje
WR61kNLuLf9fad9/15p8JSRP2Kyjp1YFb4zykRJp8HMWKqqa884NztH+I71kFHBO
0T7al6O0vhIW/MX0nfIA6BIoHwu2F8IBtXplyBqfa3xeyw7wYbh+XBeYEzqk+BmF
ZytK7fEarygpECTL4wH1zvo4y0ZZalC0CJZfaSt9Lq/Gj1EO0CYPSiCZgncNqGF1
xvCpiD4ohyJZcMz3pVr/rsxEV0U06Dyd0F5hzD3uTfUw/tZRhnerVfgX/WEc2ZuY
/aVZZIdvq22wI+BXlhVBWJPI/mQTmbY/v5pn55WPTbveX24vvkKHzOW8/nooFQh7
q4/Lt738rIyTsmT9YBmQ4/Ml+lzSuXZXfHZ/HtFupF0+/PesUXc6SbVQ2LVLB+GC
tTc0BWciIg4/l/T6b7TCRtZfmLdiYlssXea3651dY877+xyiEEH0h4o+zPdc3oh6
qi3o6kCfbIls9UGpamgnHppVZauHcyAwWnPaydyqxHT6rvMIk+Feb/jp95Zru8HA
Zq7VZ4ktDTXy5ZKjcGmUdK2AjH0jP/We/7NRtrI9t1lNCVV9Uv1K9Xu1AZARVGRC
gv2uyFe+GivPZXb1wSTVXdytSTUnU2wzdnFf67K0I7PtI/DaSJjJSO8dloSCxD34
aHTULxFuod+ggzC/Fb3sAif9K9Vx9jeRUwcjH3NC9veerDqJLZPUUnHaIqAVwMG1
zjpHBHrNZYZF63Dj7517Bn+8jbvUR5w7uMd+XpLbdBnRB3NSI+NLNVR9n79Qw8ty
jWd3AHORksQUgt19V0m8GJO4ys6I455Z+PJMtU0P7JLFxShPrBfiblxwH6XsTuWt
OP9AnwBJaDRpXoR+SEw14hj/UBrJT4UxMZgSlu2dG4EghMHv5XJQxqmU6uDSmlI3
zGDLa6/8NfA/wc0PaxW2GGKwPn+X5unXQW0h+c8qkuIL5mFC6lqQ0+UHfQFxaH0y
hzRpF3bnClWiJfxz7SFrpqFrFakW1wuHxPcn8LL6hAIbZpp8NAmFMHAtmItwD04E
AMcH/3J5h8c/asZkDvzTSrKJQttUES0ftvPX8nbjmmwxuirYLoQ1/RdwSb80VNoK
sBBCzuUcYI712YZcoU6uvdZDcaHvydJi6XNdF6g8Dn1SirZ1FXnMS2htttkF980X
F+AT0UtIdT6P4qvJMTalLtWFAtHE0WzofZgnY5SzfE5DsdhjMdtZvPfckVSLB4Um
K5i983Z6naKCIBcGJ0/FaBHdlGGMYCbj0byI6X1JEXi7sf131jvIxJPEpkxvmfSu
jWxMioZRLHVsT9VYMpC+1sLdTf/BsbR4yNR3Vzep4QKjTmSFuRNsQyUm1f+BW48E
EIY3AX+fXkEdB+hmQIU5q1baeNSORr/lf8EzqQ6zuh99bTadQ4ztstnvQvNbB8lW
cRIJ1VcVgEPAKp5facS2/iGOxMvvObcxhYJZ7BfpNU5rMUFNrSKlvCCnzstC5w5m
QznuvuPhy/3q/FNM43OXVjHmH1NTFFSNPF4cX7XM5Hbbf7PWg5KSGAqL+YJiDuYC
zzZSWh5r/k8g1zC56w4holxBwo7klnwb/zrOotZ1BcO5SuV0OtV3a0PDZFX7dJpG
mkBgGjvZjSeGte4enZdTHAlFaaapulaWUA1LkNqrMNghFclVNDuigA9KhCDK17DQ
t8pygswtfgwywuRy2XZvebJwQsKqHPxGyjkCikNdc8pubA/+ScaXivjkLeNg27qK
3TcYvz2Qgx/oudMWRu5HQo4bqpvQOZsgzOfbCRe4kJBVAlnfsekrd6JmIlt6MqFO
8fBPwCRW1qpnksqd637QQJ+O+yd79U0hqhPIwb2jVXRlifQjcxnuJVi3p+LqAIUh
WftBO5gPvNE/VauZZhIm/RfhieZ1KPFjxWVvjhUYZn1Vwmk4Ug1VEjuBOHumsupo
bPvX82tRwEEjle6LEeVKMfhdcY4BWNDaf4ijJepmGtJHKErlHU/rb1HyYOexfKUd
9qKaAXj8F2na0pE6u3zPAGQlyxWpMGFBgbwKfIGGa5q5UHwDpBDCh8o3rKPEfOZd
Q8f9T3wzXAz4+5wS1+ZlQJ5VR+LTmmpnxMxt7ZAfZks/jwJ5oWP4hgFzQ1ykXe9W
8OPlDNLb9bu8skINzDntpcJfN81f51zTV1E/lbdhXHTJ8C6F1RsQwh0Mq3ss62pc
oWFL4t4E3Z2rYt16sTmTHDexhlR/h8bcZmEuEaFLHMClJF3rvGmJtz15Qfol07Ow
ICSnPvTcjMqZdmuYjHrvjTP+gCGOmruPvaZrIepl5eRAkEMHWRMhlf1/HvdSs3Qu
3fyUytJyrrO1nfaEPK+PuQmrjc29Etx4FB1QpNRCyZqgKpott2N3tPcNE1srk+/Z
f26GA7zqJ2X8J+QzFpkGpkBauEO4+Lnpm/MevogJrXE8J50zLLXifiroD1/U4hnI
GI5RdyI0LMob44mJzsiR48WznqGs8yVg8ipnjKql63EQGWJPqtJJxcjQPUO2Y+0A
gxRV2t+N80fgs4b7YbbMBJt/JePzJjAT+2IRWeGZTOZ79jA/TewGVe9dz27Ub9Kc
VqWFtxWlZjrfFRDf7qTwDcdJLlVFakvZH2RpVoRNJcAq8fIFPD+wJfqsKkdyYzO+
vVgE8xmHWDlv/o+JKc79kUBQOo7sdcqdKNXmttiXUdE650dio9Nhdkn6QupWclhO
gcIsRC3OybtBxKRta+qZmoeppkuvD2vLc379bQDzmeurKzH5SQAq0j97AE8+Vwri
LDsEHq20y6twlrz305F36puZEL07UfQiGtd0JQ6nXKcMhKPVyKTv7dvbj+9775hg
PW6Xqp6SjWDIy9aj2A3YNQPKHWAlAVYxRWL5lS6nH6J5Eys7DwVx8DSKliaUCeLq
QZ6RcFaYZsD61EUH7TnCIfVZtBScUGzVwl/i6Bs43B27VZbyePvqZPdCo6P1UYT/
tBz/qiTvQ8/dIsdT1Yvx0kBODbc0QWJZi0CQJyFM74R0/XZHjDsamuLDSnOczszw
INgCCgmUtVKJ9MMCrpZNvnM+bKCG6mEXSckED20fCPRmzj6d7APbJ5MN3+Fcm8vC
+MxF/fLAi6Q1mWFY5o7ePB1g0xVd917K+4B+lEWK5AYRgshHRpyOJIJe5CNdzwiO
uDA+IP4glZd1BZy1E1E7zjED0WyNPXyMbgpwG7KhTSkOTsXp456pQVx0I6JTyxjn
lzMCF1LqlaUMFy48OSQlOR49tqvhRZztCu7DiplXvjp2Pfga9LcFnTDCH0mLwfF1
QxXm4B125LR2hr84A/agBxgKhvlrNWUdH2ThiPvnu9H6VWKScLzlG43eKUi65Okl
8EgFp9sIksUYYrAXlEjwrwbL/9We1nIJGXRmY4Lv7dEHcMwcLeCOpbwHL96TvCMK
CsHhpAoiPaGNpVrARxgri9ILiczh/QKXuZE1gxJYT91/koK3u5etsM69LHdGBwG2
8rRk5rVSQfyFxFU6FzqkpslBubA080Ihdm91WSzc/rNuxYlv94ipc5UOIjCauFZH
SHvzgc9qgc8ni+7XAO12LM9kgxclQh3qNuXs5cYMC3+oNgGgjwrfsYONGr9bPop+
b3+tZ6qA6Nv4Z1jbnuxgAqTfuA+8HdEVM8Lz6J7SY8FV/NAcp+OKvBibEwhHC0dD
kFZq0+Jc1OozFm130Goi9v2oJKSDTr9t7YEbwXiVLs04CMRhaZ28XlnxhR2RX1yM
qwdUxyhOhafp60DPDoSvZ7/YCBS4rsdmhbY7pASKm4/+5jTZCoz5jT9+rhspCqCW
vmBomDlNp/DHtVi+qBL9q0Zme6LzabF9DxfKNrOu/s5wY46BNPn50qaVQVsuQblU
SInPgFGI47pAbZgUxdT8S4XM890POCxTXJDRe7WXJ0rQuJWF/2q31i91B555aEfg
qLm5jdEHmGwM/qajk3HpnhqE/IOhgnYkVDE4bz5apmemIMZGNPRChHPemvda7vJA
Lw1cCzvbi/4LMKP+nQxISeXIAfKKg3cmktzvjj9ayqQDEyVIu07qymm4wt0vs379
GSnrZsVsC7lEVPoAO+NKJX7x8LsFsfrQ8S3yAF1RSxgSf0/Ko1sya7ONLXNNPNnF
7ftiOxKQbNo6/YshN65zk1ECaWBnJrGvoKj/dQmhKix1QkDZ9rwXNdY1ChfAu6iV
rCtZSBtmdwNcHtnUuUtGdprD5Q1N354ZQfc6jS7+f+0rill6LTbhSg9j+iiX0J2V
l6cglqEnHx3u/tWac83nfiPLbZgGHZ06FUBz/7t/ytH3neF5rWm4wuqxWJvJ4RUM
5BbIz/uKrBoygEPzoxpyJRAdzV8iMoA9BxAp1KtfJIyAQnlk1gZkfWL9P1YXPhUa
kDPIrfvYRKMeIfD/SCTHR/KLikvUgTYaQqYJoUKW0ymXoJ+Ej5VtMelJ8X6NkT3M
ddgWrYj8mDdE9Ai/C/OCLl09NcEZBAQY7M+ihOIU3IEXcyyuijIDiziah6hsyVii
N0LKgAh+e1mpP9iYDt7toGJkrLc1LaEYQBKELnKZg+5WO3ITbi7HwO6WBZsCQxxx
9UcPHVnFIekvAtVMNhrKcKwx2CQbc54FEK1ZduLyU+XSrUXA4a88KjbXGphL6Fcz
NchHBZwhmQyEDvDtsxUlUTHhYd3Va44PXkwjIqiwwoG0uk0JBuNHgA+ZVhdXPxrV
6OZ5IzJwb230RAnzfnnq4CP6mhCD8E91yIeyaqUu3RC1sJBAokM2yhMsujJ78KHW
NVJdJsEu/h3S3dqa+9Ns7LyS1eE7lH/eU+x1xfXCtLVkXzVlojwbwFgVAQ0WUoEl
goyUACKk8BZwRCoOXnr6z2hX4AZ13Nyjhv7MpL0owXIhh8Ru4nHpQsK4mJHv5vke
1QTJEima1STL8sKIDZUgfgWlqH8NaBsHC4NMOecK8qRzmk8E3UnJ+BbiygOB77Q9
8lGiwh1x2sqi9lDj7w5lmqFslD/YhbMazH92+b4gY3AxtQ0zJtCtxiBUWrz/5pSl
BpVWMiz9J08LRzBOfB+OO6DO2KmMtrCGQ7WOh1C0l4gTjKjHteCpQD0pFzdmlcEz
FWgcxo8jxltvvUj/nFoUeLFv/beA5LnLZHpNYbY8yfpCuAjf1NyTjXsmPBadAPLn
hnVrEsMlJeGcnmLfCn0llFqcQmzrv7QJU/64FkAk8ij+Yj8kLgv9nirbnOm2syIt
lvWdPNIK/rr8l/0u3BUemBQulq9JofIvVHbYY75ilr9jRdA/BVK1P9Qxuazjha0B
AaBPaADZF55+Ad8oVK9hciD51ywvG/qJlqy/uGZdJvlgXvtxg4TbfwCEmJ82DQtR
UwqYRfXVI3i8uksexHzYqRJSWrTWIeY+lwGblVW7Mv8hN+SFvf/sMHJ/RRDG3o57
rYNLh6xMqLzOLk171T+wwgQ+jPwehh2URbmGkWUj92OPBL1HsrOVkynedCoHJkHa
tiuj+q133B4Q5sIgYnhtXMUEYGQOc3u8tqj5cgpbDFZEFy5rMiS+PXzIlz84Pekm
sOMbwI1eGvfu6B48wZ6cfl5ZKx0TLjp3kFllIPjOI+UzWsjRp2R2sqDfKnWht4q9
IZ2fS2SmS0YNllMkk424E+1JooebrgTK1cLRZGIXMIbbbErnoWTCK2yEssRULfTt
pFQLIjxXeT0vZR54z7uUaNXMLrga5DNAJGzOvxqJUFosH29QdHrjuvobF0692VHI
I05F0Cie7yNkyboJJMo8elUrlLCG6clAHU5ijNEciYvdvkKziVYmSZFP3uIOISKA
SLnJi637uD53iHY19t6k0gB7IEIu7nES9bO/Xg2JIf4kMkiN6p9SDZL3MVxdFhCx
0jlYp8NnRn1duFP4hVhNdraXnlLqdCcIxHMJtJUH/avK48cq5YBTQzhFSeqdrwYG
3F5r98cQRneurMt7shdHUpCMWSNWx6fLzCwTKsn+j5oa/iKxvvl2PhZie78lU70s
a2shZTP0P3wCkNBT7iEB+s9KgmxNeTqgCZWqzVthoHxY5sSIhMGuHHIlvxSLqHgG
IOr22wIRkr6d1Ko6PgiALEoX31Sr5xrAPLD/uqzfpN6b4NIQU4Gho59mFr2tmxFR
yAcsjT8LsTLXmrFUsaUxIFa71UOn3JyoBmvEWRtZfyiV3k7Tf1NIs0AVZe+x4vYl
rCJBfCwsbebwfbshXbGWdFwMfxEnX5AJl+4xkEBd/VKuxfL7MxGXIaye6W14InBx
Jy05TCUFw1J9IdKNxyFMsMAxSJFcxUaFNW2il42C4hgXHrM5KRP+Bhcjzqv0JCVo
qm6L1BpDiGwlKFOxLvUtvyni2hvByhTWHhEqlcluEfX6z7jbc6W+GJ6aLF6TFbiP
o3/oMv7PXqOt8E2BcK9LCUQyxOfzxWJb1ACOAsMNhWDU8R5nYzpSAjxliYEZf1yl
5Ls33lhINqVaBdBxghOhAxIuoPENt0Juoo6HRBpjUcwXpIfLk3sd6xxKTKtYBax3
a/SdDvw3yyaHKqiS72TwVS/RU7x8dY5xoyXLEe3cxCYIj1ddjYO+15G1Ibilda1W
pK7GWg5MEWUwF821O1ZfyT2rrEsja6BuyYGbRs3QkwhKLhMJ03OJmnOHkf5rpAq/
JhVuZP1wawKtQ3HS92w597sxkl1EQbTAbF83grnTCZmi5ENXj2B/HvxdPbBjFtO0
UaoN2WsVh3VmNW/H8Bz2IWwp670+7K+5m8gDYBHPPHjS+88ysfwkSC+xSq6F88mZ
Gl1LpCekm6YERbYJl3QYg/U33rVSylVORpu2RMeh1ao0+c+WtyOL+5q7/L5A0ujo
xtW3h5bgEnh/oUa4w65kRW6yfp7JodtUHEVCSN7RKBTGQXM05C4um3h9yneI1irS
vKv1ID2J1VVRB2KcohIueC68IHoOiUl0B519Yg+GqvR0n3beuVV4AoRkjNF0yNx0
UXcz4m4aQgK8d65yNkqymeE5v6/kU484+KufhyP5XuTzCOtO+AVgLWRYRhOXFF4Y
Wt/S3+lrOAirwql8bFbteRkU+6mvxPYOpha9yXGp6y32NQfn0hhsnA4Q+AynH1Xa
7SGDsXro+wDoI0davoKcHprNLJm7DF6f5QDAwRdxZr3lAIlCYCr0fyP7y6LMbTVf
cCmhW9yfXoLuvVS9fYNbuhPko3MYKlpb4St3jpOK1J0tW12Vy9veocsIKgJgCe6D
WVr0/tm7jsitjj09DmZjZv5u2NjvbpxzR7f/orRcco/lyWB/J1mOMt24yaYQZBuy
7umxXSnx8NmzbNK78HQcMhIsDFq8kz/9HNcXK8KT4tSiZOMnnQ7gfpFvZGfxI5Tr
OHTc6aecrxuXVELyHLwRf+jookEgVp68xqin+fQcXYgH0HKGkkzkJ+niaK0Tx3P1
mMuUMdukvidQaYKoheNsjVzzVnJ8KebIgKdorD8jN7Dot364ma+ygObRQQAMPJbG
xXF9N66poSrwG4e5kIapzI5kRNe5T3u3yKqvwWSLqqipvon26wj90p+JZHfYlFL5
sVcIxBravKYlqUxoBaVVQavGigAm4w1sBuVarCB7zyw/Qg3xNVoaOF+HdttcRSgt
ZHO/46/K5vAUKYK7umRg46ngxiGFau0iSaQ9NrUuHyWgRQfGyw/EVD5AWy//XAmJ
JPSYHZZSYNzK0pttFyAOY2bpQbiUy++exmRajt1ACFR3qFi5bgfzsqP+UxpIVQ+k
4RLTyCG5MNDxltoOh0qaRHc5SbbFXRgmCM0TgVZRJ4K58gGa6kuPgdEENu4XKox/
Q3K2DNXVchN3uCT4wjbabaIR6WzDP20Ch8XmI4iKa/JqCGFbUH5PvJhnGIY0cwTN
abNcJwz3stAUKa2i6RiiKInaWEDI5Bpd/lh6eJPjZX/AiAgmCWfrobiOl4zADBTC
nnuHV6pENn/ck+NHWGVXu772vHV2Lry8ZEE6+6xdAgTwEUShNP6XeIeEc4/kq194
MfdosACPPCLxLDwbIyF6Rqe6ZRTR5v///5JC3mdG2XJNXHxCEwIBzfOhtvdGojHI
X+cE086HUoZ+SXSygKpiKlpASbnGykYFwzzaCJO7irmdhoj99URVZphxh47c3RIV
4R7uoFC+zllT7tz5okoRbp1I7SK4Sw0DjBU6e24/7WDtj1L0aCgGTEzxgqy8wuZl
EftG6Gfn9rAjrMRmArHy0QGrdY5yWL7Ox2sd5kMH1GwSfwUJTZ6vZy2b826RxrNc
FJE5xXzHBR1ldCDjuJQJalOmWlSqNbLU3LG2ZKv9XfP3fxxb8egrAP98bNgZS94S
kKUoZcR2CN4bRoLzSh5a8dsnA4rL8msx8rqUloNLgrgxKrsQtUlF32KsUBwsLanH
kpnSTM+a0K7IYReZ4nBELQa3nZkIg3M37E7y5R3r6SQUhW4IrobNMleHvnatozPz
FkzQLA6EO5YvJXy1iee7VlKOU31S2nymkt8+BHcv28f58ePB4dmqnAUupS5uw9k+
LCJmfhstUrCUPvHQZWeyNV7Kilrj5ZrawVkssNkupCYNKiOrjy/sUGjfNYLMl1yx
4gsbHVw7VMq0vQPj7jbcKHsPknFtJnQjKXPXf/zpVaasE1zVnrsbMWLDkk0ipOHv
M/6woa53qchwjI4LMj9KCwaatnSXzeVv0ETioKZM79mQO6WUNLG7e4r6CG8biJEV
+g1w3M6Vy+zK6HIqQ4amA8d9vBXLMN42MtFuMmvF+897s7caAkDzMpfKdOE/SZ0u
mT2Wy3AcI0YiYLpmJZQNHob89Z1WF9RuJ6S080XWhzfcAbwbmlROXWJkv1lLl9P0
kMNhxsJbj/NO58pK1RpkGWsvFfzxFA5Y4JwlDWGOqWTtK3N0dVdxVUeG+UF4TGSS
kUV4B7jp3PpbNq01yxsQczmW3dJrKqhYMbksbFScJ2lmYBPkPd3cJpgItGMvqfqJ
gjaAReE22kBg9vD/xGghU4R1KWRLsEt8K8x0jOIInkPyMO+ecboNTSDSm05HzGRH
MaL2fjA6cAlhx04n1UVmV+fn/zTToCXAwisDkCJmc+jvTb1lWDMGLRlvyySIiIYq
4YGyKwT+02Claw6kR5ZYtIbrYE4aLIgC4lWtI1mHektueyU4EyY20+/xVV0DvsFU
LAdV/rOHKbI4c/A35uCyPd9hIMlSbJej55XVKPhAkiOquBZ6cfpCBvVJnxNgR5/B
5HNTSjvTdVKsiCyW2LwbbBTMRzM8gGIv9ztlP9IWV6dN0YN1McDzTcGUF9G8bwHP
GWAkzCes7AHn688pG640XeAlmDtmP2dTZJ39EidTFpSyxoH6xT2lgOKrso4SOZ2E
zZAYtVT9CocGZnVjZv1/eltUNqObZueizO8ueNEwoXc/r05DhDlzp9idUVxI2+3z
9vQ5KzWDo/No8zkUbZzAGRITNbJJMhSMV+7o5VOzhL7yxW71/lOvFgidlx5LK1te
iwgPidWx7lsEq5r8vgOZfRlYvQggRCwusPBmQpdxbgF0q1/5aEPko9TCv2azwQYI
x6MzSiAqxHDnBKpQN3H3NtcBYSmrQ4yEcdfpC9qnevvNj/guilqGtTd2cYYJOuuY
qojez4BjFV5T/JG9U9XpljhG5x2TZHk9NwqT3nBV8crjgKbS//FHVrpvz7gi0UAY
LOsIvEkFPa8iUzR6yfwV4Fy9YYEPa19xNGcZP1WPIIrahMuLNgRpgYmJP3PPmD4l
0EKJoWdZkMLkBC92SM9UUEOc+Kz8pb5zn/0r4FQJkC3SncCg1bbeyy4V2YX+zWKj
c+er+ua0vYSkji9Ue7LNpprbvpoI9Dr3WAtx/PW72mlDoGWhlatFeVnIm0h/kdoD
86t7XLJPRchmui9Y2eTIp+dYx/2941vQnMXjQ4IvFPGth/liInJOZVdEKENAZEHU
Dh3qmbavhvI12heVYLupBaXr/j4Ix+5SVDdbA8pC6nJFVnE37nB9xOKMwf2rz0Y5
N15mK6AGUh5x6hlA4GVSO5/Gm6SOYDE3/V5aWcTjWMCm+13KLzBVlb2T4NomJN+1
B0zF4myA1vc9b+F39oGBlQ3lj2x9tmkH8ffSPXHecVqrHsgWdlXbi7m6n+oq1IRv
+rIy54abnrFpyHEAln/YhntwUU0RvWaqHV6csvbQW8z4MwfDkpwylG3KZdzuSUhh
TCYA+nMPpMSSN3w4xoTa2f16Dn6d/udeLVX59I/un0Ol/xKbugg8UVSSP0lku8ce
klzLK+Q9lDi1u/NZH6ZO07A2J7E53zSUSaFYMLtfBvTPsr4kswTqBnYvb3GFbmbo
5SaommfiQ1ht5ILvd0dec/eDRCvEF6jiZQ29boQs6d+mZ3m3/NcPOrXT+zVZEUM3
Ar1S0er1Y4iQ63ua3rYNLe3g87dOAzLzI57p3zMqfz+UXVkMXERKc+UlLisCpkOi
tpHu69mdCTzcLknoOpOSP0c5G2EKF4y8z3GrnVn/GV7wcevpcNslvgC09ODFGGn7
euI68N48cvU5onsDzQA0UwxHRWY3yZyngQVlK2tORqYLackX5eHd+zrzxhJM9ZRF
x35p0VtWIKOgwUYYa48uT9vbMDOVHUXQ/V1iXqxPfhVkv3ZrBHLK/qE90f4bZ8Xs
rh9A/36PNw24dlj1hZrGWxChxStK/nvGcJYzqXwOgdPx44wS0oN0+2Jc6HSrYPy5
WpRkLFlOC0pHrK1IRxiR1P0t+TmcZlPN41ZNzfvhn7wtx3LjaWG81GBf251RVdVV
xAzmB8CMw6gzMJLUXB+yQYAa1DZ74Q+3URXC4qiPcWMNB9u11cGxdY4kUyXEYGyY
ATsUzUEwihdfKzj4SrF8yi2AKeVAmPO20/6w/+la5r89RQfvclXn6nhfK6KT8jkH
bR0RXCXPiozFuSQKC2Wl8oy+d6Wl/vbsUXVg0xjjxPfSFr+JCKEOBm3UVa21KCPY
xaykgwFmIioo9daDYtKYdo/IGoxnCsJLaY/7h561oNKmRVO0KOW2DXaEojudW3T9
Xgx6KcQ7PBKkTwVYH8m+QHUHs3p4nM7RHtfRXA4GC9KdlFdPoha73xnUsI1sELVS
i4ka/zb8oMcTYj4L5fhvZX1u1u+eDmFEelZhfovlpv1ZPtBsEgEnI41UiQyAX692
T6lARlZqhe/RHm3TLOBNRAqn7R2fxNBUhPls6kWYNcE9n3vuRJ6HSLDrsZdSvu7K
nB5eZVUJ6lE7YDnnXyV+DJtpfJxwT735Hs5JnXdD36UtwdqcGtlXeMbwpuDIs9d6
BT440+eRZO2ZIFmDzxKve18B0JyyX3qGuhcZUbVulVHCuGwWnISYCXCU6YI0ptqG
ujxAYsZoxm2FI+5u7AFJVD/zFdTUQdRw3z/vbbHCWdnk/5NG9PYP6qCZiZktGInY
RXVnnOFw8QdgZ/ef0ymVoHVDVjrHrGpDQ1LZJFWJMnGywvUQ/mp2J6G95ibWoPke
MFRtVnpwHxq1jTqZ19/O3/JGZQ3LGm1kJMHLzdZcYJb94iXZU12o19VfRKqjKlsP
4i7eYEof+3SEYLNsKim2VTRkLNdzLyq6Ud9o/jpoyaKpoqt+NgJWuJ8Mx5UiKEQ1
Z7kowesWxg2W/MrEVodGwe3+W83EjJT5bIT5MewLOd5cNg6bZ5+aaE2dwPOOEfzh
aTxXZBtqaojgs9+cDOI9UGvUY2J6zTtBHA7r2EdM3BKlP4wadbvFIdNUw1L1hzl5
AWAxAiuu7HoGCzEEHfR8K3EF+hy09toZiiLGEDbMBI57zg6isKrPLoTyKYdGYsL8
bEvAiJPOmjqwXHnU06tV3RiGe3CamEjCuGB7zOFMY86EddR1PwhFjU4y2qLnMHcP
EoIPhjp/7tCVqgLTE06wFUjY/q2JaKVlvnnmzetLyrqttM25vych3c6DGLcWi9E2
E4f4NAc8zZ9us+e03frbALvgLM3mLJWENBny7X2gEIOIX6cDAlnOmbY+bvW++m0M
GPy9gi65vJ0hZ606q935gX4gJG+pGUUYZK4EKana+pGUIVXJnxnK1Dw96Cb7IsiK
T4iM5tbfwDV8Xk+tyAftk4dcP1Sai2eUo/IdnBLxDMwIQVtnt38HWemFSL8UhKTt
qhwqTVQ4LvaaVBoxSdamZxF3BJ9OupSV3XzI2mxoYVtLJby9xNBSm7MB3sWdIkKD
k+WiaYgYVuKwXJ7x1KOgrDBVnG18jzwvtnZGv0l19S/NLXbqui6+mn+JEiKZrI0D
IiJyInNyYHpCQW4GLuhdldYQmQzKBZ5x8Ksqw9yChMxnX55MSYcdOnZ9Ql388kVG
Ij8dUrpARX8seMfn0GL8s3jmBSwgg1HYbhBGM+x+DEPwbkk8qdGwwn07QyZXNkjn
eZJaiHl60Ek3Z4ueNhNcIIBl6i6Tc06NYWgd2SNnpcb0Thtlw1bky1EBbABJyxL+
/RyqAM6Df0AL92YTydlxiUUFXqo3Dfb1m/oUd7GlJuzaWCcL4i14wpb0uef5+bvz
hXf/p88icwkOxoiemAH0dLCouzQ4l0g8YC2FmDWT8WO2r0NRKltqySlaDuHstOGP
Cao7bVjKL7vZtnnpb8yTtUKCyUraSRQxqr0ETTwOZk8IMZloDqyrJ8crjc+V109A
3d8WPgYP7idNn1zpGqN7T2BpKu03mC7O/D/5lfK2EiYvbCzh3kZxHPExvLTnOB7S
r2MX4JtU3qRCnkVjXTDxOqnHpbCUUvCdcR9rr0SzZyLc4lbwv3MMzCu/Y0JXZR8M
H4r+bK0HMZkrolYmiGEDXwOgk7E8rtBT1b87wn/gP5ylsi2/6DZwY6QRrybUmJxh
MrGwdE0IEh6yac+kdE8aP9PjMu0FDnkjML7f6u/Kvlmb1tg6ujDK+ikE5o78WZBe
Wz43k7s527vUlL5xRFtHzQuDfJxiW612ycWvKK+uHIrD8U2kA2OYzcRh0hSb/dmz
IL2xj3E4ptQM/RGTg5dy0KDtWgK35iT8VjHVxbU7GW+/8tBOkCgJKRCk4PcR3lgM
b+0/mdt3e3PHBh2zE5LMbIM5DaIJ7gs+bC/Keano8YAC4sM36BptBVhNONwInyvP
38GeN2iA5IdZb22qH4Uqyj5tNiXMphbsujKWYLPB9mI3AX62eaWCZ7zB55NhpQ4R
gbvphjD/6VoW0KBD6yhwIjXkiWI3vOgp0BT2rxtXunFXETW0RivJ82a6GtAhYDTN
Tnj00JUVbu8U0rkyGKqd1cwtT18frWm/I6DykapCCUixkWmTYms7JDTk+MFpzZfj
Z5dKn9cp5pbDWz0xr+/hqKdM5ZaAn4ou0AIiIQ819+3TfG87buhTjiGcdaGdK6AP
V3b1nGxg3yromW5yEoLmh5GVzEd38gsTse3xLC8cdtsTY5VL/WxB4K9JkBHzpqyM
fuzFZIRkltdsPM+e8FuoelTL+NBrLyZ8qBokNsE+Pzi/zV1t4xwCNBTSTZ9Pfr2s
80CqsUMlubV6uHqptKh8ir6wfwleJgeU7kGmPWBKK17U8R03maIqQorrp1ck9oxL
NHSdbAG6QEzGByO+PbvHnuJe7yUw91CAFgJ1kgo9dmjsh+Y7CHkEIJUIkorJQX2x
B2fhlkE1sdLfg5INXAeW3jXgWoOHoPCPkGPJ2rN55pDs1pnzzGgS0SLw+qTlHkix
I2t12x9MHLixuAt6JZ7v1QDnL8a0VygCSbti4U9KjMSL9aCIR9L/eQOOk//EjUAZ
FyT6cf+c8DLUtz+2K7CMICvDNq1lU3SLm7xMTB1oDrykCGcsmy3veoY+wqZjbPIU
dbNaLkzxogn9I5b4cWqOFkJCnwM5NuZ2va7lpc00gKp64jDqdmW8RH21VlPgPNLq
IxEBR0z/VFKBfT2vpvIl5esHh7rsfvJkxSnHJEYOiJC3GyoukbUP1noCd8Bw/0O+
IK3f1V6P+ke1t8qkcMVogKA6sM8+vNWFD87cY7FQrJSzcjyWvESKraO/pdi8siAp
3JQCXAzTxAXBhnsNuf5S/Oqh+Y3QOLtugt5ZyjyDpFjrbYgKBtglzYYyC2sYuCCL
5OMqqHM93AjCP/F0cVwdtWxPGLAFBdcCncJCrpq3cgu+52ftN8/tWSRU54Xf51Jy
PYpgIc+0Wqgb/oEaHI6oZymjzg0QrzU/hAVaJGZyIqZ1xAuUobf/E5Cuk7cjxBO3
Lu6qJ3sfvN6SjUhHCwlws7UlY8WeIQ4Ty+haPaGYfDfg33mefKWvguHaTcwL04bi
7nRp0mRrozenUKTh422O60sxZyTyOFwCh1LBSFlSjf5unaSC02sIRd8e260LN0xW
hqf/cLAdy0oiWLynJdYpvKoupP+TktvIlY6dBXL2PTSm006H/yeZWAgbi2sVSs96
z8RrmFwKOBFQwfOjh1Wzt3FeFDsBTBetP2k0Mp9tDVO4mpTd1iDneIMY2O5XaD0W
v0QR+DG7hEQuwzJK9QUtyCCNPZTgyPgLYZMKzd1H3LZ5u1LJpx7LP5ngnIFW8YLj
6n0okwyZmxJLYKkM1NZ5K01A+YNXVnnFsvPIsb+eV7XpaEFUCtEEHrgT4Ml+RXsv
i2Tbhoi5h39gbqTpYQzik6d2bwTxBaMCXWkwdicRieCSmKUD+Xn0EnVYVza+xOCI
UELAg5JhT+bqPH2LY1lbI512N5Yu7Y29uoJ2goY6tZuf+rngsJTlnYvx0d8GJS6v
1pwiHB7gPH0GsuK+9jGf3ALjIwvUBnY82oAEcj9IZZTP7qaehowhOou7sVyBmSqY
rmEhTXlRYuBD/EGeJLXHMSzGYqLePQ80yb8t2hI6oP7FS/mdmFukKF1PMrCtTr2C
oW2bHfJ/Lr5wEeKBh/RWbHogHdgoS1a8d4kgYQwKPksaZEcKV5Z8JxhwrRLiCH5j
BuhqeXdznvzQ8eA1prkQeKRcU4xzkryy70HVi44UG741Bk7z4q75e2BhEsd08brP
joWOlWfXiC1/NT/iiYL7E6j60kfBuZsbGIyFYheIQbUkJww/ZH7CLkpNm4bFspk9
ACIcG3dPklNanl2ziZJrlxX5Qik3cpQk8VmDMMi0adI1kQoI//P969Pa/7qWknTg
CvqEYkekYWPn9FUhhtkzcGMDFxR+QrRJMGJDaPv6FVfYAK7WKvaVwlfFhGwRS10Z
/D65cLCssbXqovWzrcRejGYQhEbctP9Gc6w1WXQT3xXaLphY0WM9UrHmT3HYiFqY
vSBbOrr9e2NSQzqNFQ95xAN/3FfEFVvWvQMcm2C3rYeNULOAf8TZrhDrhqUA4fLX
JT0+FVovLlkFCag2JFYpoPh3IehZZ1Q2RfLZFTf6NTWmpfnRqFghbAy33TelxCAB
fHfJPhZE/RFyG9fWb+rxQ/5tzMCOnL9tQJaHEnS0J21vy+BGhMtOWUmGfnYyPAgF
TsSfeMLzWOv27e5sY3yzPAWvUNj36A5888LdxyYFHErPtlVZkNXrRtK9D//UnjwB
RGx245oF+EnpFSA1Ce23YgDHjvTVklwP1bRA9kWm15Zd34UM7lq1NbrHZfGqSeLZ
Wtzu0585FYdh+uMQI+I/4RVvXA1NA5dzEP4uLTMvsjMVHIed7z1tHtTu8xht5GNp
XmyDUCAmLIOT3EjQFZLcln4LfTdksHnsYKWAfoBr7x3hR0tLfD8kmYixS4gH703I
cnmiLgFUN36pnbY+36GUV92/WQ+vjaiC95HmdfXrV1fLnwrLm0mc5ZU5RXbz1mJH
9Vis7G1WFuTorNTSTOw6pcX3b3BXZpj06/lWpyZTMYvC77looFkXYxX3KxgrW+TU
BgSdzlAsp/EYIO58z5KpOdTJPwkeb5rM325lFK+67ZmA9OhqSVMBRLQigEmhzypR
hXvYKhgkyay/6mQ0smaU3Pu6zIW5hftHxfc+i0+Ctrb4Y4gLQDdufL+LjMaTDd5v
+L2MgfcDe3TOG3QTxsKMVmkC2uNx373JffI16/iPNqU6ScMeLWheSifVGz0buzDL
fL3xs+MJihdS+cPQhGf40WlDo4SZFWRcQol13iB55PO9pVbxG5Eex5bxFDhGPvLh
ivNQNSVVPJOT0yAVo08pcCPYuHtH4MzAlZ6ld+yKybqsmFM0bf4eRE/0WTuXU30w
dtXpe1tHhrxgr1pvodqrIaUBIL6MyFvPCmC2u6M+J1JAyAsB/Jo0t0+u/Sij7VUh
wqhvWBMhG3lYZR4k2wXuk5rLrruzKpEyVLLfcAG2qpfabyVjDNK6JHRTMKsbPdXG
x0wDjNG7VDImQSRNYgktNZvmxIT/zwqKADngRXY2d3U0SQllPbVzpMd/Wafd0Xdv
MthOeM4UqfB18sATJYfXj8HszziJM4ZQvP5/2CGxaIouTXNrRqZOCwRpn3V9A8Qu
PklRodUrpTGQirmPVNoLk3VvKNjX9Aqx9cwLab/LDdqsXy8McSSqAt3Ypi040zv9
af0XcjxkEWm+krJYVyY29g0e9Wmqk1i7Qfd+9Q6CyVkANaNyE0aidKq7zKJLUrFv
Ht3vkPyPJGwJ12Ot9yKbFxn1b9pwo37T0aeVzYGnaqht2Yk628XN8CTW0IkEBdcF
kTrGQGffyjpiXGh4f2fCSIzCQxoSpJBiK9eEXqVwFW/ts0kOrlp1V2/h6hg2D+yq
lTbV/kPr0ao+WKMy6B2dQ2g/eebkrTfiifzgIq7q4Z1FDtjBqUICNgPV3AdR3cMU
TnVNq6htey2ZIZwMv9VFYZMyVV++YDT1AtazfZK3jonl1S3TJwo7u24m3C+Ah35k
w3LuiiaO6NTyF7pQW9W6u8nnRdkznap92NqLN8wawPn3jNEVMvRBt0rC9rt9wXWU
+z3NggLE1/4j7aki7PS7axonlWTaECmmz9T/+IVzwgVj8qSG4S7FmTKEVTwlPTrX
NzU3zUFz7SpG3VmfGteyExeiE0QoaeolvTjCHlajy5KpZxifFEjFA9MhkK4ItJTn
C53n4ShUfb54uom3j1Ptx6eWdiiWHu6Ga6YdCo2YOwSeHZN9FJ585AG1jk+TEYfV
nN6Cm87sGHUpzHva1/4H4aShix4mIbu2iGu70g/EQqJnNmWI7hH9lsVoLKaOzvzc
O2856pv2pm9wRCfd9y34GhoDgJq4TVjNSil0815h7k+wfMqHQXrBI8UYFqM3u79u
9mePDIN/D0Jr3a/sD2DvsbgzI+ZXDkK25mQ/+f5rDJzO3zAgSqZKEAHNHiqLLD3b
yyPhihlTGtw2hKaH74VuSY92xgN+PZWHddVfRW7TrpJkwj8pUSvS0FoY+fA1lTFl
WD9HBwAKL8bG/rZvWIBgQHi6OniM4MgmI3jfu1jTxCvbLECMf2u6W43Aqf3dHQPE
/ONIL6ZwktXGs49RFxb/Jq+W++7+ZfDDe162oMeu334S3JhnJ7MW0bH0fKl4Hx2L
uGB8FxQE+VyckdY9fxqoSnnwJqbifiaDhPLuAs0BMB5Xwu/uTTutJQbdgo8hknAu
pS3R5gbDgBz8E+DI0EQ76MItzRNY26xT6faxOaWGxhuk/vEgkEZZT0b2X1wfAHte
ozJ7A7iFnsOJvUJCWe84+46qdalCpYtdEcxh7jOZOFhRKVybAE+qqSkHsy96sItb
uU+whSCNAyYHWyFMT0SjqZIIlEYGKAbOMCXamPfMZhDvnwPHZgRNtaM/ij1gCDOK
uJPQIf38QiUXvXaBNhScwfdf0JJN5Ly9mrgPLpIbQaaIK1LotxIxzJQaK1DJqj2E
J8xy43SsYyAq0Jv69aD6axjvdnZOp80Wm+ry2Qk+oMDrIFRlvXrm+uBYBPXyZRYT
Ux3XEfByrtzilPgGbb2W+dG5ktHaeY6lzGxl6XfS1hJHBYeL9djbYbUO3hLtZ/h3
639a8Ef6z7lkApC2YcfqLBasJ3N1znNmNbS4nZ8H5XQTSvs8ej8a56Q1SgslVrT7
ww0gJoxH/qXxY3b3xmt2Q5XUrxaAvsV5qzXerwW5IFqnbhbuMqSCTOp0I/jOzsxs
za4z9A1beiuqga3K0n1QpPQzkeAFTNUhBVfOtnlAaCtHQSu8sB5Xw+oRZgFKBMnS
FwTj/KiMCel3LzmR7jjNqTATs2zAaSb9R3Rac/fWb/BEgXpwfVPMT1Dr6AyTTjnm
KkqghB+Bef3xGHpkM52faB5FnQkLByn7l5Fg6g4Zw2MpoeZc8lR1/RDAZciSiq14
DZSnqNBIu1x+UgLSsFygkDUUpDTVyvWv+Oh7ajTcbHiK4w6rY1rAewzCc5PpnL/4
lZ3/LND5PEgaLOwyFeZT028aw7z3df+lPuHukDqyPLwPYSao0jZYUGwQ17a+QNC+
BJI0dKsvQQxdDODQtQfpBOSNwQKJMBl7tSAG/pX1D+EGplGEkstdhXqTe4HH3YNM
JHJlollp7IzasmNPP/Y4h9I6epXSKjBDv5Lp3LWs8m5Sek3YXMf0RtS4gPR+3lCa
ujh7itP1dGrwAocoOIknKFbgRNHCWC8f42lB+U6DQtaGPKE11nIz5M7KBiHUIlg7
66NO1CeD2U0IhmH8QhqhTxB555hgdpyxZKZrlJ84kIqjKVbSAqsuhbaL7nkASSBu
JAmwP4XfiaUT5kqwSor91fq2n0BwAQ0CD/EAIbDp8HJ/bMvDJjgPNPlVuySxKqru
8FpCXN6og9ZF1DBpZzsGU/qpCzeXHvnEQbIzbif+mtIT7n+DqeESwyiq6HULle55
8PdZvUq1R9Vhae5H9cDq4bXK0IzuL97cSHsn9QnLlLeiPIMEF69hjHaYj4I1YqQV
MUtSNR/Ul5r92lFj3LNz+Om84c0itwRt8+PpRUfD/azeIuReJLZGbeqhilXd8SaI
pyH80xsqaVjg4j/uz1NVRtwr0PL/LG9SZoSUoHbtBTmhvyGm5uXeM1KM0oBQHX5R
Wfpf36606L//QdheRBjEoM6QpaqG7+BKCixSRQyhBok5RG0gMXCQlQSvom3WcMAz
8PLcRemucwi0G6lSmczzdndxSPXPrCe9kU80SCPkzy1XsnkbzqBF7+d9R08kqNWv
CiZgmxpptC1QKRjNa+MhBBNSsPABKO+16wBwT5Gt7GrozXCyXW0u6Qk09n8uZGYC
LR6mmTQ0ZA8GAEfin2u1qICZInLUGelaNNLPi/t5PV4H/Nc77X5XlxoLb0Hyym78
d5pnXQdj1tNkBdN+1AoLy0SSD6LXS3Fy5xQoT8M5XjpFJwCguJlAL2uD7Gzk/mZa
3V7NiQeXSRNBIdzsSzX7rxNTc7U855QrLU/IP7SnFI26DzJnOfOx5R+sninGdZp/
T1yUdXGugngPyWecOgvNpaLV60qGiFQ8rL3KXIEu1YVkSnDVWe6WxEzHtUvCv2qU
5K+5TYmUrXvwEHsunjvOx9VRocRk8XD99cg/YFRNOryVReHqr0fuU9Qhd+uEJB77
VCX5fl/sGPQLIMIkcLyWKil4HfiMzGEu7Mm9avFkwR2Hd783trVffsPUEO+Iv1Rg
CXWY8uTd58/Jvz9jhxvtbX+UcKLsuXSmKyzIgQXZBOIXilY0ks42EW/j8Ey8HYBL
0Bv/i9pkqPdHTZStNz+S58nkvOIFzqzitrhtfPmbxP0aEIv8yVw6wnEe2jnaz50/
wDgPLxYgx4OwzsyEIgMNylNodwZ56czgHqanT0fNJ5PFPmIWUPV6ULQZWaef7afb
ThAHF1syL77tzeOyAvLoPGkSbymkBSnoUcAuK1x6EHgGZ/+sZBwSVtXdANRrYWeS
Rk8+eLybSXuuAaRTLFZcVH29xPeCUVWjL9rrx2gZzjMrxyQ4iqVk7mcpfBPk9MT0
qMwu2P+2RPn1snwwufEaWWLv5jSCb0r0SxWIBPeUVebUJMLnCY2vJHQuh2XjjNxR
TsIru8OUGX97AjOKxWcPZ3qnbUt9gwmHrkZG7aB6+H3i3D3ClENRwx3gYZHTuTnr
AYCI6MGrK+QnDVAxk7mewu+NLcCLyvhBUv0DDaXL5jphCXLvL49dk0H/JFsqhyLs
0xvPY/hCspAxYhSvm2FCNOTGZ+BUrBLsyBjQh021qmVe9i9SHLyo/d2xLixp6rZl
TesfjLQq7/e3xj5fKX3mFwVyKf9kb/lKzlmSsLUJx4RHcmgfOpcjZw1fm4T6gd3x
nBCr8J9n23dyoovbwJXL6z8r8hGsw6AqbV+GCXIHSUQAsFY9tbjPjhSMA5KSbLj8
cfK6mLAd+mnSrcK/FZosnRcvALnwLUzdlacq7SfJHhnMgoy5O4d4FpJRGiw/N4Ce
aixtlB6GbRJibionUBZoMEuubvOHVixBHyNlOp9qj9FIThyz0zO48IS0CjwFVUbb
jImRa+QNGnKtFb59qLwhTKx7B8zzGwnAsXjABZ7qt0YzOVsVqPMFk3xgB5p49CHr
6jSUXf3YExdh5d0iX00VhCRmTNNuzLiNE32ZPriGwTw8Im4jajTlBfScfr06i5W6
ehQRJtMu20le82y1vsDdDX8pDHO1faT5JZyktaxp7gC+f1dRC7PMJfwyifOhpGhw
7uTb+ELevc/rtGtFqusqyZPj75mEr5snRNb4KX90e6ONFnoMUtFR/fkHf8hjEqjX
Ld+CpbjuuoBoKEt1X4Cyk6HEGHYrVviqfwuSD6mAsg5zXm9FAOOJrtP9lDj4MuoL
ZhVsPNwlyF2bOJlgQ7hnkqNj/5CWEyVdC9NuM5B9QebM3wOqIGpdq3VNpJ8shJL9
XSgkrKjSQr4qUvIcVQOYJLkPESNEWLbGj5KmmKQM34ZeS5au3FQfz8xniuuuABVx
XrXvKH3qGMu+ki4iDphwShrDSHURjzPD0HsRuqbkOV8AiFWtWShciCbYkH75jGVZ
Sokm/kKpmm+Vq+zaKs+HWgqLR9N911iW2v40Lpc/+r6V907GBRcXPayWwQhUZopa
nq8fzQSJsTgUehnuY+sdiRNRtz+d4U1GlY7lyLgxZmTIquZDXB4LLzI2rnKn7hJ9
CK80nYIWSyE/3tC9xpSFdgODBRhwAoWHqmD8TK31hQiCP2CZngE7l0R6G/OXdDRw
ZovckbXM/GVi/bAZVGQ+3JH8U48krxYUriZvGoUCYQp/lm4N1URtOBugFJ7kVNjU
YRW5i4plkFZU0BFG7a3y3zatm3eVG3aHyXPjjxp4MT35b5C99OvE9p27z6Lgewvp
QRoJa3x9POZpKSm20jECybMfBrvZhsDXgoJvFlfDNWFiJbK2TMgMXkpC9Evhu0Cl
lgYlwCR23QN1rmb0mcxl1hYrQmRp5FQVL7BiYff6MaONW1z2FIGw4RmdJ75wLFXV
TMKdKuDppWH60yuRRUUm9/scLJRIQJbXlHqt7pB5IpW/4sDn3cbAy5IixNbma97E
fgkLcKkJzGzaL42V1kqsjxG/153aIbXYdJgiVjChylFUKashdybcZReiYfF7eNG1
Z/JZzKAPoJnTBbchxEaI2aV6/2H0JgA6I8aSxJApKcLWlqt4HRMBh9uWjeIGZK4o
1p4uoumy0znZr34FV6+kY2JXm1T0Vx97OibMcMNonpV/Hs8DSgC1v7i0hcx8eern
vVoIJ0pY+I8s8Am7o6vZlKrLpbRuCt2p/C/Gg7nU0N+cEzPQzIlpEUNbYJm625le
iJ5xuE/t16Tn0Qba9E4Bdct2/tyifrWr2VdIRFvxNuYfW3j+nMoo7zdKT2wgDNoR
y5flHUG/BVYy+263BFkPQypSz4SQfoSwcPKo9CMkcoMg43V02l2gmcnj6vMRQ9CP
miolPuDyM8Yf91T8wJ+52QpSGMNld4gyCY73H3lQtjCC3I8k1pBYmzqmagjN/1Ke
xd3pOaMuQe/c3uT/n2gTN13of/if6X31FLeTwxj/Sq8VY+IZb6pyLH4UG0O3fmOv
jitZppMx1IcqwUK8E/5A70JutEip/R9pePB08wy9L67i94QXhkZAaQqndt/MY1T6
uaKsB+7ci8tX+Oo9sW2HG1WoZnaRM0ALbyU3SzvT5oydF00A0eGgVNY/R0f3s6fk
B69F+b6vBiDKMV0kzLanm1r/XejD8tKIOSPNVS/U1mn22XV6PP0qaGmYc8Bhd21g
zgdSf+8ETCfF2WcpXx4gNKu5w22eCMqTd6/wS78YJpWDOzZp82MlSJeBfwVQD0sb
0luzKPCFG6evKkwV08Y5/i5mLmQh+unKPNxJEjR94BGgxvTGqzvATnJpIn/qpDrW
l284tvCkBbhCeI7B+uA+22g6Wo3nrFf9MIQtFw9PJpIfCq/P9sRr/9Z+fRiWFdX9
PnFUbN+/iD5by/yvCxkleT5fZLWJLTlqOrpOj/LGFIGtcHgQtawcxXVusstRhb9M
Q9j5vndWVLJXOKFIbGA1Emm9Pen+K5BWHYM27L6MQIfVRYK7t6dJ7KdQC/h0+c/w
dKWjiqWMru8LEIGbZFcEk7zsznlVbOdfbzKZgIXuhNatq4pR7GkwuoFyZp9jJCB2
0Z8mz6cDdSzLULF8wuh81latzVurGCx4/KgoN5+mn9dxPbg4ThFn/EftEfVVIr6h
+btjb11oaw7E7tndMFdrFfGwk+WimfyINyu6ZxijbAIbJS30f1cttn5i72TqCrdv
FQhqRld9OlQgIlx7juO8cw5iz4BnhH/b/SiQu2lnFRXP2teS+USagv6iyVpkuhIh
VLLJpaa4dsBYvts94BX+lpBFjJoF4vYhioP5jy6OspnETVt61gaY415XfLc0mOAp
Q7EYjTNrx86+kcvUFI+pc3/tsRl69wBb2JCVVEjA1xnHl5GTICi1FL3iCL8ouQF+
D6WWZiJPaD/7m9rtowdT6+njVnaBFlos3j4SArIThq3yTl+9VNowSDxEM/e7uaq+
yDoZBOqMEMCwiSr9Of7tQZ1fW26Yy+3x+1HX04VSqf8bAWrAbFQi9MJvaOYRyTzU
0JdAKpJsJsrVUXloZNmESDhKvYwgJDs59m2o67rcjteuV8ixybLemdGQ62mlKHjh
m4YDTPc8VUXpK8uiLoYnbGtjfbNCrMVft/Zdh76FuYXLizP/srWN8XzkZgeJtd8p
CBFG8wVjVRLDZ2/QtRV04QEf1mXL0ivTTij5PY8bImwsyVdsKhziilbJyProgua3
WfGITJDX+IrZvvQqou2odKnRCc3MbX/9FOR+wUSObyfIKSjd504A6lhvUUDDMMur
i0GJ3zJaV85el9jq0VmdlVHX9Nw4f3Y15Xa7NQlYCFh01XN2Uh5p7HyD8cI3ZofQ
sTKkPFR7XLDeqvHvBDrCiVo2KdrSxDEWylGxkSwR/NSxNFgkdECk17OWs0ktfLhj
pTC4FCd3WsvneHe+MitBg6lI/R8yTlJYpS7DJx01eqiYYmd0Y0FGb4c6rg2IBO4n
fBi60RggK8KoeLT5oRO2aO2x8uom18m81otBKgw9hdLPYQQTCKRXFzSIhhP7Y8vZ
FC+qbShb5FOrmCh0rQnuMkUooF1vKPj5JohQVnsTEi9EYdlgrytWCzFA6USHh/m6
NX+j+dy/bhXa/fM2PrZLiDHvktbIIHKdA1yxjnNfJK9eY/aeoYvar1e9e3pDL9DQ
4nyxlFeZtS6lqlfjyV1MrDkMhJtYK1bOdwEyjMC7HXbi9A2bm7pHx8KU1QvXp0IY
zCdBv72kZSpWxeX4Vpi4ikTnWQNPIf08/uJ24LmpMAQ9pnrrWYuhOfuroyeRtgD0
HF2siVWKXwdTptnk3kdC0XVIUi+O4j3YUQnbSuw9iNmE+TzSdPwpigi3aDRGi5wp
fvEcLRsq84PH7BDTGShfjoYvy9EdsbqhuxH1SXMw2ChfqzhpDbBFslOaL6m0t8hv
wXNXwXGKSmXoHYckwfg4Zaf3wTlmpelvalODZW5nOSptzwr9FUMG8dMWvwARFP+N
J43m3T1lQ8ZnYLBG63sscrFJWqu0BMeNUr7daK0rTfLoMUV3M2S0UH52e8gnaSla
8n7XqMsQ1QAHQXdydGrqVUARmYR8N4LZ+yjF5YIsuqMq0PI6UQBrTGLC8HJkbXL8
anW1UpNGSDt0BV5DXPRuPUgtjZI/ySA8vAdMAGK7OuoolvTCzToj3qMCfIq6JL6R
gSBMqItLRCLjVDj0lyDjksGcBJ0ZfV4BC04j8UmbhDwNXGquyT8nULZbSa+rbNMU
xkzYOlN2mXELEtUv/5zBExmoIT64mcW9lEzonwul00RBvsCKNscqyzY+PSfrYsoi
/JBRqKtW/uoXBxYq+Z4O4F7Xh4Huj9S5E9BDk9M6qzI8XiyEv/7BkroTGaMCKfSR
TbrUk5erqHO7Vktyp1INZziOp0mTo6sS17mEbaAP/N5mRN0h3GhLl7mnbf3hkSVf
p/ucJo9sppMGo3xPEUGmfcZdWjJCOwcpwMsrgceVjXEJsFI5Ss442pGU/o6+Tb+m
ezpqE/ztUMIwWIAiOgx3AbISCiCfoIKdWyEHOBaa/D2n0D9mtdpFTUn3SLovjadY
bXXLLs5hNsfz/dLRZrNfwHAu7jvjUSTWIj2z2WUkC5o48ayXr2bQ9LHCL3QTxU3L
ycLNgwm+bO9Q3KuUl/CTAFR07ZqTzplKyhnJBlOeDpLwNo1i+PSBjIf+S9mAeSIo
so5ryR0HWKLOkNvkump1dU1x0SNjw6Mwxll3KYTAHiQrnT/8btX9qDMiCIuF2eFj
GLk4czg9ZXFvYHvH0WUmEdiZtitgXvrkwNqLvm+H2Lp8Ymh4ImaHBGZOwgIR34dq
QULPFBD0SoclfG0gvcOEkRofB7Txz6UkiWAQ6sfVVkUAcMqVeKjdd9cTb40g9fPS
qao4zFQoFDq5FFJugoy1xYXAZepYYBn9w5ccsfavBMI5/7/6QThKeeSMBQetWoZT
H15oVaekVKE5TB96tAdC0pL78pALMkvPIRHmqB80Bc+NhLAM2P0pRsuvb1J227GV
2njgHceYWHqGweDhj1EWkMO56vVk2Qj5XtLBg2xx/zCJrgESBVxLp5vupJh+U4m5
qc2ghUlZoyw80e2SwHFxSwjs42uL3ViSJXUdnQtUc06ABkSTNitTo/mz3CY5woC5
9i+rUeV+4EsCMjgiatPQy6Az1azhAsjwScsLz1Ixrgry0C4GhzADWvvuoQ0RCljX
NNQEYfnLzt5H5KOFaLsI4VCSwaUeuohILeN9/NHZOs6Vd96O8yhIPZvgy6ACHNTU
C0t4Te/74NuYC/PJXa2Jl3u1X0VhPiyPht/YGB91CN7beyGLjH6lvyWeZF9V8Qp2
hRBSev2M57ODBiLRuc1NPKN3yr0I9SFk9H0GNhCRKyJKHCu1nk8Xc3qkoVnOuMTX
L+zpQ8nGhX3p0knqP5wKMJt0KsZKZ/OLfXDWfzGg5PdcP03TOQaz7xFBHJAHoSZj
fgxQ0CU8fQX2L5w3BbwNryM3SCbrSqJ1KsXovWxJPy2r6M1MljZxHeTiL6iwRNIn
oaj+huB/kfOlZIWpMg5/jw+qKBY/5F5EO6rlAB8zgj52ITNKWCpGzzPSqg6kb7YR
AKLdDQPdegVOBbLc4R0aOBCJOXUjwbBG8t4lSZhkX6yFD6X5g5HKu2VR7w06GSdF
xXJHFUrfOJEQ87GnhzTEpmsvuGoAin4EAT2Hufqs2X5z3pA/G+jpZnsKGOJ0BNyS
u2m6xr8mQrRWq2l+TlzHMa05XTbF3txlhujS9162GlbtT0hhnftJJhpwOoQEntMi
Ik/CIh6V3NV+6773Y8ELHWSZayTn0EZ7GUMP/SBLVayEswogdL20y3LPgz6DYw+X
vI4NVvqkheniJNYv67eAvzAtVh4Oa0ztigYMK3zDAKPCIhqqoOWNzXxqATWJPr6f
QgTwfwBDX/r1ZCtN1e/nwnJ+2HdOgTj4klLfcxIw1HztCrrqoWp9Nj7aWZFNTQi+
mEi8cRBcYd4eJgm2Sq6uxToS4C6+K1ZnPe6qEVUeBJOnUQzGKyk46+mFYIgLr+sV
yaftSQocP7sEUHpoEqO55s8Ux2rW0MAIcVQyytZfCo88itGRFbwzLOHNCKasoe+7
HUyI2cWs7LWNItQ1qdstowRFmOklzL1492ZgCWECacq2KtvAigVDX3M7wGgslxZI
rjHvMe+hg4myd2aGefHnvhglMI2lWNUDTBRJx+2GzpDy82W5kUVH5dMM/twUSA2q
60sF1C3QeRbXcWqQHNImSSgDqHblspTCX9S0xyktermXQjmzgCH3Jltp6E7XQ5oq
UhhtGOj2vtSomIETQDv2Bc+rLCigJavJ/HTdk407PHAELghVxz/jG98V5cooI2Lo
4U+HIuix11phyMO6ep8AnY7ZC1vHZE7bNWJQB8peCI5oXo2vhsMx20yvhK33NIc6
rkUe+dNiyi2tudcgjH6I9T08jiz+mmDNeEjiqaB9DHhoRgjGVexnfNo5nMtqXf3/
2Lqft7aGdbGDIBN3uaUOueHXwPbsiXPF6U6zIe4fkUg6hvx9vCXETYhn7gT14JIt
ggQBMxWP47+DMWflz3cGVK/HOZvOv7AfLgNqA5Ml61c/CwrpczhJk0S/r0xmxoI4
IhnHOy46lxHCl9KggGhsanOvdTqC2w3dBY/wsJQbA3ih95l4fOlSEA/PBHrKLKIb
0djveHi9+c8leohjVWvjgGCCPy/pHmXnkDHciIcVVvJXxFan+lQficwADcnO4ghY
bRvlV2DHFDoVIoLblzP3muc2gD7wNa33tqOlctDXFR4Us4zpsKNfcFf8Ou5Gb5sl
e12EiEPeBg/cJOI6kvPQiuJWT1ZxtXMZFGmijNOSlWo9VKpK1mKqls5XYYTifTJ4
rPrNInst6a3f4oHT/mVAXD5mZLc9+SweyA23JesdSu8HEWEZXIe15c6K776hTeYf
ZgWIuhhcwJKIjfUhf/raiqwqz/J2nowATsRo2KvvtT14ErI0pbmQKJOctUaV0GlM
OjtYEt07NuO8vfHM4Qy/jYicX17jg/jP/1OGCTbrpDCZ8wo01LsY+wDYGrxR6gBK
S9MVPbmgXoQ6eKaEVJixxukbDUtMKJcKRpZZWTSiKmZVpCoQvn+5hNRCi0KUQskN
ax7GiAE1aPZND+OPt3ETpXe6E+6fD2HClYl6uxY+sqb9KKR3lyZKxCvIMIroekqG
johLhWRUCOdh8Vbg4w5+WKZ+MY1ua3rP2fyDVYr53jXuIBr7DkGmmD9tZe42bK0c
6W3pr0DW9dZGzLdPBK59YFDw+dubXSMqtXP+2Xi0cDS9MaSd1nh9ZRLhga5cdExp
qUWRl2a3S+Y5l4SpoN/WtkuXoHA07oxiVBO6wsfDWwqdIaIuLHCKp1o7UkxEhwl6
gn4/RcyGgXVzufzUpZZqQBCy3lKQFQzE91eyFEKIWJuJP4I3PV6jYPPUdrlJ3P0g
ov1A+QAss4xTed8hOL/NT3HN5JGyHAGE6xVeOVlCJxQ+E/JrhKPk1yHdjRfrcqDW
EARvfqfxHRyc5yA5AmsSi80LC/nbYVOkgKGLurvs6sS+KECQxp+XgENHHMIvwC/Y
y5XcKJI4EtxtO4foB3UGpCeB8V3hFkaXUd5Ul0BAk17RswL7h96WuR3p2DKWGKx3
AI3Dy3OjBkBFj0m1Gzoetj/GIUVGjiQ2ApsskAiW8ctBGRPCEdG0WyM8SuMcdZ2f
UOCZP0sByG5sFQWpciqCO0yJGuzwctJ104W3qlR3P3RLXRw9jdfzFi9HlNpRhoD6
JrYrts7CNJgnAPLHuS/lgGltTHvcbSG9E+GkYNaixUmZOtbMfkBfPqXcx+oSPdaM
F/7l+SBE5C86J/vvScSmJjDH8NUjTIfwZtE20LXE2ftvWcwk75z9GlC1gZRjESrS
7KG9t1TvSkLd+YYE/tVcYgKZxxCq7iOqfL2CVPBhw4rs2SMcu/jEdL+PAFumrgHK
LlmTa1yHp618iqKFDp7I82z0xlD0IuhrlLowbutIoCFpOAKo1OlPf9FAQXUPcyFj
AnwfgT9GF1aWFqza0OV5fx0VK/Ml+mdtWF2kn8zk0njheZxr1a6Xm7TUDWukK6u1
tJQRpmkVgPqMG5dAe/13M3FPwBYd7R5++xbyp+grWVeS4qwzp70aUJ3v95jIB4TL
kpIqfuy5J81IW7t9jkilMvAub+Hgds49RanERySGi1O69YEmxzrPQ+ktn/k/SHZj
JJgqW6vkMOjNKM/byZkGd/G1X9Kz29imJgLpvfMNF5ulQ9JxQjn3mqQ4SJVUD2u5
hOGxi6E+jcvMCQQPmT5g/gEFVNfWi1o+Jdxv4DTe/njMEpc8x0HC8ObfFbWfpQTd
EQXlPLjqWQ8XciW1F4nCG2CpOs12GS0N4PjcnJpHNrpcILTYRDxWq/gKulN0uuo8
kBEqfwxZ+ucqUOvPh2SVnQzx3GVo3fstPhw50oWI6UN6XTbQ6DyQiACl7+YeFQKt
mNepthCb8JiJnVCEhsjudP1Zj/CSuV/BFFvHkV6urG4e2l4eUI1DFvc69hZ+j734
O8ear/TKaJcgJzQwssPBJMiL4lf/nzVR1ThBYEgUblb0y3xfOu9rdoezIv1tBYm0
o+8fnW9Ce6HPu86SUlxMlNMCWTfs24MQC8LbjEHHGT1Ge+k2eTbiTvCYpSW8pKD2
pjHblLMdZ/3yICP0vhao1vWOGozltgvLFPXNhobc6MvWuNOEPyRiRSOO46XOasFj
Xf9jAbvFrxXl8Opfngq6MaSBPHudaay5a6wLwRNirF4zY6zgU3OZti0pRlbtEyVS
0AtSlxrYhwSzJi9k24npSIV1xLtPCCePT2GqD7+UQuEeCRTOsWsEcqkSdcTYp6SY
quPsNVmCnBCE9EaP0r/rlV6o2N3Y8StcNbEVhi28+LWqZkrb0g4LzhVSdIGGSIAQ
wYc8UaJPwILx/wUgFafi9W5sL2wTa7qLKt/dYFLmXy6oabZJWlUhFgdKvV+7a3OR
gkbm8h5AzLqJxkGT48mcQ00TIK2M6zAXE62iqRcyQWxDzjSFqRJ8S2fRbApXk1Jg
iQUO6pR1xB81CEqivwdYNaB1TlueP5wn73e3Cz9OIwRa0xEYIqcN3iGlSHy3gH4T
DBt2Dy+uR9pyOw+RSO+5hWObQpsLBMC48WE/TqK0NyNqEpD674cdU6sDWweFer4j
awWSZngaZk/3UH9xKEu3jNt9fBWOYn9EExPI/rU9q0QCNCLn1L9vMSIA4pZJLe77
79SAIlovtHIzC07mx6OvGcNYwkmTMtml19S0bV+V5LzxQtl1LFZ6GxtsQfZq1Rjg
8pVOzTMKa3kA/N1Q+OVXajt7b/ECGZa4KO3OL6iSVOsgth4+4WOwUril7JlluWEl
yx7dOgwm2AoGw6xRqcqDSXjbXe7HOY1weOsK/dzwf3ke4V9i5M9vygObFxHI7RNM
lKcDuJKqAdLIrT7ttBFsfkYdRKuCoENJdtnNUFSOnxmMWodRtf60iVAmu3Ko3MfD
UqBnj9Lv4uURur1GrB8rIcG42e5SBpishkF5GBR8NwwTkEqdLWFIeIIkloKxRbnM
aM037V+TSSCc+r475k+BhOckyR0oMroPv6Nlwvgacw1ddaZ0MDQ7rTWRTJe4XlcZ
ZOglJcVXogLBVXZnRpzz1Qq8oGySmOxqqlpvhhFP1tbe1qd3H2QQSFSVnGZhmAf2
zlUnQ1+PLkPWWt3hHm6E0FbJSJu3uAk5qVm+1eqNq4wmbot9rd6Xg5TLjl08xYnM
9+mXL+T+Ec+fjd1KakWUs/jXYnptH9Kz6f2JfBKRqOhFpbe7dMEaZH7GYtUBtGM5
8/Dzg1ZkoXd4WJOvWzWMTVqfpMMHtrAv7isXPjHUz2c5/2NRW7DejPx7FkHyT3Ts
nckMvfilpij8kxsJSYPpByw0YfXxKwaeztFWa9dczC1RrY5XdZkW8j/KeuFU6aos
4DAA5XiKu8DMoDtwHUqESq2JkO9MiIxVf67hbazqFV8hDUU7EcUglwVGaihJPSgC
633+c2B6qm3MUTypojbN7oYfzxVw8/DI8pNry4J/io2Qo1Hp4l4Y71rkJQ6qN6Je
17WMPXMLWtYCE85astMNOaqy3GB0R5CLboiMPEL7OHPdyH6Z8eYdHPKrwCWzse3E
vq6GOitY6wY2WUuvO+usn+jGU/XxMRROZsCXGBUp16p0q1ssiaVwtzwJRidLaTaU
qn9TaMhmrc3ScrnPpo+Y09cQO3aMkTVStp+YU6jcLrVkK6AM3+rEofW1D94NGZp0
6eWETRzlRU42X4FayubpL5ibmaawHlozwN4bPcOCnGHWufzmbAtjmPDsUjSHQSev
s26UwV+YJ9xLHq9FiZS/xKoXIl3gEJ6yIARdSLVW6/Ddw1cYBvUdNmwVahqIByjn
FmmU4G3ed1JRqwexjHS4PNC7VfI7NHxZDDsLQ/TJ5CbFG3BWXH8SjNrzYoUC8CbI
pJ3eQw3D0cwZbSvRypTGZdPqzeAskjK9yDiJ6l+xy9sibAZyl3a5rSz31nMv+iTI
3yfqT1NM7Z96eidbIbXtGscvrYrFVoE8r++b+Vkl6X2uqdiZF/lPaUoOgGIPMpBJ
Qowke8aYyFNy+U45j+EuPhBuClG0APBJY565YpZyphqZJXSSgvwajN4lbCBKjSAK
du7a7dA6oDdRkXly20/zGCBWPYfhFUjbP7obkfAX5d8dVKuHEfmr94EehAZCRJTn
pV7XmLwWVkVww9X3ujskuLinijX2b45bPfAYkAbpdaETH2U6VAaVZMXz874Xauux
MCgVqTOniCTmro832KoL1h01HKqFQvtKGpL5HE7O+Kb1Mc0fI+Mp5x4ezOw7ed8e
ORL3c9TKpGyBMZ/IrW9RMVI0KeJLYJooU0jZrezVQwVsv9alxOrBlBWWkd7+pk9N
/ycyo/voMl0W7ju1UYUIFWWW8ubs5TnxcTtotEzh+fkMjqR3vi3aG963ImFKbT6y
3CGZ3z64bFu3mn2ZNVH3UAiUGl7Sn6r+u4vX9w5OVP6k/fW03Vjhd3kBpMQwihRZ
w5Um6LTUXPajElaCn+wMg5ud27M+mLcr0AS6uWPwwwdMsVDks1pKqXQ1kiviJIZA
2+nOIO8rYC2M4GR7eu/lC6SLl3sjC8cs8FpB2MhsrVExSnztH3IaHTeiPTXHbYbB
qlH7grN++y1VPe018hlgjjt0TfFXdA4RIZL4AokYCmeEF7Pr74BDDCUNrTrNKw6z
g3KLchRXOt06LpGFISdDfRdGgjKDt1p4y2khiKePgB6a95qiPLQZh7XC0uDTie/H
30BkbybmHqKxxIE4CZlkR5FqXRcQg9pkA2E2jTkswlIsrredS5sT8eb1z/ZdwK6o
2OIaOsLx0/VAo/jIi4CArfRv4jwdlI8e/uyRuCxZgcrjzctjPeLgLtfY/5BTp7HB
j84CkTMHacMtGqtdDwAF9/UCjuelVfnZeiPukn326a4dUG6JMlAR466/ygUNsn/c
F4X/mWYaxOrArzKXpEhXGKM1IU+nZm02xj+3Z875vsi18vREnnFitZEOvi9zYhQQ
GF7EcytFRf4nsLNiuJhZ2ARLGqW46UU+e9qfySbq3Irq4Iir31mk2epDXniPMqMw
l8BmfpCaKLRl7K1aaZVRnLIGz7l9ojgcThUHcm1ouhfeVl+3Lg3Ny+zxJjJLuc+P
9nz5qkv17SWXapkUFhxy66B/ZbUouiw6xHK6KhRYLGNkleKg35C2TwrItjBHLB1i
GELEdWRUIDoGi0FfP2hnbN8/W1cGbZ4acm+QSfhIiIlvqddcJpV1q5KuNP4m6Dkb
tSjSN2b4ivosSHVMxTl8l8Gfo2qUhZ4rHKH07gG5debl5hcZUCglimOM1Wu0z4bR
WAMNcl3wulBuwTpzv6GeVBzt8RhcLCH/L6q67xqXzOj6jLPEBJmXaNGD6oYyAYTo
AK/7xonaCai0Uugn4kXju3hTYO1EsNB5DiTCbFWR/yeSz5RIWILhr3aAFQ+UwCWH
BdZHeC2HLOtOJarV6KNAVJfpAd9l1YXJryOQuTAuEzuoCivxRBB8QutBnyKukaTT
vAfHa83x+MUD344HGdxJ9yCrHuD5YmqV4+ZIXTvHUzdCcfOBj9eGByVeCB1KGiq2
L0oP+E0hd5SO2tdXGUh68NOfeZYo8n8TnL9F0I/Ss3g789wVWg1cTSycf1EiKlXY
2tD0FCvmBFh9w+fFzHH+wsHR6PUhbfph3koDpxmSSnTmRA1p0Zwx824cDoTr3GRt
BFz5RxLyAO2X97rx9HkqldduZZ/B1sQEHchxncmuYyl4Mqz9HSdOPPeMGAd6Ca3K
siE71UkVuPztOt47lP9M9xdjB5Sjy33QIZwYtU9sUSstKxNgZCS06nvA3NGw9XCN
uDK41JVqyW0tB5aSr+NyvOCg7F3H3RzyJ2pjIFtvbhkwYI9moYKBcaPT2DNCBPew
w9pXlZGMLs9j2QJSZwbvHZu6Quc3JPpeazIzh9V4ybOWpH1HXgmOtkCn0bH3apAf
XVvTi7BDYfvXoIOQy/7Tv8pJIT/7NWQq+K7Cz5qFWq9tGxkElq32XjfxpVAYve2J
TDU0Dt75jJelAVh0dgfgYcoGCwEWw85ee3KgZ1MTt85iOA02Rhg/SObYVPgAQRpp
SgzFmSmNBbAxAHwtjYB5eQ0BisOjiF6UtmvQgVWR+awBW1PQiTKGCvz42lpBtZvp
rV4PggFna5PUadofBLzD66dMxxT2HT1GN/xyoYLpZnVY/gMDNuVMBSh8uBg+6WKQ
ikKlRwhKO4DV0XrWtti7kU46x5Hgu0s+jS5vN+qnBiyX2lBJjlvqtGQ9Y2+uJN5Q
EbBf4zS6Zdim4L0xD4J7aDlvNnVrzr2M41vUOqzkKyArqGZLYZzF+ZwBdHyyf0Qm
//6ms16ckRAKwVlLiMem1l0E5CAQcez2WfYyYsqcnAc3qrCZsihaASo5+hrc9Qmq
+f3sH8F6UHLUA/lbB2R5ArJRTelDcC11jrH5qwjKpr6vfmFtnWC+YWVA2D0XV1h0
LSzXgdJyWF6vRP20RyegCt8RLQhkxlmwe3vC/irsmWDkd2U8bVpS6YVK/pnFqFwE
3Ub1aCKhuzvpiqgbm0VwygJFwp2cJCZC4ICjyasUbe040MbbWgWvwcaxuz2Ulvoj
w5cS9ayWYSOZ3/UMKsB9Uux+WNEResGYiWIx4NvkNfD7SA/6OSLEzcOOUY0PFlq1
h7gmH6V9CHci4XrWkiCSkmOa+lm8qAnMbu0d3TB68EN9hiiY5bRwbcSHhFRjsu8p
khxJSgj/hR3ObHMhyPc4FNkq5sVe5w4LPJuxEriUDZAlv8eHGOs3nDBkfEEUt1U4
/XP4JwIUsbWq+1NcK/NflMLTWs7S8Y46dqr9k8evzPUpmebFhgT5LK7t2l6r8ARW
n6HOIoTwnfX/1cJQ9NOtC17OA1UGakoAbRkJb0VMbkb9keLg3bxZcIfk6V43Alt5
c9UCrrATEkOumUJiIK2zw3MmfVkhxgF3FnFXdOzvNJILHY+j61SVtGmTdjqpUjg2
FnVhp49jXEfy5GGA3IVYYScbJ8QEzbLvnfpxtFNdEcfKQs8XYR2lp/9XVdagiFBg
HjayDUTYAyY8qRFISZP8+u1ds8mPMZpSF1jiFPdzmu4sboq7KJ969JHxcHo7mNOm
QhK7JBHldVBG8JoESfx0cXvO4yTTMNGm/uqTEvZnz1M6aC7ncFEvDEz10EuNa4Wx
uOeXj6DfYqrMLwGamxhd0IA8rKinvIk619HPYlo6/+Eb3aPPxvs6EP+F1NGDIRk0
efx+tN/sr6PxkBa/sSdxBNWvqece5cy2PCVIM8Qr74aL2nFPBlf0guJORUNRep/T
RXIZyLh0p453dmik/2S72PSh/1o3FVBsTPcZ/m4M+FagZDCKgNNVvyTQRwOiPcPP
+xyzOu51MG1GncMJaaDqPlDd7AA/SRPVS4ynIyYNg21tEKIaZRR2+bUPXzwZJlMV
ujdf8hyaBCc4dAmqtuO4GNdIvATiHse8JuAXwGdFLF6uTSEsYQdbJN2CwE7ePB5b
adGVW2YAPygvZ/wh6/pnlhirpUbxWAG46imqLnSEWubrh+YJHBUW5wiLCXsaK8u5
S9jMGX+BxNlt4izln1noiSR8tu1XyET9bt+33QGNZ0CVzPfdJfIMw3KG/1XG43eO
vY++NEDG79dNihtDWuUwasaRXX9BCTTdOO9wnSByRPFgJXa7GpgwxLHAMnLYdpP6
zPZFD5IbwJFF0cTBW6Wv9cP4iWTbl2Q4PhGRH56OjEWysraoYWa6H9NLIGxhx4hh
cfUdTep1mWSQxMefhxUkOB/OsMQds39R7iK8mEJKXyJGxjUmUOTu/vwR21a+dFmy
Bjj0YDCOkrW0jW6TNYuL+tJ7AuYJooFiSTDmBoWFq+2WQsAJ5KmwSah2KiPVHEhK
rXxA++SlDZbkSWkdlsEmfwUA5PqgzMUoouyTlRYeh4SxbYFlkyw5OeD5byJbAbho
1I3hsvlhOs6Ji+n7ig2m1xEl/Zh30miB+hCc7EWyB7uCWzVgfitVBV3JsQQcnPoa
X+xWnwthT8JdF0ZGCNOEicbfMAxMbs1q6M+RgBepfh76SPNEMCP9/bXn4DlMapTj
GLg1oKPvApUxIEXyXdVXJZgYBLXnDLqXwmBkdZu8xTOY8Dgbi7t/usYLXipQwvia
DW/mT6tta+ndkpiirWPN0F2R74Py0ItAG+Gui5e8W1NMtSHqyWlxxlY9mG7NZTJ0
ODbj7tWRu/2TQCldwbkV5LHs5ibIEVGtvzGGyLwDxFO7JMlB7/dw0d9g/RSWktCa
MkqWm7Xvk8AVe2FiPaGEADObzkLvhXOfPX6BUKg3rk8mZKWsJp9AFMYLpQpXoPO1
HXd7Mddhu1nqMjtqR2AZHKyMRpbX9bsdxbAz/P3BtwqIicW2enod3BQOgnk4Gr+6
FkOzU5RUr7N0YDmdrxsECHDhDOGfKmEa/u8+uMmiHEm6eOSZYCXEzZnK9j02w1GW
Jd3r+Pzz9tawuQWH4l5c8s1wGHFhHiCX3B3B7mXe0umCsFRCy5OgIMnxBMv7iEBT
Lcu9XWNdy4i076TditW+MUG2KPcUPhGx1H0h8CsCGk3GEhgjHV9zI83yZEK4uomQ
8HVPP0JkW6e826FpHRf3Sm7W/8tSfhUaMNowi5uVjE472LJq8ZC1404BBMbJUlM5
9mMl5HMhaAZ42L/B3crii2cb0ARMSrdMlGqT5Yz4NnzsmzMwOt0iSC92S8qZql16
OErD+1lkUoFqkej6ZGzilndtz3cLTChx6e+K9nfeXvaxVkOCHA+v+jk+BdAKEIn9
4aBlvQGhld2/VvsDTOV2xvKtjhzXJwi0GeBC4WqWrHaaygq0NFw4BumLZTe3D1Zx
T10cdwF8B8NleC8ebt8xDiu+cdJVHkkcAzEMI6uKvGIt3mukFUlkckR8QNrDWdGL
ubhpv9MIBQ4GSzmidcMWbcyfEKIszCLHePSXvTvPjqRa0ukpqr9DjO/T1xd92KHe
IkYNu//wmOy+UqiSdZIGQNeptSoJvD9TQdaxLhPfBxQaNZc7xGxUjWFBUsJOHua3
03iSkOifHe1A/DExPyYJmxH/aNVTkFhvYR7/XOnYCbxlaCIqe60xaAcAM6cLDial
IFR60t0GVXxpRxXqe8MXkIkiAT6/lgembwSYg2DAf3SSrLMWj2Ggtc3MAchFwac+
xqddoGpFUpoJWDjDPA4JpzOtPg48gzzob6zlOADGuxlt6t0eCoUWcdydpNit1H/2
OhLwdH+hD4W2QbcD3ojISTgfeL4rabNKFhNCp7lnJVTjN+QePsLjHJH0T4aOY9QQ
XZJ20nixZpAWWLYMAb8AjPQiV+4BlW1UT380haiq3hgpjoaxGf4Cwv2gc2LoFE+X
S9KPuJJ1bQpE6fd4YA+t8tE/uh8AkAAZScEYkeahNIUxDqcd5Q92ZyPsJzTF1nsm
gmFiJOUeBcFpPS6G2L+Fk3eE78xMCqW47dpQbJkIjQH3Momk50rk1SFby03HNj1E
znkSMsb/mChRRnMuQ3+yn4sUfMG5nGQvbYVM4nvVoEg0OGcnh+whL6ewBJnms6bn
oej5xgTKN+e5qnvkPA6wK3CHQb2pti8N3BqyGx1CwpXVxFrQnbeA1Z3WDaGbYCJH
aTQX/G7QFL8hp5xoE13ASvSK9+T23U6t8d4BoAmhqZyleTBd/NnimZpxbG66IHFN
TnFOl4rIjGJntsJDo5TaRW0QUuDxsBoirigKLySu4irMCsV/xuqs+EnTF13LBzfD
ckeMG2Uuv9q0PnaW22G84V8pUSuq4wJBn+GWX19HdtEOhR/6+n1pyxgUpSuetczS
ZS5EeT7/VFnGp4AQ586i9UZbQeqk2VrJzO8RfBoDE3ybwJ2ThsxOUBZVfTcqSoLf
eeaGZsq86jNNQ7AmsYjowgPex0Ev9U4+Lzz3+TMxaU2yTyWiFJil0jFgCT8cQzDA
g/m1Bu66LtndqER0Hbk2dpNUJTYIFsp6UzjI3G5wSB1U/QwKrvwACTk4zpCcUAQ9
EBRjAcQJW1J1Qb3K/bP+6fCLpq5pxGXYTqInJ+pB8daquFnzdVWxOPMhCiaKs5A6
QYQWkMwtfOuDFJr5cY2NytZbJ7P5iFR0jTrU2xMUA1VKnF0VZ1OM7IoPMeTKjfWd
gllrM74v0WMMf1tClTUggkYRtj9WK2jt5d9ZMkiSu/PbXWwpHRLOun/QMP9GJ4bO
deHD8x70601pj0mwAbL30s+CcvURaa5I7ZLybqsZnSIOsWHg2nYRPYNwX+QGgUWx
C2bZ83wj0wTDLZ9z6tfsBm48YI3Lxwgkdn84STYvmSMt+wSAah6UEPHt7MTtsPl0
ZB21tpULdPb/zGMoT9HOO/7Z75fAFd8/wKx25eWqftRYie37toxjQW65j8pJH6ZE
alYXjGhnaSMQ5eNZVub6GU2dzsUm/o3uOKg+WgPbgtHpZx04AtysoDcPfLwhs5da
Q1BeAVf6macXhyvFPKp98QXcMaM+HqoCSr5aquwPqAOeQocr0YUghffGPbOMvfC4
XVrfmvdSY+f+A8YaQyQlqM+KOGUvi9p2Ofx5nQ4pICz8kEsdljA8j9Pfhu8C5qy5
LysG5zEy/Du8rJzzEd0e9G6RcFCCiyYsZBkK1ux9BNbQ9fFep0m6HK8i/J6q8yh4
jPrig1Cfu7MagykpMrRZXZmuMS5csFeN9QldGCRNxLyqVr33y6243tIQlRSVde2A
6aNTwvFxbGBE9DWkqaJD1c9r8EQUwTBxfvSdTXF1QeFymYUHg1tRzWLEW4AFiMby
EnU+SjiKc+lfaPC800sx2fKTeFg61QYaT2AgWSKuDDWQTUeet7QyofFiNkG4fPoU
oe1sDRwXnFBpcSLIykZUlLxB3nVSmMlR//L+RArZqKqJ8Aa2CsYUIt232ZyzFGK+
8AJzfEGMQpRY8wdkOjq8ManneyRtZYNZEgMTDIftXa7zRZCG0qKDopmmfrbJa663
LK05NRe9R7qWpA3GS8PjQZUlGDr6KY8fKDtg3G8N2mwm3MlkyDV/b7V7WygNLg6q
drRYYY9DFx+BCBEKN7Kg55o4dZfHtubuDeobJGb9avuKcVlGEaVUKnhsun7TRP+w
+V2GqysncSwGop83navUS1yMceErZEYfSKPYjIV3sGshynglCWb/z5xeLiqWTnM5
urpVQofArAd3/eRNQ69GDqKHt+4psqBag634w1MihTs+fnJ0Jd7uA7lFmpZNMpzT
0yrJRSwZggEBKYwWvO4DX4/hv3/i8YDTQdSMennzZI5foPIXsch5nS0OsXjEXQAl
oKjHSM/O2DpJZbhrkdj3wbIe9XDt/dCS0aExgR+LTjRYUxed0cLl4+79F7qPcbk+
6PIUCB5IXn4tQP3ZQGEeHx8nei1tyU+NELR0n4ZfbXt5NzenjMTirgX+nI3t7H4t
+EWGiT+0DJNaQzZoJBPZEGmEgzUjpnXOsY8G1ZSmfRn603jspp4ZqaIitkBvzC8c
gn8qtmIzChGe74vwTEMqUJ3RheeJMp9/5KKDJ/UEY5eSPRJUx2tqD+VTysQzSAEt
0eVhI7Vc1Jb3lmfhH3qnY//UoqcA85SaeSeRGYOIhSpTBE0D/paOq2VLdSWD76th
7lOA4owQkNt+BaAK+rHrYiFH/O51QLj6iAZybqh5XnULhmAPLdahRZAG/fLh8YN9
0FO8jncwFETLskqad41O2OoMIFxfotuAzO6k7p7WTVknmowrFqSmJcqw1P6tKus7
i9mp7WtBA1QJyXXxBbiXqlX42KUKJFucPpIzzJNh3nYBItZLChfS+Y2URF7HoQrf
PcuyhW75kUBX4QFF3xMmf/x54C1eooCVUfClWl4PvQO+jZM2+CsCKly9uolLE1y+
ByHSAqyu0U7eNsDkggGonwFZWwBn6WgUbhEI2Q/2SD5bqFviJutb9IWdyQJa3OAV
lWs5oFHvnGZyYtAVXncldKg2gtZPbUgOsSyw3jOG+WFSZp4NxZSEXF3AOc4Paf4J
FsY9oeHU8UuFoR5bVCctq2QgU4H4O/Tkg61ondBRbmF5PCrhiMaDe1TuCYXMzaRV
EGhJlvYa6awlEIE742nWF/yNs9tXRA/JakrziPqyEEgcyWD+jixXPTpDxn4IdOF8
g6ghxBkBR1xii5Q7QGVfF80maEYYfNdDujV6s0Si0wP66DgC0YWakO1+QGWLsNNQ
rpyfU1uRnXc7P7gIFspC7yAfl7eC6NnKSBBxDNeUg2eyaJi7OiekC+Ce1nYDKmu0
npEIllwrqCJihZJ8+efyWommEAbq5nLjTIyHG/MhvG/Bja5tzDRkHqy8TXzFulrb
NwYubORnhgDZNmEHq8CQ+9gP2DkDi4mUCiFQrhiN5koEgMpR43HNb1wYdD9EUY5m
y/VDl7Rqg7a6vFE2epSd+LchyGVUSnEMtzZJxDqD6FJvfUMrRsMJq2EZh4en7d0k
ZspBYoFdETZfE3dCveXJT7WBsERgHn2BKhPAMChD9ERPUed6eZ1D2ORhWXaKiKcx
xcaUl65PhcaNgtsrC+Hdi53znyGLICsI4XTLo/QDW3qZImBaYJTtYuG0Yv+p9H90
ZNlWeXtz8o/y9VvrZzDBhkSyftqYkZbgX+1ZGT4kTLZ6k2BGFDEMffFf2dKiVfKT
y2eePe+vWbNm9dILA7DRarNp2Ii3YTAaz2mdhn2/f8lWxi8G2vtNO0P3M2NPG0UK
PmE7cGTkqVD4T1BfEErdVk7mH+MHh3HVv0aqMDl2uxUp7nz6HQhi5xGwJa5P9kJl
MG2G8WSh37ddogaJ7lY7M97LlVtiqEWWS69HJuOBjn3th45tGSngz/aSq6Fhrgaz
guIIFTqq1Z1cJtn/ltTi+5qrbOPTNfic8Gal/lODyAQD2GW1Yx+cQcR4ybrVOB6/
Zfn6flYw1r/W8XGHpdO2Ao4Tg6mUH05x8Tkb1I3TBRC8PawJ1xYBk+zNkl8Uh/Uw
es2D1Mqkr0AvpB9V0IQMXMYOtqSAVzhZu1aOK84zTjFlFdc9lUTZXgReVYANkKUx
+8tKCfinWUZT34IRp3YD6wqX1rSsrtCvxPikCewQ3XaBK9YmbQp/RevXgHmBVFNC
VH6RP8+W1NviStN/VF/wCILK1tMRG/xHo2F9WZKHoTa5H/ZBZxxYV7BErMsMNoYR
gzXL/gQ/hHEE05pgaOjTNe8qhVgCGtuUQUEnzsw7T8AWvItreqvZlmeBiU6azKzT
H/c60hbFhejtu/4Sdz4KYlrMEOVVjWk9Wovv57WqITL2Z9psqQAipR8Ngr1Q6Zjf
f7tCH05JNyYTRmO/jWrqCBbMpp3mTGcDpqU53m/RYXkIwWWVYyaKOYwvdCzsP98e
JYs6cZecXBIjqUdkw0Tal0m0QojMaB1TTBIqN+jpXaQqxrq8EMz3Jd9MsAIoz3qJ
bzs0rdiq8b3skTRMCynJzWbNjlq/3O9bBuIvrlyBrbI3rOWD3kysDSxhaAymcdMj
GFoMn2zqaQOto4QxDn+2UQXc8N8BGailCYoaY4jT9/UOBQiaoNb5IjwBI+T22DA1
p/lzpG4BbDJHFnLArPSFXekI9HcbiMRfXpsnmmlgudUpE5F1ui6UT5OCU7a7YM2K
7wLHHDYg3qRq6pLDhgMQv2WRJwedb/yBbGY/Na2n/twhH6poD3tXjJvPN76vuG+0
khkWvS7vXERAQaMYalr1HCSN8uGu83qgLKZ0KgS0ihaPmTzwHZnaiWQdfaIKXb4O
LDqbzAEjD8aUkbRahxrVi3M1zVsLXxZ6HCfnAJGk+UqKIumHtknjTVPQUx0nnU9i
akSgxkH+uEbnoGtnwzVvlSSzkUM0I31bbn7qNo6OODOMIQUrIjFx7RxcbW7TPHZk
TmU+T6IQX7QBfpaMNonTujmiw05qS6bH0nHRe6Kr0TvW1mAi2urMid7yUHMPdgs0
VO+XmSfzc3FPhE7+cq/teqFDMFDj7KFM+C9uhH0NQb+KLeyMhOCCjSz/6OayboPV
D8LopiPqLF7aZMhFqEDTb8esVyqch4TbNlMUzwcI/nArIyqdZ0rwD2t4YMOyAHEG
cYCAG0awi19EVQ/AypzN9XKJdGUvmOwn7COshiNpjfpMy1MATvxG+//m1M5T+m1C
imqGd1KvRcqVTfUS622Ou1R3wRruqw12BwQpGZQifKkBlERbRBVyaiFfHlxurpe4
JS7sYQsNkS4SQBVQIrjT5nq9WbvxIYmIuOnr+rk5biISGrX4JUZ67EYRm1VBusSN
RDUIOt7xPfAzG/1TR+7xSj+aLmzYEZLLG9eeF+2AoxSrvDXFAtbtzqRLYCklRG+2
0G2Tq1mXyiYvIyJ8v2Xq4HXlTnsvGA9hiHwPSr8eN9gJBJ4DCJ0kCG8ZgWcLRjiO
U2pplGPFtrRRTTmFHegFuuaNM2B+MyVKLhIOdUBViOoYqrV7EPr2GGCvN1q+B3zL
9dIF8nsldkONqZ4mT+kK1H8njI96KacTKHgkBhnptsSSEMQ65YKErA3Ky8CPBkUs
FAmsKe0RUQlOlc67x6095acV9uDlPmaLI+KVDyiQLDtocYnqOL2O2y2CRZJbufme
Akb5FTa5PA3I4eKGCIpT5VqFReD5cjEC7V/mBkrUKB3U9CdQ4GMMzKEgiCyYERh8
BgrOXq9M8wb6ShFC6t4pfhdjvW60EGvU+qMHL3iawgqj89DvecG+FCjoTKYzwYIv
gLaxBVOcJPnOmPTUTdWPWXswwlyf3LN2lBa0zFaW7iWfd2r8mFkbehtv7CvG40TQ
UTQEroyFCziBtxv7VJ5SjAFaXQEftqzZ2VKZW1Vuu7GRGJFPajHsLX/V9tZvmENY
7vv250O74FuGkSij/w8Un7zPZyTZsnIx45/I7iQDHx8WB0PKPyiygjQ/rxEPE5za
VEHajCkanQoSrUXBKN3GsAEWJZEiUz8m8DYMXroqbt66sRoOWXkbSMEcBJLwGbum
Wo7rRW3QnTWDZ6XBgfNzci6/v5FCFACvdLA1cxHBFVCqAg9Q/Fgz6W7GF/94m9tq
QCmu1T97JkxKIN4my69hzoenpIW75n5pWsBmCoUKQLDnDzKKoNZux9DvaWidcO8Y
HP0Jd4cqdE1hINUl9ZIPoxUnuDpvKZrAzHzP7EBHuhofIv4Wu0sRSw76rcKzqJ9v
Zkz4/z3oXmGUzMlMue+2MtwTztZq3BU2A31l+0g9r3JYRaswqlYJJdVBE/jOMo0E
Rc4y2vyYN/m9qKx6H3DIvQxt7oxv0g0XyPNCSuqFreWMfj5yOh0Oemk2trijnlkT
7AGQ32BpqV3Ra1Zb5+wnpK0/cWkWruwXfodiJKea7cQNiDjO9wpBwgQCO2Gs6PE/
BeixYPlJWrX18O68EkVSh30uWYAdriI6UePCYMhIMIMcUbUB5b73vlwEbsXhpx4U
R3AmAB1Sp3RmdZwENEv2I5+2whV25wJJ0TIXktBgiT7SZwhpZksXqVHRLuS0uCVV
UFHMS+ZxvsNwknyktnhm89hENmel7OshaUoH6yoJZBLwhYT8db/0O5mOJoA2j32l
9+Ag/3/CP6fuVl68bOGhKZC0oNaSBXA+yY+KXk9KoJnN8CAk5mnzdkKCk8WaPo/H
Mkf8G3rZB9s0Vq0H/wZjM0kcQqosRbsRZvB/Ki124ozQNDPorLUv70jeF+sG8Lxm
LNoOik5dGyHuEtDu3/1icr0FfEKrDIuNobdame+gkDws4VUqGVWVKqjaLRS0o9p0
KAn1zHWzUt5j4VqukDDpEoILkkLCIlRSZy5rkk914f/GQqIIjrRHwh8dIAS34dNJ
0QTvQrASqaTDrsSXhsRvz62tqb5GMKizvdQF2Z5vXvnfvGDxh2tXW5dtJF29gMSj
XDB+2qxVzHmiK0V+rrlXZYs35yixki1sYfVQ+HQlvbPiVEv8ElKpQ1JUcv26Si/8
lhVV0wedt2UCELsNFY7bpW1w57qdNEtOv0Nd7kLIQ6faoNPTlqLDN+3m14atL8KS
Ke7BVMqmYcDXC8urQ1CxhDvJNqEsMhTDHncAZFCscYbFQgz4ONvOfXdo/LyaF0gZ
9LGProvkWAjZCwZPavLFSwSbiTZaY0m+73W9j+F4TPRubSOHr2FsdrJkscAw4F+E
0dQv8iXhD0L+p8lVSHphySFk7BpyYvtIgMbauIQDEE38mvktI8zUvItISKDeEQEF
RvAxrPt0a9nhelcKV7A9xM5O4EaYm1uljMZmhmNEhUxLx5Rl3wxWrXuPlW3s+Bqr
/aGRr0gGNQ7LNJsWsnoE53vMPHDyxmy1JGn2GErqVK6MGXIVzLaGLI7mNBKmLUtk
pFFXut4BFsVBx/s19oaZuAAwFf5ePuAsXRWyi2txDQWu72YXpJum1+X4+r0NhKkg
a6x1c6sA4zBmv9g6WTqW33SaiD/CZ/48DrLeNcL/hHhHgp8tiTYRNCS7v/+QWC+B
BZxL7VAi/GFPbOqt1REzsb8zZwiRC/ytAizEuBNhdQzUlewTmUiUJlFneGxA/rcW
cMM1MfLggiUtW5+i++YwcHCBxicW18EJeQkY9w6yBeTK+wQdbwtiUZupObV6D97T
cRHwBcxQFL6vUqcMKXj152bns/3dyHmiHf0VN2t8RKEcEBR0zX/L2u1bRwNoGjl9
D/VcNEP7A9iESMNSioRR2n9lUO+mtMwWYuC7xN/LVqv6e/l8jTGpDy/aa7p5NHC/
L578HBDie2jS12GjfIdYDzXfsZn9zPahH5GB7TK263WAk89dhyix1tmrbgq3HN4/
WS7UO5mA4m6uHSqYrY3xFuJ23xJIGJ3dmjG2IcLnnArtSN3zAZxbTnASm7G31DVM
gxxCKC4M2kWuj3Gp6EjQwFaojX+MHCR5jtYycqreN+04ayI242/1YH4Zd320VDkF
7FKD6VIDQOLSs/0HPufmVdNUeQV8I0fu986kYYYmcpftAgH/uEB0GkcQSSchb/B7
/jKyA9AHHKiIj74HObut4ifPOJF7wUnzG9r9OiHLf3j79ORcIIeqXq6pdusBdXjw
jBa6iEn4g4AU/Ads9VtmmWgEVklzETAAOjf4YVoOydFbf4XmEPWn/PMxabYGhOni
DZxXlmrsMPu0GxV7nsp0bpV2JxwdUVEDjRpYGc4WtNOk/fXdzGBcs+7aR1omK3KS
SWs3nxCiiZbGCKyRavSjRrOUOFhjnWvfY4lcipp9OWaVYeMW8336sD3ei6lEikrw
8SoGUUl8AuvBSf3GdP0C2OUre0MMqzIbh+CX8YrH8COORKU9VkNwFSg8L6VXVEaT
gaFE17nl2wKfQNeg0b64B7plubGDUdU7CqCjicXQQveA46UYwqjhUDV+n4lXZzqx
IrB2dFKCSbqpf1vt863QQX9WZ/IkBT8UyPk9pDCs1QsGSBXR5Kibrt+Uqh3rX2y0
50NZieWXMRpHZ4ALMbkNWJYy8AOMfB63p2GlcoKYeHEfMPEwTENWUKnRqv2X7aNh
1s9rr3cUGkGPtk8U1oKzXE6wg4Va3g/jE+E9hT6zR8YC6I/Xay6fZqilwqonU3XM
2GQJGSsJq1awtjIKZZNjozBMgtC8K9K2luU3hDxZD+ntPp2gkuhSayUlXpKS3yhz
rVsrVpGnGxXMg6bV1tTRnrvLkmzNoEo/meiHK57y6UXUy90nPslNWvTYfQcuMLL8
dl2eXJAZYL7uqtikGXkzTIpbqG+4T9Vr+YSkt6sBt+rXnpUJB5eiA6kYPdTcEqFt
Zm25eydztlT5/AahPPJaztkbIwm5PJHScri/iYFkY4+PWUQrRwVzOQBMnQupLnsM
bnYyKPEtF+JMLQb9yr43+DjVzU4Nxuj3MRs9uYbzzgagbYIkDZMmWpX/NhVOIrQi
49fh3KVHTd4D+oOXJWISrRxlYYpHG6kSRScaKhJLVn6l1gudzaWoAhM0WJhGAonG
A/io7G4pCkmRjrZgnazSpIre943m4Jtl1OxHe8MhWHQzpSdKBjbSufmFvmcsD7gS
hq+QEaDcCGc8gDZ4EWzaRS3fmniJn4mCnyzUxRUd/1RYj56nwDVi92TPtGhFWHIL
5mdKLEaL5/zsmXLB0Syad0/PqZrPef5IG8/fvEElA85XSKLWbieQIKuISLPeup74
VBMIs2FXcRJwoCQzx5anKPsCHKAVZwCqti+WSsBSLtY4QfRtPInD8wGNgU2khkHC
Ee9V7I7ZFkhntMyWUw1VDr71gx7dwV94RzMqwtpYCHDp/Q82m6C+y2RnA6j4jS/w
IGUIkqBBREoCUgoebFJMvHFANDdAdWcA8gRBklpdRzZoULji8uvx8QjqLNDApEsZ
7ZhyK9IkJmdp063TCZCNQo4ZNRIuGHkNDxirRTYAshSSsKJBF7pw0Snk7G18rvNb
6QKoNRegQ1e9O0E+nFS5ggpb/Mt/RLwgyivWctFmqB1N9qa3wlJFlDqJm1IcjH5u
dVHuasrzj2dzJMdOlj2uHlY46IaLwdmKBQ0UOYsxG+2iAmkyA436lAhiZX0/LWAg
uTroMxdK/avw7o0jjlTuKgHAqf7xivpwbYx0s9k/GwHyoUGQon/zGVU6nmjFj2Lh
rjGLH4r8XT3HHkkL2XqMxh0N5O33V5VxAXEnc42kIamMEel3MFDADBPxgRyP7sFx
LUcVyomYDIRO0LA7uQmVOd3Cxe4F/Iqz/bWSxj9Cwz5CJRYvmxoHDjmLtqZ/2eWT
Gh2S5o+rgHv23bt7R3g4fj4OKY7BLRQOz73psEukxAm2XT4cMGVIbq6qrSIPPiwN
/x6WQSp6NesIBIAzMzrKY7Zw89xuaWoYcDvBi2XToeOBjoLJgADwx4rjiLdIh7Zh
PQ5OBTAqcNG8YLZym9X329RwgK0k6RMRNtUuLy5Hov3ynNHskqmJmWijc/awlBWF
CY7hv+e7dZuLI0DF+BOjskQ4BI4YL4GbGvDTJs5gt/PwviFbJ4HAOZRW9UlKfROd
54ltLFX1tvjkOX9WOpKtw1MhM6zySGsLwaBcKf9xNO1a1GuEVUvTTUqQM9F/un/D
v9oMQrmasSceRw0vLHqTP6RUHXlyBNZlQENgLyAj62hQDBZ1ORJW4w+jQ/CqpDOG
v80PLZf43GWZwKPnbq1sUo/ENkNTtYgnuLvBQo0SBsxHYbBhAfUZHVnSxPMw3Tg7
dVdlNWc5NjzOLaFem/xVUrQgcz/Hh7RzeSrO99vtS9NcQG1bNhB5xUGgKi0yFEGC
KBNvoJXTOFzsZ9C2vsqzrahWKYgp9c1X2MtHXKlfzF+oE8bJ7MDhIhlhSSvyAc9j
eoL3pwTfhwrX9ORfVWago9gG1ISDlQOQx7Y3uyNKF6ew6IzQ6hpTAmWUW9jH8vHj
JVriG9nIFQ3dO/os7ODkXXCNQyJV/ZdUgJHyyb59KbRg9tOX2AxQijhZpsLRCbuP
IccExzfHRQMyUA0jNaIu5FiLSgRi6QVUGO02vV2ht6WtuqJE13gMcQ1Y5Lka5KbL
kD8UI/4vxxxY264IoiOf5WAlUBTGNk06+bYwTYoabXPp7/s33u0ezJTo9/Nzp6EO
wl9gWsk2/HtE60UkrAUPy7d5bF0Pu26ABwV+CgCGwzGF5WT8wDTNJzZe4zWitIPr
qOD/Y1C4z2h2fpZpqxFOcjOf8DqVoiYJnI+22hOXgh0ZfH867d3ftPxbMV4g5WWc
ePFJ1MMTDDwaHkrjx2C8wjKw+AQRxzWzqGLmQZkhjfGmF8xLeRSJCqNiYNqYBOfx
B556UUGMAeiniKWeyRjYAhh6xzmsaYgkfbxYM0C771tAESqXOoaprzMVFz2RPTJM
8mjExfLX0ei8+gBGKDBCRyWRYBOpMar8IcCxjFYKkU3cSzutjmvbi0QCO6bWPIPD
r6Kx5Jp4FtFue5aXFiHCZt8n1HikCZDUYa2mYvTYbV2hDlRZRw1YCpb0xAcEZ+1b
ubeFxCZxxHFwuolSOuDJSONqVK6lrRqWaQO7hA4Wyfk2PiQKGZKdzOdrLd9DPU46
eP/DtggBSlFkumLiTQXCpiijg6CLr8Dbbps7ArAc+dlcJww1JHncV1JCV7mkeylq
2kRaOmz6NgCmC9FTkoCvp9VxRmdqV1wi9f3xWjPhS+s9M6iENUBnMewviIhy/KUR
9OozQh2clIME7HHyWXwjQLC3iJE2jaxZYXVmhHMYwWorsnTVrHCu+RLHV3ks3Awm
VIy9ZQi8qjLxl6aoNDRjL4b0DtbaVEgOiUbf5EBPLiee3rPfw2DzyHRlkFz50TZt
ukp1kOi0rAj0py09UsDOsQxljge9h1HFYB91sxdLpfg0SpnOIhmLHOmzyuCPTBdK
MTRBQvq9U0tMNw6ot9L3J3Zt8egNengJCgxzT1UnCjZs0fZLzFnuVEUmGkYvsIpX
qhm8N1ozwMSlsyBdrNmqhKuVDgIiXuWkh9rtivDXbRn70HB+voSd7hr8qgyI6UZa
2k01B32CbYRIHF4svqB6lyBozIO0lLXZD727G4Cl+rEo11rd+WEPg8yxnifG77Di
/jnETyrnoluCULHNqYo4AhMshFkQBNnyZJJMk+bPIfs71E4zs5M7QsoRbTAOad9P
8jZiCHkcETv36LXi2hYQnnh4aU7ZS+aa/UO/xk/EqCeup5mHn5ZN8ifRLhYHtAMD
WdghKXPQGFghi+sbiCxO74Vj5gGK4Qfp/LjLnuhYsHJrUAJnHTMXzqg5ealE5G4F
7uqYYy9UmzDaOn9HvapMxP0eFMh6Ep0Jmb5KLtUF3lCwH/m1B11HaxDrztZ6I/07
aMkjZwYrKD9hhs+YqgVwEPln8WzGUdhgsTW8FpCCajL4f3TVR+G35Vc72S8cSI0m
8Gdmg+ma821eb3kQyMyiUVUPG2sYqCHn+ezlO/8fnKCM18qFjf6bqTTGpTBUIE0B
K9euHXq6NpPFMviCfQo2wz/KC0eQugUFZuCuKTok1fCjQbe3BPtRLQtgNXud3ssw
AHPAx4eIz+TFe4iPk921k6OLRcVFcfLO5ZKS/qV/bhUag+KgYEuEpStMU7LNstL3
89qdOx8D7m9/cVS8CLfiCKRcDAv9si7YzKICoD7Pq3v+y+zUWHrufkvi4QHxQkcX
SEaLrECYoEbJQk6NngWpu8za1n4JXYOng0BEr5RScEYPZAeMI1IN+XKad3CUgl7o
2+EBqOQ6RG0AUJhhnnxnhpvQ4NrBAZOrDj5/V6pN/+Uxm5iwJ5Li/p4XdTzQMEVn
E1mK2a605Fuw9G2PF7RWYIG0Gm5YWqLZA0+TqkjkSABIlx3w+0umXQDqx54P3oeg
3VVm69LGoCsAmOGUj7Kb2zYXSMnVf8YIvK0+vyH+B6aX/DJmWoMAXTyPBuWt0qAj
pkFwItPXZXtdGO8eezKpS7X1GpdJm99pZhOuyNM0Qiyw/o6OsIneWAEMSMfTPYca
q3ZbgSCKNF7WuYZ+dTp2uf6k8OSOmh+Y3kmYbRCOYxEybiuo9qI2H7caDU5kenkL
Dqh3DU6WMP62efyThqOgupKipRLtnP9ukKuYsXdSdE6uOjD/jQpiuArpZ4xLBhqS
kwJXu3yEFMb248SilEQ/h2KM4pH3v1JPbndc2EWnxgKMqZLXh3Y4Q9WkCi3LVQyk
ydsDUF5K1ZhqK9ZX90SruhaUPDKNRdZuxq3mlc0uz1Qv7cp8u8lPO5r9CoPLFtVp
VhjJuRrg2Qz1uO99umgqHFM0cusBlXMVYELc2mxBEqj/wHQ5V6iuMIDQ2SAi29gD
MgiAqQsf2Eph/k4qtzI8d7lKsVKsZSy7rVQ9CK1j0i2/G1kIkw/JJQFyay3M2mcL
hLwylfNz0f8BPh04O5+QnsTQTuTbE2QcqQzHObn1m0CJXK+tg1P8iDcTV1Ex60D/
mrkbff3XmvpKn4Y+O05C8Hrw94fQ+VYOm/U5FCyC22G+j7wJg2tGtU9xF0Z4zanE
hCiMUZlw/b6+BvEjfRtIYHI27R8Q+bPRmJhu92lNd2MTY82bR9mSry94KPzsXeli
1nBauoQuydED974fqRv+DsMhdVLERkui5EN9iK9NQgjiryuW0xdby30bw9eLkWJk
kXaJyVvrZRk5cQMNBDioMmDLFUC1+heCoEXUKocjgLsCKnmmxNsW47S7ZSKPY2rd
5TjNmmAFHpdtqcZyYYKYbA1U8gGE6LqVDZdufhIV8m9Ar4buznEwRQr8ZXwMO7Q+
6cs9pQsd3SURH4SJccoVpIc+VBSo/7BEEZciRsFmwWr4oCAhlGKEoQjLInHnWfa6
79m3F3Rft0Glo0/SbZByNPkXkjig/GTsLVCCJbTZeIJp8LzDxVlWv66AurU8JBDH
hy3wnZKU7lfBIuWYbx7owr02xpmFBDg9w4G4oyeUpsZx0p1XcyTbebKDNkzuaCJw
s90RvHm9vfmnEvom+RAutZzTkr2qOIpBdq5GkOKh7rsfyEOJ1fgx9KaFfsKp34cX
cnZkC5U65hZaqqCYRm4X2sPnCPSnFwGuoVJNNe2lTBlXR34mqtSgBiK4pep2xlIX
hWi6NuwSxHCaNYjNxvBojyjGzvCf253dvVHMsDBB7jZpOJUqJCJVx/kMnRL2YDrW
YYNN6oje/AAlGNwrcA0mysM0cqTVDcAsZ8koV8d791N3yq1FSBpbpFHrrsOu6U6l
vIh87KwCjPLtoiHG5D+4HytTuZO0MXRliJV2Af3CSl/JJLYveKAF3jZo6DCtOZNY
xR5siEEgMr2X6cJRa/kgWAFq8asQP4h9kvFQa0mFfSpgG1x0AYYss0S4kV8mqsII
0jHIJdwP61lyrufD+m9hmZqsMOtSCS4rSVqlrgKb+JPvD83krPBkueNRS9Pr1zUC
JhVVGIf+v5jOw2nOfc6WjAjaoBHpJFBkptYLRRzqhXI5uOA6TPoKfY2hvWe8ZMDo
KSkkKCONUXEWuLudQ0u03/jmW1GyXYD5rPq/ToEHrWZZq2lBOa7pdgYPIoEWV3ge
GKm5LQCIuRQdLoMF01SIzmZKneYuhe7DMODyfV6JAqXY9J+7lZHMQEHCIRhUPTv/
q37pkK6Yk8Bin+/3W+FthKFF4tycxdNMIjgCYH9u3sUMqNcgrvWHadbfQFGUZEyR
aJjLA8mqEvT45SIJZmS+cYAbSNGH0LAQz9Ba3UKorpy3JC78n15nCi4f4s7nyHvg
HYCSPXr+VdPpizM/ENcfeOq9NnTGi2xG5L9bZ4buvJoAu5vgxvAXfTAX0PCU8NGB
Rs72ecybYRR0ikhuQ3AiNXY1tB89GEr8SvVgRURWuRPCeBDqRvQP8pIGLU4tPXKE
JRyFmiTiHMxJluFwF/7QDCmQ8Jzx6JYap8hNZbj611cfa+u74Px30scq2Cu3mdIO
FFCYEUvFioiQ45Xid6d+VqKvS9h9HpGT2Hv/0eIjasiCvRMT8JA17mDcZQsjlVcS
OsfzudnjAcID6fsQq7XUq4fA+M0u8wnL6F4YPJEQ48ynl59XALnx//jia4qHp+n4
Yv2WR5xviaQ9SFnXeYPIlcXL4AEeZsg4Xx/EpY6EhijEewHMNaDh/7sbFjv4MIiI
OSQdY5UFm7PpwFSC413roQAElnaOJSTmJf0cr2MdmWU2gq+7l17RRwI/OZvzAzW6
PP5tsAkkzqeUhwL2QDjQfWvbKU/5ps3BD1OkVQur4DQf7Yc0Lf5saQEOgPYXoDMK
DS6LxakKyiatxU0xlit+b9KcpcAFQZAlv0VJeeWATVt/C8LBoZXX21KrQbU9IQlv
RLPdfB9q7VGyjAxRzOzqmUsunkfiNfm4qaswgdU3XBJqBOHd0j522jgYW1p7fJj5
45qz2MuGFi44zTpFIU2MBLlnzoKNvCZhoVOy7E8wJDjIwogzayNH8omC4CBcKLMt
YorxI3V9BuS7jQSsQaxRgKD4FMzQGi7pkyCS73QeKXKKcqlSEo6FQYvl/wQX338t
bLWnjnXFeFoWoasDPMrB34/6E2YbVaWJAS5vQ2pIgFfYFQ0GLEzN5NtuYFcDuWUY
kbunEzK+El/pjPAveYDlMTxCamsrNoX/TNnIi9hMbcjIxhNiSjnmcJDmR3E1YlCz
8NMbnSL7V7aMi0le4IUWP+hd/KwVa3DTzbxQG+7U0s3EW7SzRvHtl02PKpQXhNH8
GoTUxWaAKzqcv6Uyr2TFltzUob56ts2dz9bm1GymLU+zPh+vY6itS+kXrbVHb57c
g0QR/OXqNJn/u9FIH5mGW4TnGlCi7PEg1RE1O/MLikbGIwe2j0NaC7orc1gBmrAb
d4m5GUxviSKgmiEeDaj5i96RUk7S3qt5Ttflqu+FDCzBhilN0cTHHP4SD40n9O69
IHdqRfnLYdhz7VhtPcyPn9rvYnxm1Df1E2vtzePb5Z7GHpLF6cnJsucKnr6es+qK
b0JD0Fk8UbtwYrE3KGxgmaWhyfAPjg+SkfC+YwVUd8teX51r5PtQPVXcAlg7W9cZ
/wiLpqZOgHRyfYRxdqiTYLtXL/XjG5OasJw7/xtQPVp6+9hmAOSebaf+N5bu2leH
zHcI5FJw3E+l1zoPp/Lsb1Dec63mX0pwvZRachaxRUofoRhpGIyxt56/qcTmqfPZ
EbvT/fGo/WL+6Isc3SGWBeY6Ksoie3nNt48Ho+hN1gZGb1hR4EO8id6YxjcqVMRm
j09YJDIUdXO6lTaHgCPH6QbiUA1vnjjpI2YA8W2s6cl7AcANwJEKcpCuTiZgOeOD
B5HfoIyLEeGgOja+GlX5/YPOlbB8RtFll2taBwKvLLEweRSMM1i9e4dJN+F1+6mk
aVevXHfhwgMcPeDnXp09BaocDpoXhm/kbOfobGrfx6bL3+v0RZz/vmiA7u/he0iq
El7DtgorBIO9DU1Zq6Dih1svQmPoswR2mQvSRPj+9PqeUvqc0oAz3j/rH+X4U/+I
whRDW2SamWKYHOMvgxmmEeHlbMizHTAF1rDxxPRODVd2Ip6N/dsE9P8bfEHIZvUR
6sH1Hm4fkvbRVnmnxlzSlq9eXODFnrZSNBGDSB4k6hfY9v9Iq0y/oRCW0jDocyR4
aB1hA5cbkv+PmZ3Kf/HoyBDagp2l5YTEO3Lv1UNvsrNzooxydRnAk1g1UX3/J2jU
spr+FvjmnODLNk8ql7s6c5I0PCLrU5GeHBgo90uczJv2jaIwraWCl7fUkNwqcL5e
uq8lLeaYCOaxsRiV7aXfz4y+FDmTPZew4EfknmeugTMJxLNp09bw0ADUtM8amA+q
n93c8QVVxprUm0qJz0+tFFzgARXnMRKUBNypvF5Yw/HmB2CLwFd4yiEFEYvFnj2L
3F/3FuanKPf24UgJ9VC0U6boyjkTy+OIccbyOvO7Lnyzw/LTkEAnlUk9YuDq01i0
Yu3qzNt05UCeCECTWA7j8o+2sLQUwKffIUO5pUvpAu3wVYOnq8wC840wAkunbNtt
Yv6UuzRkmk+AtefgHOSTx+8uWoyWMqf/qVImMG8nylOJYHDKNG+OwE8B22XywC0N
cETMq1tcqccc3Zyufhv0dbzI2UjUZEfoMRqyW6DafHMyVum3LSd/9uqKp9lnYW1Z
PDlTCNOEwJRKofChqw+lDDT/8H68G1jYpoSSjp4zfBl80zEsrIZ1dQyGUwLP3ese
EreVMMvG7PnmKD7Tp0mjTPoxRP13RrIqdfYXcL5ojYgKLatFa2gfEwVxKQuuiktQ
zldBtDEUwJ3YTVhwzPnu3ZphVgLOKop9yIh4IiOBtcLbfiz+DSaAfTnjo8cfD0jU
qq2w+GVF6Dsct3MKM9JJfwePtFT5wOd4/5U4/510F+PgdxqkCmBBya0SpxVQDNYR
GVFyaX6+CJ/a6pa2avdKkaFuGOyf1dnsDSnHnvWqRTRdh4DENqNbr2qXhqqtAKT3
xdPKnVNOYpEvmOXtXxKDe4/BbWNxv9I42Z27+1VNBvqA0JNbkC57Fn24eirn5hRo
jr46pF71sdnvCD+IfbfhILIjE0wsm8FuLTxfVW9UiJ3SdWZ0LNvDhofJxfwmN701
ls4fsDuHooZkPxSaSTDswVLbHeASDLftZan6sZEdQKGqJ8BLX0i3inRSrrJORIZR
PuLnTZNy2zB8u5B6FhqdQzw0PVhWDjvIquPyVqstoVP0R4dGPEdn0iXHfzOC6jaD
ZMhssD7J+5qDKDw0F1xi4e/Q2tmbHVTtBFSSb1a7mHPEmYkmyU+B+7WU0FxL9DaX
HOvW5PgACKhvsl5Vyak3NB6lvgw/Jdl96rmjTCA0xvHVyMftqGMZ8n02DX7mdoeV
ccPsxTFr9m0M88Cs3EySvYm5XSryTVEKvMcWv9Qk0tLPm3EWC6MgD4wfpaYxSBzt
2Gjdjw1MlwtTjfjREAH0No8piZl1XJSphoKcN8S9kkopF0VE3MhirbICfjyn/iWt
4xuf+V3pxoao07zW2t/I9RSw4/lrXRlVQAXhquFE3Fb2J9vcZZ1h6ssQe3BpuzDk
AIzbpeT4GmgFCAJSoDqpGRw882e6P+cSx7aZ9QZXfup2ncW9SthwKYbyLusFCLol
rqt7XoKoCZ5F7gzymxN4+rfMmbrgfPBPtTrjehTA58m092y5nP34TlASVZtvO7Sk
uFM7U/sMSMi5GuZRDcSwrxE3esO/F5/gPvEuxJqbgexnO9XZhNMgGRPMPXJyiDMK
tl47wHeRdyvm7ja7ZmHc+gi4KiUhW4S8vzqGCt6385TRz4hWRUEvUCOGn8kSgEQT
SLo8ey2CevrPt83ixlPwLDZ7XZuQ3JVLg29aiytG7Q3SPCzecerxXtnA/W/6KlaX
E4GXRM/lOSt1QeMhJTytCmcg1Tm1gC3IygyJMIpWA9LKvyk4xDlpkLVn2mpo4VVW
FrrWeN9VwkQnalqJ6kyuvoKxkSChpoHI20V2f6fm87pz8J2Q2dNj4aWQ/x5mgpBM
S7/psDxOZTPSCGbMGNtkbViuDh+G2ImV5jPo3jYycr4BzyHZX8DYGXjDEykl+RgN
8T6SvYDM7AoPcL8+NPcYev37vr4Ll2KhUW+aKZSvCSCNrGPjysU8Y+Eh1xaJnlAc
vh61Mzdl9CbS6EjRrPL41/RG4ColWgiqsvylB1+vhaIO/5zk5mczHHsJfXJcQxMo
8Og64VDPDodNP5JUiAIyxd/UHmEl1LXnZPhr4N4POhKbFMm612JFqov7cV9BoFpR
FvVC0AsvWpRQEXjhwu5kJPFHzBRb+Nde6L9Qe+LhxwzJFAk3LjQiwLJzYhYHq2Rs
lUZXZLEsxDVvsMhcU/8stZhEfClMFfTW9YhG7Rpfi5vzr9BPzMoILujt9RzeJPCq
P4U5sr1HdE4RTglFsHyvZxk+0lqlblVTpq/gnZwcsyTDSgPIH7TPZLmFIv3Wvcbl
9De9QmlKtX19S4dnxlhLngYn/xMwVTogYtj4Ji6f8GntRlrR8k9MhcEepGvKOxR7
umL+VLY+mJCbQj93NpfhAZjje7cUUNsbjsgvaaqmJ6Zx5XPInU4GEi//9awLVzEw
WAQ+yTKytMT7pBp+IFVZm+g0MzP1Ik6/MI7Vr3Kn77SyndwwD/yy7aPzzaWBYGIq
YNwDExQJu4n8LC/FCtdTsrY2FBHzqpY3Igxx29dUNVh5fzZBPfKcamX8nKPulrpd
vsRW6uwaWLfv/RVwxFCUWxWbc5FyeKswYyNhrNrOj/6FsOE9gUes+C3/mKBa8Y/n
jWWR9p2r75bzmMwrHnvTL+qNUE4ShD7OxEp61kTSgGuKOCH8ky1G+AgNRJ+wERIL
WqPIB2G5Nt17EcD4dJDm+Sk3zZnYYtwR5OBpPrRLzT0uCsa0LM2GT3qnFqrjtldF
fsSbONz2qEEIyCh0QoP29v7vy2i2pjjlZXs+TL1HkoR0B0drJ8IzjZOaF2gDzxDW
+pkghhEIPQLiXRxiphFiGj0BSczfeV3qn4/n2eKf7pb5iXyphsulNKm6CF8RQq+i
6kVNp3J9aYjMScNwPh+8uaO6kkdlKq1r3qk9j7Lkt6GEU7h6Bd8AEoT7LquMRZqJ
m4NL/U3g7CDD5hg+D2w5KHpLae6wZ+wDVQoB946ClJJmcX/Ayavqxb0DfGxUgGYi
ilD8P6Vzc4j6K/2AKBHY3CD0vrQv+FIVAfNDRSDzx+/3SGEjObrt0VanTPQu6Qrt
By18FHU3QzBvjYRIp/5qrl55SEz2R5BAjPHRxILDVODgNKoiMzTLPXSsZjXPS5Te
X+Wx3NIiqhGjT4JZkIYJSYiwtwKbCNObhfVBqIqEEuOMx0JRblIj56quFmZH5bN2
5egh/97S0tZPFYjk4aHGmrFHi385N0X8G6TrIGjb6Bi1gA9LE775xYzPeCnYuBJu
Y0X+aZbGx7WFk7zymCUFpwi9ID1iRdpmv8OdxFE8n6dIg+Ue9XFV6C4ZgsdAxNwX
URKWp8v9fNxyNsrk/jigu3Fnx2htxIUtJRo6yCeOEjcP4l/DU7DNfz2FSuI6D2GS
MnYMcWB4w0OI9ePG5bT+fGho11AL4S23FRo3qHRVjnHBVoflbo/pzJsfG1+mXINq
hVCFqLiD78dUnbELAJC/wJKAtIqstmR+uK9GItTKNe+o9e7Cia7OKrSCHtCIxxU0
Z6eguFRsrEKhfBcpXluekXLPiy6Yrb1VAY9oK9BGZSor8yXgcqxAhg2aNGEgAXEI
uKjjV5JBJYwNutkJ4KrSQhEGoRDgzNiJV+Ne9aTjWG1UOBoUFNJN+ZeeY4neFvQP
eQLfQkV1oG2AEVDSYHgoto7LxnfPb33o/yLmYFJx+MaEAgk861fjLydbqQimmsgu
z8Sig4UIkKlYmeM8foOxS1LOp7kxtHq0/ldprips83cFg6P/y2RvZeGZGTN+X+bz
gKzxbg/KO0PQSn8wFwRW8eZWugsBXnNXuOlW9hGIyLXT8n7ZOjw8TGFpssrzNDZt
AtHW08bTcqLOadtBc97r9ZqDTDk1LgZPFdTjWIoEfN2TeUimgfZ8m1QK30eAMZsK
v1RZO9YLXRO8VJ/YHJN79gkTK/03berzDFM98BQqaMLSZi14rjVgmHLWzlh1zJnb
/OP1v1aICxI9SNCu2UQg2dRPnl1ISmxtdj95fiof3nNtMnSzFKKdGr+42SDastJE
UZUolxidFU1wDmBZIffNWj4hinza07qab5QanMzzwZPT/Bmd3Kig1BNyV30Gjtyu
z1sMBmqvvKYzeToMP956Q1AGVfk1asXzrErKoX2HzvqCdDu2eVkMIz6ICDjNov8b
wGFxoIBMrqET+dCnDmdF92poSBLkJECTjbCVChZi8kBO0rb+Vbc4HlQC7Ug1uRh/
c0Muv3KewD9s/4Mvynd1uH+/wHlvIBlu1JKGNzGHQaK4rGHOXvqwlo4vJwdRNpir
L5P3yaGrCys71XdxbXKBebyQDoVwVsV2JUQikTMzrblI/fQykrn56ZdAmRgMk0dT
xpwuF/+t6wv3Hv3jG+7PhO+tob+rCDkYIedkD8ruOh97r7kE1kLXiUiMKJYxpHNs
OnkWoAgtrbbAQaimLo5Z1d7wu1GKClkvfOXHu035reH7LRdPTjO3b4PEP5rt1I8v
L2hm64B2yeocyQRoY8IL74C0u33yCAGsdsTqQ5b/XoXTOKT+A1HOkHrYOHZWFrr7
sLu8/VQ0kFCxDm1xFjeo3rnmJZFQXXAbZ4s4rbB2m3bHxnf8Uj65itVSQrsosNTx
vaVJQEVGFR7BTHuCyPDeK03SZaGeKoF0oCKcDOUHT/6fD04bi+59LisLOdtVhZno
KThS9L9XriyAurbdcOkSDLYrysnUqWDbMkx918xfiU1oCb7ehDfwbB/tkEsp2ud/
wHzaV+wchh8zYUEcv1pcia/6CooQtnrc5BNP7HoQl7WRSK4y6H4ewH0eVfSCUp8c
Jaf8cNSd4zSD/MgZVf7iYwouIaweIdyyUKo3wSZvx8GS6Truwo63DqGTmlagBc8G
l+MonHfukvsf12UvsCcHTNAITylJWa2FKe+CYGm+23qNpGxrpTBSzv1L6TdOo3v2
HLmQSd7ZMzb2ZgS8z+ZzrBFbPwp9NwL3Nw3X/wTJAutCjw4A3oughVsOqH+cN8Sg
X0Kx2nPt/ef8zim04OEjrP0T8Eromp4uREYYcPZs5gFafQHsVESjBI1uBjSQ2k4O
A3ko8xmFqAIU2y+kMbZfNR03DhIH/k88TUcHNWoHKYwYJKVl/02j0Q1cN17ULtNF
rzAv+HMEeB+lXU5zwgR72SGz+o8TgB/OQ5LZqlokspxzhGO59FwpmzQ3ytSn8Dm4
yZD7McLzM6WMCmXIY3QN9CyscLdvA/VAsxbX6rR0Qq9kl6905ff0BxJcdvqVMs+Q
nfDYpik8QRWdFLLzd8Oz8szcoDDbuNiWj0yUjj9JT2QZiqQ6AzUVqw8kRfd4bWD/
CcmKvqQLJE68Cd69G4PHk99azAia0i9JlzGTm5LdZtEdHdYYzxgnI+EueWBHznqw
rlZJicJDGYIF3rSt7jPkCjbtn/EAydzG0rMhEVnuMiXrOCKJQHWJ7b5UqICdM/+e
vk+HMNGULrgwG+n+/KvxwZJVm+csvlIN20mOri3lMtVELyl/I6Ns1410sZ2C+/w4
nxakt/CdFs+LEDCSWPxom7297zI2DTpPn0DL46tnGYTt1dPpm8vI7ygHCJKAWhgN
hFMt8yCHS13+hrpZckW9bVKa7m48MdMbOxAyJM1k/1+KBoRKVpm8iJ+yh4vNR6yW
Qwdwl7hRdqmXmZY2Rqt2zp7kIG49oALJIV7WWaEg1ZN1O6V9O6vBApig3j3xBLE+
EpL1DyvF7CvT/hzWIGEsTPY0m49GHxF2scI/pp/NySDtZbrTct4x0ciBkpGwN3ZD
WQsRIORr7JRQvYkZkEnKGP35MeiFEhoVOocJRwjHibj8E5ghPyKYxs9YF8ooE0nu
MN6yFddeanTUp3jd2DZqz3gLT/lfDyRXcLg77SwntEmuPX2wTf9RqJFqIZVTKmLz
GOaK05ncmcOsHssdsY9O7wUqWKHnz7LFa1U1NqD+hbfFdpWf5R1aWkqHTMuZEL2C
yV6yqdFmtxV6PqLbChusf6q9U31PGFqgcyISPmuipMA+mu8zXBIANS5bbGK91FcQ
DwsplfveVIGuNQMr/W5SY/YQM9Nv+4+haEe5O6UP2z+afqXdsmfcySmM2hWu9lgP
iVXi3WKf/OSDaFP6Ly3WkYAnLCH6DOE78f3Cy6elhUklDLr5ogvIy2Ug7jTuvEoq
YnUBSHJy5f0Hvqq4R/Y6rm7/uB7kjFRrulrKGLR0XeesYlsZAHGvCL+oHBXBx7Wk
pBXHQNt1Y16MQkapAEmMI1PtBr07g8T3L+uxhJ7eDClU/hS4KfM2co8LuUHuClIt
yLnwWF4aOBseb9lIYpvHWnAj6Rrw0PEDmrn/tq6OzFgoLc8sL+BClU+w4pFo0JlM
4aIzjHWpv0bqKuef3nVANWFmCn5qQdyLNOz1pcHJzLPMTDoKYQ9ElVkH3bDVTX6B
4hGb0Hm7hTvMrhXGlV85IU7phW2FtDDD/d6zUkhpA6F7Sb48RIFJLgmQKQviiTpS
7Ye2aWzncEcrqrUOTYWA9fqtWl9Y9kUYJO+SF7IOsVXmGvYj2lg0MD3VQd46L+uV
x8qcCf/kSLM1r6p36jttD58M1ManpF4cZJbu4kr4Kw/CkDLrK5bBz3yYaY/nwk7A
vLVlIRg25n8rBxB062+jZ5THK5ryrIPKey2Su+APRKwjvxZ/tmqrCHTzax1Z2DVx
GTD8xUy1CVYKE2DUobBxj84NZPi3zHUawVrq7Oe44mtti5p8Q4h0UNXJGlakudLD
wNVf6eohY3fjvwv4hsFNhOXBu4SnTgXXBy9sa+S/xRNTWjqdpWQPdRatNkRBn4Ap
vs8fYMbTZ7rpUZtvSqQ7ocVbw0fRSgIzn4Dxs+bYRkqm2VkVYDO9+Yrfpda0iqdl
Ej28PjRyu1a9DPQwEYN4yy1tj59effMjp3hc7qKrU3wyNoUhcV9YWW/xfYu6kEHk
VLxfY/a6+GH8bjufi2ltSOODtnHmaECo87+x2OK2q72yJc2LD9yJPValxJ1axmCJ
uARIe2IhxxjsT35mN/8UxljnWyC1X4Lwu4GXVJ91/yoNTbG5ouozSL4WZ2LKhcZL
wr9FGwri5wNHBqIa3RADrn0t0kttXQPfrUjonv8JsGK1dGt42cYCNiNd8ztdq3hW
FpxkBjbX0Iv7r2foc9w14vp+YhR35Fe6wGv7co3oocKjYo2YDj1ZarETYyT0uar6
kOa/c+G6XjdNENEn0Z8OAhbkRHaR06JFi/L6ZuZzpDuc74R285rc8Ckj4qkKdZol
KncVGIZYFjAJD4acfg8pUjOIQiZq+PmUBDyRV+TnjenOU7Wlgh1mipjX0sAaC7Nd
t2TeFmF6E/FhtrOE1GcCPaZVt3JET4FH09HU9B+33xQHCC1gdvv71w+CHmmGuTZa
XXkt9g84yZE6MlUUbux5gAonkiiItKY1JaAkRqGIx9QCCB/zWT0kl32Y7XJ5jQRm
jRqlhosLA7YGpvvQpO2qbv5nkQT5tMXPcJ/GmolOjUZg8pod6HNJttPV6aJzZ8Eg
VdAeJ3S9tOqjX6pLbkI6CChUc1onwlrjj1OhdbKe5N8cr2OjeuYdX7tJX6MQmRc5
JU+vbwadG/W/o/UVVRUcvwNk2SXQzPgyH0sLjs6FFmSzxq/g7zhIW/me6NmQiJhq
GuG8OwBB/gyePkMt0itqm92ReJzpgruuzcPO3EFPZ8QHI10f9tneWyWPVMsD9MRw
Sg/8yKEWXdB97HRep/TNMhCN/1daq4WlXHGkT9YfjqeCknxEqtfKXoAnJTgZSlfg
B3Ymrx8txCpeokgBEFsbQvLU+ZPtWkvsSNNRC6QFS3BxHIGsFIZ4k/gkqdBoDcPT
WGzYLhtaIxzplLLcxwqLTOjUH7IUn6V0CM2YCGxGkubv2iRGFSev5FvyGsGPmM2q
G2GblbOXa223k9cPWRQ/GMV81STC+5OIXxk68/YvrhPjB2OeYNGlmQMJjIIESapR
es71WYPwS+ob1F3pV+37bg/jiQNQfTQ7uHe4Y9UwMSFRRx/R1mNosZ8/ICadGcW+
YxGzeyPJcfgorRBLq4pPylSZSeD0j33r0J/8uLXb5czH769j4oexpAvO1wp5SQr+
s64StaQkxjlLsydQrpMg9i2/JHHPiSz5N6UInMod3EsuPMSfqm1OpAsBzLsv8rzm
ntvREtpiMZy0Kkh3PXncgRDf0CfwSN4oH8VahBIcG9afKz98KZz3CyxSHwKv0rqb
cbT8Hi6OWa67H1zOC38zbHvAVwm7EKRh4fRx0zNjTRrkaGBJBUr5BGqfBMPN7/h5
BfxXZj1wn3zOoBTO4cxAYhthbTnutbFhzDMKMdI34fq7v+UXqolMj8ZnrIY6yc3J
VK4/wNGstPscX550sJa1wRuMJXo/Zg2I4wI6T+Iq2gpIRH13NVAa8lgUfyE6Psq8
8hfrFMs4kN6uZrh2C5t3hSpLkvtI2/v2Js+jzwMCOKnxWZoXT1rkpKkI8Me0qxlO
k4XEIHnrP+NX1PXtKvfGtwd3pUhMqdHr+9ih3rXsA94F2FuUzPWFwWz0jEkjGnSQ
99XlbO/8sj121+mptLq4CPXFUt9yuqpR30ymaVqPeeuXvQqRxbyQksj233td6otE
Qxq0+Dc8ngwNZ2kGG9g63Y111ybn0VFqNMYSeHHtB1bApJEINJX362DJECyFVxW6
JLvLr0r0te93TcSGgbBLJrBZdc37sWM93x9niAqqHgBZXqSdPgfnoCnW9aP2pS6H
q/eGHhx+ZTqQXWo8WXufxKTLVDnhXYxHwyzrwroUVg0rzd/zyOGPKH8iT2PUz6Nn
/YoyqJ8B0eW/YAsVCyYbcIjnevO3TS6VRRwtW74JAtCwswx8W6IZ3n/KX3OFqseC
1+WIKPuRZJtCfRzBx2WSCdT/qAyLKDAvwY0s2lnENUP89KWY06RwuPR5cJiInoBb
fHVNADHvZ+/wbDB01b9sG/XbYanIn7Gr9Vds39FDwjj0hfh+8XByStA9KNpV2Leb
h0tR6ZIjxod30oWKx6A0YJ+fgvsB9ve8rjMi09+8JSDkGwIyePUC3nv9k5uZdTOw
2BKuwmN8YV8x1jd/lW0I5o/bktAx6rPUzXyROMvBfiAd39BOk59MV2CTr+Kn+eiI
Vtj+3omNHd3GSMNgiBTVLKdggsiab95Z4RVWpBRGpjUFAaLdcZjsTf4eYedsTrKS
8Y59oV2z4ijLeKlo6l8t91aMyZfVzohGnOopvgmjT0ST9x2RgtwezuQyqYPPMdwD
Ok7wEuQx1K/NrsUa/wtSQ51J+s1R1zPLaIyQRr9OShMBE8HbhwAoxSM4OIhvSl0j
BIF/wRgwWHs5SUxLwZl5bmfsLXvolimPdxwnd3DnzmwROmXOvsQv37AXyaz6c4Ii
FFBwlOGIVgd8maZ4ySTTStuGNDA8CRwzD4nAUfGnrba7jJK4qhacq5VecBQ+V5IC
yGQiTpxCdRHbPi4NTweRRwGt9o4B75ycymcTPr19xteyaLeXxG0b/Kt7E/GzNKG+
uXnZ2+kZ6r/b3Z+Qx391OLXWfTehqvGncaR1Yu6vW/L0tGl2mLUBAD8Nbkn51tmJ
G3mQ/gs/lIqCFGdTvzlSj6oxBf7YSYi9CdsHqyYpbwrdA8KJyHXmoRAXxIbDS0PC
Fbk6fio+P9JdWXySaf7dqVnk6f/pkuaa7rwcfynYhHwHFof3OQtknVflRwXmOOCZ
YUIJOC1ekTpCQ2Ztw8QiTvFyUJYkjoynhFOdJkTIKnqNEdZHFuq1qfwswgymbMUV
iotxoh1JioBF/1hderP9Fvo8NCkiNKm5Y4+E5qi3bGP2tWuRY3dga3g9CdQXE402
IJo9ymhjbQsig+pGgueUWqRtJruT4F32rrL2m/TO/QuA0p4oFIMZ324Qxdk1iFUp
seWTFm2TSI+eT2qbFHUuyBJYe9QwY+fNr0nsw/Y6QPMMo8Ghziny52YGU1qh/grt
Q+D+1Dk901GST7Q5pNR2Xt+XKMDWQOAI7ENEv+nHSJnvuOCGaCX0MW5VaeMJ0bzF
zZuBeupHlvMBydSXgCA8bOAL9TFAfjaVGskr8wcdZA3rlX+eIrUoOiILZ3g8XPVn
VXgDo82WMsUBYMVa/t4ibaGupA2MZ1o2KXMTMVk55ndxHkEpH8IBXZpIjY6JoavT
I0fnxzPMLFv+URUwYw6tgx8Fso3YanLZVYVzE+N0OhyNnU1mFnynXALHkVJFmsGF
FIQvH95KSOxAP5XURyIRvX8xjqA3MPhxW2cy3N1Y+POC/t+9prVjHD3kWAg25wgs
0L6L7vOo7W0vLI8PNSU808aSYOb21oazR3P7nREjGP68JevNRyW8h4telLs24ZSk
wkZmzGv3OtnxDBsVGLarXF+0J+uyx1JXvkeHMc+jt1MRvoj/e+a1C4zHCPE/8On5
0A+MKhHYR5fhWM6Q6/0nhPCE1zMEUO36CgfoDOO7ikoMc3GZQImn8Vntk+P+qI2k
6PV+M3UpaYFuwOCS7Qzsce+zB4RZiYvs1OIMCd3/D2hE+22vMy/h2zY9H35WyUpC
PRlf22fi11uYGKULUp1jKBjKilwQORn0BwCZwk3amgudKjQm046I3pFMZrHhJQAJ
ltnQa6joE+1RPVAnjN7HUkKcF3/ZtGFZdWE167bhLiMTNaRu52+eGcWWW8ocJ8zx
qJr48dQbkhpOL1bZb27rMdU4GnAIhWAfECrh5LTgiaVNHwC6kSu2LY2u99khiCay
HDNCQWTRLgHWAJXSUDZ5ZksFtlFHSIllUHZBo+5Aj+61lSwx219spkN9I9HxbQV+
BwU68jhorfIdO9IQnWIIAcXlO1gHg6Nhz+M5p+wtv9JQaarZroPqzkDae1cGAxJC
3ev4Us0fzqk0txPzo8Qxyk8pTW4cy9hjtZy+o+/FLGXmHRhimRTqSqCovf2Dxakn
XAIKHnMyCLl0WKhnEwqJvqbHaIu81xuq84nE7Hj4Oha9luBkudFsCLXj1Nk2mSeE
5a7Dm3drPkykrClru4GE6bt7FoKgfZHTYDLQpSggLKhVoZGuAPVIUVym9KgJt1qR
ANnGqlggJwbkXyiTHhWdaTQq0StowVlhGvYXCuXaDtIthL9Eka8Kfubla9nnH5PM
jJbqpK8egDlcRn2IeFjRsC2zddWrAi4o/ZS9SKHJpQlUf6RfyMDT6RhDXyxlEIU3
4tmS9T0qfKHwvaQBxQyMEGctYiSkzQDF4IwVfP52rm6Njo9SH6OTl5sP2qFKp64j
4DMxM6V4FvMF64GhO0Gicx/06c8YXQJVxb9zm8sJXoX9hyGYStWMk3CJ4ZgyjXrk
jD6gyHUvWVhrTDComSqPlOq9A3UIhiiUq7ty6oSezosltD4jbX7esxM6aEUk9Czv
mBIg0b23CDYqcpQIIph7hz4REeLXyDqxshX0rKFlxYGOuKEZ++cCzCB3pcwDPLJa
n6nnya6rdEf+H9ti96TGbwZ3cJhlgMqphl9fO84FaqTN0NVA85ZzLFF1gDCN8i/l
PSLQkeOZBSCazj3lYDkztIzAQz1k9hAO0U14RqggvCCgQ8CXppzqvQU/MtAcFD2D
NVUn5/qlSnoQ8kY49DzoZZmjs2BCdmJ0KDRhp68/qBhQWfyENknojO8TkeNYe7XJ
gTytWWtLox8lS5wOealhhppTRvOpsfCZmQ1LkSNH+hWyE8OEGrx6whKAZ/BQMAno
I9arKcmebW1YrWe5MryKXVj3DYqvGFD8YNCPBjOv27fmMMgmaH0+bB9qYHg5+j9o
jEh/SfG8drc5Q42w4XWLwIsmNZKxb/oCCLkoQM21v37mWLAtZP0ZcXtUAZLHrjUr
oafr7AukZZM1H4POY3WBNhGt6ReZfPrw2qhr7up9nBzC9eTt8yUzKjo5zjKotIgO
4IaEQyecncqGhHP2yXT03n6snA9Cz7CkLo10q95ifqJNINcz0m6GqarizfPVgxIR
zyOk/Zh79E4B3jIvRSn3b1eaoC10gP0meBww18r19t2HtPNZaItNTib90Oc/mQTw
WPqh/rLxDWVZo8UB97rRH2/jzH6ABGqCobuut7xU6LStGfRnHLLenXtca6zsh34g
/scgRM5B2+QjPvuEI+fW5qokKOHw0CTADqDk0TvpvpJ0fw/Bh0ZHckHo9HfaVbeH
y/YeNoIa8MlUDPzbxZTxa+vjPCUh1ZbiFQ6BJHhxIw4X7tHlS2V8h8JesiXcrDOo
LsXoep9SCDgEtyeT6X9/gUZugpdydZuRg1fLnRtdOvN0Y9n80hvPI/yzI7BtqCvM
vUQRnm6L0lzF2kw/FAtTlsyYHS5DhsvmPiOUK9luDwhPZj5iNZxqohg+n4gQKMu/
vOjH+4XXyNYF24pf6F7xSjCJsgah7iUMKIaLz7oFoFgdnWlwxVXpSJMpcXGDBuIT
PcbhaFY5nDkzdP3I+Z54Wm4zWBRbMtIhD/1Qlo6J/WExSKu5AbP/BK0KH7M/GQjH
WovwIn87VXDebLOArB04L7GObb+RZjKlMMRHRcJ4hq14/gpUAn1uCUK+pbs6mnRB
WyjDdH6pbQdhgJ5pnDAIp8zbr9cqCq+Q4jVdRkQYwFxNptXbhaxScnmpk9UhbBZA
gTpTXZ4/qCf6bf5UcJq7+fYAU3UjaRxsI8vSE6UcrWQyjND4F6trFGzwyQxwJbX0
sBNGRpNG8jaxrsqi/WoOFpHMm3LIfjSvWlFPE3IbMgOl5DCE8Y7OTSUWC223YRpw
tx6LAk+QS6wwbjTznOjcC7xJ6BkldbPdkOVQjPBlq4JXZNcyaWXe+/7zmDTL4eHG
XxYRa0DNpcYt1jFOlHYQ349zQvJcdazFIzXlZnj/jdFupM6uKzgDnatQZdKArlgd
D73mcvVeHpRyQOmWhiSta+XRpsOO0Q1n4vebs8TdQzyqLi7D9dQMW9RWhrhX4ncT
KZULoYpidg59Y4qsgly0Vn1gd0WGCcjtUuuhmjyUZ9aESlHzs3pjz+Dpl6jWUVR6
XvwOUcSZuJZd0aiqrYpHZJ1KlQewaiE52kXKP2dkE4DAZiKwF0azeKqLjRsRCz9K
f1zjjxL5zvoLSA5AB9zEXDZa6oycXTazrvpyQwcCzsYlTjRd0oxlG7gDRxyPVoxR
6UbbAE6ApFws0UjmhcYuhO4iXrK7JpwC0E4vyGfD9rTEOYjZT93PU1KFI7mraIg7
tkplX8vU948Nz/hSqXPzcxIFkKKQfgnuCZ1g9mJHo9NCKWyvKRJwg7ivkTIRolQd
zkbpVQciH02gqES4Tb05Fy9plnAAn9xNZdf0RsLj6i7ciKqe4KViOKQBB+7kvdo8
e1QjHksOe4IofOaHwcyFG/xKKP4fz40o8sn5UNvBdsV+417R2c0N04L+y0v18kBD
Fx64qNErjVfeBlm3RVm+spFt+fVNkDVRU/hepTzsnDOvgH/VzqiYcn5hRqnLCpTw
G9b246bhwhbYyxd2iK/+c80mwHC87/hr7ip2RNyIxKyDHdynWK0H67OBa6ZE3PfF
skHtK3//nWbib640xgKF8qXN01ViZqtjwKSyu/nXR1Okfbj0yWvOgr3zPG1yt9dW
5XuPmFJ3BGUHpwI30+tuzzxaB7l/Vu+NbxJqi2wLZX4komvho5QUnrfGUkgu2Cut
yT8whTTOUcrFI6Z4OlqfazixMl6vg0stKTGc1gBl8fGZxCDrlKg2q7yucn/Iujty
Qsm5QpdPVYGlav2LWOwlVWWYK90hJ6+n+jsNCPyuvrzB3ri3euXTLO8IuBncLYeF
UCaZ9HOJy9qjR7CkWabnN035ihd3OFUqT0FTdYhZQVOKjzCdmP/AytVSwzgxnw4c
d2E1F+TNKCWABnGq5BqxagPDBq/4hmTB7Yoy4wYcPC7UErdV7rPeZpGcaH5WrtQW
R+zqZK8NBwgyKAlRVcrS+ZNVScn1MdlnYU2tAOha4wcbglooQ3ewJoPXYypaxJDO
8/URRDVZaKqQIeqhbr6fQBE+Ofyeu8LZEC6NDbUlho3wIfY6xsDBMs3Nm+NW9YwF
FEEpLpYoce4xd/XScCXaNPpAqe6U7u3w44YuVvIcoBqv6SwSz3d0hLPMfPxopcZ5
mv067Ytf/OPGtntySpRSoSbu12ElsMTXKLJLg27I80HgluCy8UKqPiFNfRxrqLCT
fbu/5rSZ21Wl21SINkpMyjsfZvR2+XCOtUFzt1o9nkJNpiVBturRTAMfZ86sIsOc
s9iftvoSTlOfORqPw4XX3Xus7eaOs5j4hNlcDZfom9rUXn5lqEijEpWNU252jMBE
hFjkmGPj2436umYRpNZOE5gZ6HgP2AHv9oz5h3M984+rr2EfQ/L4WE9+5ESZUSfo
qeHJWgxkqqE402ywfXPni82ROmXy8v/QOeMMYP3B71V/PkEe/OwJQcQqT8iGxOTr
fhDKyZ3gF4zRZ38sK9lwBJUtI2DFmcrq0xlq0uSGM2V7IpK1THKH7cBy1VKtJHV3
bgX+TBmkyMgss5y9u363Mmg/vA74cwyZlefZFhe45oPTaxRdSvV21tyBff67pOOJ
mT9SpYm4jMd6S3GpToBSOBKYCFDV2DBxfgIhhGVGA3EkTymnZ1Zx1sS1JxV04Vd5
7BW+jFUoAdEsWJ6GTVToaTaf6F0cpl1GvFGbMJ5B7prVbuy3T59O/3mtxPvTb6O8
vcY2xkjx7QnxHHPgNggtkC247IvmaJ6ERXqw+9NKfANkwcUvx/M66kurKi+hCCZI
JJnpNCPFngZbadh8hGZyAmEL5g8m2WTxzMvCnAPBF5Z51atadxmuRGenKE2nJbOP
NSuuvqcfz/pU+KfDjnZzN+X5TpCku3U3VNIH+mgmo4byFr6Ej0Z4+bBlXtbrUnaS
XwSBE5fEdwQQPibmfq2YKOUU4JF66QQqNsciBL5ACs8Lmu3iqBSqqFQa4v701Fr7
5wpCGimogLnIC/lt4Z/IytTlWOpMPPwZPPrmH9uruVNqhVhAXaLcJdBoqGSG1J9m
hA4RmTgJJtd27NsZ0BBmR99+6dY6en1pIh8JX/4kXuWfosp99NrGRfb6tU9Nt6bF
LaoUITkBX9wH6ozViqfihRb/Yg/u3zUf0XKVtET/8kQdd0WcfKWGDgvRduCBphlR
/8P72iGhY0lCx3ENh6FbEiUiIDY+Zd1vP3ohq+v9e47i916i6mXlyRMguxgwo3x9
Ij0x0yN+HGOvvp02kE6+vvyjxJvV9KFNzmymlZE8iSmSCcMRKKAId1ebtKVN2Vde
ZO0EOxdgHd+E696ZmlT0Lq+3lwBjqJkriX7iFUIVyVPNYhNiQG0eUd0PhtbHx+jJ
VrJBPBv8f+lywZOnioejet9Y5cKUkD4IJgRF/xYZzseYdON57WslTpRUPjo28DIl
qviCg75c4WYVoxkShEH01SuYI1otRyw1482t0DX6mnFHAWf43VPOQUj6bi1tRnyy
FK4a9VGJ2I8+ulvbqAUCa+d5xFuoLA0+4UN8OblzculMkIKmPn2sjibvmvEBVdq4
PRGD+PZqkbMFKOsvJi4E9qOmmPtW/iQhJdDsesG+MFuSUO3/cJg3fnbRG1seippO
sz1QDNTY19CErnsPw5owZ6fN99+rUpIwHQ5lJtpm2/ksz/YOnwNKbh4vJe9X6DMV
UxRg0wX1wf/MWj8ypXpFi1pkGtSOyWemXZLEaSut+Zoo3LI0n6nOc7ecGB3Y82hH
8BH3WZEj1iJzA1eyqLWB8rUl1r65Wd8Q2Xznl67iNSfWODKexyf9BXzjFpdC+UiF
XwLnCjmfkrXHRERbTxCXUrI8K68WIQ1axmZhIDuVlxtIYrnj0933c1AFPTKN9ETw
bObYRus9FPH8dY8Q50GqrPywA7A8iWpPx2RIyy4X9pPKq+N/MqbuTFooAeYPK9t9
9IRBP13eJosNj29QNfSji32KJwGkgAv0MXgPylNJZfBvSHMEhBalPMF1VQiY288o
w1Rzfzqt0/TT9jT9p6FAxtsnL+OsO6+3zbugkaTjjQESFs9vXFnMzZJ3frv29T6g
D0pSwyehi0b3l4iqv4rb7L9lVTqpsOsRiLwD6IrYUngqFo7oee+51eWa2bCZ2E75
tjqmi3YASMDCazfCoWGmsZHovpor+Z/ZMPyxBBrvBM1JtLUKi4sMOxD1d0TaRR6b
8MIVBIjb6wYY5oI9QuGctyy3spsycMvBHJxFSKfE4/MOf+c1bcxp2b4qUtXIyXFB
AdoG9lPCtgZht3Bgfm4fiyuKV4MANbMuhGarEvQRb7+p6HMZywDE6eCNgYj7XikV
DaJFtwB7GruG25zi0xNl4JmFhOjCbzdC9Si43rpubEdLgJfWLZzn9ywtqxLvpZvl
KJ4bzF6EPjQNZs4A9o1pYwT6s1cM1lH7I7KYDbVnZq7IEkZhH7SlVKrVjq9oVPv9
Ux8SI9SqolLXmLWjW3qVZnXnnOK3SmzF951H4hj1R74V79+KHCSuogMlPFhKeORP
FOLiIHe4P3guB6CkMnsUZLcEF/ERdFD5HDtyC50meVwzt5VyK2DtWCB8FIDnHvs6
TNSegi48vkUuPVjZ6noG8kXkbMkxnjPxv5tBO0FxmZJ9SQG5/0Oxon94Dz4wWG6B
PpGrbe5e3wc+9gVKac14zvfb9gpE0UAq+tCObmftiINzrL9xom3NEYHT0PbYenzY
fVhAjOoYlWOX/kYeqYH0HZEMnwEAiQVFx7/MHj5f/ybuU9xJEvkckpdOtF3hNlo+
3+FvLDOuKDYL/fG05KA8xr9WLp7Tu8BKQesDCAU/iQpv1OLI1kfgva+TPDHKlwFz
fMv1FErI2goGek+zJ6vnU8JkZb7JTJizu6o9urL/mwShKI7ycWsc1Unu7eGuswoS
sGuHhgOBuEvbYD5e5xhrr7WbpMrOUPnK6pZ89uGfrQSlRBNgB25ltdcXn7XLE8ye
cqQnVhman6uR9qNlcOadwHTHuIjfMBh6Rf2Xz+Ad9utaMrUv0HnZ6n4wGLjoKGjw
ihncdtS4AvfLZV10EAwtucTpsY7BUa0atv3Hfp91+UVfK+h063+fbL1oXdNwyQIl
hGOaeKMbviJQsE99yTThEP9CJJ9s2969mu/Zg9N1SSuxefKGvnlpxTEdv6o3uZVE
+80v7U614M1CLfK1yUnpD+nYVxyWfqQqgPm6E0Tdie1621unTgoavuI/kfWoZoZj
m+Jm2ezOSZ8vcqlR9Aa0qzMK/x6xjmTUv3dh5nq40CPpSbABx3ADnAKA2H7ErBup
qfyUB604M2JyReRFglDcvRvxVthYzCb46LzcJOLHQE1DPv6z43YLouYLCYQZFyjM
dhVWrJp8uCbHbJW8V2kqypYx+jo7Bx7Zz3ljADh7ZByrbBGBF4ZCzdxu4gdEs+rI
n2jeDBTUN8MWOV7mpWXht3CY4C5k+506Kniq8RkfQ1PIXViNO6MIIC75e4Y+dVtO
aONIfosoF07WSmpucUqNyQl/QEfrShpBdnL9lVQajf7KNlYvn5dFrr4VkfZ5bUL5
95XWABWWQ5Mshp7vucZEUFSjLBeDlLb0lwiweEpzyvIBi51txORAkrMSDgtPg0Tj
49lJKy0sYbII36vCT2OnElpTX98X1x9KMFPSiWcd53HVb8/33VoVncOqnmNMrQqq
FAfzASMMLdCMGP6nC7HJCTrtwGk0klGHRTcBg0EQ6xEZGVOOxs6GVK+SrGbeLqvX
2u3PGSsvsGC75lE5LGVSVbxBOyMdIE44Yd+NgaxXIvdOVztlItirEBEoOLyWabS6
Y+43HUCabH+IjVKmGOa0MMAlTMYy7DLAC56g5MlBCRxdE78l33Qo2wSYPncENoL3
Th3K4rLboK25nf7EkMyPBaaJ7VUXygl+5VeZF6/Rxwg2X0dmaYkLnLiHEpKYeHyt
B4G/i4K0GG6Mk11fDDzGTgSUO01wJDImsXm8NIcoMiP4zEmY38Bob0UEIAPjKcMr
/bwFb8LY1gtuBbrcC34zkWfhNxYgQ/0oI2l7rmQhCXNsj/aKmHxq/YvL8wSX1n0i
W1GxbiF0JwCghU0FEnzkpDtcDOphqVaNhx7K9IV4XPIXpHXSjup0frSd0JjP8VnI
BWj9dIKatfqEmp74fnIaMijWHGcZDHpHgPuuioQI5k1TfclmBScAiv00cbPK67z1
cjBAfIPoVDypel8TMEyrE66TggSRfrheVEGBxV+tXHMYKAwiAE+D7Ow+8OGfJE5W
lTLyRUdWDGeV9eMFPc1+k/IekSEZT3RJqGktjyaPu+sRTC23bw8aMREJyM707pt3
3F5KusQOA/PAVUK4xkNaBmbV2YDjjgxLkN0De+tW8Iuj1q4Qd7oFmmFpHshSriIi
j1NcJDEIOlb/bAh35HnYq1W/sHjyM6hSepZJMrW8o/gzmGudDC9f5lsh9QgrYTn2
FsewQ4tMZDs8TJwVAQrXq3UofJPdTZh+OYrfkqbUZHBmpbs9wTMzzqBAqD/ZC0N3
tB23gsMtVTvANO4ablmBSy/JTNpCBZEgQYWbB50LjaRKFAmo+l0zGJG/3L9CjUmW
MNGHVwbyz4T6mrvD4kzvu7ah0jbZCz780SVAsRKugIiZmOUTa7FaElNhss/xnJzs
zEgxk7dwzfbRDJPd49YZRJeFPjgRMu/5G4ADCrrzu4NLRV0/kDr3+4kN9MSUtY98
zj78L47UAfQSbM3F8B9D5miP0WNJAOAuvoMSf9uTMpudypSg9YYqH2vvMHC71aHT
AsUqTfE1JtAEi/UF2EOnSbdi3J72F8VvX9AbduIKbtBQSyp941DeBg51ln3IBxQ0
aT9dBSNVt/LF4URx/EH3NzGI5383GD7V7J1kVnKLEw2e4tKGCXJJwGjqIlUNh6dg
x4tyM8dNpXEU1O/lrqSy4Dde58iY4KTcPh6Cval31BRh/gM2TS52xoCTLZf/3oUe
ufq2p4rqKyisNAebfhJTioIZhQ3NfNXsGzN59f5pfNiBfWHXKMF8qaw+cIT7XSyA
L8q1aw4GnZs7vHgPOfnWBd7oE20h2VFrpW2YX0DAJCo+4PqqTl6L3mrl6PImzqPu
q0vsHJ8MTvePMAJ5JQ1IV7YfM4bIAzZOZ8HFlXKp/WN+4pCJIHVrx0oaqeUMuFH8
yCNL8AFH0jlA5KYfz1ybFMy2cyvyj3n1lA61MHQ8r6n1bT33rLfY1p/vMUrc9Ofo
MQIZ6BKp/eo/+LREcF598KKXy+6T28OAdyRofEPdeHzdVvzIYe0gBhpWEEz57ZWf
0dNMzUgSYp9hOZwzDYAVjgwLfiS7F/u3gpF/mNRq32hA3SZ9vas0kEq3eA9KZabz
cKIwLvUfXBBz4eoMZn+8pu8WWGUrWPrO7L4BLDrGQXieUJ3T2znim24sr2Zpcytv
7Lx151w+2z+avgaQh8lZV6Eo1ltxwRoteUNsT0x2F6wbRBOkQArtIyFuwFiHwNY9
NMZ+5OriBArXYscJjpCtvmrn4iAXaHJS/vAT67iKLyFkUd+tI3l7AOLiZZjzZjnA
1rf+lB42dPAsqfGeH+d3D9e6kdSoEFX4j2+O6EWagU96v2eRvZlfNpFR6yNblqlo
l6LjGesqVdo4/6A6bR344QMAs/8fXHspRhoqzaRbk4AW7jqgXjEX6L4WoUm117S3
LGVbyLeIu5j3zH4OSX+R8HLQsWppj2UFBxQniSFTwH2AmXI+4XXvkSLE0rkouhFi
onq+sKQ1IdL3AvTdaMKPW7nofjW7LBzLwEG2XCOCRnDSw5CV8bPSITuWYRiw4mnN
Bb8MnMICoxfOHCB++o4mT2oNKWThqyzR5s5frODk7h6YpPIPxgw+yFHKXOk1wEN2
/p5xpC6ckOzR/IvmNJ+v0E2VIJy0kTUlytbdvYLlQkHltBv9mCsUb1kz91mAsMSp
dQrlPvHASUJZjlL4LIL8TPayq6cVlbyU+09HFPW5mYrL87tEPE38jgghwpImuSiT
0Yi531Ml64gvVw0e5oJXT2T8czKzLdTTpYW+daj3lUTpbfS2KTggrvnPaYTgo0tW
ZP/ZwZvkS2qotFxFHPF3qGmq+Y/KGk7yp5GSbI2Dj0VC/UxbxDr07zL5SMDRRnAT
PK2udrek/6yysyCvoQxlLwmY/N1g1VHnA5gvZPQLEM1aUgpcjL2axDByES1ZV5v7
S7UbcWAlKOT4K3t0jCYCnryuYnxq1O/wqo8KLl8iGZrLvNCp0iamstFfcmgnHYNk
8QwKYWynaeZjA89jl+mRdiG4nhgCwUm5CvVJK4ghk/RVGx7oAXg084BKKyxe7Qt4
oGItdF8fKAQfev4OVPI2OAXErv3I6UudXmel/jxp2NqB+pqdLatLD0kmDD260K+J
Sc/kpziJPoL8j1TkDvDSON4nJtUzh02UVPeQyJfBCihc46oSibtPzJ/S/UNU3jkv
suSp48S/l5lYRVZTWbBN3cK7Ro8cgIxd3rA/DaRrVvxcredt6/Vgq4A8A0+deOAH
I8HE93Ndbj2GWDP2O1P9+ggo+yw16KoJx/DefXq7Pm1bLKfqPH3OrC8pbXFsAr0/
nkmSSydgaw/W/bsdl+QkFcOYi6Cgi7N8GwtDc7zmsh1ymhiXbXTJSKzUracZ3abw
YUme0AbUdNDI8LBx1inLDHZtzHh8lUI6t9I9osho/DQoO1BLHQdGu4anQv1ek80U
BGbqptRvAA9o5A7ODgT1b9igxFs7WRs9258sBY9xPLM4wx5NHVhWXTg0l25epVK7
6I3vwaMyJb/8/v5zNNH1bypEZmJKFMNEoeD9SZv+R1YpqjFzhufP+6OlyBkjOVNZ
VgbQIbKPPt7dtBr1OkMa8QvGCZdux8CQ5tyV/HxWsS6urk68iNy+qhHgZerBaLai
Q2IuFFf4B3trWXy0LarAxV8CtaDE1kzfb6PgNSEZ4aJZyt6nBZ1GLziMFHmIh0PJ
Ci9yNuQ2WjQhxtcDDi8qBu3subJAyYrUfJkkf3F6wTfr8909Mk4l5sCJV/gwm+A0
Dgrkw0cvCadFo9pfhWwjkVC3la4I63qQltdhGK/chRmGxl0yaetq188oL+sXz7kz
AMX3CAs8zUur9/+QxAfLc6LitwdzuY2EwRa6gbqgUEC5QRx05/3aPI3oU16eELA4
O0+MB4S45SQW244Whqpj153O7WNxRRl/R80okGXClhw4c5iWeFPQ8E2tEv1l4TAH
cApFD2pF7/3CBsublrboRDk5SbySOUwp1PCmZzba0fndI1EfDeeBrFlcxFV2KMQF
aWwVIdWbFpgSu1QKMpY/J/9/2UOepWDPn6Qr0qy84NhAH07fUVeAqc1/pNAk3/fR
/RmF7CKTlm0Qolsph3i7sK68Estn/fwXw6istM6aqlwQVfg6VWXRU77YshpqxfAq
xsffY4dqpOqtE0z9NBep2upMPFQuagTjZfUAKphPDD01pCmWEv53ZhOauQiBS22B
h4xMPGfrrR4jwTZtpJWLhVPKx7+tF5JyBQXGHaZaYJgQuqTXN1mkbXuUXwVzRiEQ
XkCI46L2LgDBHGmBCJHlXvbsuGM+thEwqIYdFjELB540ufrbMPEt9x8OOHrP118q
KeXpqaFtou1zYbwNhpIKThRFVSpU4qxFCN5ocfOei24DQRopFoCa6lsHJijnR5R9
TlZvv6i6qYOyFdMe+Q6doDgijWuNbleuHd7lzlZkNAmFsztzHWRAaOlYxAgyZXPR
1SQU3uOfGOkHpxUbljbpDN3cvOyUO2K93BLszpJ+h0fc7EN/wQ/7/t8xUsBWme8b
7ALMyw4pm7dcRwP8a3OLYvuSFuHo8sxDXkCzQKdonfXk8tRm2WvEB0ilJucoVUq+
S6BgpEq1dG3eWD6Dp4mSMvcc7NJIgEFr43KLtJs+TArSdf9Az0rL0MWkHRnqYqGT
VQmHkqjBwef3W8sEyUV9o9wItlzrOC3vI/d5kC1vH7TANdpNowRag7QCBKEvhY94
IzfiX8YUIF+j5hLOJbD+6rwubRKy9Vy642r7e6FOXKQECs3M8AkNlTL9zMjXN5G0
ENLXqLcFUHM+OJJ4jO0m/NPwleBaQ97BR4gHr9Wk6O1A4X9V/RWMRGvvQaqTe1q3
dWqD6vJsoAr+FASr4rcvZo6WTIjdQ7e+OIc9eYZBYRWf7KeAv2iwLW01Y18NC1Hu
NK4AGp4NGk5owU5upC6JNtU2yD0jKYVqtK5HGKJz5gGlLtaCtOUeDuhF0DDcEUn1
SpFruKGZu5I6itz6T4p0/2SKQnOehFbxd7mrP6nFaHei/StuMemhRccwBzi9dNYv
MmstcmBRLUvnw/AO/b5NrBNz+WQIK9QVngI926D4bwgGh536PlcQPXkGA3GuGRrt
oFhpkuvT2+B825xWZBubJkjnOiBj0uBOH2lJ89Ei7c5AQZfRsz8tuvD3Jwo1/Nji
uGzD48XBNzdusAT8P5p4V3XUEvtzTlgipKLZlVK54/hIOdZdV6UGxLirXFOJHq6u
s2eC2OYN6owkklNeywbsiTTGmwDf92uCYC9pGtvyv2pu3TKPHzJW4gXaEoI+qRiV
OEjNdciQsG4R8pc2yHPj4QMib/R7ZRk/taBoqy7jqwiJx4L+Bkk5nHYBMKoEp5c7
7pRRE3LcZGjXdA6POmRFWp6eaQ3K50w4oBB+QJdC5nmt3G30Q3ksNkG70Hskb0gg
bufikKp6pFTxfYoRfbu8seTdwZUUHhgAQfLpyl1lEeekGdUTwLM/vGcnJmQWuG4q
g5fzr+aMC6O/GIew10Z1MMnF2oEerkOCe4vFHs3Wei5rAbF7SaQ7oVKWjst/G/eX
n7uDbaAH6IasCRrKlGrhJeTwCFXP615kBiRxaBtMnj9Si8q+asPuCiP0aNilROWB
XKXI0gzSrMXoLAEdDKm++t/+r0Kn2claSohwKX2xV6D4SYFUTHvp9X6dt6QFYAxU
Ca01E90Gj04YX1BukEtnvBRgbHUQmh3KUVOx8VrWp5dG3PvyLBKNSEBGb6GJgD/I
MiExTdobULx49aJSP0Ubx/km/fzJy2sFFC5oe14LbUsJqb23b2lNgAy7VEdgut8G
6i8FIsxTzEqDBdxiUCIq7PGjhKSEjQ4Ud4DZS75eR8KSxYypKWh06UmjtdpRordU
w292K9o/RZX/0eqM9AADmqZPJhMtcMqKtogRGG1JFJ8ZKnjCCaGNL7yBQy5AuFwf
+7sjsJTlRyW/hSiWUEohyd7TXxqzM/6lCJVdEVL6edgjlEpMXW4+449KlGt1mkws
i4BFAtbxFGvn+Ts7HGPWjjhbVL6eFivNJUMEFiXXg2WSMtUpd3M8FFhG4kIsq+o0
DgD7nGOAW60tdW8UNHktZUiC5V8GB5Ud1sPWjo+HKCDXw1Qn2RfYJD7hwC6Rn6yG
h7ri3XeEnWVwguDxvxexQSYSnSPHGGggtMRXgdg8X4vY52hsOEyuvsiMeJhPN6bw
s9HqpXrToQYZxvZSJOLjljOz78hNFU5LtNKrY/gWH+cRVckdvt9/Uhp7L5hlxzv6
8Fs9vGk5aNs/IBh2Lk0eWc96J8wrfTjSinH2Z29bQVS8icNWW3B+iO2LBYbQtf0G
zU2ZsWgG/UdsWROoEiONG8ebb26JtkAXQYPeWUnAi4xT0L2oQJK5X8lGA3Wuimr1
YyHkkkORee8+3hL8ggBvWSUeoSqw56+tC1bJaaPw/vXcUNzMA/gyset6KTWfzDqj
gp8Dj2iDTpTbr1Us2snLEw+d53x7IYVtBbnVvJgAfiLrAMiJtTGxw7J8e3stjEhb
BexmrKdzEaTXKw9hnL6Va3idms2Siu6mS6XU8rsYTL+BPA0e/yA8lutH22cMkox/
+RguGGtYHk5b20R3epeDUDTKBUKOqQg4agkeLEgOCuJmamueDY0+M+kZUxSD73B0
JSOFW5n3eV5/N2AsqnVI8STRDySGeI6xWEXVsLc1VQo2FrsBhpb1p9hDHVQCKZ1g
rLi4FQLQGeR4lRHMC6St2GTD3W85cLr5q2kBPyHdBnueTrSqvbz7KuefzLdSm2pD
rEnrIsBSq5slMveV/hgHVSmrBuGsODU2tghi4EARMnkunTLyZ7XnOSjVdwmKikDV
6gq7Em9GOUFqAf1hk4TTPVMCiROCnak5DGzVDlr8/d4AcNzf38Rh4aEZoCDBxbiE
QTLwypn6boEpJVpkPXmv1q3YO6DqZw8hejXMQQDiqbT/miQjYoATj7Qa46QMvoEy
05ws0gttffeLY8MO7xBp7Oohf0M9RojmdTgplqpxN2smhYFcCsqiKTWXZ6Jvy+/z
s5eeyADfc9WTd1zRLPHxaxOXwzGGYvmLiGzQeCoeQmFqQEDWaQVv++yl4PqFKpiM
gJRbMKk3L/r5dpruydd5SNKGXkGDPpv61BNqB3MbJfBdx+2Z5Z9sb/mxlytYZWtO
eVteLfOpb90T033JZ3Yxa0lJOy1w4UAS1jmkX1pMZigQXabIPJOeVAkBh+bsNCtb
n0W0P5YtQCsmS7WsmOA6FV8PqSfVbtR5f3gSDVicWqf0gU0cgjDsGzUVOdpKdP7q
rtxnvtBLVhxeibdWXnWx1fd8gZDMcYy3oxrJuTA+PKDOyosxluZyCwue7eVyL5rZ
jWhaO6CX7fDCneFTNPQ/PHbFX/b3JQy3YIZNmbk4PUcdm74cxPfEt9Z5q/M5slxO
+s6COxqz9WvJYUQZIeOuXKwc5kOKLnU0aQ5SWE8dUWyEYyCzngxizs5U0/DA3YXN
mkh9xweog367/E/+F58d8axsEr9gyFag/qfvyzLafNdbF2GCXyDdzoUT+LQioxks
riNCUjpXGOjHLwaHGyzr6+SaFYECReRwyRSnHm0BoMdL4U2j2zRKmxVHpSesEdKM
P/gBW2NiZI0ylaU6A67pJ2dH3GqY9onUaODPKSR2Hb6taxkvpoeYNcu9Yf0QiUvO
KcUHreIYOhZULuElsJE9HP0QoFAAFpWaQy2b479iXDLDMJF7g3TDi3pbt459MQCl
ZbMaVotjOkDZyMJQ35ISf/aUc6Yk69162fCrhpSf+p7R0yB3UJk3EFkj75V+j83W
slL4Yp5FFARU8z5uv8c6U3VA8L84zGYunDMAAPlIpMkb4DDM/gKvmx0s7DKSiht+
ZlcEcaN+PzU2WhsanOMWZJbu1r84pljwx1EXkkd2SapHwI3De6BpA6oe6pYUYNeb
Ie42Y8pcKh37JClIooqAGBHRCRcDhjDVOo6RpIi71lQjf4bqHms+Jho6Cz8jTwPK
Z771L6BjfQ7V/siO6KKuX7hej6G7XmMkKpFMH71BwDHb25YM5gmsX+iOqy50agcc
AkBNUoHKq5sUK5xdTrshGhe47xiame17nMjLCb0Fy2T2EK6yhICB/gUvpaDQbgNC
mTN4h6VOpvYIsEiVf0fNjsPCoC0Ja2U0BzI4Ixj9zuyALq4WGf3tgHCV3vA4VsIc
F0XWDJkvObCgcXZpFh0gWi1iyC7VvxIMaDzcVIQwuP9Y+oHmEWVXJTKPUU79SbZA
y8cijTE3HDnCI7ojAd+wRksPP1qUP6AlvRWRulVjd9XZ8MfWxLikKeBQ/MSXtWJT
O/zax8o4O7Rf5XplgokdTZy3kkq9uKpBaOhjwBI6cf83N7BRvaphdsTKjdGORtEc
vTPBlnUV46vCSyv2RYlT0gTeKVTXcvNtBC+w/3Q+GRPkfMYZ7tVavR4LgvBh/h/T
MU5j6TgUc6Zkx5cZ317ASS2+BE+FrgVGgC1vDwcIpuKnsfL0+D0N7h8ayHoZuAai
aPW36FACo5XoUNSWHWbSLDnofXyqMORX0oPaJMIj7PKUQiglY443HrG9m0nvzLPy
NW45+1xhmlUbE7yuqX0wB5USj4ukSYCM79W6WvRg/yAivAnMSebPOP7tcHkjblo9
gGhDvxPn1xT1wzsaf0tgJRsR/fmXXWfbrdRmgqYkoRb905o8K9QP4mZp44WxnufS
ehGRcN7uJBLRxVG3l54DjShay8KffK4jJlpJAnuWBRV4w2+dNOapD1dJ77VzBOxy
zf0cqdrzILiFBfT40R5iH8AnCSeNG0M6cmcIpactwxf2olL81BsfrSEblBwIbN0v
jZ3NVniTMEM45ehPKyELRp8XOW2BDtM3TpCswl2uTL4JFAH0xzRY4ub5DzXqXyec
nOX3IYI5gjFI/Jw+TWJMUsyCdFtuV2d3YyLw/F5mmZtPCsfJtNFgYR5lJQ9nljdc
yoNPCgTY+B2HM1sNymKNpe3lCPPnAy1pWCPWHnPMkBSSiQkBqIZ55hq8xJO0gjLv
wo6SluGwj6uDB2YymOwmDchLvr4Hk0WgfO3IsqkxEtLerTK5uJA85SUxnzoSAXUB
jR5zuBa1xjdVdx0Q7yJW/Cwaw9NBr+yXWu2kgTog9Oqw/UvVlu4SExxxlOHtm7fT
2ZMmJiCjzXz8zwMYtWMb5BHgSuylq6WAlUyD+GNyIoOZdtzbFE2dk3vYtjoteWh7
rYJAjxJ0fYH0RRXKEWIK/I7HbJ2OXpSE8g0eD0nYD9VDIY+3MSjAQwVAs9pGJke/
OqSu4MTWl3ERlz5fIg4Vh2l/RkN8cm5PBaIgZMESNumPtcYYrXkVWlCm0gFvZzMv
bKHl4x7oBRSMS5cbOWlXO5uw5UL832fQ2eh9kRciGqWvHMTcXdWpLmRBB+NQBUwR
KVxZSfyxBok2UYSuD4CEQQxZEyg4ld7SBnIqXJM+uUH7z0WuYpR3C7BwJ3xX5TDP
G1uwLmdjl/1fDEL6BXlFfmW9aeJRzMEWwkOiGMpKOtAH/9G1ODt4TYPHzjqtK+3V
S87yexTxSvNUHAlH7jg5Z+f7bhvZtmmm8LbLUY+HEP+U5fCveNP92DvBv+DiPk2P
zC2nfKkBjS3UrtLzwfcZhAmYaEOU+FKNlGwEi2REd+F62SH7MGv0OjjN8ZkF1jxd
IAKyC8YV4OYoH4h/Rq4zs5Bgt5hp6rggNlg6FOnIuFdknzr9dMmj7j3fqHj+5xju
nwx/HPwVXnMZqRLN4t6aI6Qm+Dvhb8dn/JkrHwxCySuNMtoYfEt04r2Z5Mv/0JQd
04q07aMqyJpL3Vkr1cbmy8YzrrsXt5tfnGYj6UDiDbvC0rdynDFyXJxmb8aIOWRt
Z+INbc+/IcsM3+trSgsDq3gWyx3UsKw5pBozSnVnJtIxz4TlsnLoFO19UEpGpPs7
c/9uF8iVajiUCdb3UKQFZFv+yy1We4VfccbAdCt9kVQYVnI/8UWqwJmAkSkt9wEW
rGd5FfeTUWC9Bmc4khv75+VkX0wZgN6qZMeifOtTU/IYtPMgZPQmD3qxGfbCRxCk
m1toZz/yqGxjSUN0+mlzYvtwsNpPRdRcsBglvohlk1Xz+4kHSAg/y2SUU/X5Nd0n
RRWCqVFWgzbBDPt5pmoMdmBQ1rBcAKGhJj4uJY4xrOn2LAzjICLukNEMsbYHhePg
Y1B4vjiqHCDacQ1mwx4JOiWEBGtmeTR3zi44T4FqaKPpkr9qIDq1JWTL/mizM2dk
OjFETKUxKt3HTwRE65IFQUYvHzXInay4+np/i0kexlCCnSeD4zNg238eCRh74Vm8
h7/FILfwTdOxhNKseFXLc+ZceGKW9tpxQa1hXp+uFC2vkHV8/HK/XLNh597nsemT
lhX41/2t4JaIyTgzGthNSkFx3rMGFSKJck8SwO2I39LhD5wTczeSjXxDI2ibtn+u
gE0ia+BVE907w9KHpg3dBzUF2vLd7DGHjD1FEqC/0MfLD0YF5+7knrSCWX4+s2/4
1niMDrZ7qAFmtayv5LO1/cbzizW23QHw+z6VtqfCadxfft9teacZG7rfgiq0a0tJ
KPNfOze5TcJbss4MVJV3oZaV5lrLLzNCMbq95mvvTGufwY7KJFuzjtvbRSBj+tTg
5uKILfQ9SQacgUDXtAuLqxZ0v7+KzdhJ1ZSjAT6tkMD3yvIj5xVOhVttfr+2fzYT
8WYXusWo54DnflRvbx02ZTejDsAUbaqGnhpkLnqvYPkxmnhp7SNZWTVimyNuLslQ
HVxGZ0k4U8i+TNpo9sKrN/faT/zOEF0CUlSSeWu9Pr7hxAfO0Um2g3ahZZm4Fy6u
uRCEwkDEBftMeLM2oVU3Q2wO0vJ0EaR0TxvwQmEgvdXAR5314I49gEQ/Q/qQYw3Z
Paj/vDN1Oplz+JAZnehNXUlm7znC2lZ65BgnOsRdLudDlLg/XIYEnXwRymQZ5U38
YPJGhqcgBRj0IathaYCYMyHN8pVHi85Jkf94SX4+FdmuCoE655lxEF6r2N8wo8Kj
c1ZNwHN3YLnwgratGnxbWLrSgp4RlBl6Yg4iqGLye+CPguh5j1r7VaQx8bxzeApq
1onZ+1FOyxK+5A7QNVvTIAnRfXUDP8SVJs9VryawYvXSvMdkev7xlSd8WLcY/1vn
hIBGAVrjL55fm1igi+drkaI+7b2nlrcimT4Tf5nySc5j2w2ILB+aD6XLwumtxwBq
10SoCQtNQUCmjMNEQh/Ua4HotsiHaMJbJV6NL7hmygtGqfciIInYl30hjpiq6yV4
wwPEXoydp0ibNExCWJvDGfP4a49YC+wTUF5qrSTXPqirfi9ToLNrIy/BL0aGtNK7
xRXWiFVke+Pr0XZ7lW4U7BfjUPVfRUok3cu3fq0FzG1r9qs0pgcblHLY5T3VI5Pm
LSscvVoMN8XowMBoCehaRtjZejmBysScKbl9oGKoIW0ojkOV66cThnZhFWL7vSJV
FdaMn9SrSu43ir9JBmUnTMMSB5ryCvI6nQ3p5y7ceUFkI3nRpUT83R/oaQS2LSnk
c2QO/jl6KXTM4hbSTQLGL319HKTZhMAr6VUzvvuyDErvL0Rmu1PDQT81S9q1mNe8
6erv830pIJQcGTRrHDZBlH0dLBt/QD7UTX8De3TUsUsC5ue8MdkU+OORXiPw/yFw
VC5wEN3NrZkErH5OS33rk8TY4JbKBTnXoXIrGv2wB5CVHDK//u+Jr3q2VDnERKxh
GSXK/cEPKd2OazqU5jPDAJ0AziRIkjw/2Jm1nl9G7jBwGDIl80AbmsabaCJrZb70
7y1BAf8eX9gocklTgZasODgNmVDAh0LvlDH6KzhBMLdztfpvdwK0jEkmBOfQNqLO
0EX08tkx20GnZwfMLs6VsEjdJ/k+pmzBwJPVt0eUT6r7/wgvzAzMFmHsIp4e17CE
e9eBTyizQ3pHN3CaSOSHUZgFRzwezvQukTH9eMr6v4iUuqYczTMZqUPhd5lP6fPX
dnxvFz0O2a9OwSNBMVnGUFnd97RPqltRHfdz6EUcE2jpF4m7MWNd4aeweCACrHoD
XniDnXZotjTitCuH0XQVH1wehJ0p0MgHB5FBJ2G0vDu5HT8cAQzx+6TP0rMmGQ3o
j1iOVkFq3e+AeO+yG0ZinsEzSmvMgPMzmyQusuQO5oPUoqudA0JKBvwLO4X2muwx
JlOQTh3gw1gRU+wwqW3bo5BGYtgBmwc7LXiH4Xu+DQs55jLkrKLVsNi/IZc+z5Xp
4UXZ2SJUf83sQWrf8UP7raM6lRSZJu0MBMc5DnFO0DXGI1dYx3jLd0Im1yJdkFi+
onOKz37WDRp2dtl9wqOT5Mxy2ym1ZraPdpTph4OFfmhjI4BabYnZ7WAlnOVZ8+rL
Nvra5wbxoof3tZw7Kqyb/DJ6xz61auCeMZduLcKfcOLlV4+WAvNArBTfLp/Sktvb
Sl6t/cQ/ITllyCmrfE+G+ARnxZj9aucLCXZ7xr/DWOC8DwSzToxBzucLOSB7CDU0
Ec0RnV1ik3OtuIxptuPJGe+WTgofccLP5A0DEbWLjse9kSr1I+BJn7w8B6IyIRDh
VBwqNgfBBeqSC7plL55yW9GDTWpsFamrQy6VcSToY4vSp15GUhxra+8f7hllNIPD
zb3/dP68i3PeeXqCOC6prpRAUqW5/CAjXmzlqDV1JKFE1Med41K1x93K5vpt2frz
fG5jCOTEIZcIgVtfw926Dj+s/apL4n+UGs3dTTw8BLRUVUIWBo19cOKSxz9mFFub
nN1zy+lBkgGYL7x24auMoa0DSRaVo9S5yl7QbzZdnLdGHv3Wmljt+pPv2DRIafpr
WS5gx7ZC0oLBLJZyy4aYbbJVzcuYXXPKgt1Kf1tCBp9kL5a/prBlmaVsdFlHRlop
WweSch5hIS0HLwYUFdGQjE0bTAS1PtR8jVSEWnpoTrZEXZ0EQLDhw9KcNwEGz8Sa
IiB0sspVkFPkdifnlVEk0nYbC97IAW0tUYFJ3rVWzylcPiLJG6+qyKcP3R0Eq1Kf
Tpk4sQzZgogZ7AxMd9/vhaHdvBrZp8+Y++q7gfqwCABS6IAWA9TedJUGwMkjNjzi
mPQXk8kHFncHH8LeDXkdHjHZsiCXE0sanRlmBJ6xog/wbg45o6trF6IE+hnS1JHt
Xh0Xl5Kmagf/2RzS6UDlSnC3eMSEm295PVm2RLH7eD8tsQT4WRqXR+vduEKlrPD/
cncIXmITeOakybAgycuTnlvO22ahWAsXPsoB2rsQRnoegolNJq8TthburzrqzmY6
GpGGlYKwggve20gEWFwjD7iPAYr5z9rpY4OPEZ2O6aDXPAUZvZ/BUJ4kioH4258M
Kv8YeeEszWQpKN+nvHJI/YGmoVkL+IGkR1O6o2c4fHHewzQdD2Vgbb6vRQxcEGXE
0iOetG+Tb46rlGIToYJUNxtFCsTbI1jceJE5lw6+IBTmLV2lncf5sHhqdlCOIpVp
rzEucEMMlM6rM+DH4k21CIT6ngZMbLBQZ+IA0meO0Xv3iye4vg3z2qeisx5Qfg+j
OVN9z1GBCY4wHqio/3lwycB5+JTSli64jV5uCl2tJxqULm46CcJOLJoVkCQRPSqV
gNMJxD2A0oRibcFy1B5PkrA5VNjQhtU2Cqur2QlSFrckfCklog7Xed0Kn9o+GqjZ
Ik0t4X7xtfwE5HQzVj690FKlqi1AXQS+Ggj6C1EtGY13b0VfC9XhKLVHMyegErVw
OSvviLLWadMImfCEWpxAPg0OzCdvPuXaCbp4haB6xjc6MlFoKjnDEgueJ5Wuryuz
UuhhoV+63vtN8lcU/syi9COPuKEtfISxQTRB1TKx+DiyBqeqRrzDzEkxxenblYj1
RGJ9Wle3NFOQ5A4qLWd3S26r+OZfN7JXlgD8QmJJXRtDv/HkK7UzoiLB7gKZeNnK
SZCS1pMwiYxkaBwN3c28j7Rd8OAgQuHG+4KPf2ZxMOwSLA1SJuLMs0+rg2S/RS43
jYGKaE3feP+AZChApVkV21BCpNWReoS5plxiLMYL2NXMIbIsjFx4iKG9PvTX5nod
hlhGApOyPtFD5Gn/0dnbqPwbCBthJ/QDei5WuE0yEmM6xr4INYHNNMKH08U5xjHG
5diyxAdpnnmvmSodTgbxXdLTUxnJwVbsoa98HYLQZlFGuepzSMjGFvI38CDetDoC
hJfwCnem1GmsXnZiluHzzzZ8WUAHmE4dv7u0XXBA9MmpCRSVQAxDXgECNbG2oa7V
lcuHlWHICYbO6JQcnchFGHng2JumEcIeHMhibfRuj0Xc9LoBv3JYPbwMPD5tyWWo
IL0ZSzNVVZ/PaCvYR+gaq9fgQUKwo6ddtrGXxKE8DOqmvCjl5McXfo/LMteVJ1Xa
3d5O+Uxu0Mo0v0owzesvhaDdsR6ahBbE5rAE/Wb9nX9fkqg5VSS0KL4Lr4H5wIoJ
nS+S+60G6LSbRjCdoiBGFvylPtL5cqAlrz+9s7EUbx+lso+lXQ8xjT1G0SFlzgnD
PgZVMNrnmwDjGK3v3l8CQEtAu3PqL5fwIRfIzVPAMJxcVEW3bf/lrsxN2bgDNpXN
li300+CeMFrizjOsrhvhQ0rEyzm23qk/FqPrAEBW1ICLYz1Lfwlig6BRnQexxTCn
ui/UqHpMqRKMvPHWCYambweAP6mi2ueN25cq3ClXGRdNzS8W5EVUH2GtNaVmLzFk
pvPgXd70JmyzachD2FCY8PlcJyOmlo1nC0q8GUd73zRQFXa1W00Ai4njfJXF1WVQ
OZ/PWgYADS9T9g7WSSNsFId6/b+3texBaBIOJhLfO3S2sEfURMuu2qpOyLhavwH0
e+z6YrXN3ghCfc12btK/cZEgnlN/gsKQ1LVvuN/lds9QJ7p8EDautHRUM5Wh7GBH
aifgQaJ0w1v6eg16EuN1tiCi6PmtaKPIJa8P0NdlRsfuf3eTy6xqv7v0+NpkOWv8
LHeLO0cxbXv6uHzQyfRJnpCQWUlYd5DzXBbwu2xGOx+adhxOjB5UikRZtsdWxwow
KboARx8SbuI9LV3Z9SfxdL1PJ6fcPqHnai2/sCpd6HODr+N0NelFjkJQCEykbsde
LktxugXLddxM7UZ2hzx8hbZByUGcGKaLXW8CG/XFzeJJiR/w3y9D/fqvQ4aBCiIm
Gi3ihbWly0605L0G7sctSWNTbWTepuiESfaoXi1F5c+skeq07lJSp1az7h1G3fPl
kKpj+n8N+x4C6UOtE0O4tfpMqD0s5OTyLt3MdAdoUM+42IDrWdRjF3TTMRK6+4kE
U3c6aQJ4xuK9rcsq0rnbXfCYwywAUENR5HVV8hHlUXvByKw7Ch6BiwqsgAT4bpTY
QG0dlYgPZ9MqqNWd/l7NzmoHa4cV4fs8VD3r0WswYwlqF+B5TKOOps9jaJsgSV1z
X2G7eCEIMYlQdfPeRxxyFl68TxZJBluSL72m0PQ0Qugq8FNzWCGyK1qXBY2vSr/N
F2axeTDYdOl+36DXnG3iVwPrqHa7IWQ57rZFUWmbv5YZRdGv3aetOx+4GWzPs/8s
o+lMqErIbOQJ5Wsia3AkgKYVXOUqP2RHmWoFCRQ+0v2o5djjl+u+tqPL+AK0onMn
cfC9jiYjoB/6hLFpwKpKQ5X0XpYD1AYRseVUvC6/J2EOh3aIs3g7eVSXMqN0PIUp
zY1wFvHhYBn0WtD0RF1Jg0dkb4RMhU/RtoeYMLjbNrkIUxzD+Ek+qfD68WtH1SEu
TcwgnJUharG3tLXegNGjY8qfAPd2WWnBlX5kqDHmT0/I+T4oWvYKd+UmCyzwJ3VF
EQoJtzKsKFLZomxgKVECgVwGj7fmJSxcYEHZHJ+w4Ba/fVcGrnj/KJNSsS+i3C15
63f2zAoOyl7pFKGPdFlUfJR0nr7/fQ+fLqM4cvdAlmvriqzOzf5OKQ1VZUkD+ZLj
Dx3UGc1ia+Aog+rUfI8whsvQ4F1g3fO6zKqkKSY1OAS7y2zYhXnbvWMRcgOVds5i
uDk0W/xy1BQq1kIDEKXJ69DynqTRdryDmbNvVX/BOfZmzX/jaDX2fouqHXIdOwW0
XcNugNUKveIw5S8WlguGK8UYUseyznTtcxUJ+Zd/YdayPePXaazW7hnfqBks9R85
m4yr/KYu/mvLTuoA9zRbe6VX2Pov0FChkjPM/gzvb3xrsLl3DjgRWKI72v0uF7hB
2MyXfLr0VeuXi+BdsxzFRQUIO7rsCi8+QkPYQkJKWO3tUrt6wkNnxhID2dHPoj9m
GxDr8M7ylqS5odpJppmdISE6o0KACE0PO/0C+ERZ0V5v8IOaGkYcnGBRrusLNx+T
EfcbSRKg4brfvZEFTwC2Ohf7w3xSLmOLal4LuJtfG7Pjx7y+BrH4ENeZiarU0nYP
kqgGBO4/M1FCDAkVzaq1Frz9hsW8dLnEAl4EwMnbpd2hZ8H6LC8vj7ihmbEP4ztO
yVrcr0r6p/LdLP2VfVJ9o/PSPy5qfGvQwpfWPnaGG22sE2Gi0r9JoNXMfiIDfDMP
ZSW4hbrm5oRljEukJwu/d1EMT21zvyyaQ3OCVkojD0IryfU3DQfv8IhL1tIjnu2w
fjbh3INdgoqi7SqHMvsmUhl/uexYOjMcClR9XSIi5chKJta5QgSc9Dbl/DBGIDAh
nQF5xBpmGqI1lXLCDDG5PVYTGf44rwPpl6XMXrrCN6+1Layl09e9yaWl21zYR4TL
xamGEpaulJdobxIho/jYvefb2MgV3zb2OyPk6pYFVinNCuAEK9Zb4bAn1CJdeupp
aKtUXlUFh0+zqUWc0gO13rBLpkerfwgJmXGRfXW+bHLTk+QnxK18KwE5AxqHS8V3
x1FLfRWGBkKNZ9bP9XqhHwWdDgzuIeOvQSZzZGbQCyd444yX4k9NlDi12QbKvLkV
RM63KpC1YYewgL1yZOU9vZPyB24oVoByEHPbudd1DW2OiWY/wphkm/9p+8m/EVv2
sX5G8+W8nS72Pjxin4XyLDlNoiAgItXeegsYqsQ1+X1Ac7kvgfnOw/grth9RvU6H
Uo3AvKIHM7zjxYxV0MIFFjNtHuWrbhcmH/Da3KHCIIuSt0GGhTlvByNpp/PVeQmA
szPOSL5Htn5ZyAvUJmUxmJBjOnC/OP+Hig/3EGK2l8Xz+DrG+k4ErMLBCelBm+Z5
U1m+mFj6UBWBp006+CoT4qRxLXdeOIvWao1KceZJ3eLb1BIzhzRSl1u+oJSZZ4v2
vV5YG4pqReSpzCNjlJACuc5S+1Zcl/qZo6Si3co4geBlaTWH10DzODImsRkAevrd
Bahi6Gq//txDuiR62N2ZkpvjGbYrD/vg7wOYMykq+O0tB6RfXTMbBXFp8/Q2mtvv
7fOooqf2W+SGCr1wcHbI+zAP5ZX3K+FjE/SHG2Xk2x0dyV/g1ik57eu5hvCVi1dN
5ApgS4wriB5IhBxpmqSvYcAEe/O+s3DxRQnZcSYUOF0cQUz9+vqMgK3XpztaRC4I
VNi37bmkJHNiIF1oekJqPIYsWKV/IcwXFP/HQtlyBl+UUS2HGaYs9CsQAAHZOCsv
eN+u8BWFkwuS2YBxQg4ER32JTmDWrCpqxx+KVDcI7GEMO24gs3ZHQjN3PWQ6AIN2
6ztQvZ8cdkwZZSukQWnsRsTL3nv4Knqwp5FVV+Ikc9fvcGG76PO+ZkNhh8RJCdPO
PmTD6j+hLSkoCJKBt/mlrq09bVCIST4GDVRa6eVr6FGT9IujUBwPn/1b5je+KBnb
1Lzy18eNMcuTHYlzyJMFK/hBT43kQdLZL2Q7o+NxPuRwISAXEJHK/knylbljsu8Z
zQFJi9pnXER3kNx9Tfe4rkPBj8XeXTaMVAGyYqwX3MAAapR+/VFtB+4H4EXufn1f
TeKRJh6M/tnxamRZMRLWoeM39s5idaSEdDKy3qJfaNoyDgLoJPsqHdsYcrtWeTvI
+AqQoX3plzehKBREJZyjg9a9CRiTibweDE62zaiDJK9RvjqGzghCHyZ4BQF7Senk
NW/tLE59vWnVUDSHwQcZ7/HfCYw5IEUo08iRFNanE3wn675a8bE5r5x7GhdaSkey
KSkvRvMSMbpxdxCtgXxNvYvDQTI4KmLabShQmJGLhqeLOwWysIVCqbN/0cfYvmvn
VrdPPzGreXuDJitMzW27juPea1Bb1Svq8ha87W72/HIe1Nkjr69KAVibgmhfA6tg
9fkc8YiaEiTV8QDu0s9FWFUsUnzXHHqNvwAL7g9AnyLv6bPZdPaOsTC2jTwNKREw
qFxG3gyW9oeVw74R/vsAzXdIIRRHXmaP0v+9uZ7E/n9aegN0ddDQYjLjY7X+TnGE
5eXNJsrKoYlaUlUbQoD5OKUy+CXJe3p9ixGN3WhXB5UcqKXFz6leubrhlwTnNEuq
LjzJ1ewdac7cHuB7l0BINPhUrv9AzdvqJpgQ9cJTWJTsHfCaASEa+TezVJhVHZAq
x0uq86f7Z8QXoY2A19YhE1wTLdst+cHQ6u+Wf4BGsSAxHsqM1ghw0mezDmx7vIpw
oDD8agbvvND4Ef64VVSlUQcqLiQH14oSai5nmNYqnyPIecpkCtO2wObe7Oh7oghX
0GKZjhUcVRuvoSx2mTpwr1REQoMrLCBYD/F75NVHsrMjs4gC7wZXjM1k8fEbKKcq
FoAfWYf2CHpc69lLiko7NC3IAzU6lHMUaOPN9N7XnvCw9JZ3LzrtHonhkz3UzR0X
uo6QWVULvrnBEEEOKxWCVWJdSZMQ7lYI7Ffco7G4eYUkmhvgM8nTCki+Y+iV8XlH
PKPdqCQXB6UwRl35nUkmLb5lSER6uvBZCB9kKcyj0ieedsAqdy8NU2lmcKWw49KK
dCKim6BCKxris0IbST22BvShagF1ug7uKSQg3ZdtcivvbfIhXf6Hcl/EKGQ5U11m
xH8gJyNCdGZgHwJC4ii4/vUBAB5HhLOnQfMkz1RuyKbk+Pnw85Hi/6qSCbPMqW/G
3GvBsAy6B96vLuxFu+nKIlcsS19GScPZQgrsEQxIWDrjsXNHBnf83TvUKJhecuZ4
w6ycl/K7q9BlCMK7DV3CDL+ztD7OyPMh+tsDjllPPgg0QzZncIbP3y54if8kjJMm
6k9ucuToRjWMvf3d/71zlStUmHu4WmF7L4lgffTXf1nK7swi6fh/xosKDuzD2Jwp
xWHa0Ql4nRmhAXWycbUHWH6x5878pWY/RRJcazK7M77U8HVHQMQGydi9jNA5G1jt
y6SU65IxoQJQwphFsvjg8DLCigzXi6+PLjTFE+SPf2IMT8YytcVAl9g/pdis95za
hJt/Nz5g1UYFYh0pitE+oGwP4AUQ6NF9HqmUx/XSAVW729BRL3n91Awvb2w7MYxj
0I7e1BkkP5cO8eYpAGoDVBXZpSvTUIlmFJ4I6wMTX93AytDSregknJGI/Q2z1UC5
wG5/lagNihVBTwrHOxEFS05NFBe5R/tQmb4VcA9yPWeSxVvaTCZT1N0gnxHWVUi3
kn25TL8VcWSf0P7wE6rX4QYC694l4xizxOsg84dXLe4/dg54CWMOxQI5iwgU0t8k
1hf9FSQdXjqZegQ099O6v44UmJf+fo3mpJEUSbkGKE96OG3T4vSEkCeSTulmCV1v
TfxndSLyczTEGkYV8kfpS89IWX7QsIWWReGNqyG98ypVaevWBf0ZYxlY8vXCGSJQ
k9ldOxbceTCQPPGxz2DqFYHGUiCL1G9ulNN3OwokE+r34qiuiOjTVwp7vYtkEw6n
IQnZnQ5yXHjW8Ld2Eobmrx0dbTbykA5Vl7bhca0q4qMButfZ0Ec7DHAQGIW8MfVb
ixAcExQGe9UgRCz8QccWq/oJyfqc/coREA4SxVCODpivfuhaaCqT1BHrkUxuLgO9
a0S0QpNraXdtmxFNL4DIvv3t3OE/FpNJJiiQu8cr40TktMMXYSIiLG1vZ9yxxpL7
ItjM4tvNFyVva5GsZGPyZJ3UdY8ReFUq1l1jAe6uWF19MpPAe7nueIqvR3VXBMQS
waePJ/UUv2pmGnXhF4kF/06Hsc8ExgAq5AwwIcNZJgpK9TRP8gBQzmMReCFB1BWc
Zjp1i85LBEniGFzKTgsGLwmQ/SyxqWomJqwjqwYZwq3OHsl/KEtle9Pvb3a+ozpt
Ewo3iR87F4g6xmtOmK4EzhbuQzXCKB/qujBeQn05yk+UmEFygSC/wjz2RoFSL0C0
lodPz7YKprAUapvCs9ett7m2XNqg0Wq/ii8LKS+K1HRO+ZJmPQPf/+DF36RulFUl
O5eK/J1NxQQG2vqC1a16J2kWXHgdf9hJuKWX2+vE5V2/5d2yU9VJrnwxDBzu/XC+
dRSIvXVigDRAmOpDsiERI70IS+w1nNRXzh/YGzUqioRqNV33YD6o8yOUSce13mSC
eNymisjBj4XZDgnTwStY/iOGDNAdvLUs/s6lP8O/PtCtz1bPsEQB96QlfNYv0o1W
+bF8e0+Idrt4Y+lPKtifjzfeUIZhy3ewTCqih2AxxXt1YXuwzfJpa3C1/kQknCnh
dFU+9TRGjzn8ULjh5Z79M6SzwgU3YnemBN5dPBR+gadzLwHaucl407R4AIvG2md9
zG5MZIEMpvTufd+autqqidT4s0qZa3TEcifxKPYZZw9eR1JkOYJoTEDxy6uZ/7oH
1dKUBhbdF9Rbu14Izerl7xjlrmInXhPAJzO+QlbPHtCJ3sSPHasdxzRFREDOAp+W
X6bYTwOjOCnHXZ155B48EWO2gnHgV9afopQImKBK3brWEntSzTZBYVoCi+Qs/hYF
YfMBaqNrPuATDuHWO8yehxqkKzUQwHnw2cG9leL7PRPHrP5qag2eh1c3IwxM+zVJ
G763Nxa0vpZgUuM2YgUfww/DUZYFv1GRqJa2KCbKi55Qj2+OCog3fv95Vo5nS/vd
cks61Ip49FG8tqv38bRnLJzMKyzMfRG7gEPOVxQsRB2OT+WbyWSnaI/sVJTDW2Eo
JRPg7lHrrgPjmslbcPNRFKBtfPg4IQNj3WCoo5zquIPAfkUoy5hv4C+2WIjzfmYR
4t32D8adezjTKzfLXSBeMYn/bfzQKc7OKJX7EdcGwzA7afo+TSVNaEYOfThUT19N
vCyQZE3e/vZWKXvSqTaBXIRdV4MYMlD/HeCN1lCqJ23/fcBN672uetGTlzj63rtY
WWJ1oJdHoKiltR62RfgkgkEbdBgEKRLN5gXNaQ6fP5KF0Vw2d1ZfpC4EyQ+6WhJx
qLmq3pvCqTGi4uJNiDPO5ksynP2d3KawDbpq7WMNesS7YHl7Go6OCNU6dxvli1Z0
akPJTWUq6XWrHDyNP6396YXX1fxAxu7vvAOUN3MdASHOZhsFVpBjhfxvl7iFmcm0
JIKnhKqtxGxTs267ipP8s8r6GUH0v4DtEgnjeN1NUZv1Jp7+TZUW8sJRiq8PjmRe
EtifhFUTINykzaBn/8Iis+4KIUNBs1D3HtuvucMXYesBU1oYo4YH212qDMPyiZun
Et8Re2iKpKQTc6rlArud7/xfmxHFG5TWuva+bNFusMlP0ztO3pHF5hC3ZjjZLq6A
4UncijaO0OuKC7p8Po0OcNHzsePaMhRi1YRZGaPez4VnxSeDU4uVrZG81EJrJZuo
qcIw+ulgYHIUCF6Qeslx7pZzXOlUf4XYy7wSMHiDLdiQQAYRbVp2HRY8BbdRZkhR
d5uBSx/R/9Y0AK/UvplchPTaQyHjJERutoq4pwNpEjOe2yKg+r/DtXq968OjgY5Z
v3q7jE2B9rqcpCj5ytpI3F2vmX5zrFse21HlGaxBKyn+JU+bJqN2+6ApiBOqGV/7
i+f9wA4j9Zv7QpMFdHdlfvTwtLEoHVihTbKg8PCs0oHtkxg0ZVDv+p8vC/jUptxf
VqCvgx1H/ectUsdv/V0lDLDoS47/UjMD8aCnGEsFiBbLXokz4BfwEp9LYtRBgo4R
8LSSWBJmFcg2LF5gEbcdktOgmYcgMBcqFmvKLVy+WUuVihVpfjWQM5CpRrAjb5Nw
0SAsXTgqitTHMyIb4bnjSORGVZwk6/jxWh1YPkfBvwxZoA600u0tqRHW1nyppdt6
MX/aokQviX29jzg29VGG71fN9ISN9BDPWeQOnn3q2r89rz11YvBQG32fqMItJHjX
CKv5+kg4J/FO1h1hARQImeZ2LX0CKHWcfzAT2MPMGR6K7o51JVjf3kI4mSE4gJtA
61Ttuc1WTpM3QZ/WRg/mde6GfEIlK5MNPd9NPmObMOsLwQqPRyzE736OkyjhepGA
pqQUAhbY+JZE+UUV2+QUmebjHCrzZPwwpOLqd+gDQFiuZApRG/4qusdEIyvz3LHD
6A854QjJNP55f4j9/S8PgQDe6tuE8M8TJX5KzP5/eUl2k6PrmElAhbO03ZNQTcAM
dyZYvINLeqIE/HD8XsvwILNks+mkOSacroywOefibhhefBMmo5ibGFe84hWEpfqF
X2W5HKQGsHxRh/SdjJHbivL3K8A9bmZZFnCRbDwr3wAlrpXxe4Mx3/4Xc8atcv7e
dnEsDizxHgzLropKZgq63tOjNtLJXEAkIzemY+sYywpWp0GA1MZ7ylDvWj/VX51j
Ba6GeOijdsWmrp19QNoB+mvDDPTkuCTtRrNeKhzGjgZvYCcYNifhP//t8KhLBZTB
xlP39VW8xqChQrMWctNNL2SO0i9mV0cLTHtrDNjmqCZHxmIhHp/LuyyosIIoJfZ1
Qd6T5byQqpxsXUHp8mJbzjeqxEC5tXniaW5VBRP/msnxgk8PAnCn2u/zWvYjx3lQ
SUGh1otlyTafVCaTtdJWqcd0LnR2LX9LltU6cjpNOjvkIktyvj4WAZ2+EBzQDimH
eKzn098VOjlnwNCmGh9fsreW5Kt16o52uF5rbKCynGuHBPfXR6CorUsS85r03WJU
d+O65thrpj92OtycAXXkOfw8fcn4bvWluZlHfMZ5V7FIKvcOmqZBIuhf9QSs4URl
7OIhskpvp5vJmsrpObXn1pvO8jgECqQ7jo10l9Rv4WiqbD90L/eyMDB4o7RmSHkT
qbL0ZA169kdt3viVxDc1oFMN3rgzCMkD6PV4kcBhIYMvHGokHejxUQc5pZFgoufN
JjFgt/IHQCLGTWL+gDi74PhERCWhtuG+TGYqU2O00JJcJL0AmG6YnJ9Fhl+YVfgy
pJKCeuAaY4fpDTBWusPykwh7GksaskXjes037zhHGGddNchT1N03mNpS5Z9PHDEP
xh7++F4AjuKQ94kIKyCbmbJEF4cJih55ofk3RP2LGW2DBl44zfZShqvOERwzxGbF
rqSAI5xrV2yZVo9HcuaePmkYwr3q4Bk32DKYyCuBCST1lfLinJ/Zb1lbjXEoWoDg
vS4+hfnR8DnP+/gwWpE6JOLmU/TLOPZr8zT2jZdED3hWQC/enmSW9TGF1Z0jTbWG
pnYCk+ArcbEt3nUpp2GAwrS2Bp6Vv+FsAQu8JVEEgNcIMSysbHbjUcUUMffl1zfT
r9XGilLr2pdGO/l7qRS25V5FK5eaUOPoTFHiW3LkX1nBaNA0KGq28z8ibRgEEUSp
WmqVUimeOzPxu/x91utt/D/b6sf6nRHK1cgzLXV6XotTxiAx92RA1mBNMzocRY70
ClHYRUJ2HQyDfExWuyaEqFSVc17yXlEZOtfE5bK3l31rHzMpJXrXmorGOt0jxv1J
r189Be/O+JiwpMlbOz9zKs9D8WzH/KV46l0OHoaGTW6ZZc13glUorp5y/UapDozg
kRKo44XmFHPal4z0ik3HYKSkxlko6c4PbWdBXUPV6sSUmr4aT9lxxlQpq//1P1qK
cNf6Q5On/7ZJx9ReevNJNn2K7bOK3E24ufdMFJRe+bD8dGX0vJ7lyh7M/lXEIR/O
/pg4tOECmEqokx/+66bzUiunY6zKYHezmUHsOj6TF/4iS1zYVPD4htXPWfzKMPKt
1pcJOsKR6S89SNO6QS6y9QZbwi6kRPWdpDNYcZSGOh44nhHUSc7xs2RxUwG7mHeP
CRBXUU4Zb6aeCq2VSS3vkbe6ZLu3xd9nViTzbY5dTI7+STgjx6/IvLs3cIg3zx8O
05+i9bJEkv+vTskhcHMkHLhGUU+4hjpBSiNBs3tXdfEg+eEMJNBWJQVh2/v2HYYn
l8zmgHEJW2DeGELJkSEG+DauNK83/aa27Mc8HRJvwbHy9be3rRoo4EMD3Jl5nOzf
ROSxF68AubbF8mFlFnbcx4xUQ34Sl0FgtzZxS6XBuEVAuNfeUdcTsnzWiQxiL5AX
WgpKP2GNbBELBXJc+2jlh5G5AyujbiWNybAH2tqHdj+zWxinHpfO/3h7l8F2HScy
5WCCG2KxHLppD/FDCj8TT0A0etAhNMSRF7jNPj55llIYMAD6d8EAum3Akwjv1zlX
w7NwjRRyhXpc2ZI/b454vTYc6K6cPz3moWApT9F+o6HhJ6Yeywt6TwUPcymG3rU3
ALjacQ0mSKEKiV1Q/3R/il93UYZAv9VGF7JhcQraWaKn2RHTHCo1WmO/ZNnqD8a+
QwITrzgnvVkuRNN1ect6gpnsej5QBtyuhHplRCHq2B6+al6ASQq6jDplEoFGJ+3I
InwyFwwu/NKbXVwaNzVSZmZHWIfKxvw3xYAUPchQIRv9QBR0MtOy14q2nW2POIjh
drcrYyLHreDOe/NZxQdqh7IQFQmicExd7OgC5UxW0+2bSnefA8DADGWXr35klhMH
hxw3+jmCILGKYANr12WKySG3CesDPE8iPpphV+QcUwqSaT4ReIblGdLMzGzPwOm9
0K+zGDmHgUtWkG+Bp4rGGbE1hjUXJ9v9Oxesj+2r+pIpHGrlTUF7gPmGiagg69IJ
NittqnuB3+s+H8Q1eBF3eaFy78dGA84OOEpPtLcxbBmzL5oigasysmx2SOXn3isK
xP2hv7OMkv0X/C88zHCK9oi8iBYQPhQQD/vbl18u+HGTaOTr3mVmOCIUI36X69vN
TqI+FPJZojCAi2NBSew3B4BjZtveNaBlBSEOPVmj5oVdsar9LrrONgScGXLxRqyd
udB8cH9yD0GBK68hY8Se2/WniXRO0hxGiUbrpjLOaGhREO2FZ9/bw8T7B6hsBUjZ
5KdtZGRqN4QlP08IDz6n43we63VgzbuHDnO4zhigyCigt/1w1IcjTZ1GISy/Na2D
p870MiTLYPmqJkT/tcvXLmhMNItilzqA08gS4Lw4d/9t/JfxmGU3R0hKIbesjIXP
C9+PWaSmW56KtQZouaojUa6fq4TtElbnwXjOJNNmTr/pbdrZn6EFaeTZAFkDBpyV
DRjh14JsA0GN4BGGj0ArWZx6fbaVve9fuQyBYsWyBJ/pHK/NQ6N75s/7lA9XS0Vo
A4nVR0pKAxUflk2QCqKqP8qUbeyCg928e+gWj2YSCaYLZ92VSEptD8ALkxe0syY1
t5WWsiEc+Qyv8QMvfbf99x8OpxVG1av0beFbPpF5ZlI4vpbBKhXu5thPN36EI+Tq
KF3phlRbYh99hOKKjkwA+8BMyMvZpJY+PqCutFUc6c7wGDaY5bu/Ntkh2RYd9ccr
Rw/B0/oyjTMFZF5FJbq3ree2Wqi6QDYyFfZ/9YCEf6cTAc3b/+sRTvXjo1kckaXR
79cn5HZo62qTPKGXLR1ksHgztF4eAJ6sd4fFhXcbcpy37LmxEG1KhcMie3m0ATgR
PsMF0T6ZLC4zVw3rIIg5CDd1C88rTJBqlCiiw/DxcBr0pzaQVQDHAMIPDzkipJnI
RODXgplwXQiby1kO4lDLJMTFL6axwyHTnf6TfvQV5ZVaVGDiNDwqS/kRzlsqbb0Y
/crcyMQIUvmKtY2WAQloK9+NxraiYdVPS4MkXfWpmJAbi/UPMGoOK2kgChsxD0kt
yJUJMhF/+COdSDfRDJxFNU/VoplczdUiSDQdj1PGRHQwdfXf/YB0xcZ48hHM7Nxg
wTgFM/54AXwYgLDtvncD1M2Dnfac48p6p3fbYMwg/14aIWcc5WpK/jzsJ+E+/MYS
pBGRhP5KZY4f2r47v42YfN6R1LKpX2BZRwsEO0UwYWYH/U/l7eSKMeWz+Z2ZRMpk
IqIgj0jNmXxP1aUMR9F9eJlIDU9EoZAhLG1oPis8cBUP3MfJboVTGm2LyhS189BQ
GFwHruGBTsZ8wR3NMk71LGqoQZ1ELW3OrHwyaJeTRptBsMuKO7eu6c1DPMWnYVCU
exVnjp/KMaRniHiyDug6Y4uln0X8Y3NiXObdFQelFsdqkgoNP9jRM4fRFNzsQcSx
L4iD2KrkAjR+EmjR3+YsfV+DGueFMC6bm4Lyq3jqDNaI2ECwRyDg2nIbr7tdMzuY
d/eDSoG9vmpjfJgWCytjxki1BGQ0BtXk41x+AztNvLxtT12jcSEHu+YBN+PEmJWd
5Va2CC2cdcUKJzondJwkcQ/vCRyW9LJpPyh7keUUZprGb+iXdMd3V1FR0Iarmxcf
WZYdWdvB/yal3gXQ2OFi1N/1EUKC2B6yYVA/UJGDJ7aLgSBbncrCfZeDwHV1UVad
CuO0BVgXuzTjQZGm1UG4VLlb8/IBPZjYRAJliSU12vEvdHA0A5BufgsDNFreHMUp
BGoU2DlgAJ3bPTWHfRELqvJiuKtlz0KkmwliooqrZ6b/p5af+D5Dr/eW4v1TdiMb
JGkz/tPM67IlvMAQ8787bgsxQgSL2aLCTrcWALOjFlxsVLQuXdAxscxssLcuJ/8N
DQJjVRROFaVZl8XLkKKs6UU271T7vKtoU5gT0Ke+aLCNsYiwHlPrSdPWSa6MgNqC
nSE2lTNeX/XTqOfc98EYNFbkbSXTySd8vxkGY7II56DCYEkiBx9Zs/9kGCDvYUeu
jKR5Mu9IKWpoKYx6hwXJHF9dTj64NCQq8qIh/HAKiycCTBggikZDA/c3zz8W4u/F
D2leEfPRM1dLG0gUHb6UipUbGKaJfmnmnOtiM4iYo0ILf9GlzgHhQHirf3SJDeiY
yjB6w3irA+Y+OYFw0XcgW/cfE6eZLVcg9NuSu8Hd/uZqR+tJ2YOztRKPNyO9KzBI
1wLJDM4zjUGwyMeslY3mR6zvy9Ee2R1+qnRphOLavllum55EPw749YcHxR489x18
WoXIwmBZD19NLoKqms4cB/uGvywZuPg9k47sEyqpCmhFvRs439fwXIMCe5NraSGB
dadtoRG3a2gmQ2LK5mPjkWJLLRATps6zqfa8fEXsC2meVUTqkRXhNjDAt11/kHoZ
6P+epGJC6pSI7eyvpeHYQEyh/e7bRHk+mtnpV7mSQka9kLtgx0g24QVFx4rb7a0C
MnYD1IZ+fSjuQqSHYLkaklcTvJxcTk9ciF6qv/Oo4eA0ykyrkmwXKXpzTGuaUu6N
Nv+50dzUIFXlzAVDwdtD98WhBcn7sVWGhft4PgvJrJALYRB2mR/3CukfRxcu723B
Hatzq6OHmu06KkRiPRFpiv39EpyxjgRpnnOlbwmvDCRF8MCUMYBLHTvEsjtF6Qbt
YVuqGNbtEyFuGsHF8801DfDPuILvmck7aXJniT2Y9szcIZe5eDzzJn+4mzRiagV9
Q3H/R0CZxKi3BvRsuGnvguBGrBn4e6wplCPA64uNSBlkngs65w8ny2atZ0Qg8JSh
HOCYKrP8YzCkwBZner0CF/PR3dWtXtqJt4jvevX0e5xoBFkI48PZbyc47mEqDmZQ
L8XK28e/PC/3PHEC6efRtb3ZQbvJQUNKft0LTUK0P2VnrAvUd1ssBf+I3r4+w/uF
jk5uhM0BZ610ROijGt59NxfI2LaQm3bEBvlwm8glQwbnJf9rcE1/G9pcJepzlAwW
HGSJlU2c9TukyM7dXHNKQlFIGeeP8j2r+/Ux4H/Tt5HsjGFqhZHQtYtajxFv4Mwb
NwbqeDzFQoly4Zcfmw8QtKuTihC3xL8h6FkK4Rj0i3GeidCfPJXHDEmgGj8Pzcbd
pecQJbSa7faOVOf0dZmwFj7542Z8DRoI2BpPghnx501uII9VNMwRe4mhlM8M+mXI
IVvLzSDEkCeaDWthimTTrPCb04ypC/b8WGiy458n7N0ZHMCUJyyEgtd08pwneMy2
gkSYYehcLCfya5zBxBYt+88gUmYWwosRAWY9YBaHa2EgI3eMIawAghFfqbOuauSC
18210HDhfJGikRZMFuHjz6PSdVmzCd1k4Yzf4wkI8jjVnYMXhL+vsb8LrMQc/6Om
kaPQmkxvn4gzaRhIGr71z3lWlDBboskLOIaz7Qp5fuilCh260fu7G3mJDqBEI7uO
FR2x0s4FoCn/7iA735jjSIpJ2U856O5HZTYhwqNz0o3jdEcjHsJiUr8xsPWc19h9
K52ZKqiPyu/Lz9ib13yQcFlwdeRJ6Y7EVkMD+/DArK1SwB432zjcC7zqtR3kFm5e
kxk2nx1/0PTZxavyay6GzvRLvF+ZLKyjK083qP52y7OwwkBzEqmuX+KdbZbCGHgJ
v7uJnRL0P5sbH5l2YdGIuNwtWdYnzIBgHZLpwiDmOWgHLG5EZLOkRCRmCrlAne6S
8DePnp6kExn/kPUo7B9J/Q4sWG8QQT4TIRrPRt/MKlodURicG+L7DPFOksqBrPB4
wSgXOQ+ysvtTTNYupWlJlJykYbPel06Fii+wMZGEeZDoOgrFL1YW2pUOTaeWTUmA
YGccCtrbL5xtGfsCahZFzh86hSGS+IQgSxPLL1pbnBotzm5T1TUDlPJVkmFDrc0T
te+osHGJgzFC+IYRUVOBR5cGKO3bsPVannsPNYgQ7X1KLFsYgm9niq9LAcGkXmvt
+R4N2thul/EL/RRM+ocy9n/4AciSbUawwChOlhSH+WRIX8HUTrxUYRfNl/wj7BUu
BdJDquublNlLwtxz0/EJ+zrKQZw9IAM46q0EO3gY/bN6Y0xvjhkAmsF9vXxFOkL4
t93DOOe64Pdjhce8/Tud8oPGlN43CiPO7KQ1P9HcujgBb7pWebqnkzwVy5G7uNsF
kcofTn6V6sEynRAvKZikrOcUZKT6wqRURQGxT2UCFZoh3ZX1060alRbT5MK+4/gO
cZnv1YSR8a7pruuAhw62rH/aU0KvbcB0KJq+ACRCW6kPOP1q9l1L46CPpFkS6Jdz
bmnn5w5XwWdt1M96HrrlMjh/QI+cfaTxUDSmBSrxLEI+QJZ9Ydm7toCsJv8mtWka
1i0xPnRvYVkZqsgxUOQ0LkaNsxGDpBKeDm//N4VK9Fln7JHuXkGNncdiaaXs7Hs9
DiGY0rBk6QEa7upsc8VM1fKIMLu4ebdR6olvujY46BvVCV+zqEqyoTonrSa/HRcP
GZ71oF5u9264UQYvYgKHP+V/pV83cBROIGR0yhIV6cp7iX0iUqKefW/DcAKIvDBf
a4edyo6Lin68ZIy73jJ2zrkidxfpsDM03b3gFc+QteVTCga/lxZ1QYa+59XVixPB
wSlzhCBRLBF3rYcnrXHDgqKaBULMWsXam9a7LTsJI5/5HsNH3nIQtRzlU9DRKL6Y
NBuq/Ye2tnWrjOTcA81q7N5z8jb4Z5rppreHyqX6kGMWfHY6dZwBucB/tuvXPCWX
ZyU3MTORd1khZRQdwXhELzjrx8DbxK+ZOSKUFGzMJTsfuIKWJNfkTalSk8Bo8bns
ya5iLkLGKpaniCC7+ryCEA807bZOTDG7R6sE3524luwn9ltLbl/EZeGsRQMU6Z9m
tRGeHTFIU8NTczQwZxo2BfvhsrpWuF3xhOu+xHOs436ACRIPFFHmVimSIMtL/F6p
Xey49cyVEebTBY5kHdmT3Amh9+dtbfA5d7jYHfQQkrIlp3DffptsI1sd8r1JONQX
A1ZiKQKiX2HjIg7lQkbN70WzgFifXVAGgLZRiqrwmwjgrErbr7dxobugAMGbrA+D
XLA6RnCdcqH2k+F3c6Q0sqk68MpKyupeoEGFhBxeBua0dxOl1bf3mli8X7IF/9k3
GGwzwVm+ltKLrAe23clESgAA/wjaHHooCHVpPodGFIR+E9UFGuTBAo4TtfCwdCiO
hS8ci+Mw+qDw9a4LuoZIWWnt5zD7XBaTP5DfOPAqb2QedpGdrQDx8hE+KdZQMCjk
59dyizWkwKc7sJYkuZDLfkt10NkD2IiSPmiw7KIZMWJIrSitvYKbLWkxoo/dmUWY
B/vEVS6l/2aSbnNzCQSSvCBJaXh0WEIQaD/RNGv4Mi5TG5nwawwA/68ytTDkUXt/
q71uoIc1TIn3P3AF1pw4F4R4te0XhAWHammqZTdTDLtkMuIumCru1ByqWQ/qZmDM
YTOKIbRC58ompG7gyh18NyQkSseg+yEwlDgRBL8Igv+zTUbDFVAt9Jf2NKlyac1a
YwTwFirH96iR65CQhbvZ9hnSTxHZxwpqMvDAvqX48IZGEuq7o0KGIYAzQxE2F0Ug
xzy4q/jWhg85pg1hE0o2UWM4I4gdCwf8CA3SUbvlHJqD2NBQpmGSxhxgOTpACfMG
9UXYmKRxsjLA2oPyiFf3dSWLLofV5PmV3wCd3Yk1r4hMKku3v1NTflj7YtKdnKqU
Cws0nciwgN/tQlPOiGvWQ2ZfRrh36yPeBfonNDp12aqJ9bEjqx1ff1JSZpcYhtN7
EZfi+PrAIfFFjzjcM8aPQkgoY6UIvzRnMR2Qh7RBD/eKgeUs9gi4UH8vE0cHWEIE
qaw9fdjf7Fd+a1lVgfXkTvb1Rf1QA+vXFNX1b6a+wYAFdLcXYStrgDjnIsY1XW5b
Od4L4/PZ+UipPkLO0/7z3txpEYhf+SbyGgYOI1HYsi+t1Eu6LI1nNltGtbK/byBY
DyhHhBYBX+f45Zf4iMtE1x/71vEKmwCx1uQZZuyzZOr64jsQWUgRO4exqcYKWbwV
buEtrpN1KTiXlsTlz45tDzeStChwCFj9bf2HW9TjY8oGMgGwJMAoXcfcjHU0W+3X
amG8HM3mnr0NE99MTFQOgmKWVUgszoBSMzErqcMAnnjvJYVJwjcgjFhNa1lba8Se
LONCvw+CG+AVvja/7Z4T4bvq43wdNwIjiCZxe2D9BeaIWLRzHpdczFFf3tPduust
d+LU02UfA/FnH8hxYim0Hsf1HAPGgMf14fLErWaniqHS8AyrY+3RcYupYe1H6xUw
qlt7iEmw5Z7K8ZOrbevgIRBAPtBCYvS3asGgi7mfxnkTbNnmuq86OGtmgxOiEtWo
nLCivwFr5+zhDWumUHvOlYOz1gzeRJ1RA/iby+J3aly6ScQrCAhUJ1YWBG1bz2xn
dXSMa1CwICARo0Y8PhBxsQFmArjfpYLWWI+SvKI3LEVUBtao7UEr4JentbRbZa9L
GKUkbacCZ8v4JEI1Qx35/j/XzYxTd4i3GTCerVeRHErBIqE+IoexnJXajcoWAF/H
17UbQOdz5vavKGq0vbw+hyBVj2TrFLGwLYAzdLS9jG/SAxVdaVn2JqIhm4eAZjFB
3JCTMDhIEsj6QHCBUDW83R67wL+x3K5hywGKRrVsLy060Dtk1mXywEzF+didSHLH
S0BCmTw79JnSoySwgG6d+tcgvAVIVN9VN+3cIDXsO6G3oZrdnm2AiMgT6JQhKs/Z
eouNoYMRrLVenmjNaWppKLQKXSmPuclBGX6+Is/B5jKVRoiAXtrSjjxxoiux5HS/
8v/t+TTpgrAiNQrVpQuP4dX0FNxzAoiUw6jxcbFSNiIl1ViGrm7bwpoPl4xkdtSX
fD3CpmrbvAhb48teSDT7iaOvnyhycduZ+3hv6WkgLm+8MLP5fOfZtodm56BVBZHz
7sQA6IReRC4Ee6rmjKID96k0UITThQufnyZSFv2JuDYyrbQqGgEm625J30pFIkIF
8fNbTbEmzB4uVhy4J5RfX+cLjIDTGUXtzkDx7f/YZ0GPJr4IfypVsqeKPsPeFwri
NIlQW7Fil9hSyclrTWu0dwyAWQPsUWzfuCoGCQpqtlj6jH+eZSFF+xco+Q9G3kIe
HazATqYe16sQZa3ts5KHqOH1TCvpy4iBmu+V3XV1oz10J57VtJIFRFbbS/Rg05QY
AFM4i7xmAQEyzc8FmyR3bQe/jd4N3wXXC/R4SJHYMzjEiDoaoROsJr+dRlmfn9wy
qBmbPF08WGkHE4rbjKk9zq909MClSnDnBMjjIIY9yaViojjk7Z0sCaei+wciDzKV
KPzqwgayRGRBG2JM4snx/gHyCj/VuClZk0dG9Pf/ZLEE81GEzFCzIKw8XqYC1yQy
FDzWRtDabrNI6axfmnwaXnjRH6Vg2dOfe5hGQLupWK3eBLeWJOFdDBZHyv9EfJvP
Ta3rNCAir0TdAbIyq5Yz2ITXM7JWkJa87JaoQgazhDqnZGdk2UuKOcTiLh/ITjSJ
LEl+lyF+FPNwtLXajSVmCHggxa+UR1rUJP4zWaUGDF/T5CP/pYUyx8+/taTNsXnu
OdsfYdG2eAn2R+xuilwOpzFqXHciw9ctwntZ2YNcDDioGoLM7QILl0u3cL+NNHfs
2/2zNjWdTg/G5pu7HDnb79Ua+mZ6/grRcEw3SrU0Shb5cbNkzcqxi831raOy2xrl
qcGWCw8RTGc3N88ehqi0B18pmb3G8LJkhEn2NFE1gSTTHbuV3CpPfPfajWXpiGHd
PAAzzmbPgV2LNyrgzdq0V1vXas6QaIljJQrDgsvIh3hMQLmL52aK2oqL+tdRfVp0
tk2V/SNbHCQbuM+3Z2SfQviwCJUTTkSzhwvnTN3qM0F/0iDGNpiA2+lgbvbmjPz7
wXOF4jiOWOllTlGy4baMb+Gx0QYSGRZQ1UMdIfcWqCs+79/LCoO6kufVgsNQRlIl
hHpiBmoEgiglWufHOmLlq8bz2/83L2leT8O20NzyNp/0oxT1gMMA0x2xvRRAr8Gp
Knh7DPJvOKh2U5vMOzpJHLCnrzEL9aKN1xDxeZX9u0xBHvBjgoEnrMQtyD/oxgOU
3O8PEiQx2/WNuHuDZZQhFP58/+fQer6yiBuVGd/NGCq0J6hqaz7TG/Kn+sIQRLJa
s/KYi9fJzB5mfhd+grInxPJDYAdW3MtumK3EIUn3dZgvzukiII/S+/RfBNBj5NLX
vulEOjdPX0mydGBryT3rZ/ecAvKVWB8Vz+/6bXuO/yJ/oElQwXYd/WLlLTjSr+qU
If1v64Sd8MbRrVgkiPpWo6EYdinDz6GhsXhztA1SGmEDW2QEX9TN1Q6HTPhGiqWp
Cv297q2NQECudCPe2efvmoc2J6uLsye3EMFN8Y4dKfT5P9vBvml1wnehNCeqz/a6
2in9ipvHL9rFJoQdHGX/V9mxYyK165mY82Q4yVYBfKbMVrt+3VUTkStGJKgf6ozB
uCjKhDhjCKdAdLHPEfuigXfIMJ3YdL+krlFjRwCJYI2CFyi6URB0iPcrXYW/illj
zpQPn7P8Wn18clYzfg91oOaQmqAbJT70GLROw29T/xRYCBxwLkaC4EkqVcs+Tqvq
DnPyaQR/gfEq5y6CfkHMBowmUgJFQnWhto5o//xa4wLedanYHzKeKZci8/S4X5bI
MXvni7swf2aNLfrt+ONjpaRwCyou48OcYvn6PJjuhKOViDJEvEoBGVybmdjorP0g
OoUHeJfG97p4mRBxjuk6NeYTw9bHAaJUFrNERYSrqPbvq5EWYenYocitqE+0eoji
OxzjgnWvHkkyIDTnsDUo4np2BwrWiObAvHMK07mdLIXmZd77w/jNiBveJSfm/a1c
7uibV5nFjd6qoUQ6lkFcvY4FQW65CDw4xMlzXGEiGglwM8f9rcpdsiXjv1xYkoAa
Zek0yPWlYrLQqwSpVtMG0XZKx6OYsCQTmuH+SNnNZjMNl1Nh3h0gPfBVaf2H9H/3
9ha1HPfz++s969lQ7njmZyZIZWAf9JAxTW93cMG1t6ptQMUJV5xCfXYSVw8zLD9n
Itv6uHhJCRREKTXoS/Qm8Z6jtUlKuQ5nm22BHHCArqnMSA80pmO3K3fpfMPOPT0m
ikWTXOtLKmwWJW8y4O9H1UBxIW5Zl3RcR8WC+6ak7eWPzcx+Md38oYEfV7/MMHlF
/57nOXa+s/n31eWvy69m/vo34q46y5m0wjY/X4KHwu4KiAMawOZJe7/Lhc1442eW
kb3nCm0lVxqgISK/HJJ83I9sVgjyyRcRkx5XWiMQhM3dBskZfHADxoihRRbdl86f
DfXImld4zBVtCGz2BL9iLv9yaL5Yiji2A1sj/rwwFK+hygkcEbkdGhThxC1cS0QE
tQmiBJCwvurjwe3Yd+Y2YN70QrkbwSVDa1WxE9lywQzYY+CXNfsXLkexdk/pvCxS
Jnps6IfFjOZvqj0J2JCOvVJZzPhwIfc3D635ZgdGQXaITVXAR1ple8oOmXxjtJq8
cOlKLBKT5IMePFtCMvXHVqoXe/dzsLqLp/QVvr5KqaJTaKOE4K32T2Bkpjk3G7WK
+jes6RfC4rWAhRs1GiDHmqGm/KL3qcvO34W2iqN1vQp3v86bbtEideb0Wr3ROig9
jiDo1DBOZycyDV+dez5AP39aQOOmWx1NaL67NeVHfksLvQ7v7QJAX3fxbO3Ksrwr
DHJEH46eDSySEtTVhGH20AN5CWzAwploaGbhYJmarNAKLZqJE/Kp9jXDGHDEV9nT
vDjt0jrWjHgI5GLe9JDETCdT0f+cLBzhuOxqzjWv3j7VRzkFNW36iFVA66OW1Uir
xKsFbseTnONgfoxlQCAdx3Aa0jV7TKZsvrCSIXfwODoPpS0bODKw6xF5tjqGo60e
YT3OEZuXBItaUjDh1xc2LIgOe9nMC8fNth0lMPy0co7WJ/uUnBPGtatMjW4wpwDI
idLfSeB+80QKPnyNrxr/wN03e7DuhPPZeTulwtKqFSuDbUX7v13et8tSI53uCDG5
zTlK9GVTFicUdH7HZCsJARFnQ8xbUZrlOgVjhIG3gJMvb4FWV4ml3Qj7Uc3C/Ys5
WavzyxuRcax1Sy7UkpRa/SRivq8SC7gM6m/FVmY1+L+d/Zv7noHTqwDzH3Nec3k8
1qs7aVB4i2yD2GP836bGeEGK2/S1uqnWUFRMJpwNTCIe4c6KAaJD734an18BZki5
/1O2KlfV0+HpGdhoQdCkeFz117v+fgPdxa6FRQLBUFczwpGhi+hp3EWcCDmx5Ut+
m3lLDRx1d/NbFHXFPDYBgioqioHR84v7ABZVpVXR8Tx1YHVXqxMkh14qCNGs2oPr
uD6a6aSYHld1Qz0V12AIJ+vQed/UkBVdXUef2DdUbRxaMyPq9754g7LiEgE85HpC
pSDNkjs7BT1LxbO0B2Z0phd24K8WLoxKBkuEs5yOnmhRGcdPpW07r/RsWWcH4UlX
pI6ufic1CiFacRgkG409ICbPjAkSAvYTJ6HBaDOn1lVPTjPo7klBR9Pl5/NclLnK
ksD8zYHqGZGEAN1XVsy7uYq8w4LOtm61O0mU5SbpQIlpQJPNe57NVS7HZ9ceF4xE
j1oqSVu2cFju0wec26gf2o7gsrHKgRKDZaJ9JUU3XeHDlpUZPNSkCg98w6Vvkt9C
3D7V6ojbHnDh/c3mygqs/wXgWqsGO6umCHyLjEPrRQdoL6vBkQ0CoP5WQCDOJFSl
5TlcD17xkDvViG61jWaBWJtCITEn508sls3kE5bLI0HXBCKqyKuHBtMveVuOvIpv
z6e3Og0oCUQhQr7119MMYAxupM20XRRfcFU41UCmjQC9OV8zzoxXy52Tw5ltQPmi
kW4gMhIw/FLluFAd/ZEYl7A3XYy5jEmEH0KJgRU7/x8whayfLUipsySNC9UT30aj
KbL9tJD8RNLDMtuRCejMSdSpwpIXm5eCLRglqtoJ3hzC5sN9Zs4wc6tPs+k4L3zl
63JQ7JaJ8qbwPWh9VOr7Az+1rhvVKd32qE4aZ49R4VXoM89dY7ean/53gP2paThR
JO6ydQWhqLuNPKeuoX8MvW4Er0h6mETpkiRooz86YKwjtMNs0Jms9NEWaT007F49
SwkfJJ9pwv6olQSMleXIUqwi3qUyl1NOEF2EK0FTtMpOEw7a7TNOMDNhWzDzn3Lf
+xJqsZjxQ+wqfZpceLnS5oc/XLGUP0idNG8nopCdAQCo9AY0e8gU5JE2Hl1mjKCz
bzWaws/nFHN2p2GsVB24Kr8GSxxyQObfCWiKc8kw2ARrnLtTHdgQZF4WgeJF2rCP
zIlqdLSceZqLSHKeeKb6sNYJT/LdHQBRjJhbjwSwu8EA+eTGLJDNkjnXMRXUda0Y
4mK6di8b/rNBpQE7MHv3KDdqwEEPdJ7bJi3ThQVfgPhGNK2uiJCu99aDv7Mzhcjc
KsPyz+LmyQ+Ncx02p4m6v+QZskEXxcQO/U/jcRSB1mCnVnPh6jZSlIntHVpcn3Ns
SMeqtVOccZx+eiamavtqMU6Ox19N+jDSX11RQgGP+GrsMijo/cpccrd0C/SaccVz
7mZ2+kl02QrmjYPkI/Rx3sYWd5hpedJcPGfs6vfMdbdPZL6S0PBvzlcS/niMhddj
lI5IbEWYIYTJqlgDoFqW2syGoGWr/oXsZiXBPNbUMLYtWn9I9cAXesW1BnFN7xk0
O54pm/h5xUDadONrsqb+k1W4VvL6oViUoudf15rSkNNDXFr2MNKL8XqdKYjkQYNI
yWvyucs789lWtflipDaivgNxmXttLHEx8C8uGEiAXvmKMgWnmxl4hPZPPKRW/x+G
Y9uoUVHdDrvglRuafE4t4Nlx4p+ZvKH8oyx6Y3W2X0FAA8275WXhEaSCRVzNnLwj
pRyKh2czqBGHiWpMh2+zB8wxrrgHaXrOEgKkRG6EINTB6lFXVuDzk76KcgkqUN1i
1+fMt66HZpnqHO4clYdzzQ5fdJRmGUUfcDunhBRR8Z4bF2n53E9HHixdApys8/di
/kjamaai32WjQpzgDqMqf+JWBnrEwZiLdVALCXczxv3xU6yra0URjR3cbMH/FzOB
JcNwc1vVqvWTVcLeTos+E1oX9xjy72BOjZtEzkVwK/N2vnWOO4jo3kQBGUssTPvG
V1YpC5C8ngNM3fgucYSVwe8D+pJdpYHvke1OTvTXadE/LX/48ZVOClVQ6na/o5Gw
kNHPdlphlMKnTxZXEH2gWws5YNz8Dbh7QKuwiXiCPIUw11e43rw0JVuQaPgIwylI
CNWtv4dQd/cV6qvCt7pj1cpu2kN1uJsj7zTbk9iYLvhA6IVOKnva0I6N7OMFih+o
7fwNVWZl5DYQ/1lg8eUZPySKvihZNUF5LibV6kCVCrCjVsU09ZyJYxpccnkorF3j
HbtqDQiAT0u6Ye35WrqJpmynmIMa6uHdrq3F0xNomEANgyWdo9z9uxuZijLTvqLw
d2kHGSbojRMvDSm/hOhZ7Ugn6jER6IVnXnFCgN2lXjK9FzJLRxkiOgOPLUCegY22
+4b+M0kCNgQFfGRYYyAvFLpihO1E/UJipsBzWn3vXg06If5OxTjNXAefRuu40Lgr
1pGqZm2qperf2F9AHHAsdZNS5GGAkp50sjdJ9nasrMWFrqBtWE+n/GphjtfX239N
7EGkboCnzZ39TtWR2ECnVPg+r1Q4x67oQPZJwoVA4grSW1BJf8eI0bpAZsVdvfr4
4WvFiMjlWpsGBHJY7ZC6npHJkgTEhbMiG7T+pgxH3igCvNCMiS1gpo3mspN21aHg
XThlboznGp8T3LKnva9iY8KRoLeONrsOfFq4FMGSVVA7Toa27D0C5GoV2KKl1f/i
EPsv7+JQj5ODRuHoq2HqVsED5vQEA6bbhSs8bZm5IiXIGbkajWxZKRfEEDHJrrEy
aCqD+qu6vRlSkxQUaeLyLNFCs2EZBPrGFwdLuofUZri/RXtpgK1LxfNLgRCAsTtC
+7Yj2V6KwO0R17EpLszfSK6HbjUIoHUdDra5KKuATAUm/fakd7ZmT32bsYZD6i7F
6GhseCFqH20kOW7gE+tysMGiltUCkyVo0BVDtYO6GnjmTojL2um/ct1ypecmEnGJ
l1FbqtXGUTe7uR85vH3b0bMIQM5p5tQ2emqNu5EUzgUgr1tvegfxHLSKeDlSCMSi
RNDw4JlzROhrIJ6yBqP15AhDDlNQq+OJBf6xBA9IC5tpto2NQFR5AreDRgnERHyQ
DmGWfZf+avNTTbgNWc+ZiaInqS2bzIxXrbvPdfDboFd+uqkUN/nZ+2+0/Iur+xiK
+1NKjYC5qn2RO/CNddy8/caEUN5qRtzRbWUU0aLB2RKpfX0yQ3Kygq+yThGWC1ce
uEB0w9v1rqK0k20WlGmEAwNpLfe5PKplptDjjlr1pyXkazA6gp7WIVeLADMyJIO4
99cz2N0eVixqEj4n6S6eMC4mGnnpV3Zd3UijteBjuCWwuDYmx1N5W9Bj/EVVv7eF
MvI8ixZR3F8F7EXTDK8WXTgLY+VbVVB2TGSfH1hFL2hZ/pu3fQujF4SjU57Of3yF
LaNdnGBPtqq5WWbUFqQfDK1Dcuwecwf6HPLf4clcvkbQKEXBeUywe+Rq5Ed6GKnI
stVAiOyhYw2aKWsWOvn6zHAOa8tfdsUJIufE3+dUHz8C6kzKJCyozP2iP7Yupuw1
eNWqoDdaErNYbdxBMea8i28FH437Hu70Q3IyesL1a5W0Ptkh/aWDEWAU7LPbryOM
//PBZHmJMNyEiKseslArpkSCZL0OMwxbn8u1APpY19eSNSASdNpI0K5EKVewq/CB
dCelGjd4nXa2l3Bpqw2l/j3HpF7wrpX3m5AeKXrifthY1l90Y3l8PwFUHIVQvPQ0
L34gJhVdG054nm11SzjXvc5RtB5QxRNPLWB2j1uYhn06l1bAmdhZK0CUJPeEMqHQ
g56R0eo5B9C0SQQ9J3kxtvGkwvBqeil+hdr2XvBMEUfC5hpB6qPYYrJc7yIESt9R
hLPYNLOKF6IVrfzf0t0ARZ+Sja72XZNCPLZ9t4as1A1zU8tcVsDKUT9KeeUWWov/
pTKpPcmuPl1LbX34w6IgNDP1vluUkp2WeHv397sxET7WEIbkcjtAy96K1uBgMMLN
jV5ocqUIQz5ttgPBlyn6DZuJLasEPgQyeKtEWN3ZQOFAyl+QY8OdlHJSaXVVjEKK
W9ixxLR+R39dyztcn6pa+jzsWkdNrPaBY416ZEu9RspOmZX8Ezsv6hPZySuUUpoQ
xdasRhdjWuiG8CfjgwqOu1bw6iR3NEfEdLLd5srPpgSpGfQez4vO510fjkDYf4PO
p8OnTaB7Aqmxhds2RGyHfDSUSk4/TZFDEzsU0dgYSbPeO/2HAaV1whRsbnGcbot0
1DG6NYdZkjJeBfqCL27ixB1DJGt/nMTUo1487EwNyFsi3Cf72kjwcd1BZPR2jowg
okwdKKqjb+ddIsElyoRpv4trA239nhsWQecT8G/3dTEz9aFD778G54RbAX9GN9bR
kffQCPyfBCxsxlsZxPpS2cs3LcP3KQYAPJ8+n8iqh8jg/MVkRpa33MvDCSxF0bKz
6mhfs+yWozu1cSmw83i826f7CQqyE3UtRDeBWU/jv9jEpgpehsw8iTrtFHHJqRoD
Qo5L3fVBIk+Jrkz8G4xwciBIW5dXsHaJFmgmZHLMZAKceJ59PNYU0LODC5VKtf+T
LJ4qbcyRHIHPOo4QUNh/rlrAJ4IaQweHfsgYj7Aat9WbokodqnXPrzcAF7q7sPGV
muYBCksKllE3/dLLG8NkdOR5Q+jNnwywmWkfmqJWB/rBApzutsXu8UAV6d1Hx4UY
530L4zBXQ2sfZrUMtxGdh1UlIalkEfb//8XaZ7vWxhos3td5KvGVSltAneJg6nKK
brxUKbBJqKVra9diwNzBMgj1XM1S16hzSxG7wzqsnm0XVGXt46BwIwtIFOCQ6gmU
GmrXmhK2UGuGd3GGStZ6ShsmZs4MQBsGzfpQtyCCpjNRBBwo07EqE16CAGDv/9j7
p77m/qGJ9mYyzFRB5A/FlgLaWdmL22sPH6PmLuJKVKTmD2pCeOevhmcDfN3UeR6j
BdDKG4Qy1Vp9UAsj2XZxCCGOhTL00VSgUyNDfxSXXXzWaqg6DMcU8DKmCD0hr801
3e3i+zpbouogoGQveVRy/hApD5coMzu7+TQQLZ9+V1YxJ1k8QhNZB+bvy3I+4l/1
SfLbQCuen6aw2gU927+nn12r88VtGN0UckmuKRb7VxuB/yr5g26nCKJNL0OicbFY
J/ZdAbZ0QUduk+DUoPgmueXEiyDaJV3scIdQSdmRqYpM4DOO46cH5p8MgXad9j4u
sgtRnpME1X3CkNXu0X8saDEeKdt7THV/RUadRw+tetm0ShEPEE+c4MGssSYB1u7a
AMxMgXGm8NReoRaV+0t7l9uQ6i18dSHm++GfZaQu9aIQ2WvS5gDjvMN+dd+xcMFo
XwKdVeErUAupB2lskyxIeeL5SRVTnI9ZtQIHXTfHN58OQK31Dp7+P/hRMD2zwZsq
+HQistpUkIjoAQVoAqx4rgXMC4xs37Fl+AfyQGxZp5JhGf51RqsxSCegklBKDstq
tXVZqIqke35nRP91MFZ8RdJQbklmNE2cjxPPwz0l3sPn8AcSnki8Rv3mRdypo9FU
xliyXoYSFe17l5Cw12GuxSHSzQ/KOwuOBne+OdtfRuDpsfa34YfzaKtFb5ACTj0l
ol3+QC0nG22p64nzJCNyun96ySuFrGK3yOVKe+kiA8rM9MPrcFsWe4HQnYzyg7b2
M6K+Vnyp8SncN1YdQ1Sh3pv1q++/ZMTqo93gQHYHQEKk3M6b6bJWUH84X2dG0gPr
m02qkQ7BH7NPSXhSsI/Gt9ylsrg3ort0MhQUP6aubMeTvRYSeKPH+mqqYoFT62c9
QBND1wo4a3iw2k2sFVWViUxs4M/RZMXu/SW6MICU/4iQtCWi7VY//V/DJghvE9F9
f2Iez28jGASW4f/Wt9E0ACjl9DMKpnyJJDqOgArkDdrnYoPXcejRb3xTToTjqmxG
rM9AnsFwsAII9ETKkQBkQIrSp6MqZFMmo9WPElVtGZLiyK55zzCWw4lEXigWxMSN
dr4VXcI1Z9A181t+pF7ePwS+HZX11BXUlcDN2HMXYsibRF5B4DDMFeLgPoDMH/gK
AunC9UFbkVVchh9xkIDuy5ueh6TQGCyxl1eiOpEEM0X3iHr5E6zseXTnD9bhHP4L
3M/yYQvqYeVqat/0XLuwKQQO+uN4eGfbz15sNCHg6sG56dc1GIu5a7nWAo6NdmZE
OT7OOyLGKaBi52532EZlorwO5xbC/wUv7RRbmu4PEhOqoSFA4PEk5eS2/cu7pb0L
0zQQkb0VI76WvEsxGLCeiOg2vGlH2g2MfTp/aeBRibszyB58XgtOsCriQjSMr38M
ty9y3J7unI3YAonnMZgVh/0IA+EkF3uEGfovtZZxOi2W4nKGZ/p+EzwTPoclqrCc
vnduGIWcGngtkkewrrnyhKyo/h+A7fVpVaeYYuepiiEnnmob4Pqj/kBIBBqN72NX
3oDjDqPRq3amWoWLpvYkuL4/aM0sfa2mQeGh+gVdCvnUpOUzfMSw2DFo8B4AHfwm
kiMR+BFUCfTHvW2Xs4aFajkcTYUaYUMBgpNVK9QZWaRaNeq5JNpHARMt4N0hEEb3
sn8lDyJqgAijuPQnQBqDhTbEmoLeI1SGHvPH2rAuVmOe/RFeXDV2LHvENeDSZeIr
+cR5uHgsVAUDw4cszgMsdV3iXFDDZj3Ex+46PesTyEicm/ihCjdvz+syWIGbbSGX
BdpYtthA8AgkB1xfNUcMAiJ/D9c+w6pH5HkFG0CBMNYwcThGFLRD2QGCUqqCYIVa
BuaXUQkEP6oApjDaMlj54QeAl9OiNiqHJ9ZP0wTS5BKdvV269ZvH+PhHnYfNuJgj
4MMDWurUYDD2GdEQQ/w72kL4uhclokuo2zFoH7lIb/m9AyRVKJDZFoVUp50qYLy8
2uhPMJTxvK3v/M79hAIhiSytLGd1rQkFcl9MulG9C32xDOVbgLDudh5SNX6ip43k
LBDdenCm5XYJ0reNp0M1nPQ9eOnL/1ta9tFaUv5pVummS0i8CgZabnCCmDoQzRi3
9GK2dVW8TCzu6DzKQQ1K7vZWM/m8w8ZV3dabasCgUM5H6HpdJMFiZGizhR+aKHyg
asfYxdqZhvQhEQyskW+3NrhupGWEQJ0/KZ6yiyeDuMyUBZYdMy0o7XxhmLSHdnT4
edOQX9PllB1S9OQc7CqGEVIEJIV3kJnwsHdz3/SlMs6247wv/V/igiWmj/dbRP3O
WtIj+XNAHB4aygRu5bNbG1ru7439UzSb8Bg9+oTjxDxds9E5J+3PM/mnkisUZPDw
o4dRGR4F1XknZEWy+OrCt4x8U7QdPsnIvp3HfeGpsr7NOUCKrdEQq161LosL/Dbt
Vqc2WRvsCpciCoov4zDUjN32+r4Cm+KPofsuauvf2pIXjvPEjILvBaDfSjTrCBUB
a5unKpCy0HFBVhNaP+oCFPSnVZdYrmTXGACJwg4+maY8B5lTaBCPcYzYZTjTgocA
95RzprzjERyMN+fx5dGXOpprPwP4H6OUm2fC1xNSD4FeziO9qhJPLdbcduBVbFmo
Y4Wa/saxvJqfghaKmI+gbWtKhnrp/pKcwWufyz+hAS11nShxbotlTmf/cep1TIXZ
UrJNu8nShgOfoaUOWaOe7qWGmuyRpVaW6xEk35a1zSxx+P7EbQygJRDCuYyC/JoN
//QnnwWxTe4F83EeRLKMttxbnMWngEcR5BEDdt62oSWA+i2/ruP763/mQNG+VNTl
+ezx+GNXTA8C1IKoc4lhb6ytDaVQHhyC7Fo363fXADUvvgeIjGGWZYfU6EgSw5EP
lXhuSl9rYUghdIJqahBHETV3sbCw48q4w//ZfRSpoWNQoF6SQ/pQKLI5iRAXWHjy
3OsRUBdAJOizMYRejgRklwanfzzope3cmNavExTD4PkRqDVSfexp+dkvmJ/KB+RV
AQN2E8/t+FrrtpzooHsVuq1SS3g+QDhc2CuAGipTR+TQj5l3efHN00nN2WFWPv6o
4ytRVaqG5afcn8cqv/p8Cuz0G8UBDUhfP+eOTxacJ5PGzDKU11PZYMCDsEDQHQRT
4Q0roBYIIvelAmXtD02Ne8jCwaZD4ODfn2r3yW9FlZfbdtBrALYylE/Ii7BDVEOs
a9rSprIkoV9uVmsM8lOpjDrFXBdvgnLd62aTukJoRcVNjnzLh3uzsdPhCo4mcXLC
BPsiJHmDM2teK0kNFILusM0cYVcw2e006bnxHDdB7QO2Rh1IktAP+VoBw2S+TrbA
E1X71X7nCVqKgzd+gntW16hUL1CIXYozXVtg3rXN5t4SxWiILfXsm0QStfbP/gzg
v5Qzu4MoTFUC3z/N6qJtDRPm13qhuhHM9m+5MUR7qrWC9FdxkwU07p0tS11r6SEU
bNWP3n4LRxvQ7pOqPTc6GMGE1T6ivTvghG2W8bDNALUHoM5CYbbEYApiWHNAM2zf
kgVWVCggR6+IrtZ91pa0gzF7CmOhM9MKx2+Ci/E3mGmeuKcxSDJwRmAHHcTLcYeo
0hrHLYRSgFyYAlDewuPs7acvAca9StsEpeGQyvTN4NrKPTFWue+mTJZL1aRQjeXI
0awjBUpKoGT5QXTkyp8kEhVEhmNeUSK8w1pNl25I4+iHR5WnOZgGhEBBkWRELgHH
/GhQoAxSu79LT5TvVoN8PBItephToBjKf7WSFST6hHgMQd7QxV2A8o5UWLdkcxw3
PLK7XlP+KVzEPFKw5DAv9NfvHiV74t/rDh4YDSshJP9Eh+JbzWXtiQRSlwS2epKK
imjHec+bmAZ6g1jqRqTRAdh9UJ1oGmvJRTZeWrl8udL6Twdugz6SR3flFXh4UF/5
t/6OgVunmN1ec0nHwKpjzKDvgTzX56YCBI4VwUC78oG0/Ir1Dmlb050eBF45Zhni
9O63l8n++U5FPLJgvkoCKvYfAjg5gdo1xBgJm1HTg6Z4a2z8+I8doEMJV6BlYj1o
EBJaecef2naJUG2GL1iNafuLiTXw6kt2PgYeqm+cYPFJLhi3cJ652ltH451vrA02
9afxS0Cz8qVFXnLvLfCpubv3/FNrce8/MTeFH2cEXtK04bkle8GrD/uahaKheO51
mabIjufqb2sR6neiAVs8qkAok1ApVx/CDzQy3ToosEQQDkHgBh46I/f7fQaKh+1h
gmLQUFNJqV46gEN9nhjbQ9wQzOt314zjVKgPcg9YXlEz49kANEtk91rsyWX4tNRO
EI5ZwJJuHYBFtCL+p1zuy53Pup129P3/nHYYIYzatIoDWXitaffaMHBexCfpxaG/
tKqTyHdD3lVlDOsHzVhK5qCGBDqcWW+2jHnetvW4ppUXLtj2koqD1bLNcQcwBI3G
UeVPG5I0egbkZi/kIYEOz/FZTNYy0t2dEA5mw93Gyx9K2yAnNZxb42ykfuEvyWzD
UNRSIEDH8r3d3t7LcWobt6YJ4ZV2loBctuqG3br+9V7k+YYh3+oBdtJJkmAQfqbb
UzDRMm//K6L7IPeF5t3WPewZqie+MNZkIWblMlIdIbhvL/9ebcBm5hR+dLxz0FT7
puz/OXh0seR35x27MNGIaJOs3RibWOhmCoFVuJgSSOZBXtVBHXX1ZSGPZmUVFSbf
DKE58qoT0noodV5mSV6rnDKhxiRjECsVl7PP7oPH9Qs5gNujzFYp1mBigIm8DTwW
K3I1Hk8zQndMdthzYIqM5iIpSiSVkux3FXLH5/EBSZd16mjL0ogx9Qv9F+bkhJKd
ZzAd/xiVz1u7KZF9a5Q1/1yS0Ps7U4gGbKG0kbNI9RROzzeP1sZxJ7f1hPNAYPFh
ls7RVbulUZILmeA/YIPecAfZYgWT7RSJ10FBLuJBvi9TU+kcQy3knr9POY9O5mwK
fjmNKH3ht86T3uSKoecw1vHsUozntJAWtEOfl98Q2cm1dV6TmqSC06fIv7dmcHJk
y6j4Y778IzGTJ6t9+Vd4K1/XQTTn0jreBTwT2SPuy35FVutvHifOD+hzs42tkBYu
CJpIkFy9LO5ORe8VpVvSC4/+wyzL6PufFbj/gD6Bww961Ddi9mTfEZc3KKMb/UfP
CpYG3Hd+O3zNyecwbLqye75pErN2yik600sTBDK5tnAPg/8LeQbRUdpXVL9iWQMp
eGxnDj4SyL0NLxrkGEZKaCh+HqdQYFkvzuwtB0Ja2oKbrjmKOu7aFVZHeAx403uy
/I9pRkWanto3/tnesOoOUspMeTathjoUfbbCsw6B2517fUTQQtUivgpz4JsQN16X
LjZV0QvIYFO0cBvt4ZCAa9MCy4QhJqkej2V+85h80xaOevaP/1npFLcUCKCnmgM3
r+NqbNHlfKyli1Qt8gGxcKABUh+q2wdFkYdiVYT5KXU7Co4k6EVOJtxeFOqUu3oB
i4oXNkirht3zicbcUSjSfov2jHrDVmloWAorpoY+ugkp5pCuc8snEQ/VNueQ9Mdq
Damix9SRnR37V4Yi3N8zNhuBv7KtWAWFpC23lyqYRCqIddiW/U9+1lRtpoBEVy6x
AWNlxN77voIH34uylfxSaD7SIMErR1kFAECT8/1q8O6cMgX3v0nIAYU+x4pxm2Xe
oOYtvV4K7OMjpEkvzafgG10LhVpmwzYrP6Yu/bL0QsFlewtFNFdGr6zKLe8+S6yx
7s9fCD5YQPaFEXb2mGCfmnz/xK2v+/TlVyAxiIlWJ7Q8VTNg29z2kYnfvYGaDjhT
7UzZt31hLMcyBam/i/v4JrZXVVtjXEZd2kFO5VChdTxbrjwkEbdbNX7MSm1crnw5
NMXLR7GTtJi1awIc0JnVIplSU13NuHEV3oOrAOAjM/7FUTdt3UWFOVPWFOc0uAAi
0Gy6nKFkZquMnIt4CvtBIx5n6m7adDNzFwUq142dsOuB2gQw4V/bKcEujbN6nLZp
xTZpzfoI+lpgj1LVfl/ovD91mNB5O71UU49f3OPxYgSnsrcHnTsQHjKzZYWLmAvs
6K1HtpgkUAMLOtrNBNk90chW7RrW1fFSGuqmMcAQIYa6r9IjJN0rGnpcshoE2e9+
dBGGcslWwWPeJrFGfbAd81bIeTALFQ48cg8bKem5rGZxO6otVA+NpKlihJnYqPRs
6gCzQ9Eqti8e+DW//MbAjkC0L3f3j154Gqy18j3ThwAkPV0xzItdz6GRiotoqjFP
HlEDNuUy99u+/Cky7YJo4JzJJ2MoL1nU3t60WcnjFmuttMYhhS/u3+VQH5feXYYq
sknIcAa1udzeFQEFlv6dJ4Z0Jz6AI/de8dmaZBOYW/zklutXxztfmBVrvVblTBk2
TGsmld6sYhp/nJ/tRjbyrSdXpAwSXr46jw1QJgsN668xa3LtJdTOOSuXMv84saRX
7k9ge2CGOz7ERGcoSZytIcZr73Y1urjKupOgZt9lgTUEKAEi/rR0+1tSkj2QKXHY
jIrgfdlqRxHl9JGzK+rQ++YQ2BLyLrshbp2hMLFh3KRyOoGjPDoOEi0pOvJFENq2
x5X7E5kpmR/ROiHzaorHnozIjtOotudxBMjRU5v8bpet8TASHXQ5kwUHBZo6kvfT
wmJXmu3U8xk5x/r/in/A2dZMW+leaHXQVDxgTuzq7SN88L9rl3rTKjv5hiPI4W42
HhDsNySieDR/8Xyox0GkE5cFkYnnqZS2lIpRG0woZOKPmjAENP2CaFz8bio0+J6G
/iSXkxOu4lEzhhbxJQG8xbiJ4lTKT91NBSFja/8fa0AOZvShL5xrmgfmJsN8NeAO
FBI42kYea3pghqkjsa9H4sMDD/26X5DIWj/NOhkldm03sa1LV2EtO8rSOpDVmXPI
y5gBjFOoako3unYTLD5vu/VqQCH7iRQe3yMV+dKa5P5Jfr6c3ggZpdDlwnreQLdB
XV/z5UR0ycicIL4GSnvAJiERXRZyc2hVySjtDTtPOBCsXA30DxMJdJ4tlP3pd68r
oFaycdXnGY9jMhazz9p26lb5cRO7ispZIwR8LTe3iAneDHSk9pR+9PJNW18HuLOE
6XPxDKvESbyK57tYcOODBWnMC2kBE5HFdKja3vzgn/oeTmMDk8EfHdmDCNwYuV7m
D5FZR7NQ4x0LnUDDRGfiky97GquTlmSgnzS+DoeJ/1GNAtyLQgQq+5sP45x1Fudy
KpaY0+l4G8n1J+MTeOQRp8lkd25LJ+FDPZfE/5BZxwyLwhaf27CdD8yqUiEjS7dI
IiUt6Yhf1TbKijSZqRACOwL7ho7Ret/+E6Ok0EoBR0+/eGbDPV1UpKLecRA6CXPc
rFhOJYbBJRaaxXH7yKUNjZadujVdEPbzwwLyHmbTxdXZx4/DY+znUsDPfj2AOTbg
lDZcrQJ7p4uREtAocFaZqATe0u7irsZIgcoyPUxKZedWOGFzEtXbbiu+uhlEnvvP
dHFbD+n0+Az6usDRJNJi2P1xDdq9i2mylvn4AIXldMlPl961IdrOJ7V/5ngb5RdV
T1+J6uLaZnFJFobBm+DRMCHKMDg0r3VKoQ887PCyNjSQZoj9oIFhmpz9536vy6k6
hULCWz7Xg2uEZT+61zr14cJOcSpJNJdJq1D6Jvh7YU2GyfbjNkHnlTcaQGlHK9gL
3HgKsUffMa5KhT84bAjTAVLkG/R1h0uuQ+eT7nh0AVl9PaXVIXX/xSv5VLOuyVe2
9baqdlt7zbw9p3qxhTDA3W/znLa09YBwFghkjJdFU6HZANq96HjJHYqrlic2BfxG
yRhXPbkVeeu3d6hUmA9o5SJpfjab3cH9tbI70npdjbRjVUDXEG6wrU0ox5Ga3FbD
9+FP0JCplIpgXE4TYSrSyH8ZQGMITi5nJASGYKpfO+Wp7lt2Qr6mh1EU/Aux1dku
pm4gFcy+WqiYAHtxEsiPk75UXgyqG4sJgOw7VkXt3bTkBGgI1TICem2SuoeO7HIP
Cdk+YoV/XU1Ns93cVU1MW4TmgCDVmN+sx15cxpeiTJBqlnVjvBIM1EZtZNQsWS+H
XxUipnasQqpmOANlLQpv4cqJ1w69sV2PhZmhY1aOr5kfuLehJKP6vRKX1x2tPFP5
Re5Vrn+DDoAylG+EQNz2TVW/AR9uDPnoM0bmVaw6NsdU3R2/x1B0yWlL4WfUVveO
kWGfT8LGG2+UOgk+fMAwr0OslBrhyNx+rnpnRCBOQROIjQFhME6tux7cHYWLfGyy
ExQ1PX+6XN3Z/3+Jhn8NFdmV881sg4j5vkq0/2r8GnwjOXilQL9VZXFzQQ+z2NfC
hoch1FIMxsG59nERaApuHPFShfQu5FsUKTmmywG/2n+Hzz1tSLLdDzpxQ6iFnrCA
Yq5FgKqgdn9Y6dY0XRbZF1XF5+0RMy+/BLBU+I8AWfCPgkF9NH3lsHPOyhIf+jFD
WlxYXaS/kPBAAFpr4n//9tddhIKaot3pRA7q3w+3QOQfRnf89RTeT1+9cbhAN41x
CjMzwnsxvmasCl+Pb6g+Y0LtRP1NvsrO+FeBcaeC1dhN4vIhdxVeWQVAdWPV9Jk3
H7yn3Di7t1hBN/bFSJtNHliVDbAtJwfFNmbS9OJR7lxJSx//sHxxdwnA1qJGLMQR
l2QqBLQvLAFmSfUHy6xREisvKmb9bPP9lfMZloJd6+OQLAsSETU7NadU2nH4MYmD
Wco3VVmZcksLL/R7ZoZT2YHyfxg+w5yOZu+g6Ptf3PwP2E+bfN5UGU20gZPYtYt8
gAaFzbNQFZE0568ihz15hIDfhyJbDhplGNxvLtW6G3WsEzT85kyPk72WPSmZfl+N
7n4woMSdBKK2xJziL6y/rkMZ6RoFhOsVCPq/KNzlOqq4Mx3LkSX0RrBJGVpflS0w
HgVfxz7eh7vRqPNoX4cXVOce0L3AOsgacPCRWOISbsStCpgDXz1tvGNnG4BONedW
Zbjdp7BTvNiiNfZMNsQEGj2auFTmQeDZZxm5DkUNmbLUcSpzi2QRQxOqdqLQ33Tx
jg1BNuT87pVrsmISTjdjC5iw2DOELk+xbDc3si/PSUTafvbBJlAi2e9S1PVIvsjU
rGPV9a07fJT9OiJwjsF3/ursyjJFg9d5J7njMS7afTsae5QxFRxVeHJOCNPrj4Ht
UvMg8MwffBOLj9tl3/tZVMY0V2MobK2OthOHp2ZqcCDfYuoO0QW7EHO+lYwCwfV+
sIg1ASD8ufmhFtCRbjbufAveo/JBIwRt2cLytO3h6RGC5Oegn0rAsB+jpdaQR+Gl
SqGWS94t6YXY3RC5CNXt5pjEFk/xLokhXU/Sy/9vsT/JdRXGLatlg+6K5/Fe2kfa
Usju+9ejXlGVsJraEOFuG+hxeKKCkTGGNUFqa5DvQNdEhRZxRPotcSvjYK9XQNN0
Ioohdy9jbkMNlbotwksKWi8Do94D9gAfUbfyhtLz9nT4k+mUUTf+imvsQ2NKN3oM
RnCTOcIix9YzJPZfJ8MOQgejkfnOzUI08+Jh0Q+3OW2n+GBdYZ9qR4RTNwE/kit8
rUN7U+hY/S5fyF792krYFeJeJuRL+tPD2o/6ZuS44C9NjaMYbWR/OdFx/qhswslr
NWVfvZSreeBy8hm05cCDqu9E7mW/RFOSpnmkJMPCCHIb8vRmq2tVjnnxwSN6gfWM
GbFt6StJulsgQr1ADB4b8Wick9UKsUz6uIpWN3uabmz2uZLnfA/fZU/OhLtSkrGF
mtIKRgaCUdF36+0oY5G9/r9iD12jWUTsHTGBb9e4eMCQHOJS+H+hEWSIR1l1Ad9T
VaDR05aKQOU2CQ1Lh8/K8npzEFgEvTn4HOyCxd5Dse60ISua25gLQZJ5Psp8fbHp
pkhuxplTKNw/OzTJCsLIxrVGu/Ltr/ljYik78yKjyZq4F0cGFjjvVGuUbYNRyZ7O
60GyTnb4U3/Jtao5tOfxs85g2FBCjED9Co5icBYBW27fBQtPvuwzomqP8HaWIS5S
q4zyrO0w+nk5h3uDzORgzQv0Tp3e8jwHu7MQ7gzcwIB0QMMskTDB0pFgjxGaqGjY
c6QGGV90umVKfmdOGz+WzYsHFN7qBvdm7CLFQPUxWUp3U337hEvPsqDNtVDEH3UT
quAS6FM83QbZPT3IsPrGCGGUObu1mVrndZBaDGH5GVtUyd7yHcGI/u+UTJ0OKToa
SNObMcOirzRox1S+FIadGw1YTGQwYY9UnIApaF54ql3q0uNqxupbtnREQuwAJvjr
oIPiFxnfN1sDhoqytrdrwDI7yXcgSyrnZoWdgKEQObjoJShNEEZ5D+9jF+h+OYkL
hiZ8W0TDrFkngo+fo20O+Vn6/sCUD2CyeK3rUdpyjQkQ3cfhRaxldQ0iVUWTUeqo
cloP5m7zLnJ+OypG0yFrzgdFXR9NALtDmaEKYeImepDWZOT440GMgJ/QOtqi525I
5mZkoC9ymfs1Zb8TICJCNhCO0bx0kyST9JlfwwvaAg6M97buQ5pWTjgif3pMGssK
jt9Ea7FOK7Oa2ZTl2KmchxpqnGO5O1YOAiT4boSEDMVgXjJNw/yOP/tsYBeZ7WiQ
L8ajKI8Q8PJPP2vBEuNI0TLP7Pwq8jEmGWNhhGmW7NJoZbV05/spDzik7VmLUp6T
rF+VMyQZugGMC4uxjGmOjfiFnhblCJks0RX7Y5/yvSrsgvA1oR1QQYTzefxm8QWa
qcQTD8hKKeByyzYN6KUh2N7hwZFhmVV5NHDVvjUU7t2ZSwzJSHY2UVQ5NL05K7DA
UUBC856jvFsdO9p2CPOuCr72zVO9QuqZZcwZDY2T8gGhQxcg5kz8xwQESk5sulYz
kxBxNdt3TFhcp7ANSHokoCrknZVrIUva8lilKY8NLcL/AFgvVdP2u7cFnacdsjvS
K0rlBrxUxx9efcvvndb1IxeIQb7zGpnkIUoqlZQ/37Cq3gDw2WMqkYYeI5FsJ4Km
Ol/jtDjJflwv1kisQbO8w+m3ue/Yl/10t8MvqS3ZajnWo3zBePt0kzKsg4BXTuAQ
G2kYZbzp3ybkdlfy+pJP4RB9qBEKbTvr9sWcOrmd6D4XsYZpV0+B9lWdBEwUGKIn
4N/bbX+1nj+NnaFCFfm1ScU1KVTvmo2/FtVTDBQdxX0nbdW6un9Ki28/ZwfgnpPU
Qnx0pWD3GItphvrQwQGS/8gXggojo6SjvRk7fzQXPS+nuxN1NfUfAzr9K5iWJszb
eqvb1WjCnzW+89YLV5ldFgMpp1yKBoINToEChOKn6ldQOGIRkNO7hsWcsWOgJlfH
h3xJFLctfctn1Gt4jnXwou2jZk4vRqtkGCSEmGLRZ7Hgq26QU2cjKq2LjsYreuWi
xVpSemTf+p5UNAWumBbeYSnox+NB70iCHHAIutK9GjgTsSNDUhFh3NOqmNO/De4X
ovliWDlrI3kGg8TqS+URxOYgU7nZnBm4n+erL1xy7U+sB4XMpjEGabevLDhlWcfa
SdRD0y9ZUA3Me5SQZ0IRHoJamvSaoowdfCJ1CLyPCfjbnys3sr7FgWzIFInb1BKU
kNxEjBb9rVUxz+v00jh3iVq9PUAdRTaTb91L7wNUcA/FUcRT61Y3RsoIzfVhqtsE
+QQDZwKat7Jwtb1u9oMCnPp1X3gU5IoBG/24NDHirBCbLlB8S5VWxH1jCe8R9qZD
mt9qOLtBAb2YkgKMT58fLVyuavwCCrPfm+Uc+wRFOKV/9m2amTaPO1CfYSlaWdhr
YKbK02Ks8zgBa/ccpYjYIp3wwiNjSn9f7W3ePLDvjHgOBjinjwYLTHfxExaSTv2Z
XEsdTFyE0qk+PhQ8aDGj8zIsTHKA51GtNATXa0DAILNTHjIgk5KEqHhKkNlJVJfD
1GhapZmbtkbJr4QvXmMAlAntFkhtrAhfyjWJICWsASk9Fb73e6yIYjYP/3pG5y7Z
GaGyQAQ1+FFIB8eaJlaNtf6P3BJHoid9v0mT5FaFK8WNMsbmTLYnGw7LS4J4wC3m
9riKTS/yNVBClpTJ7VUKPru22w6ZI9ltuRj8MYaWsGOtIRL4LEGvj+zuipUux4PN
fbrgsOT1L/DJT6UDVm4d5IRrK7ceY3QLXyz4l+s3Vo1ga5V7uX+vx0v7dZElfya8
GiRkhRfQDff4f+HAEFvvcosJA/GXYnXzmKdMv+eTggUuXCZHIYKQ7DSOLmOSKK4B
xIIfuIXhBYanZZJZsE4YlCpondpiHDIpnFBuQnDGC16rAShbNVTbPsneWrI1glJW
neS8hMrv3gTcN45JnVOXi/2UU6ro9wyb/hQFpHB8WCVSkzrixiY118duyhGozXjM
tI9mXpoqc9h7IeQz3hFfQpbuCyvwhlhOj9wLsls34o7GFSEDkxKzCzcCS1S0Zi1Y
IjcDCZw94Qla2dGfoMwHMsf4T2OTWK1PYwqccydZYDdY8YsPtEsK6RVlgcpPlmHm
8AipzR6HkXyASyZTCqcQvVEVXY6F8L9ZRTbH6WrMn7/ttuyBZVdJv6eqZRp2X23L
TXut2KA8E+LBTU8tTlmWBij22M40QaJ1coXq+3QliM/u8fuAfWD1AZ9LvoAgAnRR
dbt0xsOw10V4FieSm00rfe7leI6RrIzgElcNZPAQBdgezUfrVP+BqU2SB2q5yrAo
tJR4FGbiwvztFXlBKfbyzOxmxHbRNr1SLEBwFRboXs9pFBTAqJVc3IiUXzxaAd1T
Fu7gKvofNLSBs6LbSFOPb4a6UP67QwB2TtKRpJgyC5yjsWbfup+UiPukJFGE6H4h
DUflGnwIe42YtjOT2K4k+tGy7EdfQho85s+qeItoLFJ3ttIievIlKhijzYMz8AX0
KkBTJPHIzHMixjijL3HrAMDgj28tJcVTHpzJ2KUdIgrU7OCO1RXKl1QOT+CrPES1
FYtT0mJHmxaEZLyCBX900cD7vuxLsFk8ySkX58/XZby6mQSY2a9Uza17s0A/rNsY
izw6SIVxLlr5uSdwSxibRpkbTLc33zlrdLXoYgcJNG2aFh7pwAgo9O7ef1UtnAIK
I8qNInCPZmt0SHy3jOG82mSbKN2sN4XpLsNmz1jkIrOPQO6S0nkiLZCjoaLN/adH
oCM7+fi+u7/caVqcZIHbNYRc4rjtPrOoTijjN7LzYL+qDEf23+ItOfnr0k11dsG6
SeQ+xEvYMpWp9Pg2Ygkj34iNiOSwdNjzY7lYOV7r3XW8b3NQxKAd+Ds0bJ/Ymwq2
R3ImmMzjWzPWiKB45xxB1312A8wovnoRnmLI2kr+ryW72e9/UHSyBa1/6Z2qJkwX
/dGxEr7xe9BQpsQ9RISyrbMlP8MUjGzd2mhLaQSZw7TvQOgi0AFfT8XJ6IpjoV2g
8tPpnlJwybEeIB+/fP4+4fsosU75SdkmtOMITjhtAWU3K4eXnL7qCD/s1B1SCsAz
kCuf+M+wHmIEpMdzdHDbkTxvy0NqwrbS4IraEc+tFiUxZELjBpTjsUky5rFxVgtF
LzCIPsRpMMaWX10nkybLsQ/IcRKzDb1V5cXXHZqr2aHwjzHWhEwx/8acFFKxwoYS
kb/CsqwKojtEyt/bobW6DkGZSj7U5wF47Siq4JiapX+TykTUg0x1zvEWb9kpZvTi
q3gDWl3TjLRQQ7A8tNzaNbbFDYvD0CdAZGa276Lxg9YYr+cPWf1rIE2dOfIehCQk
9OGeyo9t0ocD1my8RxQMU0EOYuj9dZPA/d083j+bLqB70fZf1W8xCZFDH3E0xUTH
f9rPVK1r+5YWixEyFjh1NtrSNKk4LBXKjHOYUpSdku/8hkq7br02DtL53H78CpJ5
/S8BYT56bV2sVDQ7I0yE4rLX3oRM/zT9ZAzf+NWGPIQ5DkD7oCRc5ufT9aD+7ukt
JCsUlEa3zEAjYyWpENATlQYUHRTWwB/T8GzHJ+y8mgDvW2mBMO0f5QJrcODccrSk
t5uGAb2N5JuN+QiIUIfyRo30dbhBLOHUuZ6qbSks3kg6IAzb0vaRPKb2yMbbz1MF
OTIW8AlH9BXD/2bjpZhwIlsMwnNzVAKS3qXZ5scu+vTLVLUHaXN9w9rMk3o1u3T0
Lb0+t6+qlow5xCor20mjw762J57y3exv/HYbgRwJOifQUdwnd/0jmCKyxfARWSdo
2eYD/ISYpbwCfU/NqojKuLOjbTylt9r8UZfYRJheLiNAob9LSqdXaP/mW7XkZ+O8
Y4i6elDudxVYkgyoYvrNimeriMOUm932XqZJvETt1AW610d137xjc4+bCtbnRc+z
4C+gfTZJDajGdHTSD6eqygsV55Z0mpXkwgbGI1tONxbhxqeexTa1XpK70SvEP59l
hOskzuGXSPjRvM2h3hkNee7xyF2FQPbNgMFk2Zi42S9OJvBRHkrmaIhp6RaR5kX5
jB8Ttus6YktAMlmP6i8IaPUfvxIE0nXnii95xudpkeyy5cbVnbI9M53GDmGDRWw2
V8bdK/YxWTVw8MYV7VPy0djqgXICViaT7Bj8lVzCNn8uWi7lr0069QmLa188OVGH
HNKUBYtoDpKg1FZK7yEo3mZKFGjeEoRAizSLhInDuo6MYwJphr1gFJQ9+pZ4Txx3
K4TSVRnC40sFu8qsbcxLH/4aCcQzy0HAUUxHiRMc6Bz8F9v4LHz4pahv701NJK4t
3wSU5eIDR+xR5B7fPymI+3K4jciZJSYCylXEAvNJ2aNfrMJ77T/p8bjLCZ5mBg4f
MVQObUnUGx7amn9Cp/5n/kWs2aekWLiZW8N9Xkcke91RrbUtiX8iNWxPQM65Y7tj
hIOYutgjIYkROJMjZmoJMSnw2ZsGqa7pk0Fzf3oH4e5f/c7LTl0zUxxLFvYcts6d
BGkBdgjuykRwpwVBfJUXXjcgdX9zn3vC8MbmZul6TSAm7NYU56o99s5c//mgI4Oq
40OLuSyIHK5CaSDle2SwthIqDmv8QEAyUQM2j36h4Zh1zqzqLk3h3tgSwVHV4c6l
5Ia9zmSyw7cl3os/+aSLCBrxd/n63O+78gLUsY9b3+UDsKerpJzEvc43e9Y8+fl7
l3uHGv/msrzsLJ+gzVGKQTm9GoVq6AIEe+8ruDdgKQdZh1+2JyX7gCDxMB1aVt0y
WWsQ9JAZsEOU6zBywo5DBwKsQeFKfSkjf/fXAhmZ2WwGyl7pqP0lyGzCQrqQJ1Ra
Y5J3rX3QS3kT+n55Mmg7oxOrUwhbn8nHWZKLzPUqWifFmXYClv5n/pRe+GYOIXIN
gX3RDD9y9CrxuoOt4DELepMaZp6uCdnHP5OylcKyDbIXC/XH2tZDczmyXYXeyRBO
v8bEbr0uY5Cq6MYNdycyRKAgb86W+qJE+NSmfHgMRcq4RcFdoN6KXiBVZUQ3y1O0
W2snNRuQo7VlZ2aVY9z7xbOi8bMfMQX8I2BK1noAKvYQc+WDBav9pEXgE/krfzDt
S0vBnUDOuXJIn36nI1ieMl1p8SuaCOdOwd7FVsKqt++DnDdJQ+/NEx93RbOBck/j
9rhvGmnInzwMyNKltBfoAZh2KfUNQBJ/okxOYK8ZST61zEjAbHs/s34HLdjsp7Wl
Ik8Y4NSIpv85RIgkUCmTor9qR2R5lNP6iU8GD2vKZ0z8lu9Icjv8H3xanI79vnf1
N3HBdqnDA9J8wAlH0uqp9XG4OLjBvXSxooyOUpaScioamV2MzvjJmnR1yVMZ4mOJ
uGTzEKlSNev+tjY76POxw4nTsxY00zLBTNYyO94PsQdjYeKEadbStTBnRQDgoTHN
glM0cyuCSm07vP3xSa9RvicCJRaTIhVcU0SMmi49KtFm082tuYS4dEw4yyVj9Ka9
x2WVZtgQt7Mw6pIBZOj60vIyOrFv60moYqxWabYK/Bh5EAkVwP03fOLeYKgEIYjq
cYjHReh6OHfMopr7EdmIPYlYzR6nLDBnP4otnImHHgtAh44AP3PZaMZ3sTrlcJYm
KGxauJQbxljOs9gWHX5QlJeGZ+ixnJOBIH1peSsezSPZhKDoCy11AOtNnxKtrUPM
g/IdBfkuv8wUSm8h5mNKnoVKf2nfCZ4y9HxL37uxXLIXdOSgvXf8tcDshjLwNjvN
XqVuPP1aj/AQF5JdDHaFqwfCqJT7RautvAlVB+McUc9iVD3D4ni94qbc6asrIxOl
J/HocR6pQVNltUD1osx4QtaZxkvIosf3bC6TbXh1cHw1dqyeXUtcPGW0OV/YYGMq
jwV3XlUFgzrulNrKbvwyinKNXB8FpJztL2inbJKMNLjB+av5G1KI9w6Ax+fw/utn
hRRH1vQzR2rbT7CjEBcdFQ+bLUkHZ4P+hxTDsugxQARi3PMATVN8UQftBoLMeKnJ
ZMSYtpndnD8OU/9qP3sbZiTnYXLq62p5V5737u4dNKQGBRb4DdnM+15e/daaBHaT
1ipNAoxBZrZ5oYkzwdn04Vc6xPSCnWCDFhh2zSZRmZlJAfCUK+FqhIxqLJSiApXX
IN91w3C/HPJDS2o+XNW7IMtOYy3LJ2VifkPa97Zqaz3o+Mp1AOr6M/mannx9A8mk
NrCJCpqjtXGwmaqzcKCAeEE1vM0U+Y6IIl1DwSQRRxI2pGB07aPHoB9YTFwZChhL
KvSRBnkBvSztdt0mFTdNWr9zAn4IHFMiB68iL5zYJyjEr3gOmeW4ZjxnbnjwdT8/
SPJVRloTab/GG2jygd3ik5bJGd676kR1J1VrV5tueQuRAkAVREoxCca3YeEVjqTG
JXrMYNti5/2bCpYKcHp27UJG4QavbGI3JBgIlYrKawazn3+PdJX9vDOmE4tvTMh+
XfvYo0GGX9epmGE76nwlqAuS1l7UFrlkm2WE+oL7pMEXJYGqvIHMZpcCQoAPU26r
hq9AhgpKiX7uOYx9vd8dDcGfRAwRToLc/BAZDvxP4pKKurWspYXzZgi8BqIIdY1Z
cs+u4WVj7GCYSGu4fc5q4BWb1Y6aslIgaOy1wtBH0O3NWgPIP/Fcw/V1Wqc0n0fw
EUzM31CPWgfzBcmcXMK6a/DbyVxLAXc4Yw2HY9hmg83/2FE+nAuBhHbaqbUnEftu
BL5D7/qaW/xEvm3yiSgl0wZUW1Lc/l0sdlJ/Pnr5JQSw1l0/RCTTw+Mfwi+psIZX
XdXpfJWeAG2DHCGXExsJ3xKZnx4gJ9zjPGrXpF3oYU/OTAa7UFBgZvMZeQB16t0u
eEeGGmCN6BL7rYu9vyWZXtC1pJ7m9SyoYACrs9M3KEKt1PsDueO/vwSPkgTP8EGc
s2z+cGBz9kkkTbvrx8DO7HMYA+ln7+/+tGrVIdDRcKFs4CA7c7wC+eiaYlYW0jpH
VS1el3sdqhWfvtpMl5bUczAfYdDq4HRTmHN6IyENvIDeRToEyovXvkBBJgraF+fB
k5ohwKLZlRZ5HMGef6BukepWjH+j5Ig3zQTrD45+U8zo3JNvkTJM4JCG0/FEurJ1
4tmU7DS5v4m9dSxQphNiBs22MvcjRDGVS/0Sj53fnJALuCoLOD33RTKCV5qQrcoH
y7AOcRTD4qVcEHjTaiAsVGIvyXjFb6D0QZhNLdQBnUNWHXBtT+D1R8kZ3MhoskBE
5JUXxykSUzUv+4UHm/cuslAvdICBnQAMvW1Q7PG9KKlndraLftf9bxi6LmeozXiz
WsngJ+GbUa90Y3ruGfvd4H7/NRGv5Wt5sN0kBSgeuT8ZiYWc7ub7KCA2rJi0JW2D
vJVLAqQ8z+PtkzJiw7sbn0aLd2nXGclHCDbgu56UcOhiS00rNajIeQh7jcxEK7uy
nelE8CvNvExG5kxZAWTkZZixp1JKIwn7c6CC310lG7iF30IARj7Wq2cN1l/x9tZi
2r3x8DC4hUyPs4cLH047TjjkkaQHF/Ofw4dkMQhTYLXUljpeNgFewVcaDMgmnjCQ
o+Px9PSssd1IsvuiWjX5Rvna381Q49ZkKOwL8zJuv7MOV4iDYI5y5xZN0rERpiMY
QN7w9lMU82P2rV9LUhgJXmpY0eIFrUzilJuWHS/fOQK6pGfmbToH65rrYn4rIfqP
f1m+BlC0TePxKjFOuL8Kk2+ewG+zul/er6ID2mdYwAPNs6NqiStRZWzTqf7fsP85
ZhmMaRfAONwr6F9NiF1rmho1M8aA64/bJJCVj+J2ne2rFrFdRLxwhhCFTgmAXvOD
kc2cJiKn75Wg7QnGOumZYiG5YzFMqHckubfRSxeX2xoDgwt5u9+mo3X8TGKiGMYn
2Z9KDl1dOQAQ7yUIjndaLgQjZDs7L8+dIV5+Kmc4sifCL6+GxHJJ+byoMnlhpO2f
id+0wHhbzpw2lYR76GZaB5clmA/5dU9GxQo7Y8hEwvPmf6rSw3VtjbhumeIeZsns
CHYhlJQ4v5cERWNA7lNh+3D8Q7I4z+o9Epc+GXEPyrWe7nMga4yT+EJmvcZt/4UE
j1GzvEjtcUULHnowUeJYlNIKCb8D6+js12wCLhlCZxWhvuFLA34qpf5hwDm/JwAe
9HF0ydQQ1RfO/Kr9HyX3NP8t1QBfeGuC90IkYfBncFpQVvHyPLr/RKtnlZWjOCHc
vMpZHhM46KRZQagjNgccfT2vyIPvyyf3g8Yo+Vo/fRIkiTVx9qFKMCSKGXJJ0pLJ
Uk50sj4kXUMQtverC3JRa88gjTtTsIIpVjq7QpcmXrbccIkycVOHF5E9eBsYRpK/
VnXzgKBE/yA0y2yTpnDR+gXg+4XxnXv+KxJFz14d7zcXGPjXch4w0ha+Thcjwt2G
YK1mvi9GokxwNhpc8gpxEd9JCLtnc8ae7ClEogeWhyuFyZ8ZCUqBpAKlnuZ4fMNq
uV8J2IcDUwvn4U6MlQB114OTFVUrs8n1ADpegXOGX/ZGi/oiB52KeyhPDVmgWfHY
p1VJb5UD575E47/orqAVj7mbYgUVNbg6zA17WkYVsh583V4jhDTNbmwNIq89m7NQ
GM/Iw4zCkmJsKaUhQgCa6k+hnv2G3s2oEO7PQuuiSbB3FYywbg0g4uau9sLvB2c0
NsZgpCDfQkpd4eh43EXrJCJhRFhX+rtmLyAAChiwLDyReraiq4YhetJdIwoJataY
1aojDlDHEePCKAqiX7kdtdcI5dbIg6BInVpNXIvlJv+wqZo6+Yi4sb9aS8My5Cd9
qk6tADIK2wlS1y6jbfh7KLE2iBeErWRreLnWc9GAJdJ/WvqQpjUoMZEFJnC9SFL5
sJcEMHzh79bSGKyOZDUuDLTQKSrj7pXx382izkdN29ooXGb9fgUc0mxLPU5LNjD5
H7Pq3Ojskl3sNNRCJYhsTXiIoqnfbAzRRcbWbbvC+IM82NXN2Bdv7zJ3IQbxRjq+
wbyUVu3dfqEjh8Rk5owdw2bSGXAocfSqymMCa0OPyhy1JDhIHVyCs47nIyXu/2c5
7w9S6BXl134Oglu47tsRXe6fsswsuyI8mPUsWBUECDdqtYfL6Qb2+mOW8arkWcXx
ZfP/eudxOPBlC0kO2wCejSkJgdoWsj61XlDNPjABNC69BjVSS08Xy5aFYWHudhlr
55hDUEpHUaA3gY2Beb+KJJUhE04cSNTwDJeBKSRlDdosqz+lZin09ELO6oNeTu9K
stROyJzHukMUseN/fDYRhmgNbHJJur5phjh9/swDHM41hwMivqOHOJ9HqVcJdkN8
qr4I+OS9D26XogIO18KijapsAsE+CMdXBkrgELRXsuhKc51cejkZlRsz/7uBJcjg
+yTFhPy/nVsYGXM6R257jshvz3H3dw3TZ9oKXZaqkGv8a+gIKCDxb0Rf/hwuG9uw
3YSviDLPhqvi2L8DjjzapnEDNmlXBoVyWTUYZjDEtJATW+4pFAqASMHdJTmx9nSx
+SJFi4g1y0VlpPCK340e92f4cIUv+zzQ3IaY+ngDaaFVpIWtMM89/H3hKhnsNmhA
0wmzVj1BwkUnyubAngmp2XPNtYTmOsHd2fcJDqJrWKdM+q4iFEUgEBc+CCVjHisK
6w8hik2prP0qY4MnRZ8VVENOvL1BiS+spKntYfoZMFQZrqw9bVjMEPaRmlUWOdut
ZgOhwtmzQcErw1HqMFU4Wg2yyR+2jNLXNQo3I+f2WtL+A5R76VSRkOvSwNvUOI9e
+PGXiw9TcKVWGiaER2BVDwYi6bckQFIygQ5XkzyFX3jjPzFnPmBElZoq2B1wLy5P
VkTtA7TRlE1GF89cbVC8+UML9qyB5Mfh0Iyzzh5S8JnBcwmHqSs3DsRfo06ne+Hq
iLA30/vVszVBq6qZC1Dn5DgThsnJk7O+WMj6KSttRa90Wy3bSAKSfjRVEEPg7Jga
iqkbwEXpA9/GXr0vBwPNBcE9tN0FFgESjr+XJlbF7hkQhSdOWvcauVIagqSPc1qn
O51pFB5GyGKmF+O3GYWR6PNuzcU1R56YeV84f7TiBj0IzB4CwFbRzTA19CkmH6gR
zpJbYr3yFHqCeH/NVTeb1PkrWrvul5/DDjeKjYVCounnwCpwRwdEC911va995E8L
d4Ej5VS669w49jaq4mNzjWOuShThKIeZS28gNcfp5s6LuWgqXjt/bYon3gR5qODF
bgrzKdUhW6peWJu6dv837EfyWa3kHZN/68B6CqfOf+p5amkAGiNbIe08mPOhbdJz
vW1ZeFEGg6RB27ghXFVnNgAIL2ktQWpB1pAGcdofSTbvsncHgaGniC9xBScXrk3p
VcrUAnwXsKUvFYW/m5kcxMgWVJNP6hJg+Nc1goZ3I1pPIu6nfBXdcdJgCJpbDzck
hbFBPKn/fzslWwVKHqwjtFCpvgLoXrabqkWjDaTxTNSveGp95IQa9W3TyIBR4H8T
XbSihc8w3HP0G+D4JdGSGQUi2Sxnj7+Jk1yGnueYlgqEZBwfJoLci39I9tmeNoak
nB8P43zEYIPdZEBUS/uLztyOwtdqFOShqerWkzFuuCBH1vHLBmv9ZG61tqa3l0e7
2/43R0ljKaXa6+3hwYh8cZLOty7Dw5sVzmjuAfgiE/OuWEVKPh38QzjdFvNmWCDm
/T0rL5xQ27DPS7V2sZKMhY2x2seFUcgylFqrTXsSnuK5DHHWyzkoBAvG48z2vD6W
pF6nQviyAK2SVMMO+uDLp9F4PATaVvZnu+MEmyjx77i3kGW7F4uHdF19iUnTc30i
e/2Y99ZlNheoEz3Xb9j1Qx4psboSYmuWWiD7yVXs16k7EnK4plKXMn9T7zue/HYQ
B0xHEBAXkWIsAAmZgazH8Nuai8Rr7rtMVyztPreo5ibDJi2AewvrptdP9Nm6W20B
ua4+pue41rG31FQbZzpbkrZ/fCh6XbafG8ufGAhtpMV6O86xgRZJlULmoh8dQTz7
3TpjjjNkvZum31YcV/uIC8RqbLqJjptxTLdcYex9i068ACD5omGCfTk9NH9Q1Jhw
HpC0vcLxjRZN1OIlScncgFxkzr3qCyvVQ/Z2OXdTY5YqE2yZJ91skkUJ13eJRkL0
QYBFve9jDYQ9GmLL47erj8M6jpvYW9roErZNfwnkWrJU7pHJHDJo6e2kVZ7Qz9YA
SB+czpxIbIH4+IhOaZZLivEKBuwSAJK5xTAytHXau9/TH9JNRCOlq/ufBh7jL8E2
cduNln07CtkNdd6YtqY8mQYD4LCuFEp4FFw/yr6md3AcDaup9ZX9qdkI48P6QpbE
isxEP5MTBIfybPDbkG2flhas5T8BNLr74Wo2BBch1tFMN9Va5LqIcuX0X2+i/Qln
yVPRRA7vXdRHpzMPMmIuKBz+l0uPZp6BO2DyPUocy2Fm+L0H5yMHucLgDWwmp/6a
fpC+tUMU03GZFa7Nru6tFMd6c2HAznpfo9ptQAyEpTJfXCjD/hfD2BO/d2hjzWO9
/F+g/4yFKt5Y4IkTldebSv9wl7Ks60thjgfZanKrpW52dns8/tGZtkMtWOz4hryT
isEM3JsiQwJypCV8BfaflqINvmHZX3Q3gBirU8ct16Of8AP8vqGDk49sNbcnsQbl
HnkTjU+n8JSed2wYgLKc/YzaoSlZ2iUFkhkw6W3ZKUM7sU/DUJexsA2jE/ME6Bbf
OhebSv4xB1TlYNGku/xqMUNKcNqha7Zadbja5pGJyskQyT2B639Qk7vR6MQDdSzK
cgJdAG0C/iaYHVdqUG4M2phxs9X82SZJkje6uw4FgQPp8BkuHMaUZsDkAaMtSSmk
9d7EmuQRNQBUJyNcZ98YwUwc3S6+cZhaENakmYuT+2jOsrRMD28/MTmsUVdtY3DZ
U3ejDQPox3o0Ml520drel9Wf09fQKOBYe93Ssi5TqPfE3mUSRHFsi3PIW5Wkk6L9
oRaxEliAv7EEbceCcWSWmvKjseM9AIeviKGOlTTG1SGqAQbrfMrR3MEjy1NcwdZR
o/Tcp5mnZ4lrR1MA4jpTXi+ye3kA9tNAhfds2nDzUkH5zYjCa4NCfIEKzoII2ICZ
6/5LIipglB74axYD4y5IPgtDCE94oIT6HOTcLTpWOOa6FlpPP5ustj6IKJKOSyC7
VTfgCwZqVzqg3p1tKp7c8jNo9VPpX+hvBm1wrW63PWx6wmQBXOg8kZpyW8YdSQCJ
MPesG6O3xp3s+rbcQegoPiBMKwE1/A6hf8uIb3HFZpqHSH2izXn3SUYD6Yr/jhmN
ALfWkXpSRL4cevyg/p5Xi3ZhbApSyONStGtYEpshcLsImHtjvHtkcVU4wMd8XBhx
UOQO95y5FYYEIUYtH7aaPCXV+wIdVginUuqYrr1zgrWtR0h7bATRqUFMTuEYgc+1
R7i1Y5jFtvWOhHAZ9+163zSHF5Jm4j4LLMOKA/H0UHW1kM82Ix+AyoWKlZEGfYj0
LTdaD5fxAFJcS/KTl9/yglNy0WAKgxW3w0FuRg2ppa/ZUXXfHY23PK9iu8m1u0FB
QzpKv0acwdB6du+fL6D2o5lZf9W6U7vKnG2q8ow5mo64mRCPKDNOUPIvncJW/AL9
j+5IJDIt+/kbVlONZA4SV6h1sS6whEHLAcP2PJAdeI33tkJ4ZbIngWOhdPAzeYKh
IVqAEtiBZXOnT0uLV8sF2paVfLy4EApQATqwWh+kqJNg5agkCfivM8RwvAEO7uDc
ESlAd4fzSU+6h20ZUL+HVrFV1lBl484Ab/xOmgpUZHC9f3m5LK8bSbO+usanvFZG
ieLI+PRZY0oOuoM9fvxOcTTY9z4ybxQsWURr4kkgvjmCk/NsBpfo/q7RxPXr7ZPc
RKutx8g4UM2MgsSTrJl6RZp5WGsMUm/YLrsqTFRyeRJOCf7UuefASLgzufurAbuR
SeE/Y7vVjNO7MeuQ8c7r9V3DFGj42UIQ49CuG2X15+P5EMpIYwKfuy4j1WVTeUA0
la9swyK55ONHsDzQklQapMzAhegWtNJLAboXURHSCcIHkTLozx5CfuQsp6aAOCeR
rWcgoSRjEckXdWfQ89Iwpq4s0z8s8Gm8OUJuVVKM8SBXzAJ/pvuFHeemuErnbrZq
mVtg8Z+DzciHYgxg5KmOBR0GY/FsapF+XNlgaX2Jd0wSjSOrrXSZVxGvnRlv+rul
tnBYeAxMSrKFjHIA5c9nUJkaMGZ9sP8DLQEdgyJ1tH0FtQUwhJ1Kc5yscpIcsqCj
0YK+nH2HNEaniYY6flkUJQ7B8+wvdYIJjtuU0Hx0AZ/aSsPMUi94pfGlnWe8fH9m
CHrblbCO8pFB7qcbOhFHecKDT1Ws4JsHCd6WmTRJJJ+KmndYBYKbAv1LAemcAZld
1IU4p73VQrApbX2IgHZtHz/lU2dH0td0OUGXZvI3jnrQSw3zt4TbznjjG9PYKp4K
atNS31h0NXc8xRpVV2bOasodab3pT4J+7A6rfD64oZxUYSdRCQnwvOAvgVHOo31t
wsa6Xtl9rZK7s8vM2bY18GNc4tbWZx5mcYyqJ80mKf7nkgQcJ0ODAFVQz2oh4Om3
9ScfUkclomgLhB2QZqPt5v0hGXoXxw6DWpoDp9ty9z17TIzw5DI1nSmdAdc7DR7J
ejvytgzx1G2ZOjCOc15S7oS/3xafbSPwmMRpeb3FXuRejrfv5DCGwzgZqSVG91Ux
nHgdJyaLxWIgUDiEnVr+Pf4wlKO7vYGVZrKIkGR98j9/FpIkRxQdTxqPcRa4Sswc
CgOxbTLISevxx28KrJJ9sxp9GxhCxFPx68iH9nifc/NmuYlxJNCMooERm/p74yD0
N5gJOrgSVPjmu7TfY2L9aqwjd4OfkvLa+bXSZcfNwY84un2gvaCmSK3ERIZL0h0W
xSPSuxb0s8PS9UABVmPRD3xYs72NYvlsHWCR2US+YBzQ7GXzalxJYns5keyeEK3b
3Jc4aMYhEn+uzckVKzuMm3T/YI0a7vkMCZwQPFE68CT6tTEnY66xezGBEDckEaJ3
5Y0eXBCVJFklV140UTYJsNSCWA9QJEMmghrAUfKZuVMhWWA8ryLvzoSnvtuojeBE
PaUdRLFi0VOWNJAeU+j4OHd4wy1HPc5nmlV8/8nihBLyNhumA85Pj7SHIvhE6jtV
nkn2LrjabvTHTXBaeaSTn6iRB7fCRWnM9Vq64iGv5l7FmfzvoPG4aja9pyT2ljqG
VHuvoeV1IcmFmMbKq0KlUfiqC3Xq3WNTqvTZqewRR38oMb+fYqi7bdoWPgqwpeL/
02vWL9g/jFdBl6TyaZuh1VEXS5RW4nAfeRg/E60jJDtIPiELFAdT7W74/q+BYAgY
ZTLSEuve5bq9cjlsKPdrgi8hQTQxYSWyGEJHhWIeyKa1f6JcydDsscMe3WRrDNi9
vob0ZRIuWYwiwb0ftrtJ2DD/B3ExYR6w8q2fj5oCuDEpA1pVwFMoNziICk48IhDb
qClDZ1u3zINiXURFmj0qDD40UJPRcEeqA2FxXmTPTe8j//Y/hz03LJcjYp/wh6ED
ufJeKSe+quUSOoJLtLmBsPSm44k3mLKHytqCFmjXEZS05XdkZ2qQqaEqH8lzgWw6
Q9Qf1LccVw1i404LgQU+n+/0WjX+bAUK9Bs7ompXsQ3cwypq2uvMf3SX9ZM8g8II
JMt5DRXyUelphquWm7Qc2SMnu3xlSmXKV10LvajDKFr9LfHDhSCnb6VIcPWSg8Tf
LyP2AKCEAhjZNUBVrOiZBxAl9fxVM8J22I3TzB5EZwz3fCXqI74Z015Wt24TiThX
5Imh/jdKsNuQcJjww2uc/xL4EOpXWizWoQ97Q5Fcnx/VxdX8fOJZM7fXm0wMbPwI
+ZnHWnlNuyNVw8dQENB3m1ReTg+MehFM4EKWN6VZE0fgk//XDbaN6QDCBbQhIQMj
tWN8vLQae0NuluaAS41rIF16j99mvBgN1mv0OA0EyJiCejGSgnw82duIi8G+u8zW
yrVlA7Z8fQ+caKMR5msSyO/39VtM6K9vPVLs4b5MVCu86utDWJ0LuSRyOQj7orEO
JDYRnPbeTir5Xk+uh1jVXNt06tLDp6C/gvXxjgvQ2X28GaYa7hiqPoAlVLLp9B+l
1KyoMz74eXBnvnllCxoi4+mLRWVrnPhDerRW3Vug8MDkeJ/24NlOTjwwBO7zIRvB
kHSYz44lnNAVPPq67IMehheKccO76qU2hdRHLJ8+OjFISBIC86Wzzkx9SgqWTh8a
XUS7T7JOuxQv0epqjqNWnso2NYtdyyK4SHBTLyFJgEUEyoY+3LPKqnTKeshmjASm
M8++QHF6VXPHwjnct8WWbXAGAMbWeYf2ewUH9qgHG5AMl+vhEhpsFVkNrIyTTArL
h4x9m83JKhhNrzuyX4OPzO0i4RqFcYCCxdRSkbph1Rr03rTDz1qeUYYQS6bmfojQ
UWRZ1lqOFsxn+E7IuCDpv7+1XTTiFZ+gOH9m8ECCWLCPP1L3n6yfYL753e1Ymw4d
tzsgYv+vyaLSMv1C1uk5iQzhnAVBxVHr5ApghKb67mSPlEHcXWzHgmYQ5DmwmaTt
lHfmACgChODYnH1v5v+ZZ9//6XXjjOHaHNkBwgzAe5lz9izlaAhybjAChUjUWT5x
bxmJ331J3zloFuQ+Pp4g4qWDnBij0HRHfZ3CuU29D7ogLvza+Qgc+f7KhkRW2a/Z
xJEv2i8DEo2wMsGu5cG322N7unYaqGKfc22v5325FpRWLg3jQY7YU5tEETjEfMZF
XQFKiZ7pr9il7RQpG7FQTojdiJJe8Tis+elgI2UmZCoPnDCw7+my6P7caSRQtnYI
AVQhdrAB4d4TU4taa4myF42UL2FWdcAKue4kTrdw4Af+AV8RPjw9xV+IF2BZKico
FcMeVtD1BypDLH5mjaKiaYe8aibajWiixeGFKLDvtrT7ITkSlNpdFXAAB3Jla79i
EypZYlkZu7ZRAON81/IMdqP8pZKWWux7AVl5eoHnq/L59XfcyEKCxrm+Was1pTVk
Ot7VeH/oo3Zmy+XNZJn8ROtvKls/I7o3evj0zmLFEWDyJufT8gBLPHUGq00XXl7W
BkLdlpIYg0iEo9LHQtcCgfT/6uvouVv9uYaVgniLqjYnEchY+RxiEr3ZLavUcafZ
1Wk3doEbkpfxUymg5Kg66GuxBC+VBaOL7mTVhn+ou+QZeJVmKlO3bzgabzC/fYGs
tuefMiKiDFUdJOT0aSu1yLQXrRnc0UNMuymhkqR7uUpv/5QXyBnl9vx2btNpKTCn
BaTyA457JvQ4KdMnxU5UamVyRGEgqW5hYWxOWiMSysyxES+w6W34nIp6cfepLfVB
vi/QfATgqYGjzFuDSMbD692cDdcFMD9uW8L9fy8w4C+oAPpxwX7FQTfXSsfwbxzp
36Ko2Ip+RR0rcdayL+/CyHhTGkVBOJQ/ZR5VM5fXz08wzj6jkWX5wuqCqWdVJtYv
sdmTXJcq5yN7pE52usUGP2jSFJdRKgGJzoSfPH+c05V/MTwlGPvpA11Gcbhdz1vB
M/jBALQVzNDOlcNZ3GFSAUcIt01zFOXFUxBJWw5iTqCf5CpRxObabMbR4orIJr4H
vNPRjcjlR+6dHAyMOGdZ51pnQhqXPZfNdq4Y2QfRqN6kEVrH7a65od47iYq+4jPM
5y58FqUpKtieYQOv1OCCds0m99h61fOg37RvQI7gOLJfaLzBFsbKYzKywsGQ3wOy
WccpHw6UPx3WQFZslfFULjcPSAY3ED7/4t6IL9Zz+w6dUsMsHOGdH/3q/qQAD5Ee
KGB3xFJEi9pNI18i3mPhPqZ2oFMpnlJVRtbUNF/lcUKVU7yNVbs35CLqSOd9WbJ1
8rF6QUoX7A3IwqapgiYqjzkxro4PSEMwuj1jSzfliE2Zky/0E03dcj/dMs359ALm
6JCLC4w8tmx1YBJepFZGtud53wgiiXmOa686apw7o0vu0U1Y5FdZ/8dyrQRmSFAS
0/M8OtlcOo/xDokkYH1JugywxN1nDqzU3Z8z/GnPa5wITIi6K7aYEwI7ocEZ87Ss
AI4GlACsnOuqPGS8evmkyjTnUng4m8WGtwGHGXX2w9DbKsCjGia05U0KB4oGfD16
26t64sIIdOw+VYP5lpWiOzaqhgSqxr2anb4xSZqLs1refB3EmbOgw3NDVSKGnUTi
SOp8qirEqN8jV7mjlU0YDLdsMhdgw2tH+rVaj1cblHe2TOkqG8H45PuDHfNFsY9J
3TSPRObN/pATY+3Rr+7/GcBgH9DmXftHrrIPiYBqT4Qjpi4DQEB7rhAPmKfZKYJI
bZlX3DgGkRder5xIrVNOAh3I82NEgVu1/8POmA5ZtH247lmytvPoSgeuBlYmxKBQ
TSz6vom2SPWPg3TR4bGfSKs3mF0YzlOZ8nvU8gHlduKF/AFWLsGP6jBGqYZYdaKs
y0rTKr147EEQ4Sshkhrhk7b3DjqFqr2HuIXL0iVYA/a+ped2T+yr2KsDoEne6eGr
SwT4OhcZuysOM8gZwP509Sm6VOYV7Fp56bgkorAk8Bd9P8lNeVgr9zfozmMiCzqw
jbOYwRZzP48fDC4Rqpofll6ysSFtIWbXrjC1mtuATcG2H58n/pRnpcohYafRgS17
ZO28qHmIXq0YsVLR3CtEwTNgW2HeqZEAsnbIlYLQZJG0BuSb5eOWDSG5nUUJQAQ3
npaYe2HtAjZIjT/m00fp9QFkW7BmzT0P62fQYdKTZQZkHT8UeXjyq1tlb80BzfpU
0WNfTvO+vsie2vLSq4Lig0seTZin5aprAAQyCsq/zShvpZdNiaNYiTpJV/wk7ONX
QN3cb4jTGz6oEY1rvL3b/kKcOClkgX3we7b+YThm+uLPwfETiyoFVBVdQT3hu3SK
zWkvQOSIG9LK+xOpP9HBfELQvwY0cozY41hsU+BMS1pzMMfb9Yir+N+ynjbLsY8r
G7sk2p3zn38q/I8re/S7jI75GjC3FJPVR5Q5OfJvaE1+NKgpboWEQV18wRoUu2h1
yw3CTKwMXAbIO7DB1DC2Fdp8JDuexgTv3yVCsCvBxqUqfFvBz87ERiVDRwfDNXRu
iRIXoxwBu8LG8EPcOJbZteyCqYUQbTeTJJfeB/o/RCEuVfFk+ICUn7Tq0lfcnMg4
rVvvfoz7oAqyl3936qKvo9WIGPVKLHbjhVZy45dyN8H1FtlQ2Qf80uQlmpWQB7my
7P0xai7jAhHuU+Da2MMWpZTFmsvDsJpR2MSIrHlQwbMTPCRhWlgM+d3sMx8jV3GP
eT+KtsGO/DON/vxPolwU4Wy6CUuNPQE0/PbeMEJ1RO5r62h6cRqDJP0M5uYl5bnW
AzKvxwx0Sn2UPE2bMBa7v6JRPLgZW+TC9yMXObe7nDwQyWvb4W06De+nnBHJySdj
zpWwXVnwxZc6LA1FnB8WIgAZm/IwFXKQZzddhjwG+UojfPJffKi2t+ncsrbNndKg
8U2H3Vzsae+RXc4Ez/quA9NroyCCjPBX7RvgvcaBKsS3ZL2wd8zB9AjIlvB0waeQ
9Hib+o0IMJJEp+hGr7SC+w3bEB1MspmKADIsQYYlwqHuVl1xmOaBVvL07MIsz5XI
dwewPBtzo+2iBsiEZSSN1HrpQIno+SsJtKwwWmABTIBiJqKLKRAeTMnN/wyQqINk
z+0VBAXOSkjv9PVO+ym0EbY0am6RrpiHe9EkkA2gvwKafRTzR5eTKuL3VnNCOX2+
RwTBqLjfbcQ6Jz7zcSy+7CMzbuLqDtruSQ1o4qsDp07Y3jK45Bid43nDxF4P/XlN
/sF76ey5ldbNgO360qysKyxniJSphuHTC1j9DLMrjLFuCwfP1f0lmF36ZZYSqDtf
36exW+9leB6FS/sfN5de/cRy6at8lp8lqx67ier9nvTxQX/OjQA3IBdinkAhYkJ7
k5e4KDD/jWX614y/S5zyldgvzU1NNdkCzgpGK5Pi/R09XwFosEr+3zqBbJZ5HB/f
cEpRoyUaP5VtLS58qxH5DQw7yAgnHEuR1Kx/zqnewpAwCn0a8n0rXSZLOW606vGi
lsdVwpVMki5/nsEgpIuvdB9+Mz+LRMsVp+XZ2vV/GMr2BfGJYTPIR7/WV+1XU1UF
1exPSF0/9ew4fEpP2XKhnFDEPIS+/q57u0IucohCQSbt2Azqm2jO7k96LY54i7ob
uAOIoxo4YlXTQ5hM4XDgEtxi4CYSkeg7Sqe/wEWvbPRu9ZFLlT7PtnskRbwvmjJq
vrX6s6Ivzw1eZbalq+ObqPZcbAybl5/+Lbk3FaPxTxbivWtq9wWz6PSWSxRzm391
Y7+4Ml6J8g2qh13qsrMdSGOr25IMp1kkRuDH6HzMfxbtxU0OVYkZyewgEczuc++c
HABt3C/CHI+i3ATgAXw+YjXN29KAhrLM+s04ZMCcYhLusFM4LJUUzUXNbph0CPaL
SezZyUU0tY7BfJw1reIcRygYKtmR7xKT/BxtBOWRu95jcUt9N6kj7VSNzaJTBFN4
kdpkaPE33p0r14M/JfYKfPdO4HLBleKKu89ruDe7aotlSJZPavLOWZkkCa/n7z/U
X6ebpeNqSHai+DiidcER0zSRRGwXYwXRHTCRAJ9sNfvWlar5x2Z5Lr9FX+x6+Pt/
h3UW1eId/iO+itbkIbPZiisCAvBMHBepzz9p6h1T+KaUzXraPnfhgu2z9EHGe6lE
WRgD36TrlgGixpcLF78VJxra1kLQN703jp5lhlHenUcxuY34h02QDxAdwL9xu/nL
3zhK5IgLc48L+rz8pZEM8BbAeK6iaU6fP17aq5+2VOI83l7zuBzjRsNoiFpWb83k
3gJ0DHzoo6ptr34WsYLCTQJnNAM0qo6c9y8fw8IrV0EE7Kc0f9ktznrlaaS4wvdc
CBc1fCPgHBOdz6a0guLkQoUUqoIamrPQoHCWAsFjuphoAzaZRkVcm5jp4rLxlNC5
H275OFzF5gZO1tjbllZLwNond8AmMEE7MmPREotOnb2Apm6c6FAcyUYnJcl4mN7U
8k+Xbeadn7+X0LX+f1wvkzv1fxf/MElfXHCzrPhuijjuLk3/f6Yt2nM2eP9IaB0J
ZKNwmYfToWOxJrDQG5CEQ1F6PmvyXhheFTywwP8UGytnnTDHuHl1oyL10d9G7+6y
RgWzQKf/p4tRNKaRCCORpG/v6PX78wnY1apcTCu2tTPLZiQcqvvtgq4a5ZYJwwL+
kwAaq9YTxUWIfkB+kFsq7TMuk6K1A/JHMV37ntQGF4KuEfPd5G5arRH+D4/aNtvf
NBDCCm4JR7sX1rIQqhpAoj+CIxISZM6CGnQ2+t8n+T9Ia1PxYPWQMFiDyhDsDAxW
iPETrTs+Sze32/HY1khrzPcGQRUh4gdw+Y5hRf0G4gi4MLw9dzVRSH7lkoHdnZ/j
InpM2/Q0mUM8T1TglyrviKTYchNshqE7Q/4Lbb3JvtsBMYu0Iy4Si2fqD8vKVEIR
jr6DvDpZY7LKBNTDhxGvh65lGr/lI86cAYjc+/FxHszWP9bN4Ge7ek8UpCUBmkUx
stLVRXFqeIkyUDQcY1dZeSgqcOn7q0Mhy07klefTjU25AnvSuab+ueZVX8OElpZ8
Sv27zHsOHr9hXkKXgXcykjjJ308QBDSiV2/ski9adLEkqmFIOTPQwAIJwfXz9J2p
PUtjd+5n/A4Ri8ukvhl9D3WUM0FiW0cZD/u7hp1gh9hflWrvYe6SsVvyV4OHo04R
pqE85R55bhxtn5yjMT/OoEMNbuERUs+knJAL06HeKbYX64QUq7zcRFoun+BHJpqq
6mriN3VYSNdlscjxw8gzk8lXTyMFKXQ0JYBm3dDIpOSZ/nYAdwCUmCtaLKNoHiHv
lPk32c/HY589u1bDd6oAc17Am8TN/A4znp4GJb50k/UYuDvO74JAqJm4w1HttDh6
934hNrVZPLF2+IIMBL0SOOxjDvLw9OtA2ZbQ3V5sqSjCt3jg0cyyumb2FZlrjDHr
y+uVxr1dHULsv2xFMPxOU2uoycfoevEiVdlcyJUB6QSWJgS5ENOQoGqCfAy1zvXH
dYRUzT5JnqklBKOlUMThui43A4s/W1keGEU1Y7Jtzfs96pqO+SISGqTAbIhdgkTP
5xCrsUtQapD3XmtSi1KDretAoShJg+dznN1/TO96cLeNUdYgkpfmNvQs5dOsAkm0
NoN6HCAGQgr58jKUk3dfzyvO1cYleK2i1s4xwQK/E72iQ/fDsReD7j0Mn9ngHJMN
BoCS36MvM0mFZUFcIitOAz05Lcif3FObDhIA90dEIOu5yCq0hn4tw0cer5kw951j
S1tlxwvpQOnlj0wyXQsuJY3rMbZXshfjQtCjGond+JUf61POyZW5CGUza2jR9gog
Jx6mtIutYKVyOUc1XAYivjvFo0zorsD0Zx7jzlwZVB4JMDllT9gUjPX/JM19FoZR
ExYiHj0LHBOCuPV4HZ/a+zA2y4kzDzOOVpOzbYTByvaFoQJki5+SzYKUisZuP8mi
1I/eMiaDQNMgTNZFuv7OREK00/xiPDITlJGK1n4yoG8OXv09/+UCF18V2FU+5NH+
sviWxEFR9lc07fMG0ynlw583aMeh6/CYhzjir/mIkzXo7L6Ry8Oyw6VTCX3bo7HI
Ix8pWQ5qVZB1pPZVsqMgjj3b8W001pvnnlzNJfYkNkw1sI26EgN2g11nzW+4miGW
r7OIX4MOj/KPzQn6UwSmOuIvRaMyQtS1JHF5sAyoE4WnE+Si3dh3rFdexS8WW9hY
cMCUqjQSf5ylu06O0k1UNaihMfkieUUL4Q2HRBtMhHjmoSfso2m//Mi94XU7kDCp
7nagfF+noqyAits2oaOs7myuC1fdgiI4aBENaGvG02qw4A9YpctmCseToV6uKhAi
Wza0WV6bdDoejVRgrK4VYYVaTMMflWEa3S3GAwYKJ3n0gfCCHKBsBdGqjanall7U
Kb+9mB3Ebt7OK6b/H5CIcg1DOzssiYtKEcQarW84N+o9ggahzIQ/KOx6vc1Cmiu0
Dzogc6miTRZD53Yo3MOractghwPez4rrBENRjjT7auISxVN53v7c0pIvEPH0YtS2
58IiMnXbEA7cRM7mX0vK640SXE6pl4QajwpRVJdGAvfroWK+sfncCPwizmYQVkWZ
ISosbVebJHbXmyy7KGa4TpzjpvdeNblBvdwRjaxdg6ujVuiMyyijN9ArwLiUbvzz
z2dQKQCkn/BHOhM9b4h9ybLdGq5vCObzmZkDHO9QV5t+/7scG/WKIm/hoH77m9QG
AIp/bW6wtTk2e5Yf9YeZCd54QEtGxGIwnhc04b6iYGi9HJ+dgoVgxTKPdt3DmAwZ
zWrRC0qofd2YhGKuXcMrHR17m1br+hVAU1q/QlgrBQQpNNb97n1apbmpuyRgmM2d
nTJkNSWMOaQFEXdIr9QmWSkx7TTXTtEV1DS2vRJaEF+jBbMhuRUjma6cUthBUNVi
i5SlwZf9njQVVdsdKy3dL/d78vZgya161rOJ4sukXRk9e/dX44HIIFPNl0VaNqmG
+1mH6gyex5YFFJr0cZwOFASMAQFnu/32SwnCPgoogLd35IkR7MmkGAW4T4ovt/6y
N1QO+jzY3WzfTs4Gr8Xiiobi96yoX2KUj1t3mmhBLQ04vztZLoXg3h445EXtV3Us
Yvidobi+1chNZflmm7WmZnveuNwOzLHKrzGSNlBhi9wPGRdM/tVpDv1H3zlYwM45
ev/MPFp04a0m6iNzgKYpu41TfBPnCxz8u6lgbxPHkq+ucahJjJbJnC4stuigrNKh
FRcfUHdW6s1fhAJnkHJuNr2LvXFGk7POsNfwlnF0q3mHCisBG5eqIgyTBNu+x0Te
hTqyJAbxsYRUXzAaFt3OAag4Ym72isIXWtDXlsajIIaMbJ+CWeCmlGVHL+VuvyqO
UnJvtXWtQ8eSV0Vp1p7Qk2odnQgfbB6JgVmeKmbIOr5osgFMpUmj3YYOM5tQNHOZ
aVbTUM3J28OMtMOxdcMxu1QEYlhpkK+3YXyPV/Ukgsi3Z8E4hl1E0LvfXeiw/iVc
wYj9650LAhTszJGJ7vr0T0tQ6JyhMVuRB6rKgILyyt5VR2pZ4/8I14X05lZ1WiJy
a4qxeACyHqCsOyk6gejrRa0iL5H/x7twASTJEfgWAPoT0P+uF4ZE3rqC/8cuFI8i
JK6H0Hh4Uot4lsJvbhCi4VMIz4/A2gJc9LNwI0tkgrDdW0vdeMnQrMANzprBcY1i
QOYqEL2do0+26SJMFw8necvTkFw36+cG607Z6/mDWkn5r+ObRpQGWyji52f55tKQ
TRwp6j9TR4tCq9oJmQ9VPMBCplJmte4iBcRyCB917+1ydiXvFEJmyMb5X+VZF/rx
JgNSVv615EAQDLD54bvbKMVux05Sh/+J8cAmxYyof2xmWU/yBd2eIBkeQZ7GnrIE
qXp3YgVbyvK7U1EHPB44jNVL8HjVYx8R9cwit8gP0edFbGHK9ZBpdC9StlO+PQST
RXo5L+nCDX2pA80ZNO5HJ9KJtBu4fGJXOKYdpgUoIW2HqxaKWhO6czukbDZHcKjk
4lQSAacObHvHz6TJPsWKHrdegs8e9Oh35Qxp3m0UlgPLJhp2P2gS9ZURwnjJXKG5
0ck/4TS4c5x2yk0rg53bY4JqsHz+KIrJVIDkUXj8c3OzNp0miKyy+DYxLLrdbH/5
R31riD4Kr0iGc5iFf6KADBXQErIH8ELTlOz7G9WR5HDeO3ZijmnEIvWLN9jdatAa
XIdKTYtqIlIkyhxRtXz25UGqNN14U8IUkSUc1QlBO2yMnH9MQVIVgVh8mvSf6vcD
DRpbX1T3aLX2R+hxUn7TFYTVnXMaYvYYkXhen7iXTabH5vnOIaeGUiCht3mI5D5h
4Qd4aJ5swYacJXtYrP1eXW5gZ45ImKAJ8vV9QgAqYAuKcATNo+d2i8k89g4TFIVU
U1Gv3fKGNMDvJempMgvDkXoRy301WQcFgmfY5IvKCKRB8NSNsYOV8AV6nH6QqNxI
h1dFwofkpdsTzse9CXHjlkfgGKLsc1VOHDEYr/HZQSJBuD28+DuC3V0azp5LF4co
bnhKax5oW974SDvlAy94iqnsG84AcSjNbIrfFxXiSVh0JVyseKqK5zFX7+bpx2xo
5dpJ+hw6lalCnri9wHSb3PO1I5cx7VU7raNbDq/Qa2S7kwqunsuw1HF06akYOK0r
UBpoh3YnUlCTQ7nMvzhdl2Pc24N+HWNckK1fj0fWBRxxRO9yNz/K/dy3h4i+ERLD
G9D7pCDeH/o+ZjBWuOkydnSXb2I00CnPUV9bnqYEn2JC8HFZkNsUghC6cXb2JDDO
ZP0Nx1R2MnAqJMoKsFQcNvDSikq09WpiSmgI23w8YREkTMmRqiFBDUWkAZ9e+www
JZwKgPFURcXKH+jKTgIrRYEw+nRLdFEZkBVC/OqvwOHnz3NVKw6PNsxuj7Z/IKx+
0EfyX5jxUzX3uknMocPYO8z6/Ekgzvvq8Ixy7udX//kY6DGS+4DlttObooAeIZPj
cExGYxkN4oVJtzKaTBxs2kmLJja2w9nHsbBEj7/2/72CTv+14SCmNJeOnD3lE/YT
XaIcm5wNRp2IYLax0qH6//IwI7a92FvGGXAGwq8z1NNgzgrPEvoNYAOOAVMgeSo/
70+DoE/FGG570SsVoLNQUjxRYmPFSmOh+IdIw0iNyzmfajPyOzIhsR83ozRZeQuu
tQZCfs20XSPor5Wy0dQOfPis/IrSILpTCbG/p7B8zHqZo9/u7jsumK/IVr+E0Vmj
0+3znQrfdgnY11Oopp1VOlm0Hl8UZXvffxkPyjE2sygFGz/as4mmHMEVLLH1aufz
+4abNsy/FyQ8mSo7sb2qmrL9MkLZ1loiXdIl/vOtR8SuD87xXdD1M6s/1dv5qHXg
sYGa2XmNUBryiuyxpyRqLFOyuoKWzMCsXRzsKR0nB2plaQJb/15q62XSTWul16F8
uafVAbhCSwZTSZnIw3dHb1WiQsNLyAS+2u98LxBvSmNtYpGDe49vL5k/aDwfur/H
/ho6Ea41yYqGvLL6Uo1FpF17ASdneo1X6zsBkN/zJTuoSXvTjpfZx8hZAWUyuEua
Wxp0O1RMwiUgLyiancHevlAykv5/lViVg8aSmv2cM0RmXUGC+k1EyH+0dC6LdHux
9q1lCWPL4Z6XQoz7QsaAg3nlpoVBYenwWMNSZJ/o2bxCoxkM29mx5ub5Qna88Rks
28BNQiFknpwY7ULvFjySdcvDgMS/FvQ+azrL35z4JzVDDrgxU4rOFEMNxF/imrEt
zBuqnr1xNE/NUPgtmn9KnHzkb148nlK2UqZItMIdPvCRmnW8lqodC4Kc1IPvR7qu
fSxDJ/zTfIvw+Sq3sUj6xtlyAqfnM0TkLYBt3o7ZIQTAo7Jqu+w6b6jxFoXOr7+/
VgxBpsvR2XicMe2lyLzq5TgpIyDIRMDO/YXUEMXxIwfyvTQllvGknr9rFHwoEaB5
yoDfzY/tKdtovjPWe6evhLbA+rvIUXKRhBaW+K3ezQNqgA1O86GJNps2trhQonqD
1Sqt7A1jy+026NuLssWWijVKxOPxLYnXp+xxK+cGTeGt80TCBJiS+7ZKeWvBcCV8
vPKqEIOmLLHv6QtHymsZhtoIvAOqHsEkJPh69KbdpVYVmW2I0DPesMBMZNiWm9Xg
RJpyiu+4F88u57IeA+t+Rdhx4mqGPso1EdS6gg/SM9vdbv5NugCqBEysZ/lUu/97
T7fbe9OdI+Nxz3Ej6rfPkpsg9AbRQFR5hb458grGaUuj43kGiI3YPWZ9uFiPc/Du
DLjv2EY7SVbRt3ykEi+mC/hQIPSL8QQWPBf18rEaVmm0Cq+zqAtCACuhZu/UG4xc
Ni1Z0m52kBPizzFd4CYUdrdzaZmgTlWHPGNQ1m55q0EoIfD4qT9yxONZzPRcop9K
QZrbvMWSgeb6jqOw9RLHvgIt2dsYwX3IpNy88+ziDEW+wPJaASwvI2Y2gr1C9WJy
ekW18WZoN2wV2wmzGpiCDCsFDNTpJqPNdMpBDcBIA0umC+6FwKcFcFYen70nKy0u
N/X38xpcVSclMfIHUwZSAQdb9XlQUmaUM8li881Ny1CQwY3vsRjmx/+Rwm1/s7CZ
PRZOS6yXr+cOWXAlKou4OQC/c3BBELzLn+PAeZM8MJ/iiC18wrhhRljg0X1oap+8
0vMoASpuIEdWGfBOM4oTze8bUQQ0x7tU3w4yuGW6kt4HPP4z65/BI3qx/ucdIASB
4UUCXuDQKzIIEkZrtMY2b1AB3G7BLxJ4qnoPFYIFuSGGTJ6issiTQarOOOaya+V8
tZVnZjgf90dumw4dn1TWmm/FGWegYYEpoTOvIOdXmrsq7Cd0fxGqh0Rv5289ulEz
hMs2zx+bgZbC2/pY2WtRm7sYMVGwLYbIVLDdB5ILPX2uEam6rgcGj+o5SnvCiEio
4IVYCGnt0XHyBjdgbrjrFvzVu6eaNvTFkh7sYHNBU8vWMXYirxII6raPeug6uu0L
YzbUI2ZJhANmMjxCoP2DGjT4KFJFjA5/Hg4qbvvjPft+zUKfgOk2ZE4KpCB3XDN/
E2yrweZpzf7i8e6BcOHzJQU0OFxNkg4Zp6WtSXXlH3NG+6kaxyyShQqCTYRALMPi
Ujdks1Ke6wZibo3ydjOK04SWfmeAYyWiiQUVjA8tIViYWrmvTNkhTuYTDA8gsY9b
pHFYemLs8muBXuWGxMynACqGKWX2ur04/cqDDHVZDY3D123qXuZMlRm2b+sPMNem
av28CKBU9Jqdty6+FBXwyk21TZSHa1ohecjm/DeFRmz89ap9cgRqcipnCFERqyCI
W2wnDJPx3ScZ238wG1EXNSvAX3FlZiQnFc1TMZTAGEKt3Bth551gPcNyz7D1ZQ74
Kuv5XtxI0D72F2n3+G/S2PPWZnXLt0VxVxFnqsKdhMQ6bDSJB45y8sK2OAzJJ8pH
unCPb6wAYE9Q6cwO1Kx+xtccaiyBZGo+uy/0TVYfUXIa7rM29SIRzlVSCrtMNbDj
4susy2NsmvedypMODadEAweqyOHmxgFd1OmK5bQGC6Flxz5DzQ109BoL+eUlhmZP
0R2IzLNAr0p7BO97cdyzvl9LvYI3Vn+IfIY3O/NynJqDo2PV3pOqApJ4pWYLaliS
7xeuf/NUrSw8dacH4CbluSLmcvxuFUYEMIpRuMVq3Q0q7huW1NSIcMCzPXVwP29Z
yopTr8vT3UaXSQk31Ij4hV8lgQIK76d4Ualu3J5TsMkS3qklqI0cz9aESll6Cc2k
Y4NX40cVnfnNCp+s+JETAeE3Wcn97uCtLmoFeTl1qBS7TaOm41IaSqAR9LKOxgwm
O7RaiQT+fL0pwWzJpHvyUYloGz1OGXMyEdMifQ5TmdBoGsvU/Eygf1b0b+KUNccs
GBzzGfzVJ8A24k93cjv9coTpMccp0g9YfA2OKfMSf7S0x3y+ViuzELMzIPLkCu66
WzArC+r+SkxeX1gbE45s1tHoMqj8//opq1s5hL3edsje7JCsXs/gj95wAYjHLFs3
ynUL6ilqwOfffBv8yDbn6gn5THMaA0y4kcOPsXp0DZvzWpxfZtX92kAOhVX9ElJ1
htsoun7+btFhs79R5/3/zEL2n0lmQI7AZXG8z5IYUj7DW7lGlTsIwa4iZFJBGoaW
AW4zXwS2LuTlahPK6Cnmc4FAX7K1FIUW2AsvA2lbkcnQoj3NaWv1yw3niCTE4+V5
1Ij6c5C2EOiof0QDWG5E18BACM57tVhVSPhPKCQPgPmWZiN0zMJ98KD5X782ohc2
CCx0nG/Rtr+lgQ23XVmJAUmsQa+49S8kbIaMYuctTEtQwtd/A86nXFuA4ch1q2ii
LAnRNm7mlg2zWbuSbyw30S82dsYlkrKUoAiXCpLa2o+pSW7w8GytKMjmr2aEZxoZ
rNCyarhcmbJs2OUricvQXXHdmM6yYZobcj3Ttq0ryN4cvs+ykYsdcdXxfY8LVBmG
4x2081iQRD2BNAmpio8mCQ05XyzbYDi+axjizzSeDa+KIG/QsZ82ob31m5f87SkE
faV5+XoSuxdnGFlPGbZoT/iZzDKF9nObswzQgNGYUAcsyufPL+5O0+dbDX4txVMF
lxCnyvwtizIS0QOmklFYHzvBgIhYyaT7sk2E6mDWQlxPF7E9DOnQ1osW7pdW5cwv
fJpdVCgGS+G5h618iLFmqQzF9jrCdAtGlDPRC3aUvMTh7KWjFRFB1ywnPJjlDdnA
osXvccXnDZP2Tvl3SZqzIlkHYCfTGXqn/LN4YaUJroOQIU4tzpT/T6LwG9u2+3Iw
VDjltM6B5bQIt72qkPHvopGqQ/bDxcGz13wdOWFagQ2IwbTR/FilbmYizsEmSAYz
15+9k5QvLXgtkOAOkQ6YSwij4VCxYpk9fx/qOCZiBSqq4kUZjdgD1cX9J9N7lo+v
ANF9lFuIFjYi/MqOWBQ6VC6zFel5BSkDTVScsVncXB5VeTiqgt/dOPTwRgy4yJxa
jZ8Jxkj7xAmLlLD0m8Zb+nzgDT1I8JM1k+A8A/8Ot3WEu5Q3jLUaRkSu2/08tZa9
MO2yfd8FU3b4kMlaA/cnnVGtth2AAJz6TRh+f7EnurEDj7Hb7YGCfxguZHG5+sf5
nkBMYwNluN2CvnyjiqCM+SdWzkln93i60vFrDdsT6/HeVr/GDTslX37zL06sXhyz
jMYrUGioVfBhHtjPlw9kXyXpcQbZ72u8ZXnqffHTMcYjpjWyxxTBoJVYfuIUuRFC
KUczvqQicQNdavuT8XO3dyhaPZwbk4D+rBa9xjteoVtkxEzKXmJMarlKs+w9+Mzi
wxcvFM6bZVQERQ4vleLHGECNU/OdpH1t37pYpLqmsan58SEgqkN8UFPTSsjHBSdR
IZl+XCRLD8uhXXwam2Q8WsiK9b3GuL+kYG3/Xo22Z0J2bGv+/kc2QdTIzA9eiq7/
s1+ibmBwxk9UO0ns7vjlHBJsYgzO2CcQSnSmc9L879UyMYpqJ0ApKRVXgQUQ6Ht/
1z4pjhloUAPoisy+DasWrWCj0U2rdniR6DjSj5NYuQH/IRRuXCchV29La+Al9jjD
lTMKvc7tQlW3rZiQ+n4FpS5nHIPfoUZdqlha9kgGHwtZNd1tHrE7aLlP8h//QICO
tCc5aeu5GGouW2BhqN9Dw2bBu9STdIUTvxtOYksWWjwioEG3K7wm0XSfld5a7Xpg
0CmAHy3KQvQXBhOv2ymJ8KO8/8c1vLJW7Pv0YC9U+FPnWaZc1YNaIcU/QF+Q6XPY
3n0BnuYP//9syQ0LAQBTDO2ecjHf8CnwE5gtIOqsuoyEk+jbrcd4kXHuVnb/fTCf
XaMP+M8p74k/vlJyDQ7E36jsPdm/kbbDphcCtSq2U7EX4dx0ZKuUniqFl3n1Pt3x
CaD0vPrHoF2rfG1RR4MrdgqxnoQokyvItajgB2MHwc1JQfKCMyjObnhkatkknItb
BSz4JM834EGLNSzKF7ErtfA+grbjbKIa2rxL2XwyV9EYTcpLvQRLIIHzwhWOxyva
4XnhWTeekzWWvHtzw+aZP814vfu4q9jH541xHaiV/N5DNDfEIpMFTNHu/M1mObCl
piwkUevFQRnJz0jsR1yROVnA1B9DDURYK6CZOYYe0OO8AGsOT9/NPQOXSfbuOIPb
x80Rh35zeZrfwCWUy//0flTwFBZlTOS0pdg91H0z1bYyf6kafAGT0SF+t0hhvAyn
nkKv45n81gT3p0XoAo8Nt1G8OoDGPz+5i30q61Y67ChVKzJhg8x+uF21xyRHVpKI
4/lsJXru5qlNnA6oiCsCTMLByj4dFfV98JxK4sZYxWjblcnH9e/EpkBR0UB0FT29
PX90vsitWI7sWDlOjn6Cu8x1wDph1Jda7NR4PDRuD/Hu571VO3QfNxi2q/teuAnM
2gSboo22rzxVD2o//lMOYe180Z27TsGOWkHVunqkyVDnw8r+hsFhaCJupgQSH7re
sj/ttYq2es2AvsvPZrwvntcJe0ymHKj/BM0CjJ3hSqVAeIOnBwgpir3PvRC7FvFk
I1AnoPub0ojWxgvGrLfVg5dI8Tknxhb3LRPUbM3jZi/5X5bZnumDzA3ZjXc4P1Wx
9uhbOtM/UPb6w25S3taZScMLZo7fSRtPXwfScBnWpb76vzM/AW3UAy0Sv3+hMry3
y2sZMEW+QI3eoeS7ZGZR+XIwHq/Of2rN98GoGThNC69GWymEsmbcFB+CmjFrUQK9
IHuTSrhoe3jvitV/HvItPX09a4JN17i483xQcAxWoDoyP4QNk7lHxvzzI2kDmhNs
YXHvmZNrIKHJ3NcEr/Ev0FkY5BGwiobEKHmQwx4UXFbWZj39Q5GCBeryRqs61Dql
I+DtPYojMMaVL5SYvnGSeeTkDvwnMVYv7L5m4fLPV5sybZ7Kw90riNPtkeNkSXLy
m2UQa5i3Up2NZY1lRejzKvtrLzlLewqvLDOHWAw6lFi8qG1Ft91LFX/M1A5z1X5R
SYtVDoImB+Oey03onDt2LgkuIz7tCjNm5qZ4J1Jc9tNBgP4jnY3SnuY6MglSrx1Q
sVD+c7iqO/G1/kWiOLMJP/hdo9sHdmF1rJ47KI9pEmtgNbh3dQE8dcIh1++vXeh1
pe0oR0sEVeaSQnw4XiPUm/uB3MqZP7JV6P4ly6wNsvyUOq12JfGFCDufosWr22G9
GaQ+GXzVUJT2nxV2QlSLGwQv05GM2QZVxrgdMo90qI6q25+C8SZBbpZxzkpXZZE6
ZKs6ylirYPF/HYx2gFQrpMxmXOw89hVnR2PpKtC+3GVG9bl0MEKOJV57v+HgLBko
PwSriVhIIS2ZhSYwN6oKO1h+PrCbA3crqHYA4sWQMwHJTbBa971gtRLDd4X1wRpV
YJc7dIWS8KGleJUqeY73zGE3DiUfjCOz6p5nqhdVYT76sW1vUHqSlGJa9JyGQNlI
IPmH/WC6rT8U79X7gbBWpZpVKc0aIJrkTA3ivk0DXwJTQiild1RtEJ7YbflIdZHi
XYQ1ZMkMJv3ccLylbeDv7N4GuD1qhV35hjbs5Bu2Twz7JoNdCzDVNWqhlAp0WY8L
X4qCkWijhXJBiCna2P16dSoVzEHqqsvPrW34GSFVC6l1gjeERh15pYGhEhst0WaI
yNgiibgDUQwpmAeJ1748v84b+c2aZhymQOtwgAGhoxP44GKFrDhhbJ0296YlLFs6
fpCvQq5/8ztf5r/I+qeSwAECcmMM/yFqSVbnfDzW7SCKfhcHJ/W0fkVWxpORmYUn
4Z58o0x3DT2+RgKe30vGLqfnZQJBL37a3goKC/FAIlXtriwF3P/Pp5f4d/XUzYnG
Z2H88ECV74d4QCKxwwi4yKMfATuNx/9x0G5OpurLQYpkEaJzSDxSqvCjIzd7oTk8
3DG1iP0PpjVF6lQvk8dOe1nDhfEcclr9FLs0zie4zwTgJvA+7yQ1Zx9uQxMrUvC9
ZVg1rMZYc3dGbbYsX2gPRyrZUbeRnNSDnGpPTwGNYiUKCRWHbGyFcA17PbxQYmge
FBltmkqvk63MqSNqz5sjYGDwounB++AlWpU5j0NhIbXXTQ9kCwBcm8dQBJKFxJrc
H2qdSGNjgc4pYDRdjIu0uKD+5GhEv/1UovhvUzFkiEmqYb4TTVON3j219yd4rcEW
R0a4C2fXyDmXs+GI/iSswiiHm1JgfyTBisDA6QnGo/XkOK7Gn6hgZAB60xV5OI9c
goJHh1u0LYJCp/Bj0NQVKh54R5KUtJqC6dYfSLGjWgQH2BZ23UboCmuS7GWUo4J+
om/McIBSyBDFJc8Wgd+FCJF/KbgH59mcLTkvx5ZoZ9zFxbt78fdCLguKTiU64SqH
RoYT0ImwPZOF3V0k3xq4HRf/m7yRZlPqmQ9Fi8bwSuGsNVsvdhruL1iPpmkOwJV3
sQaZUWE2K4+wq9NNCFHnhmAKFCBUb3gB84/keTMHynQt8mQknBA5HYyQx5wgHZr3
xAMB+1akX7ZgbBhAnnGa9r6vre7rtMsS7GkqAz+/h8t49rx8V9Y88OiqU0ejdVaK
H2OiUgG+dH5z8JLDRtuC4QkLSODCvpg5XU6iv/kmaKWFd0KCmjDJqYOIn1BUiq8B
/azQ2zlZOWexAiiaCxodj9RiSZvfiS5Ry7ZPHsA+AtiCDeozs7JNmvHBlncEIQ77
MU9y0RCSrd7mMcTx9I7Rz+VnMGQdkcaWtuo/jJKb+5e/j2g/lLORe1hEIp1FKXe2
GEa8OXo7J/1HQN1tOCak+w2X1SvzsGE2YlrE2RfCmcG132QDkQ7rVqqgtBUQqne5
EebF+VkHRSsZNSKNHSe24c6QHErPQLlHro86s/lCoqoozEharzyL8A7NozL3kDmw
WHjpT3gnO1AcqlLAQZBILtLu4Enj5xMsuVngSHGTKI9vHFz7E3GFnBLWApZ+MOWL
B8fyfie9OT1PbSwGf2P0CVmWwimg1PYR+rkpVPuCiNLX4uyHIFKJU5NZU3oYa0jx
OAMHQ0CrLaqUHnkQyxB5Mp1e6KaF/ijVJFFF8ttAmKHvC8IaVvAhfIW98G/Q+d7e
3GPI3Sbftf+3T2L44Ja17+cTWhM8QdsXBFqd9NHcqmPXtEevO84xs0zg5ceCIOMY
x8Z77oKhfxHt4iP7SSSjCofE5ufqGoLFSXOWUW3ptwyq0sKg3tIRrPy20pcMChv9
J2btD6x0r8NKI+2p0F9IyzXOvIVxUvp0GnYJ1bW68wFZbAmFMKnZvEhHebAjUQ+T
EdU9Xaq5oZkjtGFBc5g9tN5TTb5FMptupvm1qG6HUKusAn8tL82Asy12uUsQ6T9x
QFaZ8kkNK/ihUVz30LWVOLlgeCs/0+Rmc6sXrHjzssWO8W7jcNOauWau3tEWAShe
XPiDRojeyPJ2rwA9hlFC6E0mUvKWHpilK54sMZXNGCgGNd5y2NjsRzb+ROmIEADH
zgUWofGkDU/U/3TFLgtRdyk+cTIvWTlk8xNfd3r/LcVGQFAxMfr3MQa8Ox0GPY62
uuKxYpXx4uKcPWkdu+pFrx4+SE1Ibu5ZraqiPetq143C8+Zfx8o1OJvCYdospKYs
tocU5vr7F/EhX4gGDx8LTUJqmTm6gg7BCKuTYN2CIvnCSTiv32qAeIoxhmg9DjRn
UqeMydikofI8QO8/bhT7lzzhcoE6Hx9tZIu6NSLd/PZlZKvk2YBASd6mvZr3wJpr
xc7+7GGC3ZLA8anFW9uuDjYXm7CxEU3W3s0EfsLwj0LbPsKXtCsdoVO8mFD3Lshb
5MVvfDoky+pAeD+nUNXODTX94aSOZySlZfoXtjWWYm8zyUQKEQ6/zsmffRjo1cpD
3PLLZf8gHwJMNrIooNa+lcA1BnZfoAz+/t2xFMT5sotDmnD4K21VCZX6fCyzGfvp
3uFVbljkIB5+oQYelVcB4U1awIFJft/traSiD5U2lFtffALTUxzBCYaC00OU4AwQ
Ch4Zwik3nZUaWIuf2M/RbDtf4b5yi65mP/9G76RREu0nQzQ6YYoyBI6SL5h2GwLp
EcpvR7qBzqP1FvtdTLPlEG2YtVXfjIU2hjoMqM9rTK9QJIAsZKZ7rNozzpAO4PS6
03Zgu3e3+rvQhH4iGbWy8oeNzmowE3VTZQfiMlcw/ztJdiQCnfDwujHYRLtokco3
rliFIBMtR7j1n5TvHxlysiWoz5yAE0w6EjuCOCKGo/7dXdhG+dDMSMB5PlIdXZ7V
E20laGZafsP5a4fJ0HvAWwK2ZuuqFzQk1P/8YaxNTghI9B9C9hCC+120Wx3eL3Fv
P0wGGOB0MjvR6AMXpcJ7IukNOWcFgRhS33CSYyfzr9NCnT/dRIVXSbCwqnDaIT0E
peeNsSkNXSSYVgcS7ZT9aCTDsUlpP4yYZZERF4RUSG3XOZ5QRDCzGEkUmwCMQ+Mg
+as4tqY27+BF2vPHJNHZyi0ezDvwCbhxFQdGii22q/JSqIwYoh5JuGWbeSj/8D3R
D9hiuPkWIUQiOYsbXCOd5q+Y1/gakl+8YztxuMW2P6C0+v/PadhHATkmvBrquEBQ
eYerj9yhYqmx61CPCZPqQFAo4nfqdHoPXZNJrw9KH5Bbqm7wCJNHW4M61AuNMSRf
8moP7PRbRiz7vKL9Iq0Of18EelLspV+45DZ2ztjag6xp6XSq6ptjy3lZFmcIzoqe
T4hf9o9pDwTIL6sYwME0plYMEZ/OO140qQlO5Vnof0I1Iq0GqW+ucu2XeYRX0nU0
a0svDSylKr1yFzJA/tbWcjNIbbK4vSnrBU39cxw+dokjLqZo0hCU7v1WPQAnHvUs
DsqBXr0M721nYXFBwU/rwBf7emKCY3y9vGuhNyfwe+ZnzgrR4J1Nth2chC1dJfK7
gNZcGqEGcy2ZJ+GWeweZIiuTVfP2zcnJ9Red0Qz/DfrfOc28qKTfD4e1/vre+cUm
yAxPRsQo87L50INa2r2sMPDnvztnMYXTCiiUkQPtHQKavpPvLbUfE0OxPJUFl3co
JLiMp+zRP1kfNw76BxTr2I+8Y/dtco/XZmnI3648Sh/Wb/fwwtD1Yw/eJilFtx7R
ShLFsYANC2EnLOG4G3DB0vtPNsVU3BeRoRlh0ZfJPFLyvZow1oHnQVD72UM/Zt5o
JTSgzMqNBJy1GTrpPOoemXOo8DqltxWAGMwi4jusnVk0ea98s6jv9MNJ7YFYBw/I
/2kENI8OYb5hE24AHpoZx5popIOulKDqaPNaWJpKwleraNotzbypWP0ntV6t6/9y
/HT1Mgqh/mlr9DQ+rKXg5UR9qVlP39KQc5WthvsoGHG02J8+on12aJya4w6+gXZP
kQ9JuXaCOdk3m2/2Y8V6UYUBrx1o8UYigzonyhid+e15LfLMRi4807Xkyt+aSk4K
GTvVo42GdFJj+QBikF7L5E6kPPKC/P0/yAgh6HjHaNRpkKDbfWuJj6I88Stjeefm
+d2Aa1+1vJKHDBsIkIUpAuzZVHLybaiGGloxy6tn6gIbBTpWYb7eTGXefL18hM0A
148k4qFe/uPqs/7fPVogBqJwGtflW7TXnMI3WsL9K2rEWBTovbHEhpXEFv00lDed
b3NgI6A+/wJAzh3o3hLjxdyVzgmxyVVx0eEHWUk9fvy3cIDL8+mepsZwz5fjONqO
3voizqlQczyrHy/5JH+LOLbm7oa2pYzTptQW/R3huGlK8B5rWV9wLJMmWSzLKqpz
ELwEdteJp4DyoBJMmB9TvDaOqf9LWWAXyUTbDCuq70n2lIdPizNvW3q1DGl/n+hV
AOMvx8+6KTz6FGfwqE6T6NFwpNdCpdXLZdTQ48Bo/82SBESA5x1VRDDlSiyh8TyR
iSFNuRrZqbdveKGO9QjZfRv0oO7cyyL9I5ZBRjhEdYNvS81WXZB1Ns1FCcsO8X/R
GVO4DMKpELuzHRJIbDR5Mi8ACbB0Ue8anmyNEWRqH+EQV0DflSjO/G3bV1VvPSfS
NwqK0icrYmRH29NKQP0mYw/tyULnqU4f7d2d79AQaclsj0QFu0FoUi24yIw7D3by
eeyNReQnTJGtqF6RdaVPDZxBuGizF2uRNoNKW6SaDlQrXsTniPnltS7GeosmQqDf
BW2UmVrjkD79UjUHDKBk5QDYXmy38cvHar9PNMsCxSRqslg9Z+TutJql3/nDI7YA
tYXePxuGGarvCFy1eNTFC/m3Oney7v4Kg+4jseC5XwWgG5QsX1I4u2pr6Vif/QRp
fuIgmo18w3znzeVepJN6cWADLUln961D+8yoSebeylX2QZdsFqaX+/nrzf4j9jmn
FgqMmDKkuDwai9tuz1CpExHr68rFeUEflXDGl4zPU5rMKMoycRdMS8DhfrgPsBWX
V0caaNNBUn+e/Ci6zrzk4fTrYmNdzP++Y11XA2Y9PNRdz2gleRAvPV5XbbGME7bt
IEBQlzdJKlbCiyugZo33D9Jr11ilFoocBxiasXWEnPWlvjeTpJ5RFzKVmUngno2o
WTU47QpVTmI1KiFHHOyonicttUT2xp7BgmUBbZ2LWkTf24Mv5HUlGGLOoLsmZ9Jo
acfmqHU40MYIKzS2DBwJ049c6Aju2++xCt7GKRHj9wFPY6+y1WWO0NIRu/sKm22+
NRcNY6XupnYUlNgMazG5KFGYsvHW9xlYaCNRzzbDNSEH5kazwuYEKiMpx0PAanOF
NPIGhfXSv7c5qKAYPXTHMbdXSxVhVxFVxzXakXlH6CTgP+4xvwcFTg7yz47l73GD
FAqLlaVCfpwnSbTae+W/CD7jUhR4/3aCjNQplqkgyhV2UuowFd6yfoUD+87pdjhO
FdwqlqsPG+mPKy92JdlvGaFHws+fhYgU7D2kgW2KzfUJjkoQ7GDkySmW9H+rlmYb
zn3BuUuwCDzxGzBoUtkUQpzuQ8mrBUZTa3044i22Ykb5uDmTZrR0CXi4L7Gr7RFr
wUfksyb4AaTzhifo/99nlpzgoz74pYbYSlWgdEfhCW4Xq7vEOrNDnvqZ90YYuFOG
nyQtuTAPSy9BfuIYp94tZnipMBNuYDxJixwzQFB7wMHXtZ5P3YRRjkNEUWRZ+X2D
OjkcpdCphMkeKlPzFk/gULXmjDNnG7CJ/obI/GapZ+v9NJ4e61bvYwH3+rrSApJ5
35K4RqXsXU3Od4s+3nebyNilfFGQihz6UDaeBo/obGK+4U8itLl4mxG11OJq7fGD
nst58kLd3a29JXwhAS/iau7PVau8ZTZQehWjiVXeHj9n+5BJiL55vAITxydyTGyW
E7WMYqw5Lwvhu1y7ScMQd1LI1kmEH850es+jnKh1rGyAP/3NUNy0+0rdk01t4Xqb
CCoziavTiopJ0jKIJ0qwE4dZFpm1ORvaKOAQ9HF+YnUf99gqXqeg5+W5yY21X9UL
/2GPmZHz2Qjkw4dlXUx4I92ZU7GGbCFf4MrcIB2v+TVz42MGOR24S+nzn1zuF4NI
ThF90MH0hbqwWfI88B/tGMgF+IT4joOB2xhZ7MqtG2Gf5a/9KzoBvGecdv3k9ciS
l7tA4DxHKm/38/uGrcSDjDYP6Ga/nEMdhDjYCIbsICnaeC/CsZWaRAI5DQdKStiy
4j0tg2WpkDxfUvVkFLgNN0o/X6y6zMVvBGXtsTVT0bz5oOM7FrFpC7+gc+wFhf65
UwYO4sIVDI0ckTzazf82zIwuPfCVuP/nQ8aQSNQfQtod25ozeTqAJNxxmloPl50y
7Sim/nuoSZeYCFNxLUspyY5b/HTl3FuCNHO+uXplunfrsMbU0IFLXLRB3TuFik7Z
+mztohrm9J1st1IYI/jQdB6NSK19RUnJkudx93GlfL7zLaM/Wd/Qkh8zNiCUn8hU
nwdZYYcnf1duD2ojLeJmW/fy+sGKhSBSXy1PnjOaFML/o1mHk+baCbjtRmnM4GP3
Hq/RtCrTZS3nC73R6rii/foyj6XWj2iAY3dj961vCu8uak9cw631iOqlAHfVKmmn
hHiwsp54Oio/+knrMn2W1uvYmVvU4pqqA+0XufdaVRvJnuD5QVm0Pag0Q6oze4ZY
cC5oqzNb+tCy+9nm8KJwFauq+dE4q0gu4j14NAazQhgREp9QXdwySrodjGNbLDUD
LqN8j5wCFXLPJQ/+W1xMHWLayRY5gBahwAU3MGA/+mnC1AjzzLtICxY0r9C1Ke/k
Qpv14G6AFAoAk1PiAxeR8/2Dc56oZ8PO76a2/fqY99lvuO6HcDMJ195QbU7cuv3X
HVymJm4wbjwtceOT0YxXxqGE7+JdT9bCjIL3NBNTl0+VzZcnzMEp5QyrhXojK5mh
ZBlEQilIwScDccXASw5pA+HjitHxZSnt+qOjFS11p77yqlrzzXd8jnW3sNjYNPwG
+Iln/WtH7ONJY1iBSgLLk6Khsc4RQNGNsYKSw54KcGUzV0hvVNuAVpNMmx9RfNoc
CPfWk147C3xjyEiIKXHsA1UTWM4Mi38i1ncJep0bLwwd2uzQyF7H+lb1k2GrSL/Z
3sNzwaOflXMSAEF5cjyD/qYKfGCsGp0YykJZ8VqB0189HxgJWIMK0VuB0fMC4umZ
Xu7la2Lcvr1ZUK3AWgkMlx15nKwAILQeaPQ8//rVR7GMkEzLSpPJ0ADXKJd+l5gb
7DPzP+Dhw4Hb5GuBCrlkIXSTOhID7QkqNpJZnEMdArOu7kymr8gJ1e/+RoyZivm9
4IUp+e+ZFcDZnbGhaApBbAQXukhbyg5XHXbyrMq0BzMKkpDZZA2XZJbjVbWNDRIL
MSaxGs9edJPaEf/LMs7DGTV4jy6SV/IlWWx2lRpAXSBABDqA++iO+hIevMSpU9PK
/qfzVh4uzC+DB/rqRCpgG1PYYpNlgdBYQWKCSv0CQsEO0jHXAr57aio1HqAoB9uV
FI5rY1E2iVL4ugtX503FG/NpKj0gR+hGJBYDp4oMhSFbzn3lLO+rYPzBLKEqzevz
cyh1BgfFV/W47n4GUlnTjS69SCXDuvleS0ncNNNdKEwXPgvYIlF0OKEMJlQiaJsz
nah1iGYBkaAXwx1Y1YEIpDMDDbkyOnJ2uDYx6Wx9BtADBJC63wX5b3T/GxRQTHp/
Pmk9UJmS+PSEDd3MH3sy561TPOdKYS2ta3/vwt0BB4viCmta0vgxr3FMeIJ3wnIu
qB5qLEe3d21NZOmh2KkFf0U5eFPrUsYVWFspgC9AMR352WCfA3iCZzM2XltZmJBz
6gMw20DQvnXo8RLWKkhdxjrpRZ+4y6zOjE+oDjFyNNV0073PMLCgxTHrzrc8YRRT
QZAhwwSVfuUHE6irWWIG4ijvVJsBQwsprQk6F1eeHBQVo6RFwalEsEXXyGPMVSw4
c5e1VVYj2CXg10v1TXPa3rBtscRJjRiMMbjTRG4LLxlf9z6YqfbV2U8RlB+vku7P
klojZzpqbHeCkts/p7knvASgpjYndV92u8+dvmbWppqZ7oa6xBJ83KMZBXO1Yajr
XoacXHJhvczfVSk2fN9eN0Lh0bGwNTjnGU4TkHd0j2m2KTxnOoWx80q9wHEko/xz
qbf1Mi8AnEx9BwqmqpBobdRXo1FmutFa/WpYe4e3fb6zQPVZwIIOazIf3MYOX+Wx
2ZkBpZ+NtXJdbr6pghf/cvoh5ByT0PXugiGtNBcHjF/GhYdj0Yh42hP9WMgIo/Kk
kLjU3ueJxwfW0RugfarD3tUpWmvQ3R5DzYxfvy+Ny6HiXmkJ6wRH8cPzNqbYC+35
NFOMAdabl6IFtV1ds0Zuu7ScKJsfHIC2g0AhWbjdLlMmt49STK13vl9NF5ipQsHr
0SDEkWwaWJuri9So0hK/BKKUBhfmd1uVNpkJJqI6BY+5EwyItUFL1QloeIx2wYq9
ox6jSA+EW0PU/cKKnBHHrAKvqUzdwnIBIFtQDH8jNfHVB0C6kdUUjb8idNSDXuQ7
0V3vsHP49S20V5xY/nMMGZcBJs7uO7fjNndl9mSA/XGtUYsncLWb34cqivYxqA3J
OEK/F+4xmCticagnyCKX18+qm1eJMhuqqJSAD/METVpiHmcSf8V2RuWVNQSu1m9Z
Jj3NC8q8sCASpus/Ve68VFD6+QofT9VrXWuPnSoeuBQGnhiD5lD5hHBsNkb5lnwu
3Yb+YTUJpXFavaOaDWoM0mBGE6sYkb+SgY1WGXaXcDjWllhLGEQXeT9U8d9yGtAs
kMO7pP+jQDIM0OS8dOZCQD+x3z8Iu44VhhoQpgMb3DwC4naNvqKCH0vw8GHk8/2e
IZzaL1Ap3sgVkeuFNVrMn4TTgPgOx1QwoZ/INM1aviYzS9WcbopoA6qpJoOXrrSF
m17xRLjFlpIMzq9LSR8elFYxIh9+uFH1lY9n5s/B5oLbuiGRbrYE/XdFpJqZa17c
LI0prf5+bofLHONoyr8Kikm1KfGc4NM7TjHOEl5IeGJJ/hOcC5zf+7TejkRoyEN9
+to/uncMxvFogpaouflUxittCbzfffToDdW+Sco1kUhQ1CsayWiqhl9+zPFj1EAg
VLJNh2cBkAf6wzdkfQGI/7v9GKG0BY75emnNTARKdUJN4FeDBEXz+O34AtSAXUeI
yDPNwK6Yb9aB9dGjkqWiB91S5v05xyQrdOrxjA7x1nqE73kbIyGrZESZ5+obszUl
MLi/cZi8mRaTLayF8/gow2P5rmFPr/cxNuCQ23HYo1LRevkgAuEmaCJExIbjV13a
k0v8n5u7ckvZgYhv/ysadIFibW3J0HdgxrGjyC00dXd5tC1fuyHuGaArqFUJpWXp
2MyAoguWbUcpBGd2Bq4aqT78ngVvAjwWWzaeUheJ7vEVjY9ze04bkWQVo23Fl7K9
wS+k9abLNoFRA+XcqUIIcwiEVRJILhFaXrm0I0gP7zniT4rmHwKle+z5G6e6DEL8
FuVpMNtXHyznOabJ7Jh3t/ZYxNtJ87a4CffwsNSphRjdtB4+poBg+0iWf05Gc1Ol
YcpK3m2/ZRyv/pWv7jkiZocYLaduA2L+TuAeYg8jCntso6KYlt9kAL4R2iZzzNo+
zmu/dkf1DJG+ThbIIsmeIONKDaFv0xaq58odXTfU0kTKgRPrwltntBtpQo2dtxmn
B1CF7yaS8lNv2d3730MoaPmfwzS/549pnjYCEG2FjsCsH3KzpAAdU2OEH2UtUljF
n1BNCkgvV+FgY5IUlsLY/z72JzL5mJ5+cZTw1bH2FTrz/gDMN0GU1qLHkvPV80FO
0WglUQ/j5ipwNonnwV4GV7/qVIaLWH2h7jKKfsZhVd2g46ZvJROODozSuKVnWuuV
1SVe7mGMMWwSDOiCCslqlBnbZE7q6vI0vRPX9CDG4lR2jwpjXSBwLB42CzNdj0Me
ke35lYVZ8QfLg3/VCmtQim45Scrkl+OaFLdJfK+NxrEjEziGFfl0dxB6QW3A2QcW
BL7J+3W4tjmmapO3L0mZpTAChBLgz9qi1FhWNfv35QXqYNsWR3W18cfCx+XsIzvm
y7L4dwSAqhuSqql95da5gWKOqjOwUvWctfc3LbOE/f9knToMgramjvwYs1vZtWtU
EKTv/2mfiANR71XQKGOjxQjcQ3mC25lrX03ZFZ3sjGyQ4banSdZ97Ik7FaB3hzja
dRiuKaBo8diRdcfsQLaUx4MTF7cEnZi92e6LMk3Kn4Iu7fr/qgv3DPByVJJ+IDsY
MaguFiuGKHYsYNepMuI0/TdgbP7IK309k7xvx/l5UfePh9ejbAngA9fmXcxFAfEA
YeLK9WdMfZjhSz0ZOI7t4ktzRxZ1meVFPHNI8lRE4fUTNCar8P30UnIJ6oc/V+sH
8xguGhkaR5tG0pTqj14mbUuvVAtFpqpkTe1loEH/RxYZMWlOROj64ebDSQR/Nnja
VfowN5Ht9Bw7ZvpTf+SMcVtpL1Y25UUuZDQAiRATJEQMEvW/cB1cyLz1V86S8pbB
s4lEcms5vmMy9rP5WM5MEwnn2Q1vVbNEYtC+vNvZUErP90nLKstS+YTiNQKpBEhC
dxlFBfHeG5Tkce32ePui0OULv1iEwJ+7OQuS62manQYFAoZFEnK4g6OIX2l/mBzn
uWZ0ObNvqsHrX/6rnmpYP92QNa2shgnckN8/F8yaXTh9+va6bbjn81urC4XFXxhs
CxvUhq4+zhqayRnB84WJWJiTUvDPZVjxYfxs4uidmhb8zb9Vqgyjw29EEIm1lfHV
5pqb7wh3QFEn7lOBBPoOXmX4HfeEGRnXFiK8jFncGaclpSgWZF0fqKr3HFVrDDM3
N1QYGkPhbW4CYB3Qej8QEnseZyXiCGSfuTyLvzuWXpn5jqEJgI/SyKxys5T6uPRE
q2AINQU8J4aYfRVCyBRhV4G8ff0+K8NtKkODULKUv2KX0OrMnuD8w1TeiI/7uAp+
VLbA32JlLNzn88G/jJIivWPVfYwMz3TNOLVwzfIhhOSd0edXgnSNiE9Ouufd+E+d
Hst+/OtqN4hykAldl1lsK5pfjgJvxPxP8DZ8zCp6gCvLAfbCV6GDWB8zt82/JkxE
mhdQCWzdOTcXkuXr1bdaOlt8ItRhE6WOdjCg6KSmhGQAY4+tQpxq/I/kBmgOQvYG
SXVsuPRJ241vaVOOnbACdprSp3MyEz5sqCwk+82biwArBBtmhVR4zyPBrN+yI7Up
uOHdAWE6UYOuVskKJXBd6yAgixXL6T+uv54er1Y4CJV6x9BFhAWFw6/l5gFDqzQE
u/DWhNStTCSXZxiczrveQevu96099jNcWGhIuhx2clpmFqOWUzN8MLQaHjnx9EqM
G/l4/ZI2mdOTFL4vfGlJVf1akmVRQxFRkUQVfMHI5tGekfsysC9IFe4qKbY8aQ5V
ZmhKVE7e48cdsBk1RUsJenaMapn+OC4ocMsHlKi1vDQRTh80kmaZ4NuNpVhYs63i
Qp2ppLaZYAcJNezDwT5dNWzdMlpRURIcWfQxha06tZs68KINh3G+8E7KpghASkMW
jvNWkHxTTRjqgcRZV1l0TV1NdqzPSLOfTOHb5oYGHlW+FGrsle+ev+Bn1FqF1eaC
J8yNLwx1R1wm8POqSEqBOA4a800dLL9GSkTDR1Jg95V/ommmbAIIOrXzRcLK/VNh
uH4eCM+xhBTcsEos+PWmI0TBhvs/BFAXhK8PBoddSNvHllhNR9xYEjAN1LihkNu4
6iBQqT8RpJg+XzPOZjlgVwcCkFKco9Kykkx/eWFkrowB//ZjWfLAO2JD9lEGUbES
bi9tVoNm/b7y0lioBFmgfW4ebu6y1s7zTo2Tjz5crf80lN2uuvwfP0bWfJ7H9Xs0
HJUVEyqsDgBwmz3cKknFhQRpUMC0NU63PgiYnRBmVoj67ntJ/YkycFRtP8fxwtWZ
HaMgLJcLAUcHNuQAT6QwfBJcOrRXLL2i13wZzBGhLOH/wXzGl7SEF2WCumk6nszw
7DLK1hF2fF89BUVuAf7yal4cXIx8M/HZfhhJH636jTpSxhwdE2t9tmkrs3XB+w2F
MPlJLs6SPk7gOaDK1lbHwuB0/pOsc5XSodxjV45qnakTZQq5MuVeNVTouDNVWD/w
PWQU6XCy8FQYVM+bW4At5k/AsxrlPBqSbVBYzG1lkSyG7wFWyLeJN+e0VeCImhZJ
Kl9AFyid9lw6TgPIHsLRQrOMDMwoD9dnF6ItueGZwuKmVR6y1tSWwqjZEM0j1AuF
9QTM4ptjZlsnJVdsU2n1tkU3CuYp7W8XpYdDJ2CxIJkM1JeC4VZEjlVBbRtgSTn5
lAug4AOqpxPn7avLzeBDMhqoz/+dBUjd4u++MzMRbXY8oTxZ/4XndJVH19TvY9HJ
3G9TlAzNL3nDiBf1HH1m9NRlHDDPYewEEefMywL3Wpogmtrroc2wWokB7Tw2u5IZ
Fv4CskCtCd805M9xRMbWihHqidpQG3MoiYrKgvv79DBq6BqGWcQ+fkd/TDeBkbMC
DgtHlMurcBLCOBWvQM77O6W5NrCDsGIWq7HaR2Xca7TwZGL4T9gHoe6qhQnwwXm6
7H00dZ2KQnpTytyuMtLKKlY26SW7YQCgVjJYk8PN0du9nBplalxJyfTWM5DBCxvX
e3BTxTYLBeCS+oE4kSVuLVQXSSXe1mL8vDg027MMUdxwSFwa4hLV0WDeNSMpbwuA
CU2U9XaN2QECkZMAhppJHQh5vpt14V3CLVL+pzmKQc/5py7VY3mC6ed5NqgrttVv
9eEDkmdV4MHOFtxnqLSRdocAsX4WdVlNLiPdpyr9RnCAl7lUxIoSzOBDuX0yHwoS
T4N4/YN5wGFYn2QFwjClMC+e2Wtpcecr7CJhijJMYW44eKMXhkNXVpN1xBFrHGGC
zAeu3uBCpB7qdFYlNjyFX4eQxBjR1qnOy+UR/RHOcQj4j9vksD3K27ZujhTCAZZn
l0OQj6ZFVuOxtssw24EziwYLLYZ3Vyy0FPHY/2GKE1sV1Etkh9M1R972rlERFSup
A010w9Y5glO7Vr7qGhjqXaVUTaVNZqALQ8TDXxeeLcPaURkCyUOdzLM7aYHxmGsD
R4Yq9vbGAu2deo0r+Sz2gB5fRb2bmWRV4cPQclU+tphUHhvu7pezLb/hGr3f70dj
2OEGnnsvVlugzCzj8JwxNnWKyZb9JJgZuQMCj+vB3O7DN906zCW73a1YRUS9wbLK
sKUHQBwtJmpGWl7w6yAqsBaI+gNnZgQl4ydkvTSB8f72iABXGuD/J2qlOB7Iz58I
Ss7v4tQL3pYv7R16Q7t8tewzabancXuGdlRo/EU9JnF9pOyrJg6bKtU9p4ni6JDA
zmTnjFc6tHjslgGPg3lNxfnojpAAn60Ul3XRKylnGHTW7qREJSno8I8MAOyoNzix
X1ZaXycbTdMZShEVR+DSN1ZG8Lw6JaZfb22ZQ1iTKhHH1krZFxr3zw2Mu98xoo6p
HBAlTKtndl48kClPUMWSuEIfjEm9eYk146zHLakLjjpbeEU72hvcVuC4aAOwkQL7
uh0y9z0KblpJfshp8SxE8G/yN86eLRER/HPWvKl/0kppW795uCXBZEDvl1CA/Y3L
kdT7h1b08LmadFQpeehC8FC6atXr30ERXY7KtYcQYv3rFEazMGp2onyAG4Q+JEfX
MGzJSr5FMsSO7KnAK8HKVDag9hschrLMNEwwsPQx6qADcWOAPsyzFsW/C6VBbA5e
2wo3pUp9dX580RwJcJudfsFWUKY47YFquNp5nyMTdaMjcfS5XF8ZWV2A6SbynCXU
ID0YqJA3fRRL7VromFR96OGlAZLaWJwH2Zb/HNJFsSw+y1NV/5z9wzyvSNRhWHcT
/g1/QezQU247lGW7PYEjnjtFwyFE+A/4R8PjsSj0hdIXW83GTyq5Yi7cyTFjf4cT
R0ZtyPscb5mwLPqFpszV2VIrjDooF/czEbskxfkPcIGk/41dNsVaBSfvRzEEQg1o
YXxurNtaXmhLDZgS/eWxcoVDXwwOoq2th/B4b/mK67tZEYwUvml+aAlJw8iFktrb
5to627wPpM5Ux3ftfNGNfzxK40DP+4C/IRPk497Mch77c5Im8knSM+lZOhHKmI+x
6i5SDSr1n6NHk0wc1gsGqVDExejsgGVOfa/SHuLasdnUjwoxR1PpH6jpN5WhKfSq
AOpGckgrfg+Ki3G4RxswpqTAruA8r35wfBQ3kkDAmSznwnt1CZHqgO9q8ilPX4Zs
6O5JWf6zwNZUdQVmjL6cDKML4+A+vICaFEIH6SmtkFQgzoaUsm0UeD7XtK0WeLXW
Pu7KiPLbR6fTrNT9uKpc2GURDISuxU4R2Yfa+/s/BiPQQMuBy+WwodqcqWFjBlTv
PxY762h2fH4f2Yh6tBY3Av2GttkFNziosRDQ71zyswVdtrvUd4zVu506iT0Kj1DZ
UB7drctl07k3WGgaqIE3K+hq4GB+UVWneYNeqpM4YyFx73bNM5wgckf/I2dnvuAf
+23kTHp9O1r3GfpD65soHvIuSX2C2aQQD3yv2IQPayFxhghc0qLpqDYe4/xFJuCc
lIUwje8EpgpOWpslmEkE6Bdqpuudc6ydmNmg/hKunuqs4zzrJNISqrZakiPrYJQy
uKCyJOms1RZnWLivtuboif2DcmWWmSgbMJ2HVyUcQUHNRSLIY6tyxJwg2Fg9Z5c7
aXSEqA7mHmvK+5zJbHAY/I3HfcmOn69Ke1O+lOjf8sNY4S8O42dKAH0A19Uarfia
qZIT9MKBWjImro4Uu5qJfRAo9x2PQW3auCB2o4XIl6Y5TGlwAGhyNphlHaY+oUSB
PS1QKW/HkxbmhLyYNyZ40xIaZHYfMLXBnsvCObNZl2hZhBD5jz5tfX5Eh7DjNBpe
vDg7cv5USC+wfGhacjGQDoA/jQrJ8sxYVv3jpyi78dsiaLmwMzGA4Ep8sG2x9DBi
G3OArlIaACNYkGUU7O91XKX++4YGwtSd2/0PEw3S+OgKZbRIUWd4uLakyFQG/2IQ
BG/qsX58yU90iDgRbaaJQl2ILlD21bDTAfo1l/j1IZ/LjLMHGHh94o4FmBQsDyd2
1ITWUL5cWY2BZwvEa0lfsmiokxrSv5q/L+FxoQ5Z6o0I/045zbxG6hHhAFA81neq
3Wb76UETO68N4kkW6N9I3AM5fHp4QIXSYKZxzp529RjzIYFmsCz+gkIDfNfedrZs
WkxzkKcmnVTSN3U2WdzZEmkyMAKcOhav+ACV7WJLptrYnqUXylLeiSvdhrRLldgZ
0920cXKm8xeGI4Zuk0pp8PeEK5fzYp76uv3Up+XaQaUmV/sUXPsdTaKiAwVi7tFK
F5TRy425tUMbkbXuTTAqOkQQETZuEkMDxfbFcRLVhmpFpYwQjHXW9J1Oue6r9Alo
EHAVuXgn5VcdARbIPqFDD4j5Sf7kUrlxgRUMtAX7Qkrvx/3h3vIubqYkH7vpzBqJ
LH1eaxo+cEBG+v/YlG66uFtA1YU9jBGIN99vrU9+edOhbDP2HkSxwoaFhEKQN0W2
4v07uC6svtOygAecv/XOU/d+yLo4B+iJk0Iw4ek+97VZqpobcPnGRlPzQ6i6m8/j
H+At5t3tp2mEfTKIPFkrvnDtM6xUz7bktt8lJmXM3qnL9+C7dWJha321VlmmDDFA
lR4EIFvcqI1F87WlI0dfuOTdjN91+J0F9hewISKyFJUM/kajpOcD2//CrjJ12DIQ
hX3yML9wUXiAVc6ippnnMKP6naFT3i++q8w2kMwaRqn7AiCf/C1udO0mBlpaZm1H
TWawJrBzofO6UXmWJXYFln4eAP3ofw0GajCnsvaf49fRcomEVrFvWz/h9/1vBynd
Y2DJpaSQ5nU1KKKl7lHjG9s/R04b9RUxpsJHOu94cA7Z6LRCumTvvJ2KUny6EVjl
ECL5kNOXXmNBodf8K4SVosJxQb0PabKMV0ben8P3jiKhtoUk5f4DrqOoAVlIRGPY
oo05nl0GAXZQhoKpEH69acXdTZFil8MiE7v+gbWwnl6kGW2fNR2JKRy32/K1p1k+
KIC8TMKb19JwRghzIh+cQRorIZFjN0aD7nBDNzrHrpwUU1WhqYV8//+Kfa9Gs7GM
dKqP0cT+q5DEpF+iQuGM/6hzRtMpfCRjee3dx6BuyI3L6OHjjqXEMRy+Tj8Z/zdm
IHuHDSE+sFc0rkT0PXMwvtP+ubMFIDo/F27X1UDSNcTT65lST86YZdTAzLZLyoc4
/0ln6JDynhvmvv30S2H1XQaf9ThIcObaMZ0EqqOjLJRUss/ThWnaJQDUhEZNdrSp
pNmt9MxUsWNyhII7HhsigS2cKLA1HkdXbrjQF+/lvTpnPNQbz5AtE3zmkPF90kKc
DkumWmmyS0VekHUKnSOIQROYXiGq74b0ouJDuJ/yNRJwirx2oMV4u8JCZRmTPqKF
CklWW4B145XRFmSMA/npggKddPVMr5AkcnViRXyjxNlP1x1e+khDEc1dQKgYn8Na
AKevlXc7TaNbqWLqPR6XPbrB3eY4RcOSyFRkrvNje8JChE4MggEjDFq2aWiB20mJ
dw6N3H9+MZZ/TL2LyjhMmlP4ZQJ5UIWHB9C1X8rY4A04+sWA4qCDicEP+aFyK3J7
SmR/vSOhXOU0gmCjGOmxyc45kuBB3iUQWY4YVnn97rZ49s77yxoKdefDulbehFsm
A+Qjd9ts43Qo4M/6/ootoWgxfbIQ9y7OwauzCJwnrF30RgFN+OH4Ouz1IQ0dePEV
ILzatEAlMgw/ZEYNOr6tnsb9WMwDZRN4Jol6BX6/r2186bJx3TQEvHDxrXOK3+Il
FMOfYHxUuV4I3bP24By08+MmA8qlyHFtZ+HrVuspRyng7NZLYlxiOIzvMPDCUUzs
aEtK2mQxTPW144EGJr1JGg7Xk7mdVvHKirqRxOzKsco4PkogU/845dlf8MsF6IaS
kC09Utle+FAndetUYIVUu3Vx31Z7H/94ww1hvKhhOAoeXpirIYoANboMO4JkWvg6
7P2zDq6uaodSjRl1DdLMBGC2lRXQnfWqv87rdKvDir51a3/6U2iHcF0jUbXIiIkf
DH++fGshJMM32KkQrYyBdJendqZmB2SJ7DOER1CJ6PWvLKtghPyn4jRflVdG2+zw
ywWoo2fxJX3yUbrCAGUsGanUkUzl8yVNYuLlQyAlhT5BhK+FAQueI84qhauvaR0N
lBXuquruxqdtjbun1UR+elGME5DxyHxSR0jHE4R2v/OqSuSo2TFnahLuhUXccWLf
AnwAnXUCrPaHjuDkYOyDUvur856WTeNceuLMrzRrn/aNadWDa9YzHrdN6sd4QHqA
CI6Hs65Lxvg+ARx7PQ1EahrwYFtQCr+4MnTjUaQJSnhAu94/H9g42bsxaGg3rSEu
oII67PwVq6pJW98WFS4u92EfeDTzYVSmHftZf9sOw9JvPLkGTb4voOeiD5Gzxf+3
oMf3GfjF36EkfuzLslkfFWG+9Wz8OeD8Yyj0VA4THRJlZ00laszapIJBVxTBYIxC
D5PS7JBquJ6A7pExrt0x8mXJyn5fqJIJ+fGf4eFWeS+sgD1QGBLnDbYMZpQsnwS+
zuqY4iDttjNPpfyZQvCfOJWD6tejqQC7HSe9aoDfjY1jMAYi5M1pXscSQZPAn16x
0tOsQfJpr/DiE03bLZc9pP8TlmKXwGgqnXvQWX+fv9q0QEOER341RzkmyJ8RbeS8
nEVhMNLi6DlnR6T5FlcwP5h2zSVHZnDa38MzhxHaLHIe59pQjB4gdBUyc9juTw/0
bg/FGFbiN5j+bW/fwqYNtUHQ23cqnYWa7Iaivlteop7Fa9rh2hkClm2dyxsQ902C
EHU8SME8mJmvVosN8D1M2aBj3Gs/7FbQNoIxWtD2BIN3rINSPwlDVUnfebYu8DFh
eim4Kpk/qqPHpHKLzmt8hPmdV0BLvgravPPdIhtoaIeTYPpwnzPC63tFmdkWmsrE
zes0EjvO6hJeuR4mO51IFi2hveOugEk3lilCsoAkjXwxIZEIWRVCI2fOWk4/DpMO
0wQ5l5oHF9k5OaOgnka3/6l+2z3uyOuXnBBg3yFvtf/wbZ+k6VYUI25CZtxthER8
Z4XJK3kqHv2t6tDs3iBgGau1BOQ3wjNA6hWYxKTVW9VMIItYcLq8Jx8kKXDHoVbx
2cIY6pmUL0z/w1NgxBI/k/fFk4febWdxJ4LyuA3yrPEmgggDRR0i3NC5OeJAZhQZ
KI80Syt79oypqgqiIaraBSwFT4bOJ7Qh6wasor9QTZDZ7PEcANt0G0jyngcxINlM
8+NYsIiE1H2B57p7d6a0gv2Mqlhqts95jbHnDHtwsKEEdCmRfOcU4CbrseNa2p4b
ZTopWW/kWlgjFP1bM0D02+/UZo7baiGkEAToe8yOp07yhrrZAMsuEztXzGG8gaUB
9DdCpBwpxrcxX1zt6EfwinGgYZiPdvJF7EvT/M/JEtUxfDI7EXYn8wOtiG4LPyH/
WR50tU9s8BjWCV88r3TEJ+4r2mgiafLd6Cxgw9sgVOBXWlYLIRGXSfB+QBHSzhqd
El0vgwvl752TCpSmOGsrM+FRPaLk1bKYjvLvOh/V0mwO+7QQIhIq9iHNFNrCVg4w
W0CkD48jxiVyXtC8+VXhjlEHI+rsoxHpfMx7L5UZudAA+gJJDLikYrRhztBwVlBQ
9knHSM1PErpzFRbh2KgneG6ZyRoMjbCLl4PUAI+wUQoQmvHz223zdCouj5mukCpb
8UXTXOlaWnq4mPR6bKtKPz1O/IMSQf2joKXrYx/u9mDYbRF/s8arO1gXSoFmyKeK
B1V7ydUk847VOBUZHChgEXpHoYVhRStNx3DAUshULR9wvA2rUxYPNlU0l7iVfsz6
aOuvx1iPVsbaeXsZXhrSqOpxOuUsAGLXxw9uaWGlaGlUSD+YXuhEiNvvHj1ILSk7
FlSOJ5wDbmTCoJJeOKbcvnbit0pKZDQzVPNaigWZyZQcQlnurYMS2kUBqJBkv3P9
S5UoJ/mTlg7z2wpuRdJds24lNkIyblImchTwD7LDCkiZCyP782IaN8feP48AdG2Y
ScX4iV1NKP/znDPAWDsJv34FlgEcwXLI53aLfIKaa69ey2VCnPXC6gCNPi5ErcHX
5Rx+9jJXMzcMApFBkQHT5sBqpylI3JOkbUAzjjcLhEH9omMcy6FI2l68XQhpksIM
/N/GyeXxkm+ugJX+DlgG4mOYypOBRsupf7Q3yH5O6J5kxkzhz/wpdXkYdGs1EEbv
3Kf6QP6qlDxzZijxCl3WJlwJZY6WiDdQk5ME9y+kuFRfo6bEZ2zzr/PNX6n/Oo0R
YVq2FKnx9m+PWn6hbDyGAJOn0PJacKyQgzdPLDaTmMdTjs0deDxD9dTje9gUdZLl
fW3AZ213HnvED+4mVmHsjKWPu+SYouh5uf40GQKrnDSYhzEIy4rz662lvdJJeH/5
O8ogAMU4qCKs4OvwzNa9WbPaYbqoOm+gq3rLG6lOcv58h31k9X+LPScm4kfyh68o
3D9L/IyLU7szaMiM/FXlHQn4qbywjLJF6ZJQS7lC1PwJ81YweZu8xCbqVyiL5tc2
LcMHLqIVq/CCO8dW4Ds3jYe/9wDXktqzNwRQZdMi5kezZg3lVCYkaLqzLEJYhXE+
3JVgk5Hq+xGVRyl9fF9SC+7wgwaidIn2hPk7Z5rDJgXNVn8gyINUayw4RGAK+9Ee
se9GAy5j8uv7tbLk4quob/NRiuFIKFHR6eiFx+m+a6+nDLPngKPypMoqmey/Jbou
LyBUPlXY+7+J8+Lc4JpCsAqwrDVrRBR9Fzcqsa6l1B08zBrTDMQrd2v7BHOeCFlV
eV8cFWWpBhAnYM7pmJby6Tormf1W66I272l01bnfiYNdxJ10drdfnZKk+AOHW/tT
SplxdaZJr1py7xt+TmuIzmeCstBGabKioSEuny0QSDaTgUKxKWyBnJEkSbecxUym
hPNWVmjpc9kQxJe5xeCKQtt8iDMRp/xs49Iz0tDjDpjFvfyGkHSRZ0cR3IwpKyB8
10dsoOVmWV7SkKqC8IzBn+LxqveN6bO2Xz0fhY/e1udwfKe0Gb7A/9F0MdVc8FcH
GR5zkf9TM+I3UR0m7zHUtawJJfMU2dsCkdTpHJU1kQXrY95obDppyzLaCdIlnc+O
mYfmokXJJ0QW6Zfb3wtA0H2rU6wi/Y5qN0lIaAvlnd/lxVRNxKw4aNZboXW2yGGS
i4gR37s2Fyb6Jk7Vqyy3sZ7M4pve4Sk5yO4gtaajrRXjOKoEBpFi05+PX6dhLoBj
15/fOF0hvGe0CfM5ETGToLElQX9RQaBhyFBozlXXNV/8J3IDcIpH1HBAhlGMM/HO
FGtDiO7jgCY35C+o7ZedhcqVV5oQJIUAQkYYPylO/uw03zhCO2383inWhOjIKlr8
f4Byx8TLxnTyTy8DW5xu2V/1Btcuj9pQ00eAkkVuhm/ejFTyVV599HHRDPeNI4+M
AH8AZdX6egBy1gfEsXRJe6n394p+7PdF6Pr1rBxPJ32mG+peuObf1kmdc6FsJixH
voPhvs7BFD/xAgS7u6qg2OdgmqkcdFsOlTUfQiMxu15fsqJmmYZMbr0votSF9u37
o55rWZ4yFzBaE6slSOAYmZOBnIHwEhBkLt138ZVSqt78Ql/CVuMAQYn5Lb10YDe8
3k3atNOxsZHjgyVhqClFahYVji7YjC0K2TeYLf5WqfyiQRhLfd0wTJKdkqR/kTB6
YkZJNDUcjV9snFKGbM6+svM+ITGQHnkGmAIf9dFp8TX7rtLkQVvTDDqbj5LS+r0o
Fjls+9OTSSl097Q84zviGSjeBQqFN6VjRijcCXsHzS0fgGbJIo5oNl9jcJYhpB4R
0Ltm2a8KAgookaL1jREDS03HKtHobQdvj/q1lv2O8SDND+Ssx66L3wiqPITQ/dJG
HPLF0Ta1xyKxU5kUfW68sKEzvwB93RUZydTDMT1Su9CgyqdDmIP6/yXMVBqhprks
cmK197MRg/vABHkTylSHaG5rv7soyxrMSq1IZwkKf3hgzJGhB1MNpyqubGkHVD45
nQRav3uxsREW4hWe5kbFmi6fybsz6e76KciK2ZUjjX6DTyQ19vIklTBP0c+Jw7Sd
UcN2prFU6CJYrBKX4zvOiYpsLeStRbG1xhx67/9nzqjmjXoPs22AhyVJw7NuIniB
D/XJfAqgkuyHqsVb6rRIsWcv0tmHNujEhaVg//+Orcbnd1inVB9oyV/gSjUQUMrr
jbBaFhrvOlj2dBLBMhfhhFpO6UTCBwDzzVMkGkfjZIST4g427/ygskPNB1ILHsM3
At60hVx+/sL11imbUFLmZay3DhVvFzGt8MM3mpQel7hle5ksNEAfhWMa3UixiH9K
ZpHIuw02mBpmF1j4lXGFvSLHdudhIlF4T9OPjxRHxBPxAVB+rEW0mwTxuLK2Ut9R
06nEgeYgiXQheAOnt5ummEj35+q4csoIxBrdHnrO03HxvkE99OZJHk7JNKvcHifG
sHvFqRszTuEQcvd/D+4yv+mMUD6f58dk9P1SXrlrNHDmtIhcR21C/5zH0YoENopW
OA7+n7rNNKdYxUxUwmW6XdpgRkSoVsOl4k0NEkYd1LlXATY31u/OGwldf8mB21+0
+DihTHm+/bosNa6vrwT6OrSckkqmiRTndxnCRJhqhvMUAo1Sr4Hr5zqv4DwG+IvJ
c0wVR9OzNYosbO7M0o45akd5V4OBJmH5swc9PWGFporDX6DzDM3ywWozkJxeGkWg
QSwZ0VotZn30ZEOfavukZpwDhaG/BpA7c5Il0WBIK1wgwE8q9xclyMVI2SvMGqSU
r3plwxCB33an088bHZtlCJ+DSfG5NpQtj54wte8g5iZde5HwXXxxSfF6LnF8jFHl
SdUORVAjp8qLeuflD8nV8/qRT6ZF66r1coMm3baln1m/8ATTvIQvlmmFWhdegr6A
/Jcq3L23YtFKP45gGGzaxgHluopWa+LnykpkHi+kk66fhPNLr+Yn8pBO6tsjrXkW
KAUelDnon1chioNM+ET+d+pF07qnoQIwdWI6/adOW4mxASK6Rd2T0MkrKM+lY5h3
3vWQKLIe9x3ww474wQVLU3BmKWmjo6Zj2jqllLqxGlG60DC4f/1TJ8OQU/M3vo1Y
mnfsk6MY7wh1pzQdHwttbm4fBROMZ1R+JKhPBdE+mUtR1wB8JfjJDIX8Xy3MeANT
yXV/e8h6m/luyNVYJYaXSCvmbuwcRpYUvyHgx/452mE58Ix40cHmJzrfmWWKZAm9
zjtqGnB/+aSn9d1xHxhHeFCe3R6aR6f8qphQ7X9+g8bCgQ21ptRi6S7WwOWysHgI
7Ce4CNjMyda+Fyq6VqBBJp2bbtGWy6kRmCqxcKfPNiZQna5G4lt2yzUxvUEn6w+z
Np3Uapt9KABF0bZfbqW6SDl7MEKAb5XoF/GycAi00KroHFK8+vYfPglj4FoNNZrD
hJUGXld9OOWF3jxVDLrUlYXpklZzb5oHogTeXj+vjK5lY1i0JV1PCP3g2mUUgJXo
Fx1pp4qH9gqKpkHqAsPXyV/9AAixHUISXrhNyKPvfxpcLfazYAcvrNKQfmPFWLlk
rWRknX1F3nhL4sB8mimwg6mPkeW760U7TWwmn7rf4sKFNM+OboFxmhAv5j8Pr5/M
NeZ/pyeNZnv0lH6LzmVsR/RiwkR65iBRGnGAr3tOLAWT0VM3IEb0yNMdWu3nxs+k
j9uN8KGJ1sKwrEgSKQOaNu8HKz1tIA7aeQpYNps/WRERtD+e23myheoXFFWQs0mP
d4cFZ86fGB6lNMUD96ilBZS5EtMTtEnMVvizHxr8hxSPqzvq0wUd+g82jGYAQW1n
ok4FIMzYC7tY1M/vnRx+O3jwuj0a5yTvXBIQ18DUFpOwpIkZM5//o0LNClItZwka
PtIzu9eGjUQZ4QpVDkT3k3tKumj5w+KfbM9q0Mpq4Zc7F9k8kyhR7ximGXNR1BIi
cVh4ZzD/7LyzZILnNfWKWRs/NmWHgx4wMFNsSyd9jedr4z9tS2+tm+O9N23ToN/u
jtGm2B/THrpkzF4/Dq4fuT7kspaXjvK8peMtFZnlfgY/VpIWsZpRUufYrD96tX76
DHdutcvu/jZVeq8AGjpaV5Y6HemsV3vGfI483fZs6KJIPMU9xvluWQ4znnbFzdLw
5X0YR8VPNfCjdcFvmJx1cacVnzJNhAkgIosienVcjVmLG3HEa3zucT168NJl3pjc
wcvO+bwn6OzATXNUh76OJT3WDMNAXcqBOkWbT+NMxML8L4uBqPPit2GFfQ01PBng
3CCdyehYDydKd7bmC4KQZgdxCwp4vaZRKHrwvlA2ZLh7HlDJzwDdOwqZDodi0Gzm
Ka5PhwK0Cgzl1VQfF373+r+TGGIdgB0QLT2+zHzyEufVEjlIu3baqGS0XlHdnkxK
2KDVq+5rLkEuSmLGJwdRBXljD7FG2rcZixOMouDN4REfFIhEwTp6CsxIQnoTA0Jn
wcntm4T9V2Aq6eJKIiGOPeEJnzp5a/aIN625WIL0TjO9raMwSkDMGwoHHQCnmb5W
QJMGDeJAflhT07FvhLaQRhD/5QYGlUROCwZ3LZuBUAAge7cNSTvqu+vKphjfmGQ5
Kv+gq8UEKNMwAOzGEibFQ74N9IrOBxIo5pEAH6bdyqvZ0hJyKN3XSUYA/rHFJvV6
qDPpfcVy1sVk6AewbRVayu+PSlOt7NuS9TLCMXgqS17w+Y8QwvaAikOHJQ9uiUJJ
z+UdKzib8Sx00bqZRl/WNHyrl71FZxwtOpeP2kSm4EBULE+9zdQrGQKwClZ6o0Wx
NoccXfzbreNK+gGUKIOGa2u+2YzOMMjvQ5dXX4vWSQQoZwlj3Fz0NyKwEPTjvkX4
opWFQVPmJx6YcnPd3QzyL7jzQbXJkd8gg3s8+hiYZYg2UT2mYEYwKGV2rgl1nGKu
O3wTPA+zJoRmIDgpoiF/eisDXPgjr9r4Cm0EBDV2nbmW7R/YwYBaOYs3LnqXGTcE
GhNdisknP8aDuhdkmvYOucogADiLTHDwJ1iYVqM51sIp2GjsCQNORjBcczTHbkDI
lTu96aVcL05fk3BZCsDtSWKzJGj5Q5l0f7pRW4FYLBRpiEA6vmJbAYH6F3zH6IrS
eS2c9Cxf7cM3Pv0HhwL35QwQRQpPaB8ugu2mRdYXR4KETrIV+YZozj09PS1+rE5x
9im3PtQDah1Xjws4V6r3QaSc5ea7gIHsYPvBFa23m15taxm8wUVJEEUUEphhLBNU
v9ZxEHAgFicyAEpSETG8/zbe6WcbDSTl0HH7bOgwZ81gvsXfokbKqq/YZJoioMtT
FNCIbZNC/HdhQNmD2P4wCY6W/11FtI+3lta7LKPeddWlfcs1HHWBqQQ+huuIFFmW
oyA6iIHjy45q7tGzK/XOsJO2lNknY7hfZiFQ2DHW4gig4XlV7YfkNhxwX/jEq5Ue
MJgMo9mMV30ycjTZbq9hhni0/2cqMNs3JBzTURZgDRuq4sfPybDxjQcpOXPu/AQ0
A0A/iM/iepat7bIcTwcwDux4bN2JlD/sI4mpLYavAKONgleVVb8h9JYRy6aZ3vd3
ZAuc+/dpC8bNDISBs9NgqfeLNn2lKOOodzecIT+yxIc03TfSOwpCKC6HS9JaqeXc
6wmt+oPAx+0RKpgPguytSn/Ty+Qcmf5EgsodDkw1BvugS1qRoZR//VEb1cjh4fYj
raCNVs8uCbRawdCTMJ93cC6VrYwlVIBLYth4Hspn2RB/p52CwiPfpacsjnBJIz+H
c0IizaQcuP9RceEW4WEZQgBEpDrJ/bVz6ZhnAVL1Yw1d3HuF5JgO4e+K4ikc9qEO
SqbveBtdL6xzGuyUOKio/MOfxMM7CByBfbGto/n33YayjSaOd3bDjDZrZfQLJOsj
mveExwXvC2lzWEzv8Qj9ZRsM2cJeafI3oD88uE/er6korxIMq+2F6L59TzHCbz+K
EC9K0tHv3nMdfu1JQY/28eXB4KGRv2OT2Yfg7Aocx4c+OFtDnvSf/zsbNg8HduMs
BnRoxcwOW3MymJlSPB+/4rJrYKubpObTu2OfX1V+sAxCRqQSGrjYxz7naOVW/bz1
90kUbAenOt8EoEJaVkpKeqtHoONxb8zTDWl/14WO6zJeZvEgJuzCpfHpCiO4zx5w
lMX2YppVDz72BtpjoB5CZeoDUKMn77IX6UJzcIxMLY1kJ9NFDuHmrX2I/v4d6GkI
1UPieiZozzDb1JZxNoRpMd4pcoXs9zSLX3ER3BcrDsQ11S8DSYXNd161rE6bVYAc
vYOOmW1/+9DpDEVrHKG/V8KZBCzg7mPNkmCDoyMRgCM5OZD9diz2pH5GsBvd7Njc
PPp1yN/s6ZrUutHpf1QDvi+gEOH7qjmXT8FrUoFKNusny02kxhUb5xgIFOheDT/t
sNkyUYrzUhJNOazqOT7pmMMSw521EnUHScWrfyJdlgOUR3mdDGwT2yfuoc14HGmj
1w/te/Ku1RSe2JvylW4c9uaNYqrvIKaiw8nnByj3GQvS+P/oMGsuQHEzqreJJRaY
YFWiBtIXbu6U5Okiq0yBpIjMC46a/Sm7PwXeSylxD1TpnvR0LXM8tgAGSC3Z1N1+
/z2g0uA3ST1Wz4ac8jYIM7WN256XnRtZSex/BYF6NzDAqoZPXqh4ymZAAd6uCkRT
XbOoeRuZXdhiTfMR2c19iDc8JCeLtyA4qI1P2TsdEJD7TVVCsaHj1jrSL2L9gqCB
Gu/Pe6AjRRMWnq3Lui12QJL0CVmf7ehHLoXcEX/4FovjPDUA5A2AeI9V/CSsyicM
b8cu21QnzLobli9RE+og9buFBUMJcsPpSCt11OEQfrV8YbgviW2MR4n6s0EALAf+
pR3rV+ZhlXOQY1qDnFSllV9MX69gy+SuOVHVFH368b/YaENP6JbCjEsORcyGpUsR
L+8+bjXh2apGty3YZM6SR5Rcub8K0Nkp0RcPovLzIbi8uq9O1PNWXhDibF1gmehn
/HWka5hFsf8FsQ0OhE+eQAllg2JLsUWYtS1445GPR+sonGurJ4eGzwOCAFxYH6zy
xIyjrGOQmy4GcQfIriE1ygSfLxOY0J2Hffwy01aV5nAyHxKONGtH/BAZE2EF812h
by5L37ux8FMtai1f0YFV/nAwec7jMus99Z5xnkFuzEDcS3bHtxiMaBiTamRn4DgS
nGmKfLoOxSnHCGzV9k63ipUWFRCewgizEFQU7kZ0lijFnK1P9wHLBDVW23p9O+7T
2xi4E/RB3ypGBN3x8iD2lCTFrRFizflIQ2mFQRb1MXvHegnSw6Gjb/TIMXB84e6T
lyHm8KWwGp8jv/H3DunhYERl2OCC1WRzve2ElgIEEdYOv44AgTV6rpGssQ+yqGEx
iE88+DB/IaCFSj8eCdujDc30NBGfxnRy6qAPf2hvvMcFOMAFL9OFWvwlP5wrdYG6
6gJ0TN3CCHeOYiNjwH9VldqctYxcjuTA1b0/nvDkj6MBgYjhLNWO9KsvWafDk37c
/4N1Bq0j7fPS8odFIDkQfPkj1vYJFOrbtH954EtxxqjW6mq2Zvo22A0Nbpi4xmMH
nrvOnW+EefKixFlCvt9iqgfa9l+CjCu4NqXAFakAWCid4p084v6bxCAHf2YkYPAR
WfUp+dk/rOJK0i46majTJrlNN3zNSwilnaFPyl1tJ8d18DqGARDahdx0U4kWpm+8
l0Y7GNtr+epa/K9Bql+2kMuc4N50a1D60B4M+/DS+c4CTP+a6/Gb1r6/Mddx3hbs
DwKCw/2dO1z/AJkk2z/ae5YSMFyTF6tfbE58HFbdEu6msKuETaLj1wWe6Momlk+t
w352A71USuCaiTS476zx/0Yvx8R3oYy9F86e+aZRcmeKQqKOsFVrbKSxSTPpU83A
DhYuKQsi/TrkCgq7lGHCPS9DT8dwR/K5JaI3zBPuMPSX7rs1zUbBJmQDFKrdV9XA
5S97YO2ms/zTUUm6niz3ZfdytP+wNkGvz1+V4W0c08PppcCTvVWgD0L0sGnO/bKB
GQcnHKQO5N0qM91zGOG6Uguvii7Oy4D6+mmIBivwHlIZw8fbbUjn6yEO6XUUJxjn
YyzqUfXrSfAbdgcYmite56AQ2zp2zx9eLzEIp03wS+eW42rmYlCJUE8ULtdLiBCo
yIlOIC0G+6UfZkK333PZLMqsGG4i5xaIz5BP0dUirg1VAOH3+St6S2siEV3G4Qzd
4Pd6LV/yKjvCBivqXqtflbh7wHIdNyVy8CO6qMaTx6RPJ+H6kxSkXCcrhz1uOFtG
3Wi2cCGY/N1GCZXscRgw8+zBfa1drAn/8zPP3pPHgkJ+JGe30uxO1koO1pGDRske
EaohLNbLyAdDV9dLqj90zx4BXBj6+oGLj9iYiRPGzqM922J/fDmRjC8a9eN5LqMm
fzVWt+um1/AS8Zw/aVBScBUdRgVvjYV7KsVJrlbUydXhw/5kKvN/L3yomNNHBEka
J9odP2lV/iIOpDyJqcRpwtMCeP0YHG85jR/qGBBL7o5ILyT/fENRnmjcRRnUStGk
kQcvMTwuVY5qMpY1qzqyHHEliDEfyF0F8hHwtY1tz5l7XHTCtdfx6avPVv/1zHxf
uczKU1rknkDkHoaymp5Y/mo1xyVpn78HrJrNyzI0AmWfF+8V+V2LPaSdOUlpFjC/
oCHMcS1QPLbW7uYru0k2WmPbEN78ymcfszY5t7ZJ3+3GG6uV7mxxAIFIskEac/3U
L/4OElZpMYqdvRV4qAOBqkWAgK/YSCJ0ihN3I2SCnip1z8PAQ16FplnSSQr2z+a4
JVrgGcTs14AMx4alP9XdEnehwQ13JpIF3CLQquSAuW01WJj+q84mPA2pL+jRzumf
CcDHo6/snWE+KsUU195uKEfoaq6u94Yci7jlZL4a5NawSlrXL3p2X1P4yHC1RvXE
zVj/mEo3X32I/nF2hHwBjQi528Lt6t1zuNG7mrI3/rjrcf2SX5sNfC49x0tqtji2
u8hz17mejpfPofO0p7cFLzJfY14POew5yljIDUk4plJmyZKRiD4BTkdY5GFTC5l8
FDEBLB2VaDkBnpAr/vL8lfVDGVvgFrm4S2wKChHBPR7Yv7+IBiIbi4eiGH+X+Rwc
pI/5ReIxd/ekl0zRzNXs1B0Sa7MqfkoTgetwco6kEhLYE+oAKTFjBtcI5dbBTI3e
0QAYpRUj9rboG8UPKSyUgbb74oR/akmV/xNiwE1WP3NECri6eX9XYEka3Yzd4+n/
ut9scyIQU4TwIQ9YJD+7zRTTa9YhL1WUFRhEZAYcmOniOFADBTJsz6XbJ7Oq+h6y
N8tGRqwRl4o18SNqZ2evtkwjDXPwmN3tlStDMftwUzqoVwk0g7ZRPzvqN4shxTeP
StK7srlA76Zxl/Ux7+C6kXzL8RQXjlUiBfaEj92b5Crcyn+/aa8WPgA5ORVT2rVo
4U3CrL1lCrGLn+QhPV9BVjWQTtlBYiRQAeugLAIENIq7TMaubhbswl3gNM+ybJUj
Kg4jBJmwT1KF4f2RLtfnD2Qz22/rLtkcOpg8ubGncyXcRtIxH0G0wW/2FalrhRkh
sgi5kKo8FQpj65DvQQ8SZUtS2iQR2ura12IxJQGAgKSYHbum4VqN9u/GukumdU51
H+xFDBzi47B1vaYMZ7AcSrYS/8jWvE6gm8eRBKjPLPw9Zpz1SUSyOTaklNqj8n2Y
Q4fBzt2mT2kRVQHuTCSgM1NgXVgQmsZhVdNHU7YiYJT06y9GKN6q5eTbj6fvVl57
vAeK0PhptuqTQn5EZ7+yekEayhgtbQDZB1Zxv0f52FFoKWk0Qe3O49Xe7jLPkrBO
qzmY4Py8BNSYUmgp/EFlwXTE5432VArY+SvcJmDT3gfQC3u3K5jD9vy6onuzuWDC
FNAZQLNPhWzECquuF3O8rXnZ1472txaVlq4DeDJ7yRAe84qtQr0UbnVD+qTzXTSa
UrbfT44gwzS4+pG0DYL6ll8rwbj5hDlaAcwNbLuc7X80Mdb5KZiWBj2C/QB79eGs
MaBFMmsy7t8jUp/K/w1vBZFzKg54QtU8jpF+JUEzFFCMNGgZ/y4mfWswJELXWFkC
tyP1nb6O2NT/aOWwh9tjed5LWlSUJ8ZYHwOyiati5wlrnX2U971bUw8Rz4DY+fGk
9MA6taZGuerCBzUXrZ3uRU/g2VUda7bkkVDtR7f9ur/TeAFgNphMc/Uenib1Edtz
I2CIpJwUm9Dg8wkbt9zv5IV0pO348X8xXFiOQvdRrJZgLUFXBQfRdPggKWbcsrt+
np81idSaAhd0rD+qQrVCoGY0jJe9Snp+ZEzvGn9o7qOdrzH0u0vQ+ByBDfWrqqQ4
dNs15XS6CMX7Hej6mYujF31rysbdL9hkR4StEcswQEQARamY5iOtBUMvhVd0j7U/
DEbkwNklbvBBgarjOwfJzyfMkkNDQBqaX4PZDvnluOznTq//YDZ4SOPFX8eaFhDC
v90JK3SDVNDE8uXKrm2EmZeVtFTYGWht2ttH532cyagsevboSaeZsH6VnkWjp2MN
GXNsrZqeIula3JMObTZsQyzjlkfOFAU8qEqPLxTfHpBgm4TovXnvOfYRhOKGWDSe
GCPWgvDs/mWxfMilPBGbyAMY/zzQ6qPjeEItTXkCJLg4Uk8fX3qKd3gUYg2uK7QP
p+1tWeYpk5oL5XyE3QlaJbNB5/wmS1ImgCJILvD5xYnAqYnKWsS4Cn+Kb7y9i3r1
0LXrhcavq3nV1s8wgs/DvkqnZVgJAjFtCR+Cj04lhcKfqdEpqmZy/7LupEoaGj9B
LUlNsFsvZBgRYl5Oek+Y5XUvyP0fUFvuqD8v1stf4drM8YMExKMHPYeDoGmNirYS
vsEALuusv7HOkK8oRGUqaI+l7hcmDVQGtLEcCLtALc2r/B/A2MJOJN8viCPzPJD/
mOrMBWOYAtE1zT6Pq2/GFicbIbh16lyWuD5ba+pdFLRuKMc4+UHMPbffO6VTPAG4
ETb4LocfeOXHQOvfCHHYi6jzFyx5AcF6xF+ZXa5+L/Z+x7f2eZv/PoSjnYRU16KO
e2fvBuUwSmzEU/lbpuacLxUFHigV9WyYJLFt6xPLkW80sukZBPvSjqS1aoUjRz7q
nEpccqvrJyAVDol1sGe/6zQbAMdzmsCrwDoS1LMuZ+XR3Z584PAurrCyD+1xAKfV
UAGON+MKzMpWfT77xKNWXrinvBnAS6kz+YItg9iG1V+RUnMgAztwEemvvPUCUH+C
SkkPB/hCYLp7fCaXcz1CT8+FvrkFq4jfKb3s+Gqg+PtUi2S/eS5R/YebdtKt2fbS
615gGvgcNNoQdCgWl6hcciMMeWkc+60luNAZKpahkqCwakykZHLoFPeaWTej+gvc
ohwu0HI2Qn06b2laBoXz+Kgpl3K4OcyjJLAM6Bj1WFjWxpGAiWUh3gPgnGgQYSRE
424b6K3i9zsKI0KGWEHQMWby92TG6cbHS2BO/POZjVG6vXJNrHDRXGIkcgTBqigG
pg5yeW9jH65ZWz0CkvTtKcy1qqOJJIOyLkFH3ttdqYPSHXl7nJ+1QX64b+hnYmIC
J588bmN4Da/TQAidstfum2SOcpInDeqso+nHh/ztXRVr4PRXOcJ0zl9Kz2/WBOB3
oFb6Ud4PF4SFHM37XxDc09yWz8Rsu9vizguDP4ZMAGSxUDqQgmZEyk8h1ZbHQNng
vKbxURjdjX+OUCHX2c+nUbDCCMIsIC9ay9vI2c+CdpF+TQssIdtEF9vPVHcCKxHH
P1wywlOd7erj2HxvcuG7o1yApPsnJiOtgj5Eal4lMQz7WXc+tldgXnq7+JuFmuaM
4XMmkNb2tHoqssBbTk/gD6H7ZSuqc+wRUy8qEXoECW8WPg5DvZrxgDM3NMQsrHMt
v8UVIKMH83TqyJUU3R158bbKQmuAqjuLWTXTcalK/ypgf8JlPGdyVaCES5AE6K3U
oPH9ScPZaeilkPuGm28fgQI6q7ILH1FmRt2V3ZBAYEIiQozxqIHajvXMkKD17762
WrIrGv0JU2DUSvbNaF1GwcCrkAKn5DCnkS08OMmkifild0p4O8QhAxjO6IutjMz8
+ruor2R10iarvWK7/1s57ykbCZexwYv1UkDiFezY5FWCCWh9oeCVJeQdFTQuvDXo
a8fvN3gcjnRqHlNDWLBWnHK/phyTnYo4dor/jvGaBdI96oDXqu4cUdlKoxCQT5ym
IjP6OS7efRIRoFqee/QUs8KuLG76D72NafHmm79IdxFiX9UFY/uWiyobl/DBoiFm
00SocpGq3bYvp2Lbqp3STGTLN8rUNDkAr0dlmWa+KlGlA+kYqbezzJ+MhHRnYG4z
weJSR1tXyPDD+03iIiDwOLukvCXx/twqhnJPTY8NrsFjo3UDWyLkfNNH09dp9s3E
txIDiMe+30YJmN1vmTTOHNPdmF4e2hOa/9D8kU64XnatAA88wN1X+xis2qvIxtiQ
uetbHa9/gXKK1m3BiVfjv9Ht106B+LJ+oL1hmeIDNFHk2DZplFHmA7MQvNcGoXwo
ia2F5QrfbdpuSjgJ5mpjVWbiwipqNYKSY71KhHsIsG/Bkc/QZ+mE58W1yligAI8V
YIgKb3F6R0APrKM4D2szFKQIwHPud9PB0lf04kxMy1HVn7+xty/K8SnoKvDWpe89
SelyI5hfIX8TaMqX4SAP/QAqw49j1XCAKVaW896+VADug0gbDWx138shRWOYjZu5
OScL7+IZTWlbfIsXfNnULndb9WCEV7OvGt2S5STxsF8Tlw8UyuTBEqknCzvQlA1Y
qi4k2Ll7AxSRb/exX4//e4wPdldSpqSjiuBNERV5tyEx5P8wq4uyWRa94AXRsGU+
t06fPBk/A4jH3m1316w6jkVoh++h9T9E8X9Dtx53RnN355F31emoVf2p2V+TSJy7
kfLPMx47pLOFJyFVMCHy/NTTQnxvgl9biBBMBriJVkKOG5ovUpVJaND+znPIgCCL
4HAS5nc78a75+BK8yxs5lLRZ6ZLKEnh/6vseLxZmVGH2QXKiaiuH2J6rcZtPqwhB
jonQ+vzN+UjOY/xFohmy3SK8CVb6+9dYJwiGEaXdNyIdHLBE2PJMZaMIpCyY3la8
ghVI+H+xLKMaS7TrB/bS+mFoAfzzzNdR0NQdM4XGqik0R95GuePW8xnh3xABB0Mm
oerbdsl4hTIXw0u6jykgRGp8O5pRLQTsq5KEvNIVKHryIoyqrF7Siziro4ss+8aF
J7lqokYka1X7yC1o9UgDRfVVpgsMi3c4d7yKKMTQqIW+XwrDNHZgZLzjN/38imNq
X+kdYDpuTTURumRiMvgsqx9u3D9K6GlGa/O0f6wegYzfBEQNUecKxzEwUq+3fKzC
KKVPVn2k2VRO7XeA8QM6+kIKNEi6e7FR806oIQVe+ly9iPOR2ob+emfHrObjjQGk
SCJ7XugU4jBa5wXG+3kqE7pkBhsyX0Xe9cj+RutaLy8DTE8KpHgPVNKkvsFITThF
PbDXbhmVw8eBaM3Vj30eMdG5hNiMlZRjKxHA91q9RXV1n4f/4T3VzEwX4dmgzqqd
weoWgdSY9IqeNl+mgViejd7rF5umav0wBONiWX+ZS0oU0saTmvCHan1owhGNcZf8
fR7uMgILKYmJWyJZa0GhyEXDwiOTiXTnqmXMbf7uSYnfUcnb2P3O6vMmMNgOm6yh
c4EHyh1WKoKVxlD0ymTc4iUUEtqC56agM4Km3cT498810vJQ49t4WnBoMhbYxCzT
k00DcY4YBLpXEbuRbuoZxHOyV+gUiRWZOV+ps8fGLQ8P8ev4ov388qhHTeHiZFrW
Mk5y7abCsxFBLMs1M83gPySeFbhwKBERUUuJcdb1jA1JpxiJszuEco3LTR0g7oV4
xFH71b9xJrDB2X/qSNuH3s9RPiN4pMpTrmjljMUXz5GyK/h7vdgkIP4N9BHj/QpI
KxzSwsmSLOQ1egDhZ2I+blf9DD8TeCSuKrQoPpRKmlLXRaSUkseEZuUcw7hH5fP8
F8OWCfpOwl5mRWcBWaSbV4W/gfRfPZuDfkYhy59I6FGPd5yi1fTvblmbw94CmnFS
IR/WbY3GsAtnX2YfMqdBq21wGUVlZMbGdcK6cbVR4s9CTMdQ6F78m1M2WPtQRUpt
S+Net8Dgz+N/fbjoPipeyH3YNwqQeCHl7q6LZM1VbwjfweksuCKHqYaY4bj+S5+x
FVl+xyDKvBfUg+nFDYDB1sLaoQek3YDwgAeTlLsNAhiqWqSTDiZULJH72owhZTin
IBEQZnYsDAxVZpMj2P+Vb13dI1A8HAWooxuzxT4B/dJLo8AvR0Ss6/ZsaFp4m/RU
T+ab3TldG4f1+FYlwyie3XXFCPS+bVyy9xE/2Ik+5UuqPgRHJq8bQOKuIHkqUB39
LK9IWTBXUONaQXn3eUjq0wxXyEJRxI3Mg8XvJBDb/v/uYho/Y7Sc4Zm+8ptgTRtC
7VkVBr1yk9EjCl1CDxHBS2XedpHsWPYcrDdMkBIhS7QIKFzdolaG86mpe+NcJx5s
4KTEfJUO2diVx6CkROH8WwxharHf3XlzXqL6XhlLdpMlnhlWb6eM0UTBLZOOpQxv
JVG+cxD8Inik0cCWxUGtDbI5WiHuNjxhgKF/zZGa01XCFXbinzpfwMB6AFzVhIco
SUUAS2jN+TwQsaaBaHLv8uqTZoougUenER6ghjRQKspODtzNaRXO6D2xtV9EYW23
CBAKdYSzAoQUMH/8Wbyt2ltQQyks1CP4MiMrA5iHerVoZmJzWNYEnDzQFhilnau5
c4suu2+lR+ez6k6rc89+9sycWBzEsVowDvx8rfkQm4YBM0v/I1XCE0CCHf4NXX7V
OhybpuNIVi7L2ABpRcNZtqYf0/g//o4B8yXkvQA6tLx47AcNbmUti6DKNv7K53Mt
RKKka2f72HdjDPXDx5worPuPqWHC1tikBPBr9Fj5ExCupXfff9WV6batNCUhUJUU
Acnw5euxjx0EKXiN5wp0rQvmYATV9pJz2NNZ8XwikZ76KYwFvJMN3Xlbwvf/chne
VY0MaiX1wl4tbC+2OZocfqukHbuLaYo4FGraUJTtD073KjrMryctvNdO+dAUKI9V
smi+HqtmfMaDKzzSznMUFHhfawrMMv1NibKFIc3cu20fk/gug8unIwEFONul6kka
9G6CuGXQa4blU6ybPW6yjCJSxAxxfMXDUSJ5lFFbqBDDXRbHXRUtA/eEd/AbdRvO
2daAM2MIDZHqEelYKzHNNjrF7NXzCgbqKlkGC+w2BR/gMrxBgJOddlsihLAcaRCY
FYrCiAza92uJJdrn4RA9Bm4ngwzUcjIr/7CaX2XmaqYUfj530OwJh3loOX+OrQns
Crp3qKISlmoYT6vfVIm6bvEV9Gsp05EMeZZGblWNlgKxT0y8hPRYcpxStTzXoHst
qecaABpdYS8RzoRhWPfkCaUEwe5AfMmjnHSm2vDsKXkN77jALqLpeA6Kelk5cwz6
Ffr6hxbMFIPRtfU3Y0xJzfAMWzDnNT4VtNDG5ymAYigIayx9uQHLRox6c35AjR2n
6Rsw/15C77l50GDTUHhkug3UbybdTUFKDA+Yd5tNKj+GiV2Ot57cpkFP1MaRVz6M
DJbm5Q83HWhV/jyQeOC/ImPQHn5wEAkS52wM3ODJOs3UnVgzJ+fdV6u30iqvyr3s
R3WogxPT0BeKrvVpNHLWNKuJuHyhwP5tIVvpZgPja43R7MgtNW8C6ATelMhOmBW6
XBnA9OT5wjFR5azQsYr76/tIcM+VtoSvvAE9Po8hy29uf0SafQTwGumVeGwsAB+k
hB6YGlwUWodgDDih2HD7vjTkflPe8ehjRkiINI2CydhmHDJFNVBDIkJsCwghIrIf
OD06yAU/IJ0COeI6md+ker6x7hBaTgUF28HKGb+GsyfRTsIBmI50yfSgXV8r4ZeQ
PrqCM0AhjKuR0XkvBbLRze2JNQSqGLZCqF2nDDkEBsSgx6IagIJTdmP6mMrXTT25
wNjr7uFdFfA+JUJYnRtBTIfTFMSDvN9bnbHACdb6pEKG54b5fNVBtAEjZi/QFSfu
ywuYk12FgeJbjVc2pAyedRopyHedVZVMrp+zXvD9A5LYept+GnwqqRCyBSxXnsFO
c+ldnwbo2aK5KTh2WeB5z4NOIgYl2ffdd9iigwDOvBVsAii+zZ+GNh4R7/5Wk9WT
oNb3CrbERiKk7EIj9OC3JpNZwGAdxYRL0Oda7Ds5q2Dx44vvziKFYZudml8VL21g
r2QyM16EWQlDNl1RAY16pJbPf/q3muqg6YeUbRMUSTPk6QuaanoALzEKTDIMk/wJ
VvfY181B1C6t58PdQjFjaW7qe9f+9T7JUJp0m8G2PoHZ2aPjbzjYCHlG04FNf2XU
+pJfZsF9KZaOuCODC0BsLG4KViM/VPuxTeEnWUHA7spbB3CwjFnyhroPRTXC/HUu
h8I3hPxkrVqA+Z6HjdhIdIirzvh4HwZfHiyPaiTjomcfsrerDmWyVRkNbXLfpkmU
s3tJAidpzxSGjI8tvytHZjuU7jQmLBs4/fGrjGH404xqQJAyJMrsiLidfXKHfPxC
up3SApDHAposId/nFlnmV9P9M7H9LfKndixyhZXb94Wnm27X1MtyCEZ/Piwa6b8O
34DBOTHYnjmOx9udEJ2vuMc3gdArNrBlLN97WdxoEJVtEGwRnLtmG6GuJ0Mr/kkf
B1UDnKGyaWZj/R002tj1hWOyMS63iE5mVqN6DWElFigy8ZwikDi1mcD4VrJt1hnd
P1KbIlKydfrEdgPetiCWHy3baiLIqzRgyAcy2EE9W7SlSrAVRmwwfAUPy7ZU3Q4L
1qJxa0QYba1RlB6q7jVXhkf11VNik0+Hpvce3i/CbobRzXVVWznEqJ6fXjImncI+
5DYgMM/3cBJClBnpW5GgUj9FLLgiurgFimgfjx3TCckSGx8wwgEK2cKB8yayFY7B
na+LZM8RMHoaDHqRIWIfDAgAyHNhQR6LG+EpNbsLQdyiiji/GVjMUe+B/s6EPQEZ
xkEJo7WPRXdaxhtAjZnawmI3nGzpPxBeYr2gYNH3d65th22fyG33zY9o+uyJlSk/
5T52kTPmq8P3cblMPLnMONb96XstU4p3T/yesCCl4z0m9hkmhVzk4+pVABW1R5SH
dlCY54vTJ3MT6nGX441UKgb5fbtAr9mJIDxAwTZQjohZU7sPhrevVALxntJeds9+
nTiaIymNEB1dHllBIeqcjL0QiN+mG4y4Y6RQZQGbGEP0H+1sTfbCYdUkVEbZE9cf
X5TbAgBxFT9dFQv090hsO05F4cAFfN9+WI9IwOaSodY3tPpYBB0FI+vzU8rP6qm7
2R/CD4XEv0CwG6Gbi0B2IfjS9wuOjyHMFRCYbykgIkXyeCtMhAYUv0skjyTrtu36
qpc9ICNeeyq4HqJGzKl2jPDl7rIOhks/b81C8S/j0JVT7TL+7Rdh4B2f+bLS30AP
rYFL5Iy2In6BE3ts6badz6B9OfSKlpbrRgLhCmJf2cIYguaoAQbCQXcCCIpCxzFg
miHE7nyIRsP7W5M5IDZORcIhicjDwiW4jmHrDyorEI2EiE///RTB3YMih75roV/c
Z8jTNA9ChcoIv58N0Lji01n6Bh/7ZJQGLlGmej5LVN2tV65EZZdPPng0Th9Nuqqk
an9tDZrYviheKVpcVUPbETXhaZjxoCFHdMPGoZaSF0ahVDK2KdbLfJAbafYynYU/
3XGvOgldd5H53zogz9JfpT1PMRSuRxE1RpfeLwaGsQpaWpBPvhtWrz07wzhl73R1
rfhelrznVJd+zDpDCaPpjbW/hRYDT/c7aHiocxUPwK0BKzGolivAAC4jiNaq9Xew
jG4hb0RIPQeNQSlPifI6wRmlrUZE2AGc1r6FXLsWldNyOlyRJLRTx7FhwpZz0kit
DM6olLIg5H55Yv1DoacppYYASt++l8fB53o9dJDuK7kMipTA0YjUDM1FjelySXeq
FPsGAE3Lf0RpfnlzDzh8dc5X7J1Y1VuW7ifA2S/jm2l7kMRKNFsxLT3cy8mzPl1Y
MW0IvWyUZB9riEJmL4vpxJA+Wx6iqbyZatgwMMwlscRVWU+clPXE3JN9VeUJt0ii
hXZ7OtHRTqANUK2kqHkY2S7fB3cGQYmFF/2swBhp1i4s+vhePJfYwuy7e/At8IaD
/R/yvD1+Dq4JSmsN6mq+1XMD/5ulEk2BmHtgKCZ98jKyBoDgx3NmIUiYrmYYwxqG
vq9Iy9HtWOQGzIcTGATH56nLySQAmJ0WtuTn/jBkEOhvhHxQTOy4BVSudmg4Z2kE
/3qAO9fkHBBLyDRZdGZNgORmD7KSMcpoPqqaejZAZPB0tmQ2oDfqfYUvwQDWorpn
Ur6AKb0pNcPPeRTXYhYn965QzU5QZlBjr3XyoZRlph4EBMVNF0RF6jiAHfeaOK8e
xPcQqHR7bdCmism9YVvalt9mPt/zpFQnZZe27ZtOOzE1QGLdWDoNUFKUauZn1wvX
LqEaZNmohz86p32hW/fpoGEoa+JlhWIQCRNlv8bSHoqJaf912+kfK7DnLt1ihAhN
kRMjw38hczOvugxPKZqdkXEAgm+0tDQ400toNGVVV/RyRJxV79trxYfk+Jj0meHr
lSP4DjFmWb+clHBOUA2UwG5l5z5iGbZGUODrfssf2ftFaDXsBX1JcC4UbBhNSzYC
cAKxeT3l+szR1kYeAE/78gqtgzhtLSp/vsnH4PnCZExcJwXWOH19KxbjwWJEygvQ
yDmzQbUy7I2r1hbuEKsCUsTkR+f5bZLDdqL5AyXuGi7nrJxnWiHFPgkdxYBouCqt
//BgAlwP3r0tUjT5LarN8WQASRWbQr0Eu+B0K9L2flmEXi0j6fDKaTOGKN2nQJZw
MQUuKbDOxN2jnFDQB5RkGkQspgdYsKUYgl2qIANvqsCXIfWW1cEXeZJv72OuKPOe
FldTmTcv7PjbQhDDGE3gqXuCRSQEN4KjWMG1mBVd4WOy4bpeb+LiQJcRPJUBE/fZ
vLHR5h0BTtFtVAMBuDm3y9NWJ02AEzaDct2na3JTH7hmkb2H3MDulKJYu06Of6Ky
StYJ3epVG/rgm2BM0b/SnuUJWzdRa5MPg2YyVo2u3tRFRd3MI2+lZwfZTMnro34R
sxbXOnL+MiXHSQRwOopfi2Swz2HnXA0352sblvVE9hBiwugY+kwheoXcIJUCrBlz
al4HA9dEcKaSP9hFWs2MnTUmaMc1+tIYjXDZHaYl9jFHFuCOBFNYPmnnh+AcwjVf
LXPI6Jl3IHBxD0yQfqWsEhBjNArpqkDqmqw/VSUyoqtSHgqudbTM811wVm3c+biQ
5LGajJHwAuaDgFdctetmzL44mhDWX/KO6YDAJY2hh8XLWl0rIVy15E05w/fBgVOo
yvjb2nuQA1d5CxcWzLEpUi0kgoD2Voq6qSl/BEkx0VcJLWbpUIF/oHJZpd5oCQcm
5GNhApyrY6H+KNfIMAr6pTIoQcVUFHndX5MqulhACkpjmu7x5U0Ra4pqZzDbUy5i
sKIzFwqr/G6X8LiVmY0nyavGvYVkC4mM9YEC7Te87JnzaX2OJj7sDUHdCUcQ2U+z
sx4m4OB0bVdCvZGUr8dlOkcsJPIGJBOR4Nt0XGapZ8JI6/ZqOlvXxUtBYFfB1Q53
r1YY0cgSr1x4F6F/QAjjMZhZDk99KdXIVOgBh04BRGJq5c1L5iyJYZysaXcTvIzH
0k63QN/6M6xM+6bhBMiPW7z9spzU2Q/KjkQ7M/pOayDsMcyDJa4B60ypWsEtzffb
Ddugj7VyxwNTE1ZRm7KxVUHUabSImo2Qlr0bfyO6vewJqTlzljQ9mkccKe6T1sYi
/B0fOu7K+dU9fKuU3vligkHpAHO1kqHZwu61e++Upy6WflOS8M/y5VpK0pLyk30a
1GDFBAimnnL+HStZLGDqNMGiyPflQR4FLe/O8wjm/g8WFAnqCKBknj+bozJ1fTr7
x5bVus4ZJGgM9qVrcJX1Uq2cSoJJ122ZplQsTAdHBogYx4n5CBQ5aUL4tFBffkxC
cA1NFYZhxwhrVp0oxoxPZYxsdPsVCxZy7fhW638oARHFo3bIG1pSynAXC3rBBwZ7
vSnZw3xPwtOya0xJVFE2j8ygbBhnphorTihLnK+VxawC5bmo86h90w3jqm7IS8An
7yFjo702VnZGpfdBXSy/4Nsy0cNo/o3/uiIfIEaiIV4M36uYhvOooP+kU/lCPt+U
SN1ke8brD9IHAmEPUjCY2bFldBZvrhr+9+yNTb8d6SdWJLC2ZWNFwJzRr7Z6SKr6
Ln9VQhB9MO4CMFW9hUim2eHhFgizcSYUB+MaqTHgdH8dVLLBQOpHaixDIZ8/XpQH
gbN47T1QPf08flAeTHK9eiISPi31pXsh+S9TYpiqcCUk4HBuVzpmA7OJC4Ru5lxR
IpYPHTnLfcr9Y1N4FovaYc8w9Usn8ICq2aB3o1XQkdKnnb+zp/bebCGR80iH7UXS
1otwFTqkcatKhd3igG7ooMOPAJB0FTcRpina7SaPNZtW8/aZPHhPJMne9TpqREzn
WAR2PRBzRJEg32w7MoyySMjluRSqu6YWiskphipILQrmgUVwRlYO8ZQRs1WRONEy
R3sVeiNBJGcQ1C4FfI72fWVm398xP0znv3Y6X9UKjrmWtaAE0gRKXGyfgfCiiy/1
Ja9ez0Kz9mXKoM0zqA8IiNo7nHPyF4vc56ZmJXGYoZz8sNLrLwG1fCnFSQkY6SAQ
Ixb+O9tjoDKFZ0/Lnb4UIUVnRWxs2QqIuoK72FAUO/bE3rizdPXfVg5NxyZJWAfj
SZOUPszI3Bc5y4tgfON0kJBuZlk6rD1UjNEYzDk/3ivdKsCyJY1lieSPsZv9ysXl
3TJ2r8QBEhUmH6L7WXQtQ2ZUB8/HI/BFSYAy9ka6nOWQ+ecceKD/TuWcDnXgD/O/
JwC2FZr/Q2+1XOim6SzGPlWPx0jDmkS9FXAj9QqdjL1tajtS3L1c9lHne1hnrhfn
j5wF7ascM4aldxTruh9oY0V2iW7O9vC9IuFOtWmCdxj3fkAO9hVP8Zgfeb6ZRV16
dzjf09/TsYXTEBuMBvoQc73P6VTtgHu0rcmOsqKMbQnHO8eGtyFk0arBsE32lwVp
Fe0acXI4o1LIqOqhS5YMv/hjN3KBJF0r9e8kuVFYXzk7esnGJIIFS0H3k7vQAss6
+XJ2HeY2VH2yO9o0jNJM1YyVFoBaMAJE6PTXTcw6FE0EDYmIZg8qBg8aQjkvuJvi
elNbFKQiT+dNhgI+XAUwXn/ELf+qcrTEbk6gn31b6kFaj40cldbXvbJTOmPMqHK9
+gT8h/QgpmuQCtqF7OYXU9XZgZIZXx9L7lQyVii5AixuxoyLa7xZ7fEo/zV4ohAq
YZ+H+Fdp9Pip1C4LOhnxKmnbuOnH8U8+Cm7D80Ody1QxslhrpmPtIMCdz5204sr7
HAeLQK/8R7daeEk456QpTQXyJkfX1llHaTAhG0+Bj0uwAq3699YOijgHmr8v2UxU
ypN5QUhq5sg/J2BQ9ku7EXDnE3M8KmvdD5D5jBU2cOjQEBEJVyN3FHzYzOJ1HFlD
3/BjSialbk6XD3Fc1g9oK7r2pBAZlUfTCdodXr4ZR8mrldRPvKB8XCbC/56/BDvF
Zt8J1Qgo+Ho40v48zYl1jvhctYgzzLyTtX+tGUqhbijYcUTz/gAJ9kjA5sDbPWl+
IAoxUzQN8peXlUdzoTVh+03mtDSzHaDbLlT9QlZnVrfTBnkNoxwuoFF5VXZhCPn0
olL4jV4O/GzhHCoxJKoCNTnehGiNfFTk8Mxg/+tGbo+YgjWFmtgDrByEss3feWut
gfy0h5tB8tkLblaGqYCkXdwkBz348lhSLnauU6bPm7aVsGI/Tv8VBtgS95ryJViZ
rWhu47TJ6z3vmKTeKTnQCh16e5CplI//FCLS0JzgTtlIljSKZVKCSZdZvgjiz9qy
KEUS1DwFDtmWZgxi2QKi+FC/lfCG5dcwKzZZt1LvEoYEOstMpR0g2QSUh/DS114n
i9sXzZIrHrqdmjbq6z8dNRJVhNt3hE3NAnDUfPYieSfhWgFHJELvJkaBvkbXbzLr
IFgJQ3CBVmBwm5q58+lonETIOPX75if6Nu7H87JL6sCFLFCM82l17RfXC9ddPSCG
WWH142vGWycBBzK6qYWDvbORcnpUliRH6cu+1Q1NJjn6FM4OTqRHgJHkIy4QKYRe
7GaJQEfyV4PY/3wI18Kh0v4MTuXo8D0Jihx608JA8wvPdC7olvszcJvPH2ELl5SC
ZpOkNNBLjAhLyGbGRM4FT5wQQZRGe3urO2I/Ek0f94JDrfc8n2g0RvRwaVuyF8s3
nb3zWm4U3EsLQBAvx8zgp9uMlsElfmY2LEqqBkjJy4qBCYTQd5B1LyWItNcctwhw
6ziB033OoV6VfF/mMTh3mz4l8eepSSbe2sg1vbNWfJFCC2ys0QEQMRp8+KWY+Wpj
j7ADRF1zXxN6L5R1vbfVwCR+t3T0z1Vbl8PvYox3m3au/sRL0shvB7eV3l4LSm3d
NTxVaVNxGW+h0XeKiMbIxsRm0E7hiz3DKCf8CtVdHxXQ4k1ppqX4wIpMtTNlr0q4
roy4VNZQTr9/bA5Imw6XwwXrNrur3jmCsiK84QmcfjD/dWzWNl/6Vx965aWzP4p9
tGQftZ/5cpYLMizjdZPDaRYN0penUWWAPSueoY4eCjFiMRfpUsx3r9pz24U4mV7c
AKxU9cbpCK3w3ewG+sMrzbJeSWVFLor7HBqS191uGYA95SX5DEzE1/3Ldf2en6zT
xvh/5SGjB8XcNuRDdU5Zvp840xWcJ0hxdz8VX36kMTdnMV1nzZeOxEPOK80w+HFG
M1YE0xfp+PkTeFj4yEDk0qh/9fRCpZc3Goclmh5p0O3mB2/q4fNCViOZeLX9SaGM
tH6BklpjtCrbY+zFCT8vrJ8USvRrqY4+h27To6whjmc8w55dcRd4XZzrtDwvlXik
sLHQVtsJ1DYQ8Sa7ar2WolJdWiKJDfHnUsj0mMlPuatm+n7Ulo7QBDljyn8sxzmG
PFGiLOh7tfEyR6G2Lu+8mYZLISKLOMyPmbKstCYEqL9XGDHBI0aSCY5yd6gkFD74
UHhgkFkPgXnuMrpnzn3L+Ez1Xpq+qMEBPrm6BfWIV8kovPdIcwzl2c53LMinjgoi
ow0/eSgUPHraEUcF+7sEa9V8uKBAV1QlnYTxlfrblyxnbbog1BUcGWbVip4ktRzs
KOB8XogBTXUPYhQ6kLo+HOJBsa2H/7Efe/nD0+SF/yohj0Kq16tcfS/HGUDpgoeL
TnPuVS4BvpHmezuWJ1he970iF8cojJKfThpZ4ZmcHeo1vVmb/znXUzyg+oz7hlg+
EPjCTNCK1nzf+JDxOmvtmEYx98h5E2JsAi+LPUiM5gFpzonEx/f/abCBvNJnzZDM
mERSVLSIA+zu+TpN7TPx0je9IdT0HuLsQnENTwB1MiZ2o4KRTczjLN2WEP9CoPQZ
LfuVsxfG32pYQNjHMvVi9v0zmR5Vqvhx2HewEOLevUn1XacrHSDSnqPLGfDx5OJ4
93lDJhqTxbQtHdIRw+IMGCt9dNqa0l/ylETbYA5b8w1ImQPO2L6UorbFTTpiTZjR
nfk4PwlmSfCoLqRP6B5od5IN8VOnDQACRoY6xSJj1tEGr4dxvq5xMP8Nim7DyANk
O+UQvmwUrQ6LBJ1nNNx/a6/EmL7pzvQ6VN7PWIkPtgJEohuKB6SBQ0DJAOiArdpL
W21lYPFwI/joDsx9uCwM2M8f6wlBafJXkUOGah5hsEzmo3SLtyhXchR4AE3QDpyo
L8QRduHb9KOiHNQZXGWQIa9dx1PH9VhOicVuyK//2rg8G5fcTT4+3cdFvcobweWD
DPPZ8q4Emg5uI2Qn1GSUJPIdKoZjKre1LyBkBQRJ28CQ7Rfev/x/5aF3yb1X/ORJ
lXq8tCVb+3dbklQA5OQrV520c/HRoILYnepA1Cw79Z74vJNJgpOlGHFrTlklkll1
K1Ft9c8kwvmubur3SVdK/kiZSODXPOCN9wS5hV6XIoV+0RmgARa1GP2kdGOUFuZu
ygY3w0x370m6KPKeFP3sbxnQxF5W7I6JEGuCeOu3/N24TkPD9yiDLtGNyHZDSfBG
g5nIkNhETTVqFzgNtyvHvLd3AbBkl4SgXJcUjNVdnDKbGB3QCwV9Q5x7cfXHZiYS
mQxEnO044/XKgM6rACB+2gsozY75cRYF+chNdUmGtcHd7n23KC55wn1mtJUpc3Dv
s+OOGWU7lNMRkCtjGlVtFltl9uWuMcdddgsZrFWu8SxhPMX2AIRAHOwUlsmwGSzV
15G954RTeWlFv8cQ6G5QkxosUTqSFELD2BB+cQkIObhyJ5O2Y3S6oQAPl3qfj1pI
nq3+uGcHcigHcK8/QtljfF4qlG0Qz2oDscqQZhQ5Pd9H9jg69wQxtDZgZbDa6Vxt
DNVYEf2S7PZ+rxBI38SALIEWUY8XDF/6ShG9biG34Iy2HH55RCDQvPz4gpA/TBxC
8bhOZBrHnJYz9C5ZfO3kKG5s93nxx83TCABUVeX5gbvZ482FeWDE1/hHieZI+Ft1
zO9RL+umlrnec5ohPslWFPM5AAqHbfXO68dn2qH3xYFeLbZNJdeXi8wqQFs37g6X
krDYX9KaDJAykB9pBrd6J7oyeQZkCVHi61nWIa6E5aGI4mTrAPHtcSS0Znc5yK7D
Ci2NlMg7RHE4Nv5a4NVIQG/dfD3l9bIa6Wz3vXZBs900Mjgf/WpKXEO5aZdvhJnf
OweXb8vGza4G4hEBmvjV8EU0OM0fsJheX4jSmVFVhYbvce9yG1ADoYJP1VFlRpNL
wwgUySWRAdbu+v2n/hdvITaXiar4EfPCxdjuS2mfPvVeWPpA6RDWreesDHLNe5NX
i0tbMRrWS+VdnWv/ke9LNWOMQMn7RuYWKkzh5ajHeJTWXX3xIoOKj4pfT1fhe+6i
lWXUXgMjaDO7ojEhJThKqRchqTqBCAEq4j1TwHRLYwxB+6+8nddZxzGD6nuEeXw+
z11Ks4fqvwg5w1q46Altek81NLciv0+cN52nekZpb/eyh74v95TdqgS4ZWi2vmwe
dKnqdrOr99JfZa1t/w4Mp4wUstSCLOLyB/HONZGyBUfvn9ITM7KmZ6KoAQ2nWuZf
yO9ER2HgIBmYax2aTZl2b/qwhgzqY71DcsyONxUCPIoSyBh997KY5rjNdU/vHWbd
vHtuHx7exd+iOPjaozjq+71D+Mk+1jjJfzph2K8bdqoWdPEQst3sgExfFtOzKNmk
eOvCuaGwYVgRcUz451y5eXHisYqnBPq69dLTwLhWW3oNebuDuQbWoCEcTakYgD/F
/Un4iIJj0PaSmeFSuQPTVaZ8U+LZivRzuQVYoW4dXtc8YERdORWdalUpcZBrNyBb
jWnCyEAsk5pI3ayU5/ld+qklJz3srrvUBAk59dkAEPBtawhPncT0gOsVuub/tIAy
4ceWYFf3a4qRrmYHKeBcMU8cIde4scQylQM51h/xHbNX/AEjfP23zgTtDvwAi8rB
GpPJyzrdY2mxE1ZqgQgJMsDeQYmW4/ziaLZqZsWY6gEYxzbp68r5d22CVfIIj0bs
u0Fzom7uENolwijFKU7lhX3P4aAiZxai8d+twGM+iNzLC+G3NNA4S7eyv4Bwugom
LI1KxtQmPpTYLByF0IOpRIRiVD0cEpwBT+cRQuc50S60HhZ3MHGLHy7uKW2+h5BS
vFhas6jQM12/7ne5gUUczrRJ4ohEUSBZK9smcpdmbYh2uVYzEJ3RY6miQb0NfNcV
RrSbNKr1IBCzZjUcc+yMJQdmoK4TXGqdgVYn7USpkgfTB/bScU/JlhlvLtu9NCI9
DxlRb8f+W1VrzTqGVqV+70fQaasWc2GM7nVXr2a3A4eQRA2czrHj3p36wJONiTYq
abuq0EdSowr7b84hnJh4Z8ljaVEz3ZYTxlQ3JMu0k7hxg+GyjClQnz+NTRgAa4Yw
IuMese557qTl3Olu4T3J5p3gxvKfFT8K80g7jQJr482hAxBPo7TPpFWlfAWNDBEx
pi7Rl9gZ3CfI+P3MrKL/4Fv0ObMWZ739CUVlG1krEDr8UmX3heSPtFLcz6FgmPpG
UXdEcXj9SXJw+HMBafHbJEmiS20HPG2KJa7F04NgxzuLSFfi05LCBJfb8C8KqF/6
FCkavDEQeQUFy6/vVUVy1t3exZyiS1BzrUSalo6JcVIQfPAPojKHQARcdEiTlZtA
09eIu2lFh9L5WUPQl3nOy4cS8e+drHxjSSyvkeyfM7QId9utxHRwwR7ikCYg3/cL
1W8MZ6zyQSgySGT6LWg0qfCcEoHz8IPJzDUncBnqkCCAsi5OYRbbyztJwYbVwDV2
ozXmckPop2K9Mds18JmTGOZ96ldvSnhC4nu/08z+pqHivVPr4liVJMF7VLedfhgc
OEGhEmZ7ZqOcpK9925y8YyoLmL3wEvvZlU28MNw5SnKGaVC9RJ4HpTmEJMS4yZ2F
gbkZhkVocu1XafpweACiicv7pHSShGGzbKXejDRCmdgXGJUgDU709U4OzdjKUVq0
jXyJZvFr3BVCuuwFgzP5pxH+Po/chIN/rEgfb6gkTuSsfZD7rwmrJjeCfm0Ud6bg
1dq+Zz/TRNZCjzGX+dfRR8Sd+7u2yjxQ3HwuaQZlm+vGFhZjPVf8UuAcC4i7f5FC
jPp9qYJx/P0/R5OsK4LJw1DzM7XP6FWLgmNrR5U23JVUYIj7n3xFOcw58ZIN4uOf
0VojKD2Xu+B6w8ctkKpudXEHYijbq/sKPZBRcDIo+qGJ7IU6XSD4xhYh/mQq8dT+
qEXj89iaIUOJMPjpku9nqKSedyVXwDB14tqihzPoqV0BIDH0LS3bpHRA/h37Qcac
jUUiqU0OY5qQkNDPAQC4nLtXVkou+woFKAerupBYbIEPFOZCA+hWzRUd4WLVfsto
gmPgpCJ0zLGzFkBbotnzLrl+bcDWQoqYwYHiVyMv89aKdzcKlUulwfA1zKB70Qpu
Z1sjgwHMzhyM0mVzeKt3u59E0WkAw+kH6tBZWNYpHMO92UTNBdu34CXYpcnLmLBU
LcZgXIH1t3d+dQ0azn+uPKH+gkMgrHngCsOh/rFknejOUqVDuXhDxsjVHEX5/is1
UkDAqE6wsGvv52fE7LaFzkt0g94dxzxHtAG6l3iNCGrJHvwAwsssXNiUScjZAffs
9wM7uQDA0KtQ4449FBZ5ldcFII6d+9GZDbI7qVJpM8INUvNZzzvidfnQfQfzh2gK
mVoatIGPbS577/+fi6isxqekJc3hdiv7mQl/3/UY5Y0uEFdNaQyP01I93toMjz0v
ez/892+fnhnimGx03kNF81i1UtK3XEOs5FJke19JlM42MdexKbse8Pg2wBC1Edj9
/0QPhYGrQ/1PopXPJGKKWdl6DYcczezhtVLPdkl3kcB0YgCwqGsP0LPDO8JgKtO6
bLfaipor5yu3B5gskYtkuNofBcFltulRix2tLzb4rSn61ytIYN9mnBLLeG/GELug
Z7rBaI2m9C2BToGx5CJDRVqV0kp2nFVGMJLrhvAVr98LBfZdRUs/71FvWsiEBMh2
i6aw9dRgY+AeUE9kU1l72BLJmORON16dz5lDsQDg9AcO5joXmCxEvIO7V/6pyDCR
JbEtUgJk2OGntlozvQ/fRQXWeK3E+Jp34vUvgC6DgzpYtkB2SiX1n/zuiEQKP64a
TAF0cWt58cSpSY+T+vMu3JzosMfcTs9Qi4WTbNsYggw693tUQFvNqRdyyXsJmpTy
imi5xLpkTTLUoWZ4aSlMtJrHaoeutOMU9v7DexE7lHQ/JmHyRQtLcbDj+J92f/On
j+NhFCLicL8OLnBfvtnecpmmxGYVXVNjwYffnRQkCP5mt6qlmTkf5FM2vHvg4HO2
cEqBfBulggFYZaO79wQ0bQtzq9+uU5cD/mx6r3aaKbeb/JvC0V0IIT4+4Vcderhg
zlW+VlRVJXaMVUTDZj/KCOBCQ6CVWJniOIdljfmreCsoTHcjB5LRHz7hQiVTFqxT
/oyxoC9AVOXCRKIZpP5LyaybFdhQpkN1nqfNR+JNkVZQpTCst/xbl2R1uRCNbC1l
xyZPm0pxyF+2bMauYYTvxi+rBDXvsBvE5AGbNeEmNSrs0WByIoKT2MThcdFmq1oL
EneLS++lztc9kii/9Al512rNAenpwxM8GTssUkFyltEEXR3I1iTWru8AOKIj4iaT
xQGcgBQpS3sImzjMzlQ5WW4A/FoZZ9IjRkya5w7wOcdhJYqT7TyyNk20M/sihex9
Ks62owqyKCnd0C52xcn4AUqMeWOEqL64gyPKvRiD1evvyBjCB45upKQ3pWIWkjRU
Mt/sWO1NUKnG62TIdeXsodRgWsqCl0not8qv3KNjgMxQISNRZ4WQN+bq7VEcXM5p
+ct8mKdaIywVHM8GRgEqn24k5pCrVHryJj9sIGADEZDG7QLI8dj0xb9jBJi6soix
epgp1Cw81af4fPccSOHIfOaSfGexf+mz7m3fqQnoAUFhDrfN7Z2LKI4BaPVfTtLy
RSCHDrWtItXGrg0QlSngMdu0L3MJ9LhAYfvnC8scZ82fbXhEELI6sZArAwWnUNV1
XDypr8ywEtYvmqTpm02zCsxNU8IkK0O4+Fm/x7TjHxk0iXyP45GzPuRr6mfrPaYp
pSQNV/G3lBG+HmyLaMGqO3V4ug7FK7OU/H/vMwywBvU/udzbOhzSQdW4DFMyUOpz
ILKTXVpy41mYsQBCWU/gXzk1K9ovSuGBRnkQ1yOTAnsm2k6HJVfWT8Lceq3adeAW
IIjqtjBslWJaXHuZV7MLK4/5jQTdduX004EW1Uk10RmDAEfAWw0Soa9L/z9JpsVs
xB3Y7pukEBJX9O+CWXU/cdutQjhbCC1ICmXyOUD9oJRhKSWCS3Fdh6Xu7oxJw5Xf
VImgDWR7ie52DCZ0R2Yjo8wcTsqpgIAdtk+DodbD52lr4QZCppG+xqv5UbTu7udY
wl+CTh9JLXv+3wLURnaM/iC0CwNUrvnqpdPInE2RSiJvwX3OeAyk9tCJ86mwofRY
fBkt/VL/an8LV4JOm0UT7BzzG1M4qg1jWpLqsvXcYQX8DvS0ONz2OW8Yny/W9PI+
yOD35D42dd2EMxCf2aOW6PKMVTnu2ao7NEg/XZr4gkOmPe96ISxzCBrkWnMo6kHn
/7cmapzwuEsudtGIw5d5e4aW4dVgaf19xoqMPs8Gsm4I9Oie874NTE5kFuz7ZDCO
C5ZziTkUFLX3t1qykOEHiLSNakT+ukBIiTbTn7rZZgSyDDNJSXokMOcggSsC9WiU
vMqEtZU3yaYDVheyG64xsr7MihmzlOn/+qfyYuVJy5UNmrL9sFI5tNb80/AAtX7M
0CLNvrcQqcVpPJnvNoAB22ylS58Ij7o/6MpjjLHAb4QmrHNxlMkR5OUIjljp2DFO
A+XIj4twG+gRoqfP8qv51Og7yUU4pS4EtswkR1i9JcmXAJNJtaw890fRQc9WJUI5
yZ1X5/W/kMfQFJRZ9BZstjfvFfdcKgJSjqPmW9QxXVH7/NsH201OkZurOuEMKXub
5WWg1F+x+CDBOZG6X0A/B/UmucnMbOCpKTY9RcXf/2RKY+RUpPswxz+Fc7ziPihP
KSHQKVwmnl8KLn6qsdgcos1bjNorKV1/syknzIKEO0hpvfClSZDZ/PaFYEDcWsRB
/yThfSUoB2bVTZocXXo09l5TwnK5il18EzLhqwqXW9Ziu6aYWN7kSmoRaCNllX8L
yR3S8rAq59tC4IZzZVN9Mu4M3uRQDGOskHNmMMxasHedcv6pledcsMV0Je1FrsHF
w6x8pw6YDYXGixUE+/GNAVAeUsWnFS5nTtvvnSpLNjqXcYVV+SasUU8vnmZDHFPW
H01ikRtlJA+tJIdpTpbQygitA+2fkUFBX/Tj8KhFHKSvCs01RWqOC0Rdi6bdP736
nb66pGktrt+XjBSYSItdTNz+eeqI9ikG8f3xYwDy6ccPk1l5nDjJNKnBmu6KzOVk
wjV30aLlnApr+7f804VC1Hay+j+OTc0t6Jlh+q2bumZWMQSvRDiSoMSjAkkq6DsA
SAyVWoc39jM1XoBTL+z6Vv3JLa1LSfEc8RgKZT1oUZAG2GESo+1G/JaBv0dmkuR/
ujr5ddpnw1k9caEk23jM1+mgXk5br5l3G7cU1n+2f/9PH8SpeCsxhe/PFi8/dY1i
V67YxdCMduxrIahfzn66kPfYuUlR9M38XucnBTbxQm413Nga45y+iC16pgrOujAW
ASqVkKLX+36RveW9tsTMWZzheqQNwUZCPgNCAT6Z3KdUtvpJMTwztvveFFroBDfs
UPNL5PsbYfSa0qFjIIEz5sqEs8YAxPc0D1wBg+IAv8UeBoGkvwrAmQz1a/HprEsE
f4rVaEjq8T6hDKe9TJe0cmvQBV+M94y6pEebdnA1uCABoaZjRUUKdotnqqRj3jQ9
50oi5DuUM6f+3I4ZObhIUAZJkinIjyU7/2AqtMzN1QbY/SDWaFrnvkLLHJ6Yw7bZ
4Pu66aZU4P3zoZh/ve6Bkr7Up/3F9B9gNGRPdMVZ7VAR+PZ3u0vRZFEcLBu+zmmN
bx6MXT8NMvtKp4709wS+nuqTqBDdBNL2r2n8SjPHtkx9wD6aGY410NFH/XZdHUmC
MGdCMdUxQgbBQu+2HYrU4rVkCqi7AP16dEPBwATO+XruVhGlQW6gqAsnfJ4SSTj0
Extnf0DpDO4TFoiDnbQ6yHF2Wu/B/93vOB7Gj8EGTn2wPTDfqSFbsW/0Vz2bPMru
QBdGk8y7E03pfmNRfPpBIGQAfFj7zPPy+Y04+IrjKKDeuY30/NEZDLqEwKOLShzM
o1NG0VwzMsqHUijqCnjH10YsEFrP8ydVXbbiYDoNXAMGGgyLgMxm9glVnoQuhOqc
XlHnLEfv6nb2+GQlmvggj8YiL+G97bJ8m8P9SWsJp9mqoDbzUJCubFU+GL+w+i2E
UM2zHD4YoAtTA5ow0NpIxBOk8olK0t00LS+3SPYjh4vu9u1kmpyEQK0QLidrGEFZ
Z6PlcavbFGMB4znej/nMJl4KmXYoCjqIj9D30hNJrlIKw8Uu4OPej3sYJfDObUQm
buthY0zakslnuyQJozfaBYROwVh8DghtHYIynG/+aNCon6Rq6O+9uOIo0+t/XIaP
R1JszYsSoOlAjiCGISPOi2CvPghKbGM3wNE0NRGuRTquEwkWSultEMoNCTBqI4IW
F6CXtIon6T+kKb8Xh3BczTYRil8uYoVIvYvX2C4XxYcqxKFKGaKjKubEUbJ7iuBX
s+FOn75ibvqlEU/IsjxcJrO5Rbc6P1LoEDdRbKgPwqT4cu2xssDLdC33u2o1QtqY
vq5y16gyLjMP0Zon6RkFg4xHUPqUD0D1iDBb5SCWUBdnuN3rvs21pobe8IXC/H5i
niDclzuJL5J41Ny1jJ2th8FraTIwaORh67DGD0/vz7WWP1cuHG8RVCyiHC4Z9nNp
UrDWDK08kgyUI0Q4iRG+unRCne+/omYWK+qd5ScT5+/o+vLJ5UN/lpM6i5vGbNrg
U27r3t3sycSkdBSgqYNWYKsKRNLsf8+WHIwyNNbN08D+TVjcKlgE3x+DVrNYGmvM
YFMbiF8tvDOdl73cefB9oBdBgt9IAJ9NPgaLG/XWABpL9R/7KYc/YRH6it+C+Xha
A9Cxg+0YjSqBkmrs0zFZpMY+0JjonhOlLM8xwA9Yy7R2e8jH95goNUgpbNcOZTy1
d7ogvTMYyLTYeJZnspP6TJIdqi37aX/INKhEpd/BEwHY3/MiQkye0Sy/IbNdGPSI
8tBCb5shakQJTo+IGvPQycQQyK5JOdX8SvTX/CdGHC8n0R3ZMD2m+hPPVyY0Kh+V
hki2+12fmFaFK1Y6UNTWwSFI7STyOuZlDw26arD5siqqXnQ3AbDXZz2ZbKNpeI0/
KwH3yowzVFlgAWGeL5zke59Wkx9OQicRn0SfJYI2a1DBOtgQtt0au1akzDcih/S1
k9PKH6pFGQwCNm4Mrjli/mbfHBx+kW8nIiSfO30fG5+d9yGIS7eXhb/hU3nf6rix
6XncTRofbToRmpVDezd0PyrqOEXez5D8CZiItwdXpiVO18L6Oe886nIIBIbeSFrO
ZdH9BJHiWDskfBTFqu2ZZW46L6nZMOnF5BPxEo6v3ntRsuomF4K7JpK18XNnA/B5
ztRr5lX8UfF2zoMvOCNGDSiP61lgV2GObOMOEO2IQM7N0HP+fOriHTXZQLUEUFtJ
aw2+B+RYPlkZKDFkD+qKHWrKkuTOmrcEFtO2Tg4piDhzMSr4DJ5/ymhBumWHCuvx
Wdslc+55WAc8ofgXOp6KbBmUJNNzSN1YdhsGX997GZiPdFtUFpay2cqUXmV7YeMX
2/xmdFsfW8tOOX4EgixDIdiuiZyQPkANKOOUWEpqF1Bv7dM22uKV2VK7WSm3Rti5
4kE7FEcCVajQhFFcgQOQa2Pq2kf3ZZ9SSuVajQ9HgE/LVOd2InRRSRm1OkN6D3Oo
WzWNBotCew0mKG/67MlYeapzpRQQ7hvVLLKXLDP04H5NXQeQ8J8cPwSgRn18gE/b
k9ZPu2P9KQgp9KMQvnHIY8QgQibPvUUBdiCAYAZFEhK1dV8hb1YZuF2divCEPMm1
waAMMhRMt4AoVjd4TVgrdT3Ka/S/RG+zkngez7HJkn74V/gF70zwJ44FY0xFIRMp
89/NPy8PjXRzMLtxVJIneTkDgoKkGmoQH7PvB+uD6XmNjP1b3GdD6QyRsLZFVubq
wG6C+drmTB7K3wmwY0xStzKlNilffRtAtaLs+dVB893LrI5E6GLM/Ij40JlObrys
wNUn34EgmTEJmT77LfspAgpC1m+mL40sKRIs30AwqLcqkPVnvVzyR3h6/HdJyPcc
tx8YYtjSDebd2dapBtqD8hrFhtxDo6BYHuYdYojwryoVe6G+b4A3+3Ei8fISDvbD
4a7RmzmLWteshG1lWQ7CH/aIOylRgKGTEzZKot+JkSzSTGPlG1JcoYETurDSFP3F
nd6sFEsdGh91or4wo4uSwXcSFXkn8BKKHnxaO7Vz7es+iJgmNJgp5/kkCtEx3NDr
/t+K0B2AUE3lNhkES2SOGmtj4hiHrw2pHFoaM5UaeVTkCkt37TBH7sWImhW8EVi6
WU/njazwqIaCt6Spc6r39bwx+JrnNwm2h1chIBW8VF2qdL5H2ElpcVXDsDyeDW7q
nwfSmvu9xlJ573fi0U/mdCTZQejZFwP9GMwQbTJSGCA+VZBhZQUkBYzGz+VUD3R9
T4pyAtJk+aTaZyDH/w9vAgeuZxptONlpA0QP7llxyNOsqUxYHBSfGSL0da4dW0pr
x9A1dnrnTruwhmKIWzW5APWUINOlvwPYScpSuuXXrPKRQm11J1JE77slYmAK2JQM
QDK/7XLGv439iFjOvGqeqDcMUwHHq95558BFjeXSFufZApuvNUuTuCHOuFjlfyt8
VM0hQk6mxy8NIJrRn0GROqPrpr5Y+3vFSfcI45hlBo8FF2K1hk/ShsUa2qwJ1cOY
zwgIstgnp4t2pm4bsenOS48uKxjFRrYCGF2YZywLRUMOWiIqAcwrXRS+wNa1x1D2
OqMrFsX8RhJp52lPVODEjvHgqt97ydtVJxvwj5ExOvbqMpL5ej0I8VtYSmsISd3k
FHMfo1p2TB2tLMndCo9D0IOvJS9zYi4wZrOQPlflBAJ69H8f5C5xHkQj17YyivD/
a6ok1Y7ARV+Y3p20p9BEE2c8TfB8L6irt+vsoXPxxD23GWQpOMbKE9EOJTtjf5+S
GdjEnqb3DhCoPVagmMH2GFb5wDJhFy6GSg1PRJW/exbK6fzFrLCpmgy5BjNvjs/+
nDKluWq1zOR3B094+k9SFR7AwMrU1HaNeFkF5xjKsUP3/JDwPwfvH2MJURkeCOew
a3of5Io9MkqC3NBWYcYqfYY/F1iXzbt+LWlv/bBCaD/AMHm2giYuV+NNsfRL6rRk
J9Xxlp9NbEGV7aojXj7qiJF/hSP4lxwkRDoctuGn3TnRGeB/MqEo8tdO3po77WI0
7lHmvLYxj1dI/ofqbz4R2ARZ4+BfVJ92Sr/FhI3HNQfWCDWECo111ksUWUQ7ynl1
2pb6chAamtAizzuRG3yzCCje0zAAOeH5qofifoyiVxHLnJ7ImGmVRmw73/aQaRTf
HQ/ntEOM9Z35Qc7YP1Fs5p+oDHPbJ5OVbj5hltTWgBFG1V3ayy/093r0ki+qGZSW
GROqxAh2MB1jsAoqJZOIbs4Th+ISn8jxIy02EqBDB2AGlBInORbvaWLTPfAWgkv3
aYN3kukXKPzoS9toSBUvUVcAf7PV9XhzzGdL5dLSoxL0D4hF4yHIRbS1pZxhWWjx
84RUhCXwqiYm2rO+BGiuEJhgmOxtGJvqJ23bTi/WNqZ+7Q2PRacRy5WuY8uV9TIO
FKF/ToyAQEdrtlim0rRTIYLbGAgexvlebyoh++suXYT1y7/YrnyGRykx09zOeO0f
oEtZXgnA/4YS2fRuI0NAKzF8BonrdqJL3v/C9dAtq+MlmWiAesJ0OwHfJ/bljmnh
T2X7imcwQIQYdCSN8uIm7OkdDZIE3oiad5ot31yd6DuLTFdtJGnfaNtMkx0muuvr
GbUw37nYVx+Vc5Xb0LUzPw1lxI0mM8ShcrKIUIq6jb7qL50zC4+LAMgxsgX1l8g2
4L/dv+jdJWg3mzIeEEg7v1sB8bcXwcPX7x/E43amWAYoO8qRdjqDxLsZlq8uP5hm
/ILdJ8V0zzhfk/OsQrOeM0l9ydzLSVsJeRAFZAjorazQ884CvpgwCQIy2ElcaPv5
N1FgpNr7L9FyJaJu2di84LPfRYFjgp72ghKKmp+RQO/WQVHHQRwmwgdijT1DDzfp
SbI0bZx2lr3zGYA9jipKYLpeNxr2xhXMvvK7jQ0KK/Ltu7k2A37BUMoOBWxqWocN
pPHESXY9cu7jkglyN4iMZhZy/ZdonSgmwGWvl+7/4q5psZ3JN6MDSzdLU9lReXSY
7oRliydervzpgqk3WKuCCTr9zopeXlDs5N5o0+AFAwxmm1U/NeDT0IWBK1YvDxzh
DQLw8NmlYHpc8FrphtfH39enJTNPi7V+7E3/kQl93U/aDvMbKOIkmWK4nomTs9My
gy1i/YFvPqRW6va8BK3JaVkl0iZA6+kg1q9yqcRoh5DzC4+HnyFy1Ybd0FruEssD
CY5VwUsAly8AoRtYR9nLUMxfKvmGQRkXbuQiYWuaN1gap1t6hwQSgEUVQnNXK8hL
DjQQEpvrzsSuSl6eqa0yplGU4RNA8F+pgEPFTsrL9nYolwbqRO9DGpDjaC/4dY9L
AEXiO4xXrXERhMem04QOWuXCd/2svtl/w71fqUvn21bmlzUs7UAqFt+gzdVrmjTW
X5wuEw3+QwL8dlCfkRo4YEl6lHJgiema9otxF4ls+7Zx179gpgv8WMG5v+9tNNN/
BuGJAEQ9FIdJyqjE+xARX+rqOEvmqeqz166vVM+lHE+EdUhYdMSfYAEJBdi1mK4G
DvxOO7ZMXdfX/78FxB2bqRYqEnY1MSpgRQQyot1gn+kHpGifN1hsc5V3wRHeqEua
VEMLEscaOPjBRieZFEGDJp++6wee3e12mVbLhFWBfQhpbReJu2oVfhL5iaDyjihW
JLr2Ij577jvKh1GZrzs19202QmbG5hmwf5ETzpk125mTt9DX1lQ0q9c9D0SUEVrj
cdQWK55UIYfzeJe9KV46l1toio+5EnvUc95OIIvbTr0guwUP3iZ49gLmtYVsX5pw
YSDjwIGasA7UxSubhSTj11L215VCXEg31TWGLC/skBXy8Jm/KrG3eP6TilntSK7z
N7Nf8ChGieTHMcUwqzyLKvm4Ck4ygK5mPk8+L6GKo/QdA1MKjWq55XWG9baFoBI3
JHTYXJIeh0rLsoErp0mgCkpodYLpYlKTZ1H+2Mq4gO901E8iFqo1SWtnSupXZ8d0
AvjryBGSBCGcEXf30Bp0NHJEt069h2ySXlX6wouw7owNetoGNjbmwpoD2JaeFia/
uCv2VQfjav9Gi9BlbmtMJbvlOPbFJMr7MOYh9cJu0xgA087B/HMQo9k8+6EGhk2o
y89gd+wKNdaifCOaK/uiHFPRrPovfpyC70gPtWdwL5d4BDly0pbLm4LPsi6tuV9p
NRPrdpAjrHHso6ceF9RY2S1zDy2h78ZJ+yPrzU/rUlePe93Tp40qC+s3keeeBX7J
addKkbapt1Nyg4NBF+t3DHhE7SPIS+KIfvIgaDITaZ8QxEdyUH4orCnUiHRPw0q6
T9MS3X+W5XWjYB3It4CaViLwbUBJBwm2JKhofpNpCs9ph9AjoYFYJmU5uoJfVed2
dfcBmgF0N9EZukB+LJweMGXS8pJhyFuriBZczdLoJkKoDkhUxEur72K/Oe7y3DkR
Vxqknwab/aTusxr49C7pkI0Usana/vORbo23Kmsa4HnDmXoABbutFh+B5yHsktEe
NZzXtLp+COs+poNckm0AOaSpP7EHZgLPxibBMyvJtFIfeMEd36pf/HYQO06lA4x2
rGJot0kbw+jALQE1Q1OIFXdR/4Z/rKYD0CInjIYOwhqzGCW0FHqeof7gVjfJuGh1
aLK2Yd+oNJ4Zp1jAZNNREGy4s61vLvaQopmr+DMkoQnuCcV+AgN3i7XYri0PNVlY
pmnFL+nwEPpmAQ/ss5dW2/W4sbhFYtvSyYCMKdteoOZZqnINf4wDbEyYMoZt+JyT
JFaX0vPxdw20f31Dj6Gxxgyvp2Z/8iqsRx52OTlJEXdnikmLVN6AItvpT9IgpaRC
0vlG40jMfWD6jda6rQ8X0946lWy/099q21zsVihbYhmToit+ZPEwK5X+5JxZeEyd
PkP3YWmlLIGgTtqigAWrmA1W2IHx8FeLTSwKomqAB0zj1759ZKKHvOHUx9XP0LmL
46Reuu4tFRfvEwxzmhFvyn50OiDlXPqoE4ejmyOPQuofltTwKSfWYF5kCDj7CYWu
98ie8BTPEJWleQOuPlfoGE4/gCMVggvhL0zyYbLzFFIX2+xfNhYiHezFHGdvNT7Y
Eel/PxDOBNAZxziJ9uj859IlXrT4wLEhC994H6K6skOCGOa1C+XcEyX4+8o+6nly
ygQuo/DoyyRaked6QewNcq1ZZV+99JpUsvQXDYsMoxe5ezJwxWOiF5Cwaw5rhVPl
3289MMe2bzS5Ce8te9IuzapsWHEFNVILUxbkM2NACyYRy3D08i4aT/+NlsmQzjTq
lvGvf4+u/NDYoyWMSjEWcUrVL1nVtWlBQtoY9ehdb6QsNzetg1gsp6myWZ3MIOKx
6IzcOdxvHD0ZlUwfZv3VVFQLONvVkNrRwrcFvTCirrFpvoFNkB6WX4gDZa0xBKja
lZ/wbJnYqDt0bZzzGPyqeFi1dB1CMxyV37+mkW47FNfgz1h3sehZXO1RAYaeMDoR
d3S8QIhcYu8QTqEzljjN4CTbFRpdz6OjEdFTOWUHg7j9CHH+uoVYZwbjBhwtJaCv
mEBZtXovsM53lGBDJLwh16pHBw7vivyfEUXF9r8RaRn4C0nVtKFNp3KXIPfmBNfW
L0yO7ZVm6CW7AvgZeQYjAxgdOlH+EtidM1oeOCJK2fPQMASLKuod3RG5jNN9Ax97
vxxI/d2IuyJclDntR7/cJzdIAh4UUzqmoDEnOdf+h+QSi5yeFp2HviWiU+M7PKJ/
pycBI/YhO8Q1JlZT9N58QDfMkNfNXqXfIESGW9WtpRR2yuxNbtP9BRnPKnjZ/7fW
vF9hYNIPuz48eJkhK3Xcir3I+zMuOeRNRHC2gkNtt/N3fkPcpSE5W+ea55FhjP8i
uX27LbCw8OlkA4GX3IfmyYzZIJedBfgujLuIhTFFaLUJOWjDyp5OPDXrOrywBhyS
mb5vGgJniE1DjsMKBUshOgLwbX+VUlzDOEAfAmCXb9/8fMRhYbqWpINIKDJC4uw6
z07z4hzb8yxy7jKeNuWrGxWE76RyZoWO8R/pLuZFAuDJdJGC1L4aPYCoFJqAtBm5
Qmm3o9T6MIvqaljUsFvz85daHpAtBNepcrNCgt2M3+St56FXyEt37pvhjS5Lh9UW
nngKT7y1n6J3K5QlzIKrbxtCEFZw42p+O2DmUrreO161K7ItdTazlOIsIxDsbo3j
MJQdS0PSx+oZF9tHmStKdT/rw6+wsXDk9q+lEHmAMq0Gb+N8BN9IxrKxVjcdIpq3
A70/D4C3Y3eHOtKJ+wo/cWfCq/Y4+2r1yup69vP+EeHAX6rrAGNKh+ImovPnsN5p
jIaGDwYT/1c8h+n9Tf2d2Gm/HNoToWkuDL40/DzkXScazkIFCw/2g5GRIf9OoUXk
Vu+PW6gaBrfVlVc9bfjPXRH6FWkSjV2R3n0zOvbUJq29fDrgtZlqN2HXBwPFZGVY
ylur2gkACnVA4ZXjR5UvAp+SL9de0nfSIH+42xUS3MvHjjcui6a/1IU/vlJsmK8C
TvzzLHtbUqo58WzD3ZPpASADD/Dzv+uxhbnrQzta+81s67/uWuS8OHTwag+4aamz
+CX7SHuT+Xz+m1cdHk2SzlG1nQSwSEyVuHjW/D62/AqXyPCXqh14e4cWYSgpz8si
DHkYaXgZDUYtqWwaltteVDA9kXN1ryyQtFKFBFmLHuTrHq/apHAlZDNPKsXWEfCr
2HfE6dcrs4HbXBfkMCdf+RXqlopXG1kvBBu0+8iOOaMsa6wGaLWpAmxwZKlFiYI3
VlfADLiryCjN1TdzZ6CDq2KE9QoTTCY6SUwcYyw1zdBsnQiXZyg9gGCZY5cKMHtx
34djwFPwG3/UEPiNwV2yZjRYlv45VVX8KkTTYlcAx4Z2uR1uDfKUNlM1HqE5HiJB
z/CI2poMRFRLQpRBvN3WxggDz3Oopbzw5ETOdN1uatQjrm1WQ6Z9OiUuedSc8YMV
tBcj16MTrfxolJES1pprV/L2EhUbcf26pppufe/F+WQXQx8U8ow6QsrszEs6ki8c
dtdWJL0Uu8YNPykjp4h5obm6kIB3tjAfA4XXqMvsDgokY8aDNZE7UoCLw9UNBNvZ
hMFHyQyT5Xo2bXPAgV0Y3ez6LWqX+Iaru7Q/sEAPc1BdoCRiiKLnsTm8otF5bpGC
zYAukhspLsk0EjgdbxtqTMv2yST3QJLye3Qw+5oCKexfenr2WFCBKQ/NrLjHGOu9
RniTq7tMzERcvoswZkt39uhqH7UaerBzfg8Qf0vIIz9NVfFpLRVspIz1N7TYl4G4
EcD5+plRHE0pzaYtwbTlk8RwnV6nwxKwQhbxI2rsFMpxwCUHTEKEsrIdmWNVgQUm
oAfrP2mN0YT2dCJjZh7iBPn/XLFHvzGwsKCnJrlnO/+v+wG5eqxZyJjhy7q2Z3yD
XWKUw6wbad1Ej7+oPqwdyJoLFjjhsIIE6yp21x7nWQhzepNRZrASXtCHufFArHVu
P3jZpxXYMcUX3a4ZGa7BKI5ZfkeNk+4tOy1BjDkw9JufrArFhav6ik6tPm44R0BX
WojJB9GNPX2sdrc8dIjxfgi7Fah/nZwJQYGABM9MGtzYanVMz2JX0Xvh3oSqPR7I
mN8/VeM0nDJo40w4gX7SXPSuyr8L84nDYmgzhfIV/Sfd0NdeN4AxMc77lAxHtUMQ
lKA2DYe+72vArAN5He2aqpLZocUueNwu9aQQk5c1rP2mN3MfAQ31Cd+Q0BoPfQxV
V3kurSIxbXoclgcnVEUVDh3z0T5iIGSeDxBEkR90+4mnui6oO7tdD4YjEPSEt/TL
cqftM016Yufv/Ggg6bBxq8yBvlZ62lDo1ezN6Eo3HGvRM0F22wG60wLZ/o9Lw5C4
31Ne2q0kBGPKZY68XufvHXfe1cD5P6YPBISUHZzwpOpZ0mjw9IPOyeV1e6zSdLCN
FyPzsCIcWXNjkH2iR2M1aFpf+LjVMKLq4QmX2pFY7MTBf6siyQCUcjiNM+LIgBjU
cGA/YlkJ8QbXSPfTEmXLYPfFE7UcNuIhbnvbdrWUKScNxPq+nMneRc6ucm1mbx/b
xXYf7d9LleryX9HNMumcWZb5CJ0s6ziPUPQL+KjfTdmEfz4uSNDppzIrq6o5g94r
65Q8HG43paGTmcSFOwN3oXxWBvCy8HNHCNGTclDVn+g3xB5cPE54FAAF5IfzSiF6
IbLVZRoSjJ3X9f7XT0KME1AGKy7dH7LoQc4iyYeIo6eZLRS1fL11VbpiCQwZoRTq
H2yIGYKB+1mm/HT233WgLU/9l9FUDamqWjmYjR84zVROI2tUrldyV8Oy9bcF+U5p
JJyX8+xLSkiBOtQlYbx910GhPOgM9ftwMKOd3Rb0ah+lhI+JgYAZswk4eBEqK3vx
9sK/o6uOHr4tmwUSf9n7esUFbqfg7Ec0r+sSa/ut4sJ3z/6f1aW33ES4y1x7Qkrb
WrkuRxkSo2biCDMdMKu4svkegq5IUQZ+J3lHnIAwx8svG6TcB2Y4Xe6HtoBGHMXC
M0ZeMDPGy7uMYfnUsIAew6rBd39Nqw7c4ksUN1iw3iY2sMuG/Sx7X8K8ZPNyiazy
ZRHe59GNBoEQvG+QetJwm4MAa+f3gvJJzW70qbZ7fffXrS/kiuRi0Un1R64cQ5nr
3EMTiG8sIB+d5YWKDzYJXs/h0ad4y9Whp4ZQE7GNwYOREmxir3Qdi9O9Cn++iUaj
J5sXXMM1wQGwD+yoDRsBFifxlpYrmYgVCned9RsmovrbQlX9U0n9nuy5JjV1DHSQ
OOWxEO8mb76PJrDYhirCWGt4naH5HxbpdRTRPklxv2ukoPZGkhHkrypAYftJ6DcY
lk61ShHIHSBcEseESopxFtY2dK1kAcbL81/avukbSQNXXpQ1HI/v3e+YllASj8lz
dUgJA1wNe2bqMFpn9LtB/YCJnuTl/jJECP8+f0ipgmyuzKyn7fiH9TKo6tDJyGeU
L1LYmIq9oervw806q9fQVSNOWZrGblqGbvCdIHWJ1c2cRBbA+7D1jAYKo2ReVZQw
62utZ63nxvAc1kox/6S+mbwYA5wWk1WcKZa44PF/Udfj+nJctYyVfgiR78ITl+bj
is0Q3KXm7BXeVgBJbH3Wxn0699Lmr4pp48Y8V2HDF4xqgesjCfVvtI7JOmUvX+U3
WVINUxJyH82v8nnZdtqYxt9PP8tscLMdMUdRoOOh5hp0IjfPRPp48tU/YdWY2EaQ
NU0QU0J0PMCmYrhoi/hCfjm61S9rp+2vxKW709k4/kXd5JEGc1d3VBF5AQEYkGZv
SoFFrDrZ5TzRTun0Q06uGsHsD/rkPhulSk+nHCLL70zZ/CSDBPuduB+E/u/Gunvs
WlkaU0nI7Sy9GkTB6x32YgvC1EQfVSbId/9nZuwuvqNUrpbsJs50nYm3PSTJS9Ec
UWpy6MeMBuuR+3jfu1eUtD+/+G5EeOG/VO4TtLPTvP0LcRXRDN+INjtc3OGqm9Yv
Ee1uPn6f3EEAbgY7WfekpuXtiCFQlekuhXVUlwPPfm43fEdBAw4P6y6OSnE09531
t/Yx6el0TQwhKKpjv8S8NEISBoiIfRvkQLspLpbBYmin5ZbmyXNHh8YLeQLms6as
JSW1oDiadEoMqiZxi5BWZq/r5A6iWHV2zFi0o3zVdhkBzGLKz7QyA03rw16ceZQW
MnEp+F3KjcXEN2b1trMOPAXZ5bIWoGZrIQanfBd5MDbx0VNNfPoX8tMBBIlODHKe
ROq5gbWdQyAig36JpF32lR8t7I18H0sZTJoccIJjSHB9UO18pnn0iSrh4l46uqS7
pz0mXjaoYVZZN4fFlvtYmKxhPn1a1O5mFuCw7PL+k7Jo7ZAMfxme+JiuO+Adr4qd
L+8qCPqumnesrLB2T0ezMIfmpJwrBt2Xv6S/v3UIdQb2wQ03S3E4+BJsYFlQSThv
IRM6CcQ2uH0er7TK5X29GvLUzzk9g4NfQFH+ATVn9nbcI+LsnVz3R5c4vCGow+j1
WwBY9HXGOCy2k1Y9rWCFlKUOUROtOQjPAdkhDRkBR3qwXq0Z/PBl+0PHJ0KKCiVg
gpustaZSAJKxR5aD6FdJ6WWfBid/bCgc31hJ/BCdebNUu6UV4bdwJuYgvelMABOU
xU8Fmnt0B/Oh6tmL+1PShOAxEP0JJi5kAzSEvhVdW4YDLRbfj5OpZT1KhRk9n/x6
8erEd0nGzPPUMCgLoNjWf6tKjqNYvKfmgU/pd6CCH+hktZKzloSJgsZjOpacce0B
Udt7wjohYrj01sgALShCh7HdBr1EVooSed1yQ2uxiV8mlbhmQG1QVDMsEMIhdted
K991yh6JFenglFWImikWRexZ64QPAj3ebALYiBS1211U/ZZbP8BNjm/QoNQfHaFt
qHN2LcmVb9aY+IlIPpFgmGS4iNwDSURyrnUdURIVAbWDW0ikWZF3Qe0AQWSXhGEJ
YH58jL4fMFujrJRCxeh/dlNQ1T0ARurRoxYAoEKGQmXU7rXKkVgfa558kX15GKow
ab0ayFlzq//yTDUFz/ISZz6n89N6Eq6mpEXPHGBb7oBkqIxWEKh1WEQYPVS66vjn
8j4W6w28Cs5nmsZevmoMPj+GVQtoCB1lyO93IXF725rFASkzz5mjZT0LRW/Am7MI
AD9CkpYENhUuTNq7JYUIS/f0FcyXYiMa3woNOPmLrVHFuL0OpuC3lOpa40IaquNY
VlW8gROrv+OxK2Eiaa9+w9It8calZE4ZDTttzJ6SnfTw0BsfQWozCRmGv3CRQQMy
WdCeQW1BZQXcaHouxmryY84Ou0o42Hz8BlaqnC1XUf4pJ5PIIqZyTS5pe8isHQS0
XXALFJE2OUEgle//SfEAuoYDgqudLbev9QjSsw4rw5OjFTEwPybyNHk/CZZYV8NF
o7l9syAJVbM1ntAAXCvZou4V5RBPRp5uRZgpRM4L+GvLJtqyxTh4uO7SNK0JFM2d
BIvdEMocpOakhqAWdMLBKl1MyRFs68X38yxgyDI3xqcK2GrSiSKpFRKz47K7SOvW
5lnQRDT4L74A43jEAyqtUfN2OLsOeVecvj70LLKU24MO1WxsGDZABr2pSp5H2uJx
g9qPJS4CdiEDhG6CBhvY0FJhJtbe8GbEU7El46ja9Fwama0LttXv1/Kd8ZChClj3
j5+DRUGTBiUrAl9g+00/u3XVIPBEk4bwO9TDWsEMdd1567Tc8/h6bNHDYpzZCquH
OdRh6lRNPtvlSoZNiMHIV5wRg5BRS7ofsxtxVmFhcZHpaxjPxRGb+OnXsJ2a0lRU
Ks1lkV5bhqWh0xynUbmSl2FLVx0IDl9rPU/AHjNgvG/ufaLd7YJLdrN82EWPLK+E
4SZfUcDG8ew8a2+P9HAWrRUcn0kCazL349FZGacWXAryplyH9c/ZEvZS3G4HTlOg
HJ1TKF0Q7kNAAsJclhkXO9A/Qtb/igfgwEUs7r9ihMFeccH1q8rnqi6o8b5xseSv
3wSwgljG6JJdMHUBzmHw32sZxbLInEzRUB0Bm7CUKREOWLfTsE2vC4rlixubLvDt
Xj5KZ57snbs81KpFeTS8fSmAg3TCUSrPrF+hQjqBUETwYhmMA6lLIPMB5qom9EaM
88DfBi2SX4tR05/v1nOR4/2lwWivwhdoMFG2dbecvdUX/eT0GR3Ajtjj3CgHMTwi
h39v/yu+Oe5JmSFKcv/keNhNkr4BtaT3YwwZQi8DDDpZjlIaVjqNBni1Z1OzoiZL
4SssegN1jc9DIhy7mK3ytpo5ler8RekfweF/DsMVZThQ0etlt2QBC5Ox5RfG/voq
I7R76IDdibxQO6ddG9ucb2Hau4tiXVI8VComs/X4CleA75RYisfYq9+0wLDsmQYZ
cHrogedWx0DLfKZrqiB9OLabds3Wc8u2qxM7GMAjElENnkqsxKIGQnNoQOA4v0Ws
bqagwgYCk7BVCWkUN2vUnk+olqjcJcf9hEI7pzv5fk1MjNyE1vpeuLju1QsAwSfw
iII2BiuaVt38sf+HN2qurzdg3z2vgl06lNuVatG0UKbSU+sqFjMxpeFd7ngVIpGn
O6qFOyCbKhxUhfHXBKWK0s3UsCyriGRANDyvE+KqrT4ElIyAfZFBooGkLp9C6cRv
q809FyVFQCo0BmqyJ+DOv2ddhenHaTaid5uuoxiTe7SykK0/0vqYteurVcd97cAb
n9Txp+BeQMsn6xL9MajUIGCJTMjWCVtAgrbaPgn/vfxxJTZuY8SbIPSkT3xgfQOd
/oBFWaPRnQQLK1jVMZm2eOFrS3Udg+AGvtA8tB+UFQFcg2YTofIQWGJbnw2JBMNU
uzC1hc4O7bzUuBZq0e1WRZl/RTUes/jeObWkdeTxwZeWiKikiBEV4mW7nD1HQ0AB
cF+wseQuo2g+2FqgOL1Q1ML2Jg+ZSjOsgsFuIggZ4g1lVigEMXp3+/iOItCQoFXf
qTWnDDVEh3MenkphQlgzXjmlvwKLxELlKIBmA9agwVYXX61vzvDGhkdfkSmunghu
mMy3/8bHNFuOmKHnhrz0Ql7NsjW26w2pPq8cMRKmvv7cpwA1x2+sEDNokYjqKckc
RSjXAcqym1GoCFBUCQY+jsVLgsOASngkY4/H0g3/7MyVSlGy5m1Hn6zIX0IfXyR1
gseTiWRbF3d9htsQgWmRgD7lrHeA/e1zD57QaaRnmHYxJv20f8chFeH4Vim0El2D
6KqbQBTOoSh+toEO9UztykCNZ/abAOxlomhSX+ZpqvI6MCwn+1iUm/qqkJkVcxJY
gtXohKiStLlrLMkYt8xgXoQ3hNg4FHjhmg6ljX/Ojs2I8Slpy0pASv01isWrlYgR
0BKlwyDOUfF1gecVGJ3ycTAeyMquVEvLbHIKUXn3tj1YEsdUCrlHCXjevcKIZsEC
3SqP8TXDsCXap+O9D57/kbgFdqH1mofSMEOMEknSp75JPxTw0LDj0l26tgKtpQSg
2yjzem3qp3FOTm5M50dmmSMT/PhFyZOLerqhcsToAHZ6qmfc/RFLI6c4i8t37X6o
5A/rqOJ+T98T/anOzjjNvahdNiy7atEK2ha8fbOt3eSCiz73F0621csuBwKmi2s0
mB/+RzB+YNt4EPJmAnDDC1GYYGr09JDlpZIr26ckOp7mxCcvx3lGnK1hRHgqhNXK
RT8WWzkU89I2VjT7jXyOrroSvtQUwZs2gBsrGUYFYMwLK6SBgba5T+8d2akIk6b+
vdDvp5/FWMK/wXAJn6sbUQVtFOe4FPZhwsCfKM5bjkXVCyayJktxEN5H0QT/L1dK
cEslqIwUFEMkrjHNG3/y7Fa/BOPLzPfAlGfsW36c5PxkvGe9A2YTWCSodGh6qNw+
iOwI+3mszKQC4zozPv4DNy1LF0LUDTE84EVE/haeBCR/Xz6o0YDapJY/UzdJIjlW
MAcyyPwNn0hFx0qw/B4E6o1zIUjoSwUPDQpT4BiQvU/0aavvv/brkj/CwMX2xaqm
Cg8pdFTXpqgg9kGP9I++nAJNewcpNwZZQbyz1ytGY8mYF5pEJKAAexCI0nnCnDsT
uFOVI3K1DZ9LwBt8FMDhVBpCeonAu6HL+IXDM7yL/wduLDUbuchjRmX8lOA0HkIh
4DZ/3XCtEp5zTz5ozoPGLnnSuX3ryCMRjKUhKeJP3lo1TuPI09V4x3pztuQR5rcs
J8e2KY+Dfi1aCSbCHs310Idbrc5iqFPS06gSyAqpA6v9LRSKFjdy8AjvQefe/tYo
vjb6LMxKeFXvGeKUAJmgfBUq47MGvrK9VJsIMOCS21GVqSkkvwlX9DOG3rURP56b
Sl8deAq8BOdCZ526uhaDJ5Ug5MObHyCSI7fiK5caWcC8SNFvM3CJ1wTufy2M9br1
mBIlgTCHJU/qNZuOwwlFZ8DhkGOnf4/7mTKKDZ0IhxWq7Tx0Zxt6CYqp1ISpZ5PL
OMnL48l8bKjMyckEMrfCpqQ1Vpn+uecTcf7/inCcXxz55xRqPG/HRSN+OSH2T8YY
mZfVF3MuCHuf3iloeqd6CGnwDxTd6R0JGsBJtAd6kbY66gsEikqp5oBAqw5mvz0d
UtoVKga9lMsGQMoUbLy+5JB1VheDbLdodkvY5bPtlAPG6fv0N0M2Ma5YJiNaANIu
KqCWRHtRp0eBhiCWCGlWbq9rx9hchAOEt87Tg7NKeSkL9hm57y3lBYp/+5t5ZHJw
Y2SbDvZP2ui3waZLxPpSvIkcwjHSTNR3qgcKrri9E0WvVHohcSHr8RSYBoyKq9FL
MZFlInbHPP6Ijk8T6YpK5hOqaPAXABsKoJoz9KE16cBBflVKgZ4d92IaaXVhwJiD
xMaanR1p6dOTaS3Log2HngityxTcwp+1+G1d/cpY2t6EfrsrTvY8RQYo7IpFXJDj
xTY57YopGIZC3lu9d/IQOZN0KUzrOdhG9ltJbYd2a8tuG67w3AFm4Kpaj3ojQiCf
kxK7G3aZaapfy0MREqH2wiOdPDdqZ/EhwNAdnbKxZo+wBFkBBCp0qoNIFQuj41un
dJukzLjSAtaPY/Tsv3AgvUAWb1O3on349mRwEb8+IwW8EoqXOZpoBj5IbgKmJ/Rh
0v33/RCvA05QX+YGQy2YlR5jIHOObei10riIHHgAS09KMUW9J3PYEKKGCCLKkrOa
2/Zfm2RtKY/QAKVFak/ZdlzLbP2AeKgR5b1zlSQEPiHkN4zwrTmx8lqIRDJSRl6T
x3miG0P0ABuYkDJ9vzrS+9CUlesOBvoZaG7018TjPKDnClMvbHVGarzdGYcywtIM
lR5qqAjKSRCF07NtFx1Q6AC9jyUG+/u7GEs4/+a+ehDH0HEdLDXwwjltKKxwXy79
0D9r4w5RIpX8TyJTR207gOw4T3CA/JAeXW+uwnkNbXjVehCw57Jmbzra5RrwnDBO
0/gPlYDN/IzuwKOgm3125lbswDYFnZSRJotvHdEttijs/1U4zOXobcnNc2lVyx3+
JiKbp2SbdxkNKabhl802xb1JdhYXguxQ7E3UuAWvbF5g75LKXdwTk6ldhuePY1Ff
kOzfxbVrOQYWyZ/lQ63okPYcgyQl7cnqKpcXTghIofnGDt4iILJcjZ6YQntGkFh/
RtfqJJHXwxZphEb7rkq5cxmz0wNBceWxT2Sp6mBnHOpHtD183J+l4Od8pOjdDnGS
q4ad2FdqpviqYjQnWesy+1kcZv43XQj6FpJYW3U+Dy1+g8pubs4ubFGAvePSF5Q5
pS3gY0dYHCXcQdF8iSC7jIcHM7w7Ztd8hIFt+EA5uIwJk2xzTDOgu8unIsQ/qH0I
78yyASZMFYKlQUqWRLn9+zLnwDhgVkvlaGnD/90WhMVWP9B4ZZvlELJRjXaS3AI7
+4Jd4LOx3rG6gubUXz8zKrVFwzqrx1bnRB0Y+kUpf2ysKqT526Qiq2DfQ3NrF3eQ
tsy4joKAJRxQ+3D/F9sNZ3WxiJSZ6DFyilFsML5BLDqvvdflu5JjMY7K5pEFiA3y
vil6R1RZgfXXWJt1xeQx/hEhRMOp4IqlUA6bY552KlVQ15zPhW4/R8XMDQOwkqG+
FfRASM6CI+2DjR+2s0eYggVEH/Qm13ccapVK7W7gKXD3xuLgDcw4UJt+rlrgLegM
3HFdv3JFfnmk37PpBwREg5h/Q7yte9b+HWjCJHliuQSrATpcdbyFQsrDVGP+Quc9
1Oz6IxHq4s4TLGMcvXsc/bE4k73QyTQeiAGkVLrsTMJkwNZANFVhHi1uIJoTkO2t
NoHsh22HiVTunRGdldhs2C4Afyq5JCD6onS2MF4tpXR3EeJ6bIH87EEhPEfNv5OE
tppTs+/NAj25Go/gIlJgJk+4Tw/whB0croZ6/NE5EL6wwACQOCpmM9fxiLcueLpz
y/oxwKd1L2cgtKof2vJid/ebWbhieOG1+vjAFG0fHlaeNgBm5dScGxC6ZAKaE25Y
Hk7GKlL8I0fYKPnedC1C5IyvMboG/o2eeen8Wlr3gG9BEgnW/OgDI4XCEawPPUQf
tCYBpaLuMQGrkuFJiRjZRq6DmxudqWNv7OLNsLDJXZoQZEuc/OpJy/yJ7du2t9Xv
BSKHkhSVXNgMFOhoj7ylGYCsk6BfoAdKyZlj2hqidgvIcGbyqeksBsszztCdLcfz
GFfFVIGDbiXn0NZb5ArtgMZs1b9X+Ch61kmuULLpdrSrvXrnfPVbnk1uOFqJi+Ff
9nX7IGUHWneLAbcpZmbyrZNaoPiVRF7qC9dJSptfVmHci8ULO8bLnDGuY8FS2FhA
YiRIo5jD2O6PLS8mT5sVj/t3L5qhJRoTmbXQz1Hs/C1nLxZfh4oHCKHE2zbD3xVm
+mn3N7cse3OSDxOu2+pIHuPbvpXRqtXbz4Eqytd1cX6Oc76MJc3OTkmKaxAgpr4y
/Npe7kYFdePSY2PMQKKVuO6JHK5a5nc0+j/NvPJMFgRlxvn/2atNPTPidKYrapas
z9hXpaiYhcgmejTLD5Wtxo9zl9fPhBVJPxjcB7GTgxHbfaWQKjPiwU1O0Mj6xZSC
XAUjpTQBpaHn0Yj3eyg2d9lgny/Ohn7DzWgpSU6O8Le00tlF8oco5oME3BhkN3sB
omplMVEzg/eb49b97zovgmY9S5MQc+tuM/wGUI6RKFj727PBP3prGd6F0p/n8798
8qPBJ3/S2vYN9Vrnpwh1JAePVo5PviV7/hjCGXHdQVdmmz6ZKqr1ZeTrJL05bRBz
O2yBQw+qDQ0nQgv/VZrxhRFwqKF1MnV+pM4Gju0Zq9Nr2EXt3FmJtx8zClhFjGJ+
uLaxWEVPXzdEOxKLZJ2S/RKGy1jw8jWBb+amSIuSwHWC6Q77dCGI55bpDU3zsORw
HXx/8dSljYQVjDqTFOtWgL4HG+tAbXXMHady5sG5ife2yCBVP8T+IpR2jcSUDjOF
/R99ZlyHJ5IThDvVe/j0QRlo6pQgYysjD5mdO4Q3IX8PU0VReakP8QdZLKC31oqu
gou0cPKqAObPQe7PfjMFH+a44Zi0qGZi/rqTY97MLHVVRgfW9Ye+8UQY8GmqCgDK
ag/+GsEanF6eO+XsrWUxEhfawFHi8j7oruZHHRRbnyeMlDOvvtRq+E+vTxLT38nN
LtAhxPo7z/TIedAWDAqG9aX2i/5huMI8zglRg9IMKrzQS/9N3Z8W9KoVxZFOGpWU
3mcepg0zRfu/ZqyRzcOkHSlkmi/Nw1UobDwrvDx9Fjg9Ot4/MGX7VPhYNuvEMmb4
Zh7vBihWikiYNEtbLuDTrHDxHXCl5fmq8kP33Kl/K97XO3C9oSaqnLZZsEqXJHwP
8SKBh/3JRelnF9B8z7NIg9S+3Q/xQq452TKdbk2u0QsjJ3o5lsoue/GVsnI9Oz8b
pVTyC5d3KqmgodxMs/yKQf859PPIAPFirtmle8dpA0b68mWZhZU7Oj08qRKjbdWM
FtueNDsB7GVoxizQ8zTw2k8yjx3tYILEFB8CTflm4rE6Cg+hS6hLzlBEzMlcgxVi
PQWGWMZLY0unKxdX9m+I/YwwGliGWyPX50qe+K5/xAuqdWfyGqL3gQNXiy4L8YBZ
h1v4T4RQYJxGdSEatezQpFgOJXnfWpSQnkOSdoLzAcm4oPCYEltrzcC2daGqy4jm
I6OKq1t2Z+5dU6rcSeWPRkdDbXNQrK+QPX9zjdwg0AkOcyeB2rfMPy1rEhyiUd9d
mqdufPimaKPVSInewkjlWr/ijQom9vTNuefSDwtBPYTTEcWw3IjK8LgincAyxPyc
rc5G8TpjHkaJSR4CMUi1ypIhX5pB2dmNAMKU4y2MPj2k8gK0HZbG8kXcB5cS52vO
yoNpKNjuLqR07cmFFMBXNOwwxrXk2l3Vp7j8R2irkCWLJYyUrBrqffs+nnJenDTA
eNJ4bwUy9NW+h/hHmQFbpwdx2QlLizBdVCWRhEpTw3GATQCia9vJvrOn05itMql5
D2rU2qV55ha8n97FbBoj5f2w3LxNheSsdB2Aqz0UdcGXVQKch9PgUgIEhkxH2Ljh
zH8Wito8QxwPXshPI/QlNiK13fVKclVMFlTq+PqWm0jmCx50ayqesAM4ijm8yapT
p1SulWGjEMU+0Fkw4uDzbaQl56zLPJZFNTKgLyGzqiUUrvdVp1kKYCrk+X6bjEtr
ggvrnMquyoaeU/owO/st4u8R1gELOBJB/nDFPd6RXSnEIOpbw2BSl8uiA9bTvX45
uhCyHmpSLS29OrxPJrv4OneDlCapVQqXIvvbSy4Ov+eYcVOGrtpu4E19SJnDP3jJ
/yIGPd07MqTc1U8RI0hRnKaKx/v1nFDxZqeAJPcIBGWHRgKkXS6B4W/7ayaKQ3vi
QFmAbh1vDImNv3zMHmlAUiAjEnm14VB1v32yoNtRkEgq4v8sVjZItlbplwOnktTm
fQ/whbOLdqJr8IgWja+GAX5O1yEukJHdZf2nK7qQfWWKf87pyKSfyP94XcE0CpWS
U6j7Q2ATx5q3lkKsk3juOQ+WEguzw6xSb/ZZo6EmyCPMaeO+tdN5THTL595Di0+W
dplDdGkjQjLsAW93eWdjtb5DfD3z1cs4HE2K+ZLXIm6ng0WHpcenJdfyHyLbdmsb
mpbaUzkeMgOypnigQg2Htszaksv9tygjvh8HdXvj99o5ZK//88t22PSPnFJhrwkH
d1j3OofStXx8BgfyA41YGPVTpiUFwqqtr12BqmrGZBnvCCaDBQmLW+OKYKIwETRC
omtVYzzGBY88pzhGGtCY6pR6cDflTfcxnQ9jPQzJx7WpatRxOTZsmXmAjGLYWUa8
EsJgL+0BsSr4w5fT1Wmz0Vtz+Dv9+vvlNPixIfrWJaAC+xiFfTAut4HJ7y56frTn
0B/i0OSR4Ao+sZx/SYAfOofIi2WSZoDpxVz3tugRppK0/Y9CK8PmAVGMLxA63XWw
TsDp5jeWl4xLk69Klks2VH9mFq/BxbpRw03Se0UCapk9Yso5+RdVdBECSRmC2gof
wmQbnrSfQSeBgHO8Jm1CuPph2K8PggJDRDGZ+Egi1UqnvFgEBgGWoU+XNSN/eRW8
7roWdT+CFP8WHum/tVe8FiheiUmDWtfnqA90HNSs7WOhsa/eN+fEeYmob2GHhnm0
bFtyfXz5cTOEhjVjzt88bAFAFPNI6+rpyD53TlvFwduKkIS6R3vqtG9L8LnCpEnG
dQQnGJCTCRYf0Ihru5ew3+Myd/zpBfO9IOVDLkDbLW3I/LRMYFeflxqePHFN04jY
ott6KtMY/9/T8r5s+zkh9Md3yX4DwVBzvWlnoThyFykqrI/gQGEKvswMHp+GYmUw
Lu1v33M8IECNWS4Luhp9+u8m1cVDSBPT2LZw5aLiVwu9PkDT0Heo14R1tMEHN86+
sb7Krey1/7J/bbmFQbRJcVHUUtJm0uzjswRyqw8metz7suiAncdDQgFwTNUb2D3O
ko81ToBH73zthy4tssVTEXSjz5H5wB1fujR4bdYYszcloM4bYWmpbRqGxWGFM2Jm
0d3aYJywdsbouXlUCTRQDUl+vk5H/M/CDxPOT6rJkojVxPaEQDCqlctzVQmrrWjL
xA5zIpAdZPIfLvMryfIbSKs1++0nU/hsCtQE+CecWY8Zrwh3I5kNNrnkpbbNnasd
drNEQh9Co6sczbAb/hrmvlu9SnzKbCbaTUkmd12ApaMCRDmmEXNDQ4/Nwwco2ps8
CLELctTH2sR0j3pafhin8/09dJaCjB7EcK78SPAVljz/FrwIkDGWaEwxhndjcfg0
d+KFcV/kJ7RXr8GI247o+Yusn3xBrfuIgM3eWvCVwv8MyALX8g9OMtGmjdG3fdg0
rbU7Tqc0x4Q46Oyxqmzqtx27QAvL8jSLA/bJv0DCokOaNraRzILZDl5dUdSEoX13
F6Gjo/AIzu+eBLCZSLP6ChfpStE9It23SWknOzmmq6CGM+NeP/ASFoYfDy+BUy48
7c/ynVdZXIA4iKjXXYgmL63J9y77Ullwozy3ojCU+w8PQxd8n65xu87NKw591yb/
/uYDBIxrrtBRPDSJ8OW9bKQ75ePILMsUp4oWyWIM0hKjZInrrZrMav7uGKQhQXJq
gA1nPnEJ3tse8sBMrmNxhord7CdriR90oz6znWgLH7L4rwRlLOtx+9jgfbQWJs+x
RT9jUx43grUU1SW2pLO/HclhDKHnM6Sz9LxoA5bDOSutmHPPIh4C1oMLMVbAbIOv
zC3Po0CuCU383wkoL2KriIBNZqeMhB69eWRpCPI5EWYUqynl/TW0X5Wrt5tNWX9w
TzFiBEYqv8T6vR3QhpMNQz+wuhf33uTicbdZMjkNO32ic4zX5oxI/NUdNw6eRnn/
LlRmJfbcF6oLDQ9vmLsSxP8OBaY8pqWBdu9hQe4d0HlXRCpScvUIXeVd2FdySuM7
9NHW+/6PIDT2Cj6RsUnQIMhWk5Q6Q704oDot5g5d2nb8sVb5mQ0FH1CU4KohE3dx
Tiah4PqZh9/DEkUIpmjqeb0tvlSKFahhaAMdXQ9yrUhfBp3NTuGoO0mhrY5NlIAR
ptYQf1hk1x+6OReyRyNhERExLnLGvQ5TU8tK5P7Ll3PnN6JFSz0fTg/Bp/TNL6cG
buw2uZ6sdL1/hcZhY2cVcDk8Qpis+TNwFZXH6CiuemGwq03ZKhxZNuvseU8d+v32
iLXU7kOM8DsUguxMHsOfSKia2IcLyenLpwbK15xZXt37Vqa85WSWgrx4eVToHT9t
hoxEEghO9o2ngVd25OH7HQEq/isKz8soj/DucUWA49gxNfxSvCGefuCBOsi01iSD
8kNt/gWegGn/u24SRz+fZYY+MqRPHl0MIERcsapfz395dRFI+QzHfpAANhMk42Ed
jWxRB1xlX6Jh8h47AQ1XoDUbOa157MM5xYWua4jhFJNGf6/Kpqbny8S5v28iMtbU
cYWV0dKAhe9ID7KKE6JX8hKgan3P+/D/nALymtpkNthcm7AChTpKuP25mSknkPa+
SuOzXJfxmUP9McnuLpYqWnA7hwK1Yzaeu7Vyd8eVA7byCf4+qKJ4EB9sxecoTCFV
k4FF38GhzLwKiT5vHfWHe7MBPNpAqZdt/hmYMXsjWXuqkhwY24+impKu2nNPszan
z4Wq14z8hI/uV8IxurWKOyFjMGKQF7+yLa4x8BoiBO3Hc3b6lSC0LzpyyBdDUEC1
Mc8QXfTISNmd427uIfBiaAu0miu/8jBvEO44IQnw2dqEWs5npR4JB7Osf9WcuWvB
bantPUxISrjA3UpTNJr/bAl+aNcCoR67A5I8xM+1gwpMZjoVuvosXu6CCemnBeg0
1NbxxZvE0H7b7mBuagR1O9b2OgmQqk8I0neUjkJ1TBQYPNleYEg/GAd3zPZ91AAz
GHh4CJ01g3HWhF04FtjbvRXQIjP0Nqv+CA/A1ZO65FzdY2MdWQ+N4Bp4dVW9921z
//sG1xgNU12iyCf2hGt+uWrvbHi9g3divIBKfjY1SS1EhdpgaZLQX8t9Hq4YZFRk
kmZrgHFs+5EB73ClawigAlnXvileY7rAHDNSd9YG2Ih8sUw8L7za3RTngnubdEYq
72NbgSPoCtlD7mS5qNoyBuEdEl9XSLSNbf6X1+gYmwlKjzxSkYU1j463q+RX/mFP
b7LPFRiRYvP7wHYecuaHfuovAMEQxRaU2pwrla7TJ8P0eQKCWx6C9PhSxa9hp6iJ
R2wVMPdX9L7FAgLtceja+/Bq+o9Z95xALYZqVU5M8SBVlvn5w7QiwXG7F7ZwTTS4
7SqMShJ4cN5iPLLRzzNoRdeSG5kc4Rt28u+lYZAWso8wnxCdsUg6crHduvJb73Oz
nL23lJ1Rj0xe3pKN8GCBvDaj9jVvV/+dysJqTica9CtqjWJzUZxhd0JRJWTi+twx
CSYMyzsWVrBKoIkYGFKYPrPo9l14Ogf/SNK/NonrvWEblUi08+Df5b1reQkK3o3X
hIE2uAu81HERmWx1hM0UPBo+Oa9CpXH9HJ7C6XSQkkpoC+2MBb7cgl7CA0EK3W5G
W1UxKwbOryZJ7POhD+xBUrjEjtRIpN8Dof1HnRmk+rs/SMeEkwN9x1cr4rW3zwb/
CFnm7n0WbRiVvQ58t7+/PnQxaBfZqPYAvQJfXs4pSU+FutIIm6f8bBkZwgdcbAIt
ms4fsJ8iDznFk4me8RRpvCboaHNO8gLQSebvkr4DIJWkavPbdNH1A4TaQl3mRLXO
IZKZYr9d681aZ9qWqKOYW8tiBy5h1gJJ4ImQB01uJQuN9V+qnPZ+vdQBRFQ+mPoO
4H2skdcIJeq+HCy0LISeZNw59yc0I4roXY7P5l1dpzGa33uNCAUzi7jphhWisPM4
BkPUyPDaKootvcmHJfzm6+e089kryEoklZpg3cGP3woFxJHk5rYCMU6TK59tjxIt
3ttxMkHodovh8ZgoOJzIXULiwo0EiB5lLWYT3vX74jwVHuJD6oyOeoj8tVdcmv6M
jHZCUb4nF0B4NoFIA9H2KCXMxA0WMW12GdInH1PMssaMPpfO7bVknvXWk2MatsGx
DqntZKNzV/JwXI4srb4KU9VftWKdsV3aAXy29v/xapWUQoW0jB3dzxxPKCW3bOxb
G0T+S3LVTz1JjCG64xzFdlrqKol/ECoTjdXw9PglOdrPqT1FjeuTuzf6ba0J2Uor
+qfHzGRh2RVL30wXu2IqjY4g6Cl5I5Elu7r3TIznqNUezVQJQSdcj3om43dn0rl8
OnW/Qynszl3XrrZH7n99IhstjZCvBt9jYML7UJ2DafK6yySeJp3ZV/sDYbtI3JLS
kPk7xrnnKWuFcF7BU5xmeZy99/uNdgD3Jdr1QO3smrUqxvMdn7sNIFmdHC8+ZTFI
XqBDVBQyPVDgVNmkr9Y7R1Sa15TkvRxf+80+SVzZOaHXQ884X5NFJRHggYVib69O
TYYldEyzNTB8nc1GFM4QeHtk5kULem/VdipYQkZujTb+e8WRMRT8rOyvf1P9TK3w
6RwIK8HvvBxZolZcCa3K3jduBCO+mZ89Bq15gqfUP8UMjMi2ptvcV8VRZXSO1riM
DJ8L9AtPVBa3uf/f1M/jmKJss8AvhFXtt58S/B1cS99XY+m5Tt3XPLu+YceR1y5I
C2uDyFolh8m+yNeUqQsn6MgydrGjheEOJXXoaiDRtWdK1FvgWsatxwhCsAdxbAP6
aB1R9jLnvZab07Bje3kxvoyjgmJ3T+KWHN1gLx4VOTluA4gwTnyRFTJHV5LNQgFn
iD1CQA8oQtUDHmKycRMpRPcDK1FYZ/VKIRgxsK8WZ0t0lrUNoorDbiydyxOkgme5
S5HEGHBGc53aswVpXC1BTlKwLOl/zt/k5DxttxcJ8fIIevbVfm8VRcW4lhebdk2S
kZHwmRK5o9vVCeZ31rfmjJtRMfCaVgr/6d2Telkn7PCFt4tWt5ahQDJvYhvqHEpc
mwPZj+4N9nulwAtEUyZLmUXAwAntUJujbeEEfgd+9O+S1kjw0pWsAwkTku6HJzuJ
PpPq44qJHLOB/GpD75pdmzy1Sk39ZMiz61DFdsuCekEypTVC5XYbxTCK3HvUk1rP
umCyr2pHJ+s9F+KwcIEDFJ6DuEBDlArLu/AF/dCHbMtgWZjI6vQDyamytD5Z5DKN
NywSfZs7Ous0yTkv3mQd/JcLrJmUAstB/ORH8HfAi888ABkDyId0pxr6w2fGlYFe
N+LSkUQCsXXkm0GdmViNIVwhsefr5IHgyNokhViXmN9mqcL6hzrqo3D/mh/ZUdvX
PmhbsqSkoOns3b8UQQ8zJuKi3RA69eHDrt5Zfsl45+q/T5RbB9eLsx71sS+DIvn6
GwNdJO+dY+7OFctZfrLb3KNS2aVKYER6LWaC7E+M0n9D+Ka8S7kx9DTJfsiY6nD/
VgzzACuvMp+6ZUCHlGuK9XHoqv4qj+EfpHNg/+laF065TQas4CM6/Cg1Z+VI9bMH
kbQtHrfeJxwFqQZOs+CwHgBmRc0RfB8sqUsJ9UwuTWWf6YkZ5fBkJ44kw15+Qluy
o/qT9DjesiAw/jwxLqxMGZ3dIFKgJntganXx6wKl4f9TWtyVMD8pNgpfXqoOaUvA
j8x3SZ5rlh/CA9b5ocmA449R+HWZ2NVOW96eWjfPSMrFCjyDkl2VuMcSs9sDBJuT
4B7XZ56FMZehboViWi7c+tcWGvXKzjpZULQmG44dxKSwrDB8baEGspKzHrdadmOi
eFwp9ipJ2CBpRKaIPjwB1rtaBmtPDAgrbPBbxuyDc3UmYJkxU5LKindJ8A073O4H
uyqn3SwFdIHy9jz5kpIY9NoGuGwbxvp8JG8RP580VVqMCzS9ZqfkBr99K/32c3Av
frf4UYnf77NIF1aycNH4qLu5S1+dOpkbv2oBXKvA+99jmTi7SaS0Ur1+8pm3U+2P
5b8o7YHanb2r8YzJq58PJwt3e2MT/fUYUsnh28D2WdYSs/0A5KZhgeT5hY2HQVHk
XOT822KC2NX34RRs2LB29Htpedii7zmDi7JlBxz9ltGYDHk97qk3qkV05q0UqDpu
8UO+zH1pVzCMEoOur1b+x6NuFSTNZcDfhqy05HbsnprjeUbyn7HOsYUGisGcNmJm
0KT0Q/HMUlwQW59U2Q+Tms2aPtyIXIKTmAs/7CzCrff9OZlPM1Wgl6jv/blkB+32
qhre4ItcHw0i0q4G6gtp601NmV+GFSEvqwUOYe7FIw2fgti6aSDNxJd1hyvTcCqg
0jsA7kkGjt7ShEU+Z7AWAeH1w8C7ooHya8qnvHv0Tf/ean3JyCgyutug6F0py1KR
c4i/nHfvR3WYPGwrhGpFpHUh7VJlXVWPai8qHEMa/CEiM/B9dnxT6wJ6MHjvHAOX
oesCyOnJP1lkON6Lr3RRB8p08V782yU6hGDB08IgF3c2VG6DMZWh48w8LDzrlnsa
KZmmyLUE8W+kAmRyGyXO3amHyVvOrbf0+V8AX4nF0Qsfgj6yArIyd7vS1rSZVOni
ZfAze6pYljGG+GQsLJ9yrdI0NPycS8O2ajLUWEkYbFJlPDhXdm3ZMKpNaMYSsO6N
0R2hoPiwzCrTlsBHviuhtEVpaXuxX0+kPcCGJ3/J2U+11oRmwAo+YVImY7tc3LBy
drMRcdk45kHFRxFQ2sWaD6hsvVfSO1/2qrlSxVPURcbCH8hh26mjtMrlQcehoRy9
P5lx5D8tM6+QuE0uMe6xt+0gVP1u+YW4WF+nWRKaoUj9o92adjY+JKIjb0rSleAB
KlfmjCJNiulvNMZaujWDNC3tmhQUelqtGJ5xdXch3137NBJpPZinsUitYQB6ZBOV
8c39U0jrzNPVLfyyL8ZrFoQQigE79a6tGIGs2NcSJ65AjuygiT73saK+jrq+fIIK
unVSIzBuQvm0nzQT88fCvXnddaTEhN/+qUjsSSOHOMSpbaeCQGClaAw1IVuTjYx9
bVF8elUBnK7gW68HV4LqGHUO+iAEaNPGS7m2wPxtffW6CzSNtu4UP0RI2aVLhA2f
Kly/UoZmWdnSJvG2M2+yJKtix2s56QGusjIwxfP2a/194ROrZ/cd2j8dFCp+umfo
pJ4d60+l6hSFZRInrDOXMguyJ9bSNL6aZC+OimTnl4Gu3HS2sWQYqKI0WdwV2qJj
CtqINAqkWiULX0XEL1cWUNykopgBMfMpvnTZZeE7UCN0ebp9kRHvr5Gv7U7p7VAk
P1r8XHDZgdIkVSIjWh3LQl0by7EZ7pRbSQ9CRCzdPqxmYdTMA1Bk3XR0JZ23Sy0t
bghRXlQeOfeCNgdIAYPdRV96RjIIGJ2f2DS/rnlEhuqNQQvtmOeH43HHAxpxonfL
rT8HEZNUx1RrESYrLSBPC2Cb5uDA1QeV7nuaFBmLCIt8mCXqY0EmxhlAi5R7Lhc+
DZHBu8vdEtoVmwlh/CHB2NFFfWMrwqaY51xtmem2DVgbGvEOppPtOmf14NZZmJXb
woNFtRQ49sO9wEA04Hg5kA5sR22m05hsovIzKIa2wf0htK8xm8R78OwtwuD4f2pI
v7b9NM8qoO3d2NcPYN3LyLCxRJ2s/qGXo7ASI2Sacs/3B7oYNh+NdsrtdhcFbeC3
JfecWuI/S0j1lX1h7HNijVS6rRyj17xuSP90XFbPFcA1rp2qGWWoppgzVOG/qs1v
+Zz5FvqY8uEpjybSCEFMmfJsfKzwhIzc50Jjx+a01RFbe3Uvrzu1Fh94t2RTgo5j
EWAw4P9eT0jZqrhOgwqW513f/enwofNgM6bUiVJ+JRtzQYOUnpA2TBUE7Caab9zK
EIjn+NM940Lwc/w0kIDj3fuNljkzc4fYfQdErdpEdOHKsN0PnJofhu320Exz2zL2
fLZQe2f2t0Hj4sb3uSQRLzjYlelGVbxuWN3U7jcJW/b1Au53TT+Q4Ejof9Xz1s6U
wjopu2jykgwEHqMbWNSfI+Yhy4Xnz7xsJTmL9yfh21Q7zYC5uBUgrYzl6UQg8x04
yRYPGODS3VbmtUl083N9QRQ/+UyQYRaNc6t3pPP6dLyFqeY9ui5mlLctyo7z7+7g
KnVahVBmbLp0myRyLJ/Q6wUzedKqFMKVPs7ONWGiaQ/zrxIP0Zyz/L9ZZGfJE44+
/G2Rm09ziJ2MqDTB6jsQZdjhjAJzrJvyo+OAj9leJGt2rXrveYZTcJpRS38Ohe2B
nk2V/I3zZNM9LYGqNLmAR/5VhhfwYVAF3p5oeXV+uchJsqx8ovjHoVMWgHjQOgq9
j12R395h0uUwB+8kk2ahiBJbpMigYEhJS1QWAWZ+HY/U1WmKZjQzpC4kX1gd5bf2
tK4hLMmgnA/zQno/Gqhp3HE2ZQxHWVsw1cAtBDtDqYnY/CfxvGzIw6Npt/KJKGfM
HrcYugjGRzqMbA5hx2qX+FXNMhTmq5hIVNnydThmeWaLblBsvo4wmI2V+Mp2yhNa
JJwxc38iaPMjD1gFq6juhEi6fHBmw9grNOVONzmxP6HWGgEzIDqHMeKWDRv7XLdH
HsRSOkeDI1Fi0MpCSGCjgQDFmww1YJ6smt287WRLneOnNXPhVga8KqmhUCb/StsH
LkZBDEF69l4UEVqPVs7tS+CcavOjRLpLhmOCdK4U0Ez54MPKfkIPFsUFGoUAnW1g
2uL1VQGBDZNnjBwGPp0Bhma/hPCNrAKGuaqWRf0fxqVKlv/PbzdlpfleSYCl0T+I
UqjgbYIi9ldsaEy1tp0mLvzzlkoBGOKAynMX4Qq/s9hozQ+RuOU8raQmA5cJyrmg
b+1u65SDDH9FRE/wg58DJn11/YloMPImidGQ/AktIW9/VE5y0x8AwTU1uDMVFE9e
V88Sy+RZ5CQ0ChcXOhn7HewMtAoktS2fa+tGNcVlVMoWHbWnnSDtDeIPdNkEEzRD
0ZfgillXi9hmE/uxAoLVcqV1amCVzwzzn6Rvq3TEx0ocudeRktOjDezN77NRNE3j
5FkRI47g2Uhl/63RKK1alWfVks1oZzja4c3Ujm1FcNIblv5hR/5YJE/ZtRPZYQAs
Rn1raXjALrkz8l+zSA2pR4oABRymAgeR1R1CWGsQPrQxoIeEHpBTzelIaR+G+M5O
0Zla1Wak7EI2omWo8Zq49CUS5iDftxjMXUrMvoRuham+1ZIlcrV8YMeOJ338DmDB
yWSZylCoj8pPqizIqY9K1OavACb74r4c76jpznwAXbXbxmMECs6L1o0K19I26QQD
8xT3xlDLBqbtVbGAWP45KSWgG2Wf089UrKP4w5DKVWtcn2UT5DMpzwPTu53PLXLW
yMhTohEZWMW+GsEQF3r3P1a4B/Vo4P2ZK/uKEU6fFeSdOg7Xzcw8c24etNt2ZkMa
3rf/0UxMuEZygLg7BMixB2hqyXuM04MmjKMBwiNOVZZN2KglC9DAnQ4UVCBatmH3
AKivtpKLibiM5wDbEwHOl52I0Sn4hBWIq0P4vFCorVJM0osPAc27Mlj4wrqACNTL
/kiBSlUjgYF2MBY/ESpOe9Yw4kFZ8+WY2Hyq2BiOLDM4+NtcG9FpZMgWW0ENWv6E
lxaMSRxMqjf6Z9N3t3mZuAKxESuWeKmvFuynSsyCukw4mWYL9D0HiHU02VB19D0S
RbVzGXLIYeGDIgtap9F2piZvz3cAvi9qTNSnXhwki1XIWvVBNDLLqTf3dpNf0scR
NWihNUHsXxFd+Tj5G3Y09U+g/kFEwLkmvKrhxbZ0s9WAm4TxU2YPsSNd8an1I/65
1qOLhPIhJal7pJDWXNNXIr3+M3YqOG3haoBQRkS7UFrEYDerY7A/L86M4R1DgUrU
VX6oa7XpdVXJeo8t+6br8yV9uaK+guAcK1MjZn0hY3ADrXam0zXQkt7x3CdeXOAu
5xogDUE9zXiVA6uKKhYLHmGW6h+GtkKrXUMwzIVaehefGVguPyBJ+UAfqOLJOqGj
QwIa9mfIj4pMkV3EJjYzcG/G8fdLYhWMGs76Q+ZePZm1YUGirbKPEzCjaTNrkbvU
HTvoBhTfOk386Mib5gB2cqmiXg+uPkTsc0wGVyyWWWqM08kquyK6UKvH0tYPnvWg
YgH6sqlhk0NXh35gxf6XWGwewczU61JoOS36gTuSIonJ0uWm4IFYiBRzppGjaKad
XhrcvChOVwUHigJKbe08UkYUwzsjXeHbe+69dGZRxPJDBjqZeMRjLHlork7cjcY8
Wm68nSxU1ayTiefkALC1Y9xPoMdH74YYoAaW6fbUjNN6wFKANMmAxjACKhe/ZaHd
IH54lp+nKkmh54MTfJxUScbwtyI9OcLTu7SRpFsJcZ2fTADipZfRxxez5nhFhi84
adD3FQTAth4qcazve5orV56wCFGwhWAOkSU038hGJL8CXKqRwGG4cuxyRX0Tscwz
1NyKtYjNAj/KUFXsDUb6VhBLuxx9QzF0ig+51XCwKm/MbFGCKZaa9ajhabLowG/k
RXoOyn3g1MBSNzhtBnM7b5nQRFTkK0LBHYt5cxwB2EVQ47PdOH6bQ+yhQb0nMOxz
SuknNKu2vCsvR4mlxyNQT7YfnK3cIgLhDLNxkl6Z0Saiy7oe/T6dXVrTAZtUac/e
/+oshAur1TU/R/aWAxfEwrQMyf99ldxelypefHVs0Ns4m+02dZUpivx+bheuvKJ4
SoPp0VeR4BT0lUNQRuXRKvTG/I//34wy4lpJp4tXeyTtXeTtcOdHK0JZ+8S7KJ9G
9scnTMnhpGFicjG/VUwQvGAQllGWDLCKMMV3ic7oAVXS70/eHgTq+Ir7LaOUGLm5
aqqJxhbx3smi0Xt2Jer9yanQCdKJWJ5IfKUv8praOdXrpV7y+rHS42jankJuzMdN
Q7pv30oKSvpNuRvj20aEphhitBgtI7+83pTyiYh7yuQccKggHhVOqvVrUWwlJe5h
v0nIKb6HLP8bVnlWlQ0r5TQO34vBp4MQHPlP7IKHOfhO7MsVzYJ2eJwG1D6zi+TP
nRegHI76dytPuBx6GT9rgB8eEPsMwxzh5x/WCqejF2Q+dLktT95Rp3vK6Aym3azr
Z38SaC/TGvnZVN/UH1uBMGFxAEwrU+6GDsxXYnx6gVQ8P3A8A8KnBakt20C6552F
iMQbp2QttarR8UNpLD9QoXYQ30F5LtBMtkYC13/Ih3n/dMdW2E7X2TRxNaJdtqaU
LVpwdNpuWJvk2faPJZ/qC90jbMU408g+SE6CsDTlUVF8UJiGeQa4glo8scCMU8is
twG9jgoG4lwZPHHLCNuOcHG4+mPKWa3Z1xwkQHdZ3Feo1YZtAmdoca00LTGGYEmM
SEl3vLg5J+F8aTf/LH5PcUhIkrf1YLIscqS6lqVDB0CxvyAMlbsUsamKrgd+q6Jl
sO5W31C398sA/ZCo/FyFaFHrPaMdE/qe+htJUYk75F2nH4ZH6tq22Ob21OdBHbsm
5A65vf+L22GemJqWHiXUiYfVP9RAk3hROSsp7zrND1ZpRmvCIKFy7dFDp5pCPmtX
QvBzNHwfsiPAWymam03bytph92VYv8tcP6EX4eqYZWNqTgy5/Q3ACZ+EAe/7nHuH
heo4RWZ3ZUKRJPx6/zjnYCufAz7MGGcyg8YWm7l1gSwEhU3m+MSsDgs8gb2SQDQI
QrjEdn3C0Sf+twXoTKGcfZxq5MMoDHLOK5DOiB4ZiwJa2xKNBg0xITTnp1QND94V
8Mkgf6Fb7vKNjmGO3ICrLxRsXOZdFIbsHmu6kVng58qR3iM7tM7gLZZ3e9MnlMT2
TPuHWpFU/19NxrYX/W6o9zbsIgIKlyECuyAbf6OJPaTUvzRrEEYAH6WKzVsvtw+r
UY6C60yU5hwE+vEUav+rb1lmwXP3C3Z3UStBMBavpKX6ZZYXV0w4Ocb8jhdDA/CQ
gQrKWx8dsVOnwIraeI11ww+YDxeyVQEuKT63VN0r1GbgNWXhKC6Q7S8EyMpSDHN8
ZRnqwlSnvKV/0mRFFiVkO7NpZrkbkACT5KcjP1hwGKuRGh8KaFCFGqq32gT3i2p1
QSbvs3RYqjr9RITbm/Dcr4Caui4Mom6zgZ/h+M1CuRZEAdftktWq5YQ/Gt+fSmXp
xvXYSyIlNLjuyoH3DK1mMRYu1N2vIH8mpVbSycEtAtMxHDxvjjpytUbTO0j2FtKh
f9BRYqWBIejJNnZGlKadzqhoSC9KqYXXYHY2qEjNlEVUkWkd+UOm/Ra4QPn5e6nx
hnt1FqnBHu5WXSpQxv0tIAiVjxZqCy1GQooOIyTW1Y8IyLUkzwpSVXOp3F61YKJd
fWhEL5Vbu99numQ8+h6IOL7vt4hp9uUiqi/CAQ582yNdPZsKGaDQBAwI5drDfnBy
8McVcPQg7jVwdgmRPz/kGbBLo//ehfCdGE5Vx3cqr4yJdll4GDC5DKcLCOzVRJ1a
MtQd0S9iLF5WJJ150rCvPbks/tnS4ER8euV8wp7lf/w+lt+GQ01CgI3Q4csDSENl
KQAARQ5SUPojz8/hObwyb+7ViuPQuF7fucBLIA/Uldeljog5RMneIGc2GMVuO420
gnk7raAqvVA33ztk0fF3+BCHAb6mnm0mjnGBtM8myKvBbsIBJwg4fIh32tBdsT5M
KACOEdg7QguXHNEJJ1DqWsf/UgI33ID+COsDye8o8E2mPgXQGOoYWJiGVZ+rNHZb
L/i2tkhytk7ttqfJUuQQ5lgvsW0s6tnxYfySZemnG44JvEdQnM2vQbRUPz7lXbj0
MunvfnpGHnibqSdqWRtRJY308mIJL7+KsVhfzfMUn0NewwZvTIuV/sa0DYmbJLnx
0R7PbbalH4Hj9rhD3qYOOfSmDdG4zlUTXDwGYqbEWcKiWNNnXoLW1L/VquYrniNG
gvQS08uvKCCTQ9/PJOCgv8Ug9mnHp3BkMmKICHVxjr6quq3h6RYtJqvJFBOYWgHy
doBDTY/sFaH4f2mI9zd4MrJAiSz5jDXFmr57xi+F4AlJj9iTjiTHjuCaBtabfDPv
h+stpzxctqUVs5hYmDcu+UcjBpbk7Zx7n5OM4j3MahUBL9aQrQPDkbQFvYEfY5ue
N4w4+MYhloP+v3Q4SFSh5TjgUjgt9aT8xrIrk3R3LhMt9/2E/86G08JW8pggD/CF
3nJnPJBApyn0dOaDQwgzSB3q82jdo+lPTEVdSNrIybaoEZLX4LldZOi9QXMygbDw
Crl1WKUfSjfqrWb03J5X4crijks3izTW6QMDZM0cc4fv5i9tlGauE+DTDrt9tELI
R8dt8RbLrjHBb5qPmHbxmWwvbIvmRoFcZn7Sde3p9oxO7WFukQuJSVDlItlMHBZC
7yVdUrLbiBDjECScRpJs/SLv4TInhObkKLUOuekm/eUSp+Nj1k8YvDkeCukB+LxX
o/103cOIcw5sCPFgecSkSw0zOBLvrvK8cYapcOUKfB1lgwiFjHrl/BrDsqmyf2pK
CRtN6tk7LYrYR7MzPfv7AFGjHiPnNMUSia+LDvS67Gcn7g+RWfLZ2jQ43I6Q6EWt
kPu9WHYFzGhdiSsbphMZIwr95ZrunUYMzhnJlT9W7oe2yAuIuWo5xEO8tPR94fiD
UJT/jptLhRAolbqe4FO3ZnrYAotSy2grbMHnFfYV7tWdB/yAvB2r9/z1Au3BrcD6
EYj8mnhTGkUvt7B49NahNHaWpnmvDsDgzlhB63sNmgciWhGyyhp9JRHulOIo9wmK
kVvS4k92NjJO3jfOf4JquH4a/ynD7pvPbTFpOkz4Ul2ApE03OkIiXSopVAwwkEb1
p/4IjkxrNmO3Eq1sFIbt3+7DLA1IMqVdIYtZ9r7iQzIexrpMyawUdzYSrBOfQcsI
86vbEC7+Z5vwDgDEjSe1W/fpisIUgqNlGaRn+vzSvlewCo1Y1b28pRF9mQkB1okc
nTjQ+sVqS+f6QdCbBK+zbjvg8i6i/BTjlpkyaVfZjElmBGIZOAxFrGSHXvoFgWZ8
3V0H8SauFlcDHSPPRFAtYtXLyYwFRS8AWhZ2tln6hkkmV35nUtVHQdbq6sujqTdL
Z/Hjhtvb//yw7Dyz1fkR33EgxHu4/G+SMpWDpbI5J7EuSsmi5tO67dNCopGoqyWd
xXZez5QCI2dNayPz80E84hMOv48MxYnvefTvodcoKH6cUTLVTIknfm8nBFwbu+LL
pC/jP2hYkWhSA28EUL/5sg/1IRAJVZRrKKQO12MGZJbijoJyyUkfJV+Alb32kaCO
KezHadgEMVjNx/ZsrlL/iLgIXK8uTZjyh1y5IADGcOsvdX7TQUB+54z7JJiSfmaI
TpzbXaCifVZESv//3mKg5ewCyk1A1n8bi1U4XOnlAGkQlcWq6M3nZjEHTYhime1G
+dchUezJKCEQGAk6WI4CbeBmgCr4xkewCRf0ysJr0eEGhc31lKx2Z6bW9HQpwcen
mVA7GGVI2YhPHkDJEp82rRIg7jrVZv2QcJuZg6fqjyUd3GiIM6eRoTpWxe04ndTg
orOItr7Nj3QIiPBe+h8Ewid1zuAWm/TYQwPP+pPbg5PElmGTl2JNuZ5Uz4JAOhzZ
rUTGxZlKNkLwOY3gJhTerP+w3smbBcm+XwNKhz49Mezo5+9CbeQVMNk0BzevONMW
xvawVlBeIxcLpCDBlmOEzI9ntyoae6ktlGvM/yA4deDl0cQ6dv81PknIU3PJjVXd
GRSVz4tNUJNHpBdUWmvYIT/hmJT915kLzNA/CU+xcmQWWXCp6gmiCP3t/ZcqnUdb
TaJjjV6xAmcjRFlGfPJAWTAr4Vy36hFcJ0DHFEFEfSQnh2kd4wDva2NDEJgJn1bw
CYutUOEZyVpnI0eUe9epVvcU0vGl2tr6oE3cx5ZoCPxOqSyPPfun875BvDT2PUQe
LOWXbzStOTrtY98Mq3swwauEw/Y2ozr09fq0EcxZywZF9mQaFOOBf0snGoxVG4LW
p2wISGgn4GUk2bDESiYihxMLh5iyO2WAXUCZ9J0eJJplrDVd4b4nApkYgXcNsCsh
qRtmhytB+e2jAlj5oU4Rq3ZPCjLSEvbPOek0kipyDMZ70R93jXZu0at9aHDSAebE
vXNeGYfGz9wRt/vFeftGZ8Vi8jMZh6djU2VEofBOuxGndmdUpUvSCrkjDqwnkqg1
FoD9MX9yI6PBx5oCcWAVtuW/cMRn1Usx1XT+DKA75kNVaVXXGZuL6j+ZnFHY+Rjn
cDQqfrknKFtZ5jdwuVQ4+v8y2gPE4FwyAPFk9qhhlCN28E//DCc8cZ02lBAZ3Ivf
VKcb2MK5+gw3w5gSETjkG+dgZLEjq4xfJg9Cm8r4tELsNwk8xnzuUx2G5+zJdUdZ
69L+MTP9U+cwp6grWy1ApNRKO2o9XseIySx64WQzgePlr2tS7NG92MckRPVo8x1b
teMtCTh3VeZoPxBJiiQIFIT/rQnchs4iCy8VuvoyRZ1hEAIJ1TAI+XMH61j/jp+n
iY5BOs/qJvKhJbuxNti3+U44n9jMRNmehTGdI9dXeD8+HjIEPJaZ/3s+TVdIFStH
DTP8TyCxkiSppWr6li+XNbDTK3Uli3/gUbjJ7LSMNTg19ZTCDVeesb2ScKwEUK9k
r33VmbGmEQK9+69eYu136lRhkDq8uvmGKM3voEVPOExBIDw9THzJ49P1e2e398WO
2/P4yUM+nhDeYocl8T483uPVATMaEUskfxPTyS5FXFYFmKU3tk/Bdznp+EI3ygLZ
AbjRKEqZ3Xu7JDMHeGvNsas/vEPkUL1Stftd2w+GDcFyhygqRVIe4ZqGTkTiYLit
MmQWXoTQwkeOh0luaSrXk9SqtkYhDVgK6UhKd//KPmrIrNlvEDtfMeHc+env1SBK
c7QczrRAU1MHCaBiiJ+/3qFmnGibVuq1MLtZ7+caNdahh8yCus4vYB7LZzbAMJWp
5CY2y00sKhI9A0k0IIYdbQS9xh12nTl+Q2xXPKl91zLt+kJ+S8W3f0GTS+K2FEyT
Ademy+uZXNkiMq2YOM3Ac3aR7yNNDZZJipXMyU3O4Oidy4Fn7vbSGH7UtJBUZTNn
ceuKPqXp68pW9lFQuY7d3reiiTU59OtSygQyc6wnUp9zoO11IDHfABOvyAuuHX7f
BhXu/v6l6eb/9Ewf1WMJnruQKf+z2Jjcre53nstUuLod1JMMhXZhZzgsa8xuo8J2
UC4pwszVlZNu/pplNRYE3H2gzbQPl5dHdEkselowkUD0k0rUSGYIiBOTCTmKZbLA
SMH+TFLLvD4PhbVvPkGtcLqBDmbXwqSCB4o2o/8AERvY+RRDdYNkTnyGCP4w0NJX
0mJYjg+hiN+A2LdojaPyzn9Z7m/1gE4AkMHXfsQpo3YOLeqQkHjXtM7JBKWsZrCU
o+zFruhJQZxs4EvVYATWrlWj2YJt7SNx0kOkv5V32fxcqwQYdCg/2/ATRM7kBm7c
5sKJj+K557lL0K2Oxk8SITISucAZP8lSJDkwDDDPf64y8a+eP0SZodrD5dtMEJOq
tE63+YbS75plOkMNtg+GkWK2MHTR7qGl2yExdcomEMKGbGstXFXW3exUGj2aC1Il
KvQYO1YCxacGdW2qyDXHW9SX+E6mMB6Zv7WtKTLXpUn7VBeCXokFQiSsyJWwyYuO
N0PE0QNPDulMrZCtaCGVVLp3FBBmCmvj6n+CJtl816z92r9AAEWoFgMXdDQjIa68
JI93jKvJh6NUQJImeVevz++wqOo7tXvAX4HNs1P9et+XmWgHYMhhsiqoXM3FScQb
hfcdGZl9Iber2T0DIE8tnzN/biE2ZVRG4IYXyMYXr0EU+2qQkN2dCn0v37IhsFzN
L8AJ1WVE1ID0QTBDN6rDI7gplHAzb+GdNOxsFLtqRmpVBBVBPo83KHdUC2yGLi1J
lESTSCdyc6L+I/2LmP/ZuEgCsZmla24Z7Xf0iCe7WAzQmSMbAiKWBCnL1zgIr2+D
YYIVg4l63rfhPFDeK2RyicEjVP3D7ijiUDomzpzMZ5KBxgd1Mx2Uyt6oAcFQiQyD
9LHnsS4+QM1aDVNap2pCEqRVP1YWa/6G2L58n0ctLljoDxfUOIOjqaVu3ACaXs/L
OuyGq+ZOetA9X3HQpFokC4L1CdDUT8SYbTV2Ie7KZyWkWjsT02+u+4zz28JXTSny
0nj+x/UcTiFHTYl+cwlL23AbEqo7sRvSA6hRIC9IEevlWX1zB+F55SlUCJZnWn3B
7DsZZ9jMA658QSCJoF8hPu+kQZRrVN9SM0MSEU0S51fVUbrc48faDQNfmVPdRdYU
NKUnFz/8cNGc9LjTWIsmhg1IUn54kYq730Rt8Qx4fRgGD1MALIF3HWfbuCoo39aU
hRxeRlgQe8xkb5K8P6XyiQuAFLUDkGwu0s+98xPrv2hbVSzbcq8FDqahgCv9usvk
kygxeiMqL23H/NJd6T2EIsAAdU9hPjddcqAoCaNAcEoRHMW4FDk2Cg3QQFeI50sN
1QBCuvP8bIKHjjH1KCWq60pPUK1lXtPPek3HHHpuOSnsOb7E+3al27YpZvvbM32x
YYQpr/cnLOVUTzBFD9LKsbIW5tSoBVkIyl+VSR6VKiPfIrYuhkZL2muCARTyTC5p
R9D+aMG0VDLqEejewtikBcH/J8tPcLRT4ppZIfA+VXLEoaXDZgqKwU3uo8VoQEd8
0NUP1b699WkE8VIGoxNRRsPfDA6noIzB3CJHS/uY+7RmQyTq3fmnnlhUqSgFfhBa
n3LGQ2Tjjz47N5uNYHYL4frSs8BbmpJdO0Syu/Kn8j48TZhMibThqi5MEJQuE1cX
OoTLGxo1WXgen8mA46GoLRHZidKXm0uZfY5OHCRyiLRGpyqrxMM7K8fePwjW/f68
smLdhlxmWSP6pWH6BXK2S6svQp5TI61DnhQQng9AZtms7SV6C3DV0G/SzTI8kyuC
ukXGW0Hphs4vL/s/bEmKF+EOqHwsn+A1+635lZx9hP5DyO9U9xq5q2TfI6eruoC3
XgOygzTv3MZBr7e5fkhvCdIVi3mVd3iuj0t/ofkyMUsakGRf3J/fmQkfmHKySW02
TG90/M60inqnQ8A8MQVzwIpb8FwKOUODCRKkumPHfpNGFap49EXE/NdSQZUALRFa
mBH0pCypnI0lioDtMuIkU14LEzEqFoLBNxsA7gftPXY7z2EKFg+z2mqbNUYGVV7x
sT5AiSe8yyAXbyxO132YMOsY5WwaWccHNiUMcGbxz8DUmZ88+tu+LVxyH8OK7mwl
/m24GPXb3MZgW7ICFG+du/LlItKXNNx9DbCjxgeSRsQrP74r5XqGChZx3uMdh3mQ
IVrYYnRxReKMEICAKlQe+p9/bhvPRh0te2Mw0B/wtNxzbiwEWCK9kbKMpChQVb8r
4V72FpQC7S6lgiBUaVyp8MVxXhwh+WHpLsZgWTlYPfoBfpnonY/xgwhmQW8v98Mg
ruIuRJIRlXUhbNxTy3uTthFfew883hjnJeKPOCyi5UGT98RwiPVWG+Q4dhUM5jGC
yAP6/c0rZ1wo2OJSZD48t7tlemvykykKOWQ6THCSOf1Iuq0AAjzeA3RAat0r1FBb
iA7udb3pBBirG2jivmxr5TNov9EzFkvdn1p3GjtCkhgyx6rnsJHlhDS9ZKYegPvA
/rEi6iz616DvJHPbP24Iyv8HGgA77YqKzL5I88cR9lVKPo1mWJf3d6GyWN+t8ch9
cUVkHRYEgh7kyduL8bqeZ8r1F5Tl160NEz/0CWLZ43cNvCMXl5SRgFxOT7B+SNLL
WonSvTPSElVODEzDp7cHFgc76/o7xeXlmUB0C5ne8Kr8zg1EMSqXfvA00lZ0y3ox
Uvpfdeo741eSm/BBnDUx40NlT9MzpQO3YiyFlm74tqtpjl+AeOmxkmfZcctghSQN
4Wu6tURq77tSIjb0UGxW/xhrNdjnrXYXMG1s0LaQJQmw6ftGGS7CUEI9WV2YpBWu
oKgPoqaT9xnYNkc2hs7WQUlsXXlpvl/St2xx0xmt8/AeV/PDl+BV4dz/hqq3nZEE
v/+oMOcdRjObppv7YlZREG0nE8WXU9TvAMzhi3ye4JGFrsydh0ootPhlEmMnmlQV
SocWE6l4fVCDA9zuOwX+jKNJcmPIcjtei6rX6aQ/oeBNJsZd/mqT5EnmsSDZ0/VI
IBptKnaVgT5gmDwlvS1tvfZ3Gjwe72Nkc2zcIqrpBxwJhXEiQJoUaqDkGlfpEnAz
YQhWYUI1TmowrEu7xdZJWIP0UBErLIkvow2wDNjbQCYIC0vQrsHkxGtUnaqSIse3
8DD6pOFI/S5mWfJUVT7ukI7EcJRnkXIpuHqTQC0+/UaKikj/yTgPxU96f056tqlw
nNw1MimJT3USJNQXjPLquR0rt3uX2kEoNvT1JEjfUy7obfYQ09zuTXJWSInSqLVt
EiErRcJch74/PUF0IepjeUO47Bm6koE/lu98I9tqbRQHawL2ehsKsPCb+sthb5fG
wSzOfKLUYMDJzplorIcAVHMNh03plKWqUC+OQq9HE/G11dp6GShscGh/we7Uij4a
Swrz54grz5RvbNP3evGrRDLYct1jWXtrx1D2lu6InBdWZxF+xe+LP3T9AWaprkVR
OQq8kuTIDK7AtnrcPWxySnSId/dhquoDp4WM67FLo7/yk/5B70vKovy/2hDcw58t
/MEl8dRn6qt2MKN5ZssFraDDRXW03Xs6fCPM0ytP4SEUaY2QoEjiASFHZOty/Cpm
T17q98HrIItiizfe9Vq0D62b+r78SLO1Pdk82bzo6CGKFg0X3pFI6qYinXv52G2f
Fqf62WPrrTGkj2bd0PTa3eBITIONBteXfcZxFPcfk0h4I1tkjHzPOBYRxgYboXS7
DPhZx4eaf0xWlTaQLM6wvrHiAUajjNTPWJmH6YYXxV8B48fJ9NkN3ecVGfq9qRn4
iqrjPvXvNWl4/1qKi0WIdZ0UHxm2HHxY/50qGHltd7B5ryjGH8F66Wj6ZELZ3KBG
wagDQbfPH0ebqq8KnVhZKtNMkFeM26kgmCU0g7/aZkJoQr34Xj7Y8rJWNBuvE1YV
oI+tq4LcyfipsqGMPH7/Ph6NImgPLMcBLHSA8ItXGDLyFKbkNV65wzY2AZdLcUym
UQEsAAucCB9w98ig8dacpO0A2FDM6wWA+6i2egSGpKt7ZvemhO0eq+Zqc4nQxWn4
89XvLADPZKX5ZCJ/LOTNl7shmg1f3ZfZBzwpkICRCUK1YlLKaoGCguUWyMh48RCJ
6NKerJo5TQxlhP09g+Uxx/FxbSHYUzoom1VS2b1LXkjdTiGwtt4+ccEZZ1B39Zh9
t12BE/o9iJ+vDW4HanLYd6LP8VNyiRov+N6lckOLnwITlrfl6XRGlJzvOmlKJdNo
aZqt+uRHdD4RONZo7zpk8V8abm+dKyGqTx9YjwCpV5U6NgpAL56mBCJCoBWxTBfG
cm8HjoiFX/dt488SJep6jMJkpb4zww1bWxCx2GazFPkDPQ8l1IOXGkyO2bm30VF+
ZhUDmafjMkKgtQw+m3mg2c3kY37HTOMGT0F0+3ZmCuhNdNgefVHEnu/1Z3bcOfh5
Zw5TW3EI3QSpNSOFop8rNkrW9efyv+lHx8B8I5bmetyzlRhNAljwk5XxJP+Rgd9H
5B+gn0Hv1XJnt8mLPO9OJzmWdqiCLY+Sc9kgZSBeVowIcGE71fCihA28BLP/IXoS
uJXbqQbbJ2Zgjh33imi7TilHmzaMN92h7mfgnkt02dc5YKvUWwZWqyGiGYLy/oZk
O9PFLoiycG34IEb7vU6R+OiZEmQ/j89T3zZyt4ZZ1S2ZQyRE6LYkmOMpp6sI6BAX
a2ZBq0MwZ0hi6QCGGAWMvZIBQvvbnUOD4hsR452b+erNf1PP5i/xSCIA6QSGKOtD
0lCxWl04EPalH+PBDt2aBOn/Qy5c4Rv8rXbrwL2GtAHZMWw/TGW/QWjQ9bBwvCNu
rgn5OoBjfLd4eeT6NdD06noe2P7nozayRpcwbFDrn5lEq2d/CtVtqs+VAe5/l09V
z5+3PR+mgEM6pPfKeqwdzV6f89i0aWfRKGo7vNmIqBz02fU+ZIiJNuDe5RD1TPbX
iPAJTxCNsUwio3Vj04JCyLvOEF2llObPFoUNYFtT6mj3yYRO+nT02FjbgtowJsa9
aJfzeEp2yy58tgObOOE+sK3IRAbjhgAFyWHxuWgvLYxlL0qwjiK4tNYz7tuPB0zJ
xA7+7OKGdNFwQ8oU+iJQyRbIdv64hMCLcSQehQP7gHKjVC5IDpAyirg9+TKh0KYF
VCPPUivXI++VB3xkERwQ+5qDSiMM5x1gytR8p73OcdmWYI2kW5ScYdHwxSV/ncdS
gNqTaJBVEvSV7xyTM2Jl2EIb1jW/hol2tpxENy4kHs6j4t/tKCefbGHrytvs8d5U
ah8lH3wlpi+UzTgNMF/VBvVb7+Rx2SeAK2xSQSXUq7uTpk6EpIi3nyCfB6hd/sm5
079/tpaDxPHJ0E3z1D5PYZV5sMZsN1jFedAA6ujB5RUyOQAChVjmQSrrmuEkS4yv
sHHSsHv3kqnHrGKb057uddZbjRe3gKaa/hS+lK4Yn6j9RVXCHItpU5IKjARWeFYI
JUzxE6nRtcE9hIxcKs3uAUlmqTCgG9CyYEkIieKwGx0kT5KvPrJEnsjmk9AYaoll
afm/nN6qPL2c//Jb9d74unyQtGvfXewZY6wMoj48W+TPja4v5DYGHZlkG1Muf6Tk
9uHbdvy3thZXHzEXYYwYySM1rO/RgxReZ8VIGRpA1JsQd+ItSJT3PZpgPQul1fAA
gH+YcWVdWhczpAPBCAHD54pslJe8ttaBmcrzg5ognyx25g45RRwsGSFIK8pncUUU
MKgI+7O7KYZU7WuAKGxq2X8E4rBTfzC0aGoxVxRjEK9E0LmfDxWybQYWR9GKjnlD
oOnW1JQJYUzVwGODFe6vjLhVMyOGYa7lgRe4BO/P4XbJhN9SCpLwz0ylq2oiSFx8
40htZKjLiR+AFvNmtb1HDc49Et9rfxS9A5F394vQLz+042xC+wxZMgBEETgQFTQo
MS/EzHuOJNg0nDBpmoebpCBG80KD+NrD/s2QItvjob4jAgD+OLAE+dZK8fUdwp+v
bSa/QyRuRRookSWjlq78itg1qTKs+TMfRK5999AU6SYRlJsRl74kcKYFmhT5xEV7
hoFFg90kZmdl3+dTuK/9WjiuLy3FKwsq7I9ZP2F8N0rRIa7mHDJUVJN/ZY/NoiOK
OH/i9pljI398SP5o+FYF19m3/26oHKtrmteXrCFrqVJMsmqs7VZmlL4urJ7oQ++L
u3pT77nLzXeTXSNAl7ktGoxD6m+00fs7NyfMdhRbAvof9j8cuDuvDvArtFANtM2z
U65Tt3gsH+F3SCreVMb0UwpvxH+PB37OJQq7OlYNOxAuoTGrznoy9HXKkVxDi9Mn
O1ZGLgVq2Um9EOqbDAb03erkjHxSIbiTBSR4y2LQaRc+IxFIfzI9K1tn/5yr87pE
PmI1nYNX/HXc+H4UJFcuY0TLwF+eKNkfDqKLI5ybbZut4a7MoUh/gX6syF6xS+R6
0UoWSwlUbAPzLh1sy5kfBA0+JVmQLK6G1qLQzJBrE3y+IGormwSxWdMvYub+SfAB
vS9dUIQDpeU2WHPiSqA3+NTadsFmL94WTpZmGcTwj9cvlIofSp8pGFR6du9QGWSk
DiCdO4ndyZ2eiEP4FwJi50sm5xeKUiZ4q14o6GNZ6oIWGDSlZAE7yOdNb52BH2rh
XjniElUwTVvlCp4Ss/WyXmY/ED2+Tcq2ye51AxrvUnTjXY2FXPgevr2rRdDp+zln
BxfZDB6xBfVkYfCCEU294RbShYqJcfNnhs8/M13yhZSBWCE4WaZoD8jXuxg9u21d
upxpgLDPx8V68jb+uoVLV+yqIG6tAy/sY4xAYRwWaVJRqdRC03i2I+PdLG1Y83+n
ztKD2GksvODVyasye9JcGtfByaFarekYoo/r+JcnP0WraFw6uYvVsXyGquQFK2ZU
pPfdqfX6NyBp6OAx8KmZAIzKKNKKQ/TaD5JQtKKePHdXDf/WSywhqMIcitAJVvIx
Gu2YqivN/SIWqC3h/EwjMHEPa8Z7oNeVzypCykZG30JLeZgdXKjJKLYRJK0abuRT
rbamidprgW3MGFjTp6FB+NwYvi++y2qWN4Iyc6/peBYSi7f2KdGic8qCFUXqSpeB
ug+Zqwq0TgwT4jeQWB2tIwO077Mmwqtk03EmxeP1zHL8hKbyWpakkZApDGtjB9r8
eiwWiUqpTlFdC+7hBASRL5cgXEzid35FX5+iGdPMwcXlrqAyQjhOn7FJOVu4+anm
nSP7k8WWbcMLdhAKBAsyKGMpdIQTZ50ZxbY1feqDy5DiFgw3eOqUPpdlp89MvwD7
5jnvhJeGkhpL5MOWVNPZzk0SDh0dqlaz3us8Zai2LR+1Hi8GBfqVxD+xu8Y1tDnO
T8OFdbGCw2XgUfrJFVFfMLUmSD8E70GVP0YNgFqogUU7rOpwo+ssmMSvl+reOxK2
qyNbFdOrUE2Vqcervtr+IlBxAXAEEjfXu9VSnjl7t/uQLPU9xyg2XwgK24Dbjv+T
LDHo2HD2hWYMdd4Ppwtb0+k0gzGc7cw5xcHGtXQPQpf338oVjcLEAnLq/Dkynhj/
G8GLehHgfXdhjLQRJwzbQo3dQq20auQikXEEygr+puJJ4GYeXHhIKxurVJCdLXuF
1BEaVPxSG64432hZYSnAGLHw8Slb2V3vv90BDt0ydU6xz8DjWJEcrKTFJXQzu+O4
cZY6/dYsI1SwdAy3fFj+inOOw6hHec5c2hjk+7B1HWBrMgyF8tkHY2xE39WI+4E+
8h0TY3auBgQJNlYRhRWY8OQyTikDy+4FAe/CAcxZch0iNME0TASuydipfwcKVtV6
lFa6BXNcdhjJ3na1cRr4augcfzqPfjccE75lHG4TAzSlzOfTtafpASw87gmiTxv+
pqK+a20zPqZnf8HDjqdz+0m6cBe9JgYwmZHf+1huPprFPJxmIWWN0v7WBmhDEohm
QC6U9HNwOWm3iIyzfhfXM0/59ru+v4rSAbHylLrg0w0CViNo6tRb/WHD57p7ggoX
VcGGKl80BTDtPSKfJ+9eJG38ED6SW+5BGpMONLOqi6xUqFIN6RXIxe/UJf/3sVYb
RL9S9nOsZxwd/1ESW0JfR8SC3Bt302B9qOISGWXBcukIigvlx+kV10SqMrD2jaBp
BchsheIxd54V2RUdJLE81ZfAJYoAGZgbvMgp+k2BYu2Bqe8JgMO4ZFtgAcDSwNow
sExx0+VIXxZlA6uhecq5blPAEedyNZhe1zc6pQeOejEikRBLzjl37G7SNkuCxtWC
Sg+BsEJO0HwN7yINkgIOqlgw02174/Ex+2Nd5J9kbNRgoTZgXN409Wr+fuLR8P5w
uibIteCN8sEW2un132wmfoUPFw//M1A1nhHdWAbRRa9Fc9tkyBgxTkWm7opKm+Tp
cbwGR5yeRTHa9qcufsysDbnbrWqjIxKcJO3yYcFGheC9few+e9lhjh4PJO2gflq3
VQgZUvSAea4iQzy4E4Wz5f5OFTysuJyjnfvQe6gz6eRbtsTxFExOioE9aevykvRq
9nTHmv9bw0+XbgrLJPh0U1m6+fN+/aiYe28Ilhluw+YCesmJlDZRS5AtqbFJdZr0
Ak7Y2xPKJ7GzT21+tXYt0PhV2XwVpWsFLu0uHmYnWag+dMdHKCWub3CVYSD1DOjw
esNGeHBF4c6XZ2C1XUPewIGo1y4vuIcer12Onybrpnxc8xzd0hd8sJaPFHJV6Sfo
wcjiL7PdLMqpcXa94EDcZXgDPe/oYuOKLon1iRzjyy0oV+KPO/Qv8sPE+8BBeabL
NhJVrpcQEZ5xHKyW5t0LyW8ea+/2BVG181F6/W1aWgvR7tqWKnroM/An52W1MwVg
Au9qoP5XbOBw/+tpxH+WfbHFECPr+YFiktkAeKo2ylVoXAwdwzo/1YS1ZW045jgh
ccwnSqbknlPLH8jEDIaMTwF5Q91lepUpBjo1GqdbTvqHdd3rjm+Wr0eU3qPIAqDt
Cq3Footsh7498m/5nOUSx4+ihAmIas15HzCUbi56dWyoLm+B4kMuf+jyEuwWh7op
CS/976JjDlDoN58GfaAMVTM6QWOlnv9N8fusvCcRjbL4NDXGpZUN3Bk25YjFfr42
/vBj8GUHM/pE/wvMXhY1JRedW1qC7d0rlx/QQeDp+QEQp0W5G/1Y6HKGrMdgMXp6
YfO/Q/8mirxHRZ8uDGilXy18I55yepzoMMjqSmAwlgRCfeM/KJirphT+bafPKXaP
1JceQmPhEuTvCKh2qG5sCbrmC3Eul/vq5KQOljqqEiVlZPz4wPtzVlObuxhskCrk
jBJRMVEurbmWzvHXenECxYnti0a3DDLxcoTGx60Iof5i9pKc6AGXrsKw4hZFZb4h
6uM8R0jrdqQpyhPHsEbyElW5X6P3KHoIFKZ1AmwQlzjGNUT+lTvyQJ1t57Mq2kYj
TgRULxc5+fR1noMxi6cbiBBQJlkZddA1rbTCk/ReXH5Y4TNouztsquHEBETUNN7U
VmAXmZ6SWywkDbtSNSSBOKvuJDWP4x5vFTpbow7f4dNYpyLEBDwXy1WOxsLpy/zl
MvDiC/MGIZX8BOc8uhhHibOMgrDcP7UWtlA466lJKUiy5hU86NgKhh64YIqeGzUE
oUr3T0o9MD1ZQSY+pzqhwKSRZGmy3RBrlJpEAvSNQ1vsA9toXvjb3yg6kEOzEMN/
QeLpJet0qEcr1yXh3WJNCkAUtUeQ0wunHmyMHREGYh4M1rSTji0asFMGZsWiGfuw
S8eO1r3a4MsRnQazaE3M5lEqnBp8exhlS0TjDVmf2bCUiwW+Yhb0Wl7OdjWxA3t2
U+xIvqWVsJ23k32yN9X1Ak5Njq9Cj1DCOorInXnFj7RYhLeNGX0VlaF/6MZ9m4il
o3NV7gmnSwUcc8jDD3MfVfr9PwXR8LgVCtItxdWd9epccbvUQkmHFXu6kDYogRGo
NiqYKlX9EOk1y/hL+o2x4yIEtAqrE7Pc0VKtvsMGD3GDcB/DjXgjZ2RUiv7HPOiH
lmSD2Y76UBjb9nf59nab1NJmAFMeYoK0ULcUZl9DlmEtlBotm//DHaMcPL4ynXpG
iB3A0uEe6cOMBHkuKIcWFkep02oGETzYSt3eFpi4t8cIzpDNSV+MKbl5aUvxcQCQ
JFyS+i1N4rVe1vf5lmL2ZQNB3JT6LDPoiTPBUOcp+Qmoel9HuEAWCEosOV4XlFpg
ZAwL4TUXn2VNmyxTASIIhopZ7RFi/CyoE7ajutQX1bF5Y0DbbV91Xw5YBydCdneo
Xbwaidqn4p6Ka193g0+ZjTO+rZaAlegiOMbRJnR8PUWxjOjVXL4cRH+wiXpI3Jou
MIL72LgWTsdtOZXrE2J/DxT8Nvk89QwmohqVxaE96YD2vQaz1+CswMUIxBIjsb36
HquklrDtF1qS/hNdTOdPg62qr6rayHo3wBUPPNyZ5pkxnmWG2a92id/W/sVFvE66
KONWKAEfkVkCqJMJCXaJgWYfeI8DB1N8COoQowXiihtfYWPYgTe1gIi8BZroSnct
1kPUbLA4RhOSX2AIFUM6xV6G/Z/1VdrhpM7hW6u5BBc7mxq24rtT0LlMkbHHf4SB
h+9LNv9swobOsBgLGAN/sowexvgSxNiAgIXgKjYNqX21v/kAKqMTNLJ02KuQDMto
hucR8AIo6mZtas0exwMOMKC8H/ZGRcBR125LqWBZEMSEzBIqC6tNLPP6Vc7pAzmQ
Uc1ZmaxqVYiTiCV0oKes70Qx1Jg/blev5A4xNWTZ157llbJTCTbtxUXDoL+Hyn8M
XGk2nGhdfA6xFqAf7YNdK2fU180XdhN+KliWuQzEnSFgBhqRxEOQeZYvCQLV9TDe
K87Ozh1O1VWYyjUH/m4xxWiEazsvg3OW8cbSsbJkGuGrZ9jQW3tMgBk3g6IoUTqJ
Earj3bhwFtQarB2jyG/vBCE0HBIll6jSH6i7ttJxxnajr/leFsDjxCuzMXvnngta
ENR2LWqTYI0FSrdvAdKaN9Gs5rn0s9PG5aIA3f6O5IRgA54ceAFlbrQ8HyM0y2go
kC7PfhuXNSs0DqxsBsteIK9i9FlEjSDePztZp0K8+2vzhnIMCeejRViV48MlKQ3K
DsYzW728l6NXVcKkfbvshRaaHMy7VB//goKwU5R9LEfWbcGH0Sym5I8DoysXj1uB
Chk5q8HHSUkDN1m45WSmBpBFaSKphoh72GVBycAAqIozpEYg2BeEOXAWqrcGbBzb
hSBdIxNUXrJuTBaiOromaTv5jEAjnJ3QaLhhYkUT6LkpeK4KavLLMeSaXDu+1KAl
we75MH2clu1jRhM6AggsFi4YsX5+sWE14UZjZVPBi4w4qt+/8YlbqeRn9sRDJjzF
Tx/iv/Wfyu9h1QCzR3VraU3ySWBlOHohsWy/erG1yY8i02zPruGxZCMJN1paY/UM
UlGcy9fSRt5ND0AFZdzXjOjW11uTLisGErfT1koyQVwgsIi2xOyW6/EBwm4OCKRw
O7sJeSUPh7K6LJTXgsFdHCr/oWk1uVAGQnUa3g7sofhwcOtYxxBdIruSJODxCOrl
QzkTGnwPjzMhBULQnRWwXFJAUu4s55LVZSi4raj3D48kKRARKpTIyS6fBqlnJTgZ
FUjWRJLTNQhTKevVxEGKQe5waa9YF3olVRW4jCuKWK/kXUG8koEv4/cFC6TrZfa2
Pvb6lFAIpc6Mrt4R2XR35xWLbZ2iBIGxjEZVeja6KF1kldTjZQL1md67/vnEf965
zv9ypdDgVNkHMy+b2FYaC9++OKZ92OCjNqUQGVw3ooTpN1L8Wp2fft6rDIvMrh4y
l3RBw5wnXMyEjyL3v4q56bOLDOvQ9mxpIve3KPF+XlWooimgtzQJ9S1MOQVFJLOB
nPsGzymFIlnOntEXqwGVq6hC315q9IBVaE34bfYbNisTWVRS3nst8LXKdrjscV9Z
u+2P4OclvSznYQWgr8iaBvyA73JMz0ahNzWOTdBBDZ5CsJNj+l407KPReuZVMCRy
8PDiu0ShW/OePoqvkseEkCGnvWbdZNhlnX5IaUXI6Ze3F3q3zypqX6D3VemI5S9G
c9pX29jkcUdeO6OYxgjBlsxE+kciIzlIlfPnw+52drSJphbPuynwBhopi3UrBDcv
cpipB0mROTBIKLWRDV9ZjdqgKXH3f8xtv9sQxzMo/KYNjxJcgZ8ifw7xjv0nrzHS
/wnapLPEtwImIKFRbsrfc6TBXwycel8TquEqLSZlrKSrVWmL6xKS6pHOQMq87JZN
FVHLf7a9ZDXXlsShjfziJlcUKU+cp48/K5y/JonEE0G/+sKHxVWr2wJCIdwdI81R
1hwXMJjnPjNKhAhLrxW75qjJ78UQMsauPGdPQVn3NO0NP/tKsl49ELgjb2Oe01+A
Upci3CVc5YgoBqBJeMKWjXtwpCZtkDAsKZj5muSg3gCwLFE/qo13+xBa/vQAPsB1
VhW00IkEW4Bjc6yZ9V7SPY83kHBI8N7JvMOOJYUTofuy+k1sQYq8wrG4oW99bl+2
1dkC7KSr7BNpDm4X2vS7u68P9BRh1N3+XaDO/Hte+gJJFtUkoH1aSHHOMlP80Nyo
0FcQy8EI7BprzG7D47H7wOnRhz0lxWcC50+ef9OG2X1YczHRDo2KUcXy8O+UU0dc
8cWgNdr4WAEujQXDftZHJL1xNfjrwKCW7PD9JT8uO3h86nESS7qhk+vl1MCmDICv
5K1PFgLKIqDcBiUmE+bpq7RgqPOGU+KOnXFB0aAc2d+h5dgkB/0cyOK3fwEgWqZd
Ix/p2zmKsFcIxn2jhmSHqY8XAkFCLjWjSMRnr2NGFR4AOfW5kGNxoPMEv6bjrDSD
OWulQDSbnofzUz6I4hkQeS/cCYerK4lug8BmWIlI7W7wSsJFOIrW9Li5c6nK8Qo3
YlIJ3gkqKqFW4ETlw2bdUhRdWxtyoF91c8JWCnXta3zNwLLD/8pCEQPA/0W2USfa
Yklm9C0YoS2BMO7E6q5xsnV1SjZ3oqHdYw5Kf3fSQfGqnKArY8xaiBlReS3AgJKW
qy9WWCOJPU4B89XyrJjMYRYW4agwqp7mqLqfTSbVXjABqOWzvBd76hVakQAPnJ/j
AMAMoYgwmxEViGURlBR5kETWJFZ09OXUxAlraGvKaaSnKIQ+k7eTts4kfgVMbuI5
HNXMF6AuE+if8zWeradCxd68T3yjjQ8w/KvbfmvFPS4Sx7ojooGpdntAjY6WZZZI
+8dEG/n6tAy52TYmQPJc0zrMxiImaV8kRqEZxTVme3mVySX6Qfe0/8vDfhXGuvKi
rsvusWZsfHUo5KZ+lV1Z7MGZAbOYu2R3r4tNyWns7mMNCIJ/nQZX/OflZy7VQRgV
Jpnh8GxF6c+1pjF4VnlZcPbC4bW/3mW1F4XmWa990axsIBSnEipRBzSu0GMIRPzo
0h9sSyNY4GiUJBnmYuP6n3X1P9tvTjx2x94n41RPiTZPvw/beSSzYFxnjjRBjz6e
9raF+M5vSm3fEQiMX1+MNT1pW/TBHLSz70Q32E8lI2FFAuRE9JaeWuVk5HjMkEvB
Wz2WxaDz4EdVXLItzCRIfO9X6B+Ub2CdFteivGYL9fQ0/fp7bc6DpllDn9nnu0No
2kLA4wDSUozcSiizw7ML64o7Vg1rllivqsrOOx7PlS5aw6zVXn4HiqU/WSEtYEf4
JUqtop6jUaSZSq+PJExMSbxCBzEeQ2ScJGM495fCJrRMvcH/h1i4WjBxTH9/5baw
Nr4VbIuAbVp+2CK+cxpya7WK2VP3lHJBRPEWh1qNcUzKh2XfnQjBGb5V+lax/hUH
ua6Vn8ipivfSf5soTnZIRcw6u9wjzN8tvPTGb8MX1DmBngX8WNq6/lmULnwA2Eau
aR+6Do6T1PxDs0q/LHSzt1nBbWcMn4FHoJ6S3Mxcc5FTV0t81yBVSfZ4z1bOqF7N
dnQRsyOSUb+falK+DB+h+UgaIE6CZukzgtcPYQU8ojsfdkR8/j2F6TEpFd6aCeYF
TwG56JiXh0AeFjnjsDR2drVtBNpCsAAR7HEoYA4CNmdomfOPXtViBp9vv6jNGKrj
H/kQfzpCSt7padyKsXxja4inUAEylMne3CdSEwaujulQ4K+g4SQkwezBe//8/t1I
r74XOuN6KUMcT0KRkTgD7Oa+9NoYvZVMRBt05Q6tVTsQcStc9xwgEcojlnN/7IR3
HSA1LW4LKWMTyzREkxIhJulWKS52nCejzhCHqudz4hvJlz1pQTU0BdokjifDXmvw
P7aBDKwMb1vhxiuZyEqkIL1mDg3EW3c7Ll+rdbylgrLw6W73oj/RX7QJt8wGsCIj
eozZU9lBDoSTafGjWq00885qFHN0aBKd9XT57gYpFcSU7a7HhXpWB7W2PEOftVxj
rpaViBOGkCBDeEGVry6xgds1NZij9+xrxb4EWHU2hxgC0yRA0ufU8ev3y3yextue
qKGBc1ZLr7tQC0mWHfUk7BBPzdz5dcuHenNO04sENeHBbrxNqjp8BgEXj5VmttjU
Ox7EhI62d3pIbmi4Gjcen5XmBdkPTlLAkO+FN6bAMexDJYaBfJPFetlJ/vCdP45V
IpHj5CAbWWCxPkC8ZHUQ/96i1maw7XlLBBv+jbm2DQLu2ADQAP0CHiAjuBWbpu19
OAlahGRqVCcXPM3izv4a5/fQwrckDmSRXl+dP+1VdCudzIvgBF5iae4RgVQFYVN7
ZDD1PZt8Rv5NKwHj5OgsXafez+dqWo/Rx5vHViU5D6Bs0NdKp3dqa1Ce5+TvHBlp
1XPFOrvAjxSZOVBR6Wsis9TXQoivu4cl+oA+bymGUfKQ9V5Km+uyR7KDQAVC2J6d
oGfxknLMKvRXOraH7gTaxigbQCalW3701wk9FYQqN+JHJrh3rX1GuEovHfo9YgIZ
Plmto67ceMDyMn6x9pVdKrrrn7Njl783FKAP8Y0Fb499kgFsRfQgrPnHUcXytqtz
VIh2+dNi5JAecD9Q3y8rpkrGnUQo0o13Hw/dl6JKU/RVqEsxjm/Z8N/gTR4IW2X4
+vPi7VoYhLMrDnzvgrh3kaUDP0dk9ZrfzuVyIFafFIFCCcFZNcn+AisXHYenBeun
bwvKwXRhILHaYqDfvzF4cCcjKEBsCN8MidxFagF49XZuy0FHE20cTzYWu8KnR3ZM
h53kpByTi0lV7pGNG7gt1PS1lg5ICjNSnJOh3wGLPh1S46cUCXWz/9eIcKtPrRm4
7zAaVym7cT9iL5QxlfZDfvtD1jUrpi8MY+2ijRmI3mLSkB7jvCRoIrjRxoLSkO0q
d+itJF1YDQuHmYkOqpGl8T7mbCqFy6ybx7Kwxh9g8FWvzbJtqjKqdhB7FabzoHP1
XgPkczaG9kaBEv9J1PnT1mIa8HWn1d1MhvO/ixWfYmXknC+nsty0KLZ1KIBc45Ev
pO5eDqspNSFR0GA5Oi264xYyMOMlF/AF3lWtYFlT9eGcZA2APG6ueswviWO9nz6k
Z1iBPn4Cj/7kqp+KRxlhsTvkFBO41XKead3o9HXH687pKdCLzqVlPQjAdBvLjMge
P5VChVSNmOVlEihRT5yHWneK/XFe7W/6295UKwDb/tvhuyAE+nzeuSA7z8OPCvdn
hlc/zERgXtPxpUSK4+bH7jeLafRAAoDaI/8kPmUiqS0++G1+2Z+mrgkIs/V7Fl66
jX7IgC3fdeKaX7IJ0WdQWXQK0XInTWoY0uMRIneOQcCF47Ef5Ie1Q89igkpeXlIP
dkXvRFpz2BWV7p9L42I7+xzoB7+nST5rRkdzJx6gwKsBCXah6j5Ruu88Jzmi3UmF
cszCbsOePNgNYmB/q/CjEv3+jjOw5gI5DA7BHY/4qr6JnavY1pvyyI+MKUjpfvOh
/FysVoIdfdBkK6UfNoP51PXMmjOQitx3qNm53+CurkLeR6qId1fR64gpVrTAbHGs
Qym5M6sJGXHfbnplX92i+bKgenb76sNYRvslVTagBkZyHZw04Z7ddRZgElwHynsB
xlgZ+5NOy0MSE8tPli6bgWcVvivg3jMTXw+LtC3r0z24Xn0oYGY3FR9gj6mS5lYz
+HrR9AFm6irCxH/MCEQum5UHwOksWu+K0abKYbch0A6/HWj+KYCqmHQAINKmfQXr
nNruryEpSfknxJb9ByP3/kBKrnIEL/MBIdas6xybGwNffWJ1mXVNtvWj8eJtBx4m
J7tmINlCQBdobGc/YrApwZriu9bAetkGKHrOoojCKveq191lOySrjIOCMeu5qEHe
jZQTYpt18000EC1Kp3AQqnOg8/Op05fuAjyQCKVfi6e50fldRCHQFQnVK1xDOBmn
i2U0nV1xYa14Kl9O2xnJ6goJdjPuDIRFl/vrg3w60mPwZY/yLNz/aMvbN9medCIu
50UgyyfhIWmJ/6u2IefpWiXBNrdR0M5xBSEoY0W1Yyot6ruVCcBzVJC1L1B0TDTk
Ja0KXxN75qKBwUZlCy4Fgvuj/XFcXrG0+tXq8O295kv2jlLpyENLfsEYuuNLwa+x
vUT352ffkWEo78YeVwAfkmRqORYauQpGsahu/UueKiq7fxz6SSKkJ/tUDc25S3FJ
Trbe1imChOC9WpgeJJlSZZ8Vs4o2I920dlSMWwvD8ChBSJyL2PK7HuQDyBT/llGV
WNZaGXSQdhY5aQFTqmlVDNXe1J9/YYIMsuvRyyGSKRBwdE7PBvhW+tSD5jzoocoE
JYAx+ni6TqDL0NzWGS70sTptZwM6h9apTzh5GPk8Zt0TD2tgrUqNm88f4PAFni4g
c6Vvi+uzAej0AHlDjRsafwUKIHCw+UCbl2fRNh0aSPP2CnrqPyGgUCToC8CEya7t
K2fqeX0iA8Hrzke5HtyDoMceqOVVp3YKaiDga9KbQZM17txLoFiieBVXRB8EqjVb
ywL6AYJeLEPlvxA8RGThKB1iqFNapNkKuKTibsgeaCnYXNoKtIt11JINviB1oX8s
lnOwm6MKJQgZUMYf/pD9/Fh568e5grXBClBFfZKRxSNJlYiJCL7iXz09lfbaAVTv
9meDQNk95aiDzbp4PA9bJO1ULJrD5a4TGVxPvX8QfJeartOLhjrCRovgFzoGkPvl
0lZ7c+GGph8YEC9PT4xOu9ZMn7gPVIUrx3AFsQKgZTB5LcX79SmXHj3/P47YCNzl
uU4vlbwjpfdPJa+ovPNjrZyyOnrryK2EZWKvyzVxkdQjHnO7vq2wvlb+V/Q6gKU6
edVvYuBmLtGE81ixWz2643zw3BmEqSt79/Q1mT3B2KsbnJBOLadHCD0+5DK1iFsW
Wrnbg4eDOg7wPS2iXOwFmAktKOZPSWynIBmb7prPgcb7hmtA6SYex2UOuTprz1Dt
E6NMaCmLsCkoj3X8fMGMlvFFPBaizGU4cuYCTP942fy7yIHOm2iLh31NATA8WxK9
9oXRZk968KtNpNcBXmBoqlYGZHrkZS9OyLilnEmwv1WHV0FtlKAaLwipmzFWlx2G
BpKghGi9z+AabiOi+RfSCI0CiWaVLhs6LI8EvBK2I4DcL3fBaYxfHxOse7haN7xM
AWP/OaiQ4zLN4lMoah9M7dAsFe+vOpcQquJOquYYxE8Ca99IB2dEYP1E8HlT84+l
j5buOyKA83CXHW2aRAbqZR8eJrgvwaDlW62hzxOTiY166NA95XX2lN22zIYLKrkx
Yzpo86W+7DlC7Murz3BEpZm70lAxBf5qJA8BKTe/lkAofKQR7fA+P4PSQ7cuO7X9
Y936ntUNK11qwNmXYE1ywhEWKrgFCjWaRJMIcTIKtmKyZQ3c4Ily1wcQkf6A+KkQ
dBOBEoOxhE2+c8dKncXfQRUVZd/01ipkeFyQPEtXmAva8xTZXhSTxIhydHT2nV3v
Vvj8HCrRnSVSKFDt9Y8qMtH/OvGjzAtpNR+nBiXNl1nj+FNYHLWfOFyUWmESUxlq
slm9QLQ6U9ocS9HF+ClvLR5A/SKE0pUbbeuO8XR9grFGQShnrLCWur8TH6YEb0UF
3gFVvt1Bn1ASG44F5bL9z3l2gXo0NiCBailLxUeXuzeko9RQdSB5oDcCHmfR+SNj
xpNcPSHDALIEeyeNFQHte3ykEaVCv3dKQ8yM6H+1ZxDeN+kQL85PSInokmsq0dKS
jBdTsaKVFxwuo2y3bf4l7fKzsEQ4Es9pr8jroWgPhWp+idq51y2ctSmrE86Wxcqx
Aiw9Y3lKMNummtbRBdyfnWfk4Cu/yEcG0U6x4NEK3t8WUnkQeTcsDCkjoDPebA0s
X6AKpvWTTwLf8SrtULD1ydzY75rCIYAjgRIdHkwEv4IL3eey4FKE+HH0QNS2Fml7
mHWdfwRABQXlHPhAxxR2jINqyHy5KCy0cVPOWWLbdMqKedEafJVnYqYoJ728sHu8
BMkiHdLn8wxl43ZstbrjTPgoFw0QaMhS6aVehnD0bHrAPt9P8GeIEL+IOfPYONu/
kgNwImgG86XiHsQojkGxCu5o2M84V5N1mKbDY3t1QmSyLyZX7Q5dqJNpInv5QxUD
LRogpFqcv7HQymzCr2G0NN0hs6J7pDPkonLhBhecejbQJt1fdUhB9Nrnir7qQ5OH
MBHpiTY7HpmWTCBLE7BB2SNpue3NqgKt0lkQqco/mZGz7gEI5t772I6i9/DKgfPH
WVUDXmwotaFPSEPRa5ydMa4s9mTH6EEM4TynvTwGqwlnLxK71sfayj7DQPyHKDX2
ulSkMnvPiPwUH3lKUajHC+wETEVVI3O5VQ9/o7i0pD54/faBVotklJyHDqjYTvKp
U4GN+lxhXhZTTfoD7fDSL5g7hj8tPre3eeymRJyYV1pb/gsoFuUUit6Ysyky1B8K
Ocr+0x7i+T9aqRZBDGY0A6Q/KHXk8pjb6AODB459EDrm+bz05H0Gp7QzksfNgvR9
+eOoDCnph9JYPtoW9ouy88hDqr+VNP2/Uh9Q1+R0Xw/1C1NYYjkg5xBS5Tr9dJEN
CbeVYjBt8qfftD/nc0Pj+ZDu2iZE5Vmdu+v/tlhdv/eagXdVtvhVsiWwIdYn3KMM
hMsmMJv3OLzmu+7sq7zHINZ/UXyKjar3nU3UvIsyVK+AReDPbiyF8LcfvZ2pmGws
MFimBerJkhTOYMSavRBEmlxqgkMKgFIhr+5R9YKVaGxGwtB0GiYyof4LN+4A7THO
XtQQlYHWdi9ttBnzGMu28wRFglQCVdR960DIDpzicZ8g1Y0DLmym9M5gWGSzBCiq
reVgXZx1nGEasmWvyprUlM+Ql+ZVFOE3fTehgju7Pr+0jk1txuDl5zQxDnk1xSu8
Ed5O4x/7Lgrt1hSDCTGWx1sXLp/itTBF2ZnDdHHuhUHzSrIOWufHsON0L0j297Ze
8DkHZgfNvhCeAq55/SemYu3POXq+Ke3vR0g44oICewZl6tLa84mqwJfBxGkfw+zq
CjgWS3q5UvBW5RqfA93GgYWzWki7c90gARIsX8J6wjz/JmFddLtI5lhyVs/uVA3q
MsKJfMXQC+3/I2g3RDLpclHWXNj1RVZJgSVg9Pd2x6X0Cx2OqWVDC4HhmCZuR6Ch
fsrzJnL74ifhp03fm6AO+kV0Bu09cuNUxLTso1oP1iExAxcA6yvBtv/QSnkZx6RZ
t5d0/t/Gt+6VO54cjydI/ZBmFAwPRmpX6foiuHP92ioPm6fKulpUXi+N8JTxHLxh
MXREeV4t3xREmBBFwrvPw1jLyfilSxA9cSthNRfPnUnjw842Qquvi/FTF3nexQ+N
5Pu50Qi+M72xkcWon402lJAyVeyr6UjyOUE4tePDKQehv8SFgq74SDFFzo31//uX
xddHhYLQhFE3WGS8uI2wnRyLuWRzNy69KvES5TvCuBZnn+LP/sM1ygPzXAPktJW4
Ps+lG8Vq3KqLH9NjaRQtLk0liBoXlZ0QOJgmdAvne+mjb26PGjK5FXt+c2zRgzSP
HT8KhgFiEqqIO+pVpcxWR0cdLaEuSWH5+Jk15xkk7NgRlXOr51FdEbs/B5cFfFsf
I8LdBA9vGi697xOnVGThrrZPk68tIOZN5+07CHHUlyiIisF/LcyU8MtzV8RnVi9+
t/lIYXT2aqZ0IfHC9+/824BReAG+qCyAyv9RQo05ul0xVl95pGuoOc+n6pwE5M4v
X6VXdOHpSsY06i6K5nwEp131A413/MfA28w3UxQCMG2d0qBgXGaVTLam5mBkMcDL
FQ3+xXALKDwZP/7rCWwedWASPmXB87kUVUgRBev8iB3IToKIbO8zobGNOJENgnJ3
nLmWNe+/7xY1vMvrdu4qQq5EjxAYaFpuL2qWpaFzyql5IKu/ZjKrOkfYBWlK85bN
hLeZlcRcamcUuEZ4Ft9H/4aSuhXjQoY85jFQC4acczdD6+WTS2fbr/4E1RpnSX4O
3I5RsvSYKuecG4MYN0ejhgylxZNbFqhfsNXrDkgTExtMNron7fXh9BtpVeDQKpAa
aBXX70KboBvfByqOG8v8xgfppmcATTCdmty07mxSyiVsL7LmRvfugiYHH7H1NTPC
rsgeA3jJhL0jRcxiooGTv1WsI7byPScin+Sqvve1N77LFZv/YTq4fSubVDTbuAA3
eyDuh8QPYKiIaKEKH+x9ipid6uXPxTfxcEIKsgNJeaXR5JB08Wn8TGtdClDs+dv5
smKBm5X9Pmdd+3hocke9zS13nVHv3NmepkaInIlqXf0lXr3FQX6x7AawkzJB5a5W
r8gYX5xeZje5gvwU0jdDcArY38fw0t6JC1RmIB+hMtr42HZyp9fEaym6la9B8k/k
IpBPyK3KV+oC0k3G+QHuj/rI3dim0nnIkQAS8bAbSnDxDEVGb+Mj7//3Mmm/hkC9
vS1V6Pf0H4Ftq/Ol5/4IycZH4ByEur0WlyAFvhcvUCt70sLQX0yoRBi3nf0HVLja
ECOYoNRVQTVVgYdgjZvXey0PGNhcsCWahNm/1rJhI6oi/kntwY5oBPIXa2LDLGD7
N1roZtVvltxA3TNQzuJlX/yBawXtG6PFxBa7u0jnGWFE1FIcJycNgn0Ya86Vp8cZ
0kKiaLabyEu7RgCXlO5ZYNiOuDb9EwC/2W2r51Clu3ORd9bgSxmC/TUTQE5OHSgM
y91A3gAAWYKjL9IEjUVrH4DMxMbopiBAVvPYeQDCQn9jOgpceWNI508MG28b1wDZ
yRAbGwW+j1srHj2yBWXiPfghqN083n0vznHrsMimsj2fOEYN9e6JVyTlxUYCuQBj
ybyQjMsQNPcbZB8Euu885YbUcI56cH6wgwQMV/6ldvbwuc1P+Gq6LptQYbNFVmHG
hab2SjsGvbuqQrExS7SLVw4l7tWnE90UEqwXsJvkps8Syh7wwZrL/cgEMwCkv3P8
yMDpWlFo90SybWCUdZbUGlBgkpct9iYz80F1CKgeaFogCX034EokEMbeJsMaEDZ6
vGnvEx3bg2KKM4qsbIwbO35NVwWyV1aAKDyT/wdX6lAOL17LGTYxfmJMgVf1ruC2
1s0AmUwIisS4dwq4E2R3T9MZDqnQZxvcDAs2TXaRtpeZDHXFKXqyDdZw2jBIHF6P
4JfJgao1QcE92laWPpHq5C6kPc4bDgi3GDY8WyTtWtdECRPWFHdu8klDHelexgn9
eoYVP0QWao8hiebvbcb6HSpeyMUVzGtEtyxQGZNc5NEv6GqopQZl4UeIq/sbu+gt
2ZbYxVAXeDlOPVTCo+6qpN88KjcbWaO2TH/iU9Gx2/hX3bfsT6pSdbp0vEZP+iK9
5wWpmKN3AY7mT4GElFuSNoV9FPGNwVa63q3xqQOxzlza70SkyMkA+QW73/KsAgWn
CkqqfRu1F1/33PBXsbkAotj4c8h9DBazf+67ozMT8gcWtFLRR1VYFdLDK7tuSIEh
gSW1H3UOUxKBboL4d/HL9FEY+gVRyujQOeNlziduhG3Bvz2stYFD+iOud8VXuVpD
W6+C93UScxSwUEKwum8uX1B6/PzJ9bCIwfT8r4Y8pztstcqHSjk9myHq8Rnf/KWH
5+N03jGejSs9ZNzyYiFas9zDMrJ7J+ZPjejRkTpKRpsPeOKc+k6u4DxwgyEu1A2+
6FD3nbSD8stDHLrInuIxDn6Ue3yH+F39UmhiSVfuheK4VrRXsG6UUHHju9FsOCFk
srTco9peO05SZvjxsxXn8RtZ84HPfVfYt7UYUdAhsCMWgld0Dw3jloiOOmM3xdBX
pMLZYvCPqrtgYuSulKtKor2xWx7533UAOD7xbGSYneyh4ARmyNqioeaB9qJ0YReF
TJojYkwJggXPMk8nO+vCiD2jLAvNGOU5ZeU8OlWHF4gsx5YeU9GHb28KzzJhE0Uu
z4XVVL702HfJGZjycehFljIh957fn+op+GoHlsQKNG3U1AjKUKh3y3LpEKadnjRq
lF8tbKvbTzt32aQKF06+/8069zWmi1y7tInjFN9lKFHgCSNuDD84/hTLO7CLKDr9
yklPotyWcdWU8HnuzI6dlWQ5J4kwNU3J+DTD4kEwqs1SpOOzN/74wq6JdrXM92ju
bMw5RotYwg56JCsExJqAjXSpfndRbaAdP/s+pZ3mG4IVc4EfMw12uEnLLURwt2I7
6IatMXhvzKPlXd3WWWRisoUCmMylhQLH+U8oedu0yWwsSkO4uXllK9xbHQKC795J
7/jiL5eaeIrLFjcuABxTKj4XCjO1VQRlbNS3dC0yOrjgKjjnLfN8iZmYjoCBhvyK
eod2FKbcOdgvVJjlaDxG8xAeFRtRLCpy7bnW9STuECTVo/RVNvl9AmwcoYxfoRzs
FF8inWgIa6GdzLCONE7quMQM1NQ3BD5CFSmGX5XyoCeqh9wVTkiIhq7dvPYNSxL2
M2iQTwfGWHei73xw4C3gN0xLLgBhBB3qN2djx+tZLh9/P14pv3e9RB03M+i77t21
L7U3s+Pfriv/Q1YvPhNw7Y8K5eiAxLJFlL33nb+rCdXciuWtS1PLtu8UV5lB/S+Y
/VbdMj1tkTZbP2H/5+yPLlA6lLPyzyVKA9Zw/dN+dd+dwFio+bo1TRJHGjqatwtz
5S9fqS1j9wESij4jL0K/lOYrFvORNpaOKCCvgxQR37fKhqMPPAVe+c6kE94NsRuo
hSA8Jm2UiZnb02L8Hyaek15L/GQQljDMPQ5IB+0TLYAb38Ndpj2wsX7SMALmuj4o
M0FU+sqBzYx77WNSUGG9tdaNN+obpfTk6fne+rD9KgopuIkidj/9cTaeaoJctgPh
MZXXQCT9wElcNBwgl6+AVDYHgBMVNSE3+KgufKfaDsdr4VCS0cp/5eIkP21e0mOl
vhslbodj5EL72/2ohXJLBd23LSCB9BicApPJrzytaucyA6Qr1m45uQc5Z/2FVcEO
neAoWLuOBW8lQCy4IxlnrxJHDkhx6ljDrxBwVStQ9yL2hQBgt/1qmiywCTPhyLZq
+gxsYlMA12Z1e3nnKfjOBlYfloDqlc/eDxMzPeonQqN3M4TSrdRmbGjeAr39BQwS
ZlJRCBU3CYjeKQ3tD29vGZvJnWELJJbsA3BuHJBv1v26yLoOpNhADQqyizZSwjwo
Q17OZE/iqYXlcAMxuG1wL1j8hjNLpvDDVBvJI2ShdMlB7rokvZ+XxAJMtA1IAn7S
vMMzySZlTqjV5YqsXJojIyDN0hepNBhbx3fTBUgERvKvEqzTDoZ2T09107/ZuMIV
giC4PhgLiPpLw5KR5eTsj3durq21UvGReKAX48Ij88i7goyf4hZf1lWDLafW8hNd
CYVBInfwTkBmdpUJxqN+8Qpaby8ZUgLn3Y3sotHy4CdpmsahlHIm4C1cJTj22c8B
QY6a3gnwxZyTexNxRkNaj4aF8TP10mv/tuggphpQjtZBVodI7kn8HLSvTXROn8xR
sAd+0PZNHn4MiuqBnA+GDwwoeorSg3QEdt9mjc/I5ETHnHoJTs9l5ynwjDL9AA9K
2NQAUVv3QV690SGd41QW0EUFn0u9Sv4lU9GpU+wvX9UkZ975oATmD8cdCt8I49bL
0+qakSi0qK68dyXFLifff5NG0kSIOiXEcCCK7Akiq8gYiMdqPzJr/c4l38HApb8r
lSdW5V9pmk2oehDlV3OVw/L1DDMHS0H6m46DZhXm94yP9sazIUgBhdY80e9vpBwn
gkYmbfer6xRR6ZeASrQa9OeW8uFo/qROD1+1ID/MNWSE+CMvw7Ea/zb6dbBD1eLh
3VcdZjLAzLyXrEnPwXvAxatlXx2wG0kGVghCvWOvqWkdK3jxskz+dygiPGLtXuwm
RWdJaeasqeaAqtqGnnJ/es7kfwOzmkINhyvcvmcY15dXohGicxn2yfW8gx7uqCMA
3WX5wZf6419pWCPzGQwSVs3f6ODELZSPGxsOg+0crWQzom7MwSH9b+Rofh4PvhyB
I7GPjG4lsdErwrEsI8te76fgy1Th0DxFmEgtmT8ms3pGCCQPOhJBWZvvfnkNV/w5
lXXXpf4fTF8m/xuMH4h0+41cVMaqD1zB/86sSMaRCqh3Re6dRMiF1AcrsExpYI/t
vQ4TvBeiza7tDEVWYDQeHbrPRaobvtq/paB8seI6cCCkR47E3488z7wpejZiTyjy
kYzRly6e7+N/RKqNdjNOPlGXhl3WXTHm6EOwDZL4DUjKno+oru0OSr+B3H6m9gdV
KFLAs2MMPatfO8kDGLgT7V24g0IuhQL28eTU2kCWi+GYjuI2cAFSejeh+4W0hTW8
L2zuHdmL02ODu2ZG5/GuFfrK8IEkbhIbQaTq+5fGJV6RWtkg/WDFsb7EmRmjVawi
+Ya5EJoFHBoyzZ23k88/wibAAHrF8XamITqsqLZKEVM3D/U0ojYBKm7hA+Wos4cn
n9VxewhmnYwYWGP52WGWWBg6DeOxLUyNw4vj4id8YVXqXVOmVd3RWYosn0zrt9Kv
5P8R3lfaz4GxWkJAxf+d9uzuB19Zph/3VYHA7XUL3nCIcMSw/fyMMViBesQIkZOo
De3fpbSRG+3hnF+kU+4J5TN0TX/21NMdN0JL8AOJbwnXn14B+Q2qbYf0lGbjqdhy
/RLmwPcTlO4Jj2EHBQxp6/hVu5/Tyz0z8uqhylkkkUb3RKt36DoC4BXhNGAUPEqM
+mjhi5pY96jR01E2RzRlbeDBrj1J/2gSbBj55bbS31bzGaJmb8GxRZ8Y9kr0BTax
Av2gmdN4/PBii9WBnAPPu49YebMZGOL9UQP8aJrndGk8gdpHBTylSaOW99g/iiKU
4gDvaTJBZVEta4hRI0vstjg6kn1YgDsLoeHrobnWEaztHJZqD+4SpwrpCsIpuOZu
00f54CMmET3IEWcn/8wwPKH7DgA354sdSGtOkuAhQnjvjerCY83bPl8a+IhvQoyz
XXUkWDNoJhUHBsVCvRQpaldSgUGXkqOH9PYFHp0oZu856TDVha+Y8ykqT97OnqHs
sOF3dzwxf4aCS2zEz70U1Eij2AtSTJZE/nc6D6OvZhy1ChjfPtmp9vlEwXoEbwfI
BTnyIpgcyZDRnKbzFMxjxsEH4lvtTG4Lw+Sr/Tbjuw9mpP71P8l/DH1fFDi3mnTC
v3+k9ufcy786g313tRklA3TSnTGZOlZxaIBcSwz+wyhWpjsq+TzIVYj2RUbAxhzk
Uz6ASi18tnFsvtjvWx4155ctULRoz/irvtTRV2kt7V4tSS7bWTlm4nvmkoEKsAUl
v+XI+XvYD7ZAZ8RAlUuE+zw7HFdRo6E2fXi4aCkaqJ2XfKmWRfmiLYUeYA/CYBvr
0yddBT6K/DXMUUUZq2haALyA5JyP27+51gW5lLdo3rAx7sWENxwYlfH0ZV+qwnj0
b/FdERIBcYUy/cUHMjpau8cqOv3tOiE3h176Hbw8RlN3+F2YF7+w+30EY5+30lPY
IrvUStOJjHa6aZ+GrhrdaAP01iFjm7/fZWSfz14Zlv8VPdKV5jxamfKG+99Lhcue
Ka65SqBArYhEZxAY8hrQO5ggJI16PKZWmYgFqeKVv+8GbbqWCBRtWdXajULEHqU2
E81TLP4ReiP5o74Z3O1pkKTd4mLVZ+zwdoehu69Ip5Il4bu60FxRqnidfqm8lguY
aFRAuFreqeU24CBuxM36Ka4PH7E91LgoQVFu3jK+X/4trZ8yf/eYkrZ3xu3sfLtd
ToewPUM2/KrbVQsYbGPVdexFHlKKK0o3zfC8xyxxtVjpQRU5Qye3uYLZPlIqxHrl
2OYOoxJZJhgs8NlSCZOkXmYqRIplo6HMDaLPDPgXSPEEq5Rw4jucLW8OT6qP57CS
guY3AadbMuPCdxBy1yhqrt3zaXxWPs+5hwErzg/uPpK4XuERWhkXkTLE9wz9CbKY
ZUTJgywspUtuyeBg8fWKMhtmzCuculZQ5ZbCSLu7pHiGylOoEPufhfzxw+fZSRkI
91VXam8xono/hO3eeSzDvKtdw/1CZusysBAUb8Hz5dW7pTh6iWPQPdQuhMb2+l6M
5y7ulU670Y7J0IFWk5+7r3OZkhlB+c+54YjVM2RurV0O2UCbJ1jb0NoEIQADjGDp
wp9QC99a0HT/OSjmLsdqclRvXQsT2mS/28ko0B/CJtD1CtgCo8Fej6kB6kNuDCK8
9dRhUyTY+Fevx5rVVkP/M7mhICxqDmQu4/fDy4XnZ3o3oqk9wTtJ8p68HA+L9SBs
ebYfcw+38R/lQfEImW18p64W7MZBKakVw49LBXRzwR9OWMY8WColvbxVfw1b1n0+
gSjlvkmiPJ3Gv/rjS/cLXL01Zts4sks99K4zZ8YvWvu6ERoc0RUad59n6r7z1Xru
HF1/lVhqaQSskPIyM4KJVL8QF9xQsjbbzwSNRJoQQXm8NAuLTiSRtkXaq5t1v8T/
Z7I7aWicpE+7XdMF0eyL7xToI+Pq5+vODSp5nbfJfEGvYv4iYCZQXZTWGJ3/CVLo
gtefIIM5CwZhCWvqGMSzu0PJ+6/xqRUiGXVc4qJck9NMNvseZqQ+MBSYGYLEAnG/
WWeX9fNxLNifvMFz98avd7MefB36Mdr+L+fMRpUaMbkHxs/JWs/+Eg4WTy/R98t7
sZbmxwPQ4ItNh9FSmk49J9lUU7+6MjZ1ulTFNVZVpxyOPKEgtjaCPSzAGR/BNET0
2Gq26imM5qoNpBmBfT2rD33PmmMtzBQGbpELHfz5HqbBcYL77/GHGlKx8rKas1bD
7u6iXuqVf1HhbxcOPnRjimoZD46u0uRVYoqoOAHRq+gcQ73uy9M74s7Wi5WgMpiT
SrfqqTjdIftRUVIirAiUWCYRT0Gqa4ZJLhYggnl0C7WpPU2rdnLhdhWMzkviIf+Y
Q8daD1XKlBIKwCKL6YZdQX6J5UggvtTvm5185mTRxBhlLEfQIkUrMLotuVlAneto
Yjiors8FmkKK1Gy85FFMjIqtuowf30bVahGOVVMsHCy5AJ0QUcrJqa6V6q+R/P/2
3ysKbQcgmqW6TjlgysywZ0fu3YgbDJ5t+H+fV6HagX9PxaFWbEFCKRgokzQFKuFp
jjR/bD1lFQyeU9orkVUFgzdbYNylCBjzNKUoZn3ECi6GE3FmmGrA7znJRzSoQmb9
Yjff3WS+zzodxgVCEL24XORtfOxL4cj8L1ZwvWWm6E72o2BAp+Et9pO5uMnpBrO1
1BdkdQZha9qLeFIg9/jiH11KgPqp3ioaDmJZv6pJM59qAzNO15juAolhgR1T3gBe
3EnO29T++z68qqTbJNZs2MVNoVswk6SUhM+Fa8Kog4EmSXZRbUzye6w2fcXzCd/Z
RRST/zoaPfrR10MSFlKX/11ipT15d8wO0qvaPFU//RoRxYU32bxq/SsSaRFWqZGG
XuUaWlzQm8mVWbwbCiaXPOWySlRZ9Mt3OFx2Gu9Tjsk0lC57O1zZbuccCVLC03Sq
yJDjZf/KMkvb9hytO6ETfMZDZG4FOFoHOtBW2vrVzhn0tj9AIQFOlhpn4FAloAhZ
0+VKnAp9fMW/bV5lv1kxHL3WDc2HHItR0Dl5EYhcXsQSiowVc1QMgSRnxw3b3qv6
j3XnpB3VcejJeLChqGCS11hNkvFXOhT11Ddga4OUOZXhq4Wc+xHHJtRS/lWKSeZs
RM8tX5Oa657VOLJTEX4W0wkFJkOoDdwtZVDVT7F3Nu4HuRHOnJg6jDmiykCERECC
GVy6gqZAIPnJ/1lT9Dujyj93PVD7OymRRjgioi1oX8mWgR31V3P4e4aLI1/JE8gK
eRmzLkZvkasrk23rTxtzSxvdJmiAeHX4b9Hs2NGA8VrCg3+npUYrPPkdIAtiTbYT
ZQB0JoaPTRzOnc1Sy6DbBjAc8PHL4JYj6R+TVuRwkfXW7QY5ACfnFhkTWKuWq1oi
7J+XpkynT126meCKl+6skxZu/EUyBTFTiLG+d0aazZnrOxBZbahPspuxnD0Gpncu
/jqyLpeI2ZV4U0WWn/ohnZc556MpThbmzQ36Q+TM584scLGlR5FVO3OB4CgCLIwQ
FA+30gxIW6q95RME7ahvC/tmokNxLU8ZQK32L114/kLH/sopvL9gp/CiKDibx0TL
ib0ygC6PY8uwu3TEVctc6TJEHyKetheALO35H8ji1t3bRiu3iQo6t7qLzZyxp5VD
hKnyZXGMhFafBWWpPr1GHOP70gaSgUvHVSS4h0eyfF8qbeuzIsFh7B19ZqzPPwyJ
+h2Ya52UPacFR3CJ/wel2wuY9PPm7LrvRXvnBkWs8hYZctEnBcTAIGfYMTiWaWhT
djp6sxrmGpfKy3brmLp0z/JK2iFatDbxjcLFgF023b0tTjM0joRqajoLp5LlBgsh
AGib2sSjHVk2e3dTDSG4bCItdanBZwIFmVk9jOeNlRhhGSf5MITTa3AeFdSHic3i
CQuNH+zAZuvqQOfjnOMnLD9FEjOd1OUBK74nr/Peh/sjWmYKodjJYiLqXRrcZz7T
aPHg/R7wfgOAfyo2CX/7Hr/Z+7kdbkdb4brW1aT+uj3NoMrXXGrbcMs9gI/rVbKB
P9IWz8sUwVZnO1nbCDpY0cE+3c8e456LzopGpgmpkanqKWRb234Ak5rgnysKNBIu
IGGGQiIKQapHMAlR3pGZWU1z2ks+ZQuqNi0G/DSKEcJdtJnrncBr7H8bYKzAYMCX
RNp0szQgtGCn+onjpwPjzjJeCmfIk1lWGFDbeWYcy5SSDjSN5+7+AaD3QW6rmucp
XOTc1C8SKlx0P3ZebCf2vCtnig4mKTJzhtNmL8SkKrSb+fdgx3EPuZjyXGuoYkpj
AGZF5CmmAju8D6kqkVLk0du1rA3UdqP5Y43rm6vQuyNi37F6On8hAFV/G31J/BPM
t3FeHLj8NEmEszNs1/iw92DTc1OPWbInLXdnFNWuyBd3SFyQwT1YIYtCaMWEp5RQ
XSh4jDq3o8UV824vxlSr4cKirKh+FZS7ab0fb9a7XRmSTCUJVXbraWsKTzlU2ZG9
0oUfSZ1ePZXljpE2XYO4dtYXwUZvPyMKoKRLI1ejY9cHQIcOaFdZVuMAf6cYYGX6
23E7GJQe5OpCbdJldjO/ynOQ5eScyO/oKT0GXNhx0GjDF6BYoRBvS8RDwFZT2+lo
eNPMGxgwezO/cVrFmPw2GuM8rv79JcJcNC2R+ae8pEVOu6dES0GAW2Ow9BTqW00t
z3B7U6vH2oRcDXITTHdXI5CDlWRh4Xlohk3ogwM4YOZUXLZ9WAsHC19AWV7VhRYo
5j+sh/sWS4dZej4FiuYJluLtYQ/ASxW1pBn+RW9lV9NyjuUHSe7d0MPnPmgxLYqR
toYAWTzbI2n1krfGDjhnjk+tIH7QPI8xd7zmnME0r2twwEWDHTJ095PcV1AVI6l4
90h1uqr+qwcC9Q5gUO62hjiGv+cRYxQN4tGXEkpo2DSVgS5EcbqlDZHPzxJziz+Q
DfJA3vNlSN/qBg1WSdnShEIoLBtaucR/SgOC6wuLZ8Y1hYk88f3oip4Z7sTx4t2t
VdUApazS4ZLbBblgdAAThUQhLF/OxC2gUxRtWKYb3zueYXXvWedz7UQyEFqr2Z1J
ujld89h3T61HeI5MxhXgvgb/CIAzfrQKHfE7RkufebKISXzqnSTAIJeqR2qR47l4
/aRQR9LxLVvlmFOU+YNxy/Asa15652YeCApAHpYLg44O6h+alX+aGKMYLC4vY44E
y7Mpdo/TGuUhefVXYHeS8KwkAjTAX0lkM3Qj56U1Fp0vrTmYywJGIY215BMDzTUX
Vp2/V+yR+XOoJzdUxvdnKfyhpsKvQrmjQGLZX/NbjUQ0SL8hLlMVL1sd5koOeDJ3
DVKyWrnN+f7+LkUuFEZeG0pVz6Ra786ikrzp+Hlvo2Q2Q4X39aibqyVHD97TuRqc
IgctLwkmcJhp7ggR47gJUC96LLKT8jNa1O44AsAILS+Mxg9dCqgkRGDAAfo8rqhw
zd0pyxjBeNwKcAw2fIrsuMSpBBomvk8PFX/eLcE5Hc7mWL9CBsQ3+Xhb7NDk7O/C
5QBzb2A6B9hkJRWFDTmsZm0z7MvHVuBcl8H6qbBQWnUDCe0GGvbbvCOd+LG5unil
TEmR5HP4MN87wkBh5Kz95uJlsh3BBXzUvRh2ZGNh0ESZTiapMhSuptOGRxJ9RXr7
/VdIyiZZnAOwLCOp5JnFdxPELpr5B0DVjYX9IdAEF1rJt55ZrcNoCv7CVTxUT43O
AGVV9hRdsbFmPnkZxjJNbN+95yN/V5/GkNaIMgaVRbliWfJ19lUOzY9zYqHawb4m
43Z+uv8Ang5smANbt1Wdp1dmu3cu0mbcvQXvHv/gyaIGoxmp8vc2bPqb15Ka/XTq
9B/LnpcC86g61r4lJQBfhWIDgFoNB5RmFVx8MD4L6xJNr/ecSVILiYrt/SMQ4JHl
K9XVmoJcAEw/CpfZaMvQvnK66WR/X1N23XJLrJ3mNuoShPUDLNaOS5+zipB59/dA
DJIiViHHCzBQ00lF/RGiKUADKgTZYTL5T7+sRheT6tMGs6/gGmWWsPCkDpuOw19N
QJY6zf+wdO2P0GokRefkGEfbfSZcX6LMQX2DiXL2d0ncaV/H+esj26hql2RQgU+J
ifmM9FOLVsKekSDXZ+9mMY9AjS6ONH+Mye4bmr97n9P5+s9H5aY7v9DKk0LHJWO8
WR4uNUhL2hzdIG3/3UZAXpLwPIhHkvtI1qqO5HUvB/oyl/nHF6res7uAE8F43p+3
VrUJpiqB5o2VJSW0rdgKD/lNLYcTEav05daSycO4scvhSSg4AT19EoI46ACeS8xK
jBZLU+mEMeE7MATgdcNHCQNy4mibJwp3BI8Xk67PSfoiEGF6NmYgj2wY5HFmBqZU
XN5zQI3bSV6ZC8Q81dTKm0AQqIk5ydfK5ilPh6nwKNoKEntw1ctBQOItbn49dQJo
Pfr7ELVjXnSY54314rh8L73PwJ/th2txUmmPfa0guL94Mwp1EySEonwGOLmPgWiV
D4Smu1s55TnS5knreQ7t/a9xu4SmhbY4R0r1l9vZIPzpxJ0ZWL3qsJWb/u2Iil4V
KOAP7rZrarWOg/nIa19EqhDBmakY2AHKQBJi4VxuDHfKSYkpnC7WKhkK9w01A7cy
SUIkMUr/8cRh25HF8uDbA07hWe+RmEu1aNeP7S/+W8mEZPS9pamXprI4LeBRTsKD
spM22/Lew9oyrx30QCJjxlKu4mXDP2nayDpW/lnIOPBi1w73J2ZJBzZQsMuX7O9S
f7jlXLHGQzsqgvnSE3gEqfKrz5WEm8+Z7TcukfZB1VxRWEFA2t1h8jeUUEpb1Ii3
11yZ2voTLqNiNEwt+1ZsMe4Jkegkkr6AJBteQSxWHVTV1GD8Uw3AqAgqO3NON0aM
KJQ1SVQXk+SB5IpAVDAwJiXSqpP4/eWz5a6UYWozT90wC+ZMwF1StHxfHgDAZIYc
UCvWVowq8A4ko3EVtD9Bg/e0Yx38oGRh5HTryYyi52zjQzvK6AGho9bfdIzDK0tT
wUtKEtynoiEQhfBt/Rr/cZk2kGB73TJofPe/kwvLDBaR7OUuxTJQOX79qKKrzR14
YLWAQkv4XCBnDWqeozj9dyTYGvEDHVDXpB9O+yr3/uUJmhBpDc26pSLn9/YVP1dD
eZi3yzonACOlgpf66ALJHdA24jUM6Wm08wWLC07EimFROY7dR8zJUk01UcZ4aadZ
iRP/ZS2bky3ess2Y64S2W+Eo3A3W1Y8wpFcsRujS9rre3M5VckkGH2wjBBtuc4MY
gV50Ek0j4q6TiEu2JecOS89NEUh3JSa/+6YUycAlf3MnZIj4GLuJsIOPmsrXMaSN
8VPUgGM/zGft+gsJMRvE1ImjxmcQLfNSAsQb496kVRc47KRKHVMc0yj0FGNhOpbx
nACTTsJenHJ9oP71STUEoGrhHuHIiPnKuH45XCnL726xWZdHS8ya7FQgq2CYWpg+
DZrDwcmXep2aw5rpNBQhYD+8JLAtsJF/hjrasInbdfHdFMKXcwwhaAGrmNxE4+5X
qFaDY5Kv7itgXk9C0TcIRkY6XEc2FwPKgN3yU+yefmOQ417IU7KnhvobOY97UWpy
uMxbyKFf715UuyuNt71e3k2bfjxH1ttWvuHB0eAt/j4utTHjsYjCXChxfuKGZ44q
uTwUvbjngk8XiTfDqTGXFuniskAIJDDZ+Pt2ORfNDqeSFh0lWA3dulVxNPYsoEYl
9IyhBXBcjSjlHOzZCOCWObCznem29VtatHNRTo+Uf+UhhrIu1a4oWxiWjEQmuLyX
UC/v6XKGTCHJaRbKFRMZH5X388Ufj2F1FuygZiJIbgLFpduTwFDbjKU75Gbk2RXA
9gBy2EoANXXbUEgDePpR1we3ASXqd60CRVc3K7lcVF5IrpWCegZbRleW48NzS7qd
KxjqErt78J7IKLmarx/H0s1gaswxbY/rA+D43QngRM8/7oh1JPjJzhi8FuF9PpAt
mMxUqOnFvvZskIRnGMiFQSnaelHdrCEtiPOiq1VHASTj00MIsoDgI5Q7X8sfovjm
Yr1igy2Y8L2O6h+uSzwxdVAUI3c6YEX4uFE0Y8pWfqioN2LWbrP9NkffUPvpabZP
9st0/Hx9IabErJtuwe3wAstmljjQJT3B9ngPIRzKNWbSDkLDtk5T5k6xqFnRTyPq
T6IZqvn61eqWP5AUX5U/i7zu1SOS36uZU0znKYNSC/i15Ysb9mVHZw3PMpKnDPXJ
1BsJXIQjF3X64JA12Qsmz+ywK8LKzxoeh4BdTmYpalw1ZFI1ZofHf53TooHSLZgh
MPUo93SyQgGZL5h3QK6rYb4qcSJO9UzqlvtyxhP7inULfM0/DRWore6OAV//747C
VGuEQSVIqCUD9omPn6wieMY8AKvyqs4lB1R1P2ZJSeLdGfDh+8W67DGYPCy+HZyr
HmCOY2JJsZc+WhAkwh2wRHunoJuTWbLBEsGsUW54Ppb4ABKRtTaQYQ3nUehSWAs1
/f6+FN3hY6LM0r/Ibyv3WPBFKp66BbxYrJ7F7SuemhitT6n/wnE9UDQmhZADoO+y
syB5Qir6BV0M3EldGdqTBq6Kc9EeAlBvQyA4ADbM5Sb0fH/9KEs4e0C2k3CHsY0B
/CxrdadmXI5Uxr5kpLeeK2Hqb78gzYoTIlx/qP+UP1nSkJnkTG0mA9RhIpTdu/bX
all0aBebpb5GxWsqvGUpGTPpSW+Be15Bm3vsPPqdQ7YWc1TxYhFHvbX4CMZZbhi3
KO69LKf7buReiTmkg3de1IvuyYcNCr9yuDoIpssaPp3IP9otKEb42p6eucZj7YDc
1ZbMe8LVt3qBRuBhB+kA1IHz3efjIZ8cmatu++rHZ9c0PCJcKuzXCIj75je7hU4R
9VOY9wxnvhX7DVZAHkyWZNNyTjApF+vvQZw0CQKicgWWvYyVba1P8nx/OJ2m+P3N
wXDPPASc0OLMGk3A5qnED7QEUkhm7rcmfuwuTBKY5oiCvCrAHAurZKJCDQveHbi8
HAbMc6vL5rG/ctE4nzOyIK0TMC5QGSzwLYGi3MHCgaQYEAzE5NRL9Rr7IlG/nTyL
fGLzKuAnQxpn/B0rzifqbbq6DEeAeqflLI6AH3UMuxxdwElMZYZI0R8Qbo1HJqKN
ZtGgDzZv9AwR012LAr6XU7WQs1DTP2PtyTSdB6ozFxXnhiOEWA/tT4jKhj6V4aJv
OHVNpSdkUmhcYQxuLvhU24drl8zy3ufBIpJweTq/6vPsv5SEgpzCxYdUyEy8FYf9
wUIs79vv+dkwhNToSr2yoTzeg/yLcAwrBng42Ry7ZU8dQ46DW72hxtfC6llUu/sb
XTwLosXhUhVx6PWYj90YVAwiX00xdvroZrywLU73iOQSUSxfr3ll86bX+dvN4j4U
6dMODnuy2Bf8BkgToYuTUu+oaDjOfVsDQ65jppi7sgmJzP88/T78p9zRNMLHrGch
jqhP+6dab4JXkPT98zF38Duy8Ih7B3OBDeNhYRK8eHXnW22++tDOEYEKUeL8u5nu
jvqAjg4MkA3XLBMJ7MehZcJQyglXwjRm+z1Ebgw1KRdu34KL/EkubLLU0VbG9D5T
WQUX9Qznzh70Yg3XPkUfvqZ9VzJDjxUVNLWO842UUYiGmTnHGw7AccBCrpXobb+0
wUm9ig+DC1ZNQ96iw7h26i4HOwqJ+JwV8uXEYRdyr+/GZvnHl4Ojs43x9gtMuye4
oW91qfRzwLgPxg5G7wxZTcSGz4zdzJUFiRi5rSEyrmm1A1nHcFKl0qZjtgDNZkSH
dStdnzuZZoPOrsP5rmjyvA2P8uM8zA0HAVhaR1OGyMpX1vT3kOzWITkAq4gbIRxz
QSLyb9WquYETcBA01sXQ5wb9orUqiNjJgepX/Ygaw6r62gRtQbjHtri2TcbZ5WpC
cdApwaq8wXAq7rg8vaO/PQvf7+y2Rq/V7ctxu8hOaxtoOjTB8/Bnqi1Xiuhd87Vv
bxQoh4nZeDa3CKp25RMcV44EYD8JsCdavJOopWf6eThpSWxiWlox/Hk3QijfoUUb
hbamltTWdm4sT/UQX4Gb4pWM9on24+w1v1KGZoPJcVqc4KXJ+bKgYtL7NvA/oA8g
NT5lMkUUNjjNJXVL3H4Gb+C+u1dD8Fikli0una/crCiABKrscfc+2+wLF5T7A9he
vj9i0QPIQmmfXoqO4ua575wQn4R4wSVwIYRBb1XbX8WMvVd/aVzqBnWfen8D7z20
qdUXySKPvkGTJn+Osf0z6234kaXNv3oH5ticZYVk5U8U/iA4q/X7Q4GaZTIIsHwQ
62Op94tJgI1+LiD/RB8doj8YPedSYBiCyXAx97AL5P9F4uczeT05qmNZJBbYauMZ
u6KP3prAVGTRJQCnsmb3WGzsbwykC+4W366qoRc3fxijKPjNt7UigMs9jcNwXrF7
yNy7rneuxPO8UlISycJCKooRRPHYoQwQ20dF1bSrnLuGXyQVA9CQsYkOz4/23W7w
C4wrH0nevbA+q7HwZRPVHPIK5udsQ+6my2bxusfjXPxb32/HK9B/y/LCrmUqRTYM
fSGItmIiJTwCsk78nkye6ysSxPoSn5SinrrGhD7qIk9lv590yUX3eRnPf6/5tW0Y
qfN/kpbpmlRZkwKPRNnQueDbNYJy4IOy0WJUcbXRJwP25+knPUiJh73T2HoaC35J
lOa9A/G09wBBK6Oy46KAREOvwBnt8wR09ozlejzh56hiRXn9UaXlL30X5VFTt8s9
wS7fsoSGqEe8+GV2KzInu8v2dUcCrKdrTwW8RKNLVSXZePpqXA/GqPzBFYlJkw3l
icX8x7Cos+gh9LlQqsfqIIfhDysXXvM7aSFSgvt7e0sCkjqnryuofPxbAkyV+G/l
wukBQTHY1bXtTJC/FDE8Zrqp22tc+9fjRIOy6pQ0wVDdlNEIrQ6tZ0LPZKdY2B4R
qxMXQI7cDWscXPIdjUpsmeQTdnNxL6/nnoZbcgYTc425Kt6TLq6SScIYb5P6WbCH
hqKysP/Zvd5RUrTKVsq8X5HO8/LqdJe5Mwm7T5tZCu3J2aRqUnxsvizI0yccgFhE
7+v1osbbjUlFQSCc0w5QU5WpTIaRRoCTC+/Dxs8+0nyCtOp2cJ5NURxRDOcyyFCp
i1C6q/T7JUBwMfl7f5D1pdIRMERs+3RFNayAyCOPKVjDGPkxdxedMbQntf/mJa+J
od378YsMpy5mKCImlkMhkHGfNX1xJEi+wEKYL0XmDC9ZR5gW1gcVzYHPLXtBgNFY
hGp0yrjUI9Nz1jqZdt9rB9qOvRfIqN0skZgvuBAytEo8/Y4hfB0mrjvVBMQNME67
DjWflT/e17ZRQXveGB2u3hqA76Kkhp8I3JJduJ6XdvvDyR5sICBSuJN+R0lo00QF
24A0smwxhH6g07radjzp4W+FBj4vN6xIBckoa1FTmgjGyme57ejZVF4cXDR2Wq7V
vAh/BJl/3gLlaWLVPd5G7ShfAnXQOCiECBYFcIurbGgkJj5hr0gl1YG8IbJETOy8
9JPoGXdU1g6pjZ3qwviUnpVSYXd6ylC8hEl7socR+ddsUWoSfjd4wZlMcR5p0EJT
74NnUfo+KhAqkeXA3FeVRQYyhG1bz5ltGiRaw/OBbVB5os3mavPQlc1nLiBf5lC8
wZfsspgYS0squ7NvwYbf76QNUv0yGSf/YDzIAU/L9fauaBMHiJ9ZoOJQRYKdvuQr
F8RStoVm32AilmuRJyBpd9UeYePg8QxFdiiAmzojLJoLDgDFYK/xYV/E97snfNj0
XuffA5ilQfxHE86ZhT3J125CKdhp0FYWE2oqm0dSZPJg4yhdgBZd8GSAvhAWnZsG
vzM0/h3YioH/lA76e7Q07kLWoAVTlmzFbZjrDxJ3pX51irp9qnb3jayIbWA6pQ0Z
gEIHnuY+LvR+QVNXBvJk8oPZ5O8S3quwBe9q5e5c/BsKhrWz68lk6/K7nmbfmtOM
/zVp1X5oQCc7UDPbGrh8MKj92xtQHWtmwPcOQJf1R2XGhqA3GCf2aB5WOAL2za9F
4qVWbUmU2ueGXwIavkowtQ+QjxFh2Mmv7Yxq9ZfZdwenjHPNTwI6fdBdoS1wldIc
io+nO4RsUSvY0vjoIqGz7rRfeaPXjURcV2+K/Rq5l3EPG6e6f41sgGFJyCzIlhr3
7EjWw7UEhgMUC7pr3JTboWr1exeSK0ocmTjEkrL7VVrCaih6WUVoloZhBouzUO3q
zzCRh5NSSZk6yfOhOqq5+5CsQf3tw37qG1mcQtTq/IMJpxnMJJjXjZQJ44Ip0PuN
ipMOz8f2PuLHzRQMgyIvxGh/H0otL7UTHt4ZEgWRc8QlZvZMXTS44u+ZxXhGd3HW
YhHwMRvBDor1Ik/t3e7NJmVGj7LVi6wdilxQaxQKhpzJBB/s4eDx3aW81eSlvRlW
BgK/JEfoHrP80fuwGYJsqCDTt6Vd4kSBpQH9ttAdMnpuL8iOy+jZGvH8qr8vCeNR
4khA9+fF9A+V1SYw2VWwD+f/X8NzSNifTdDunsZc6r47Q5KpQb9op7I+7XPWr5dg
I9cQHkVTfNr8ryAqWjUUoCINai6tbt3kL18U4HaWI5+qb3Z5QoS9gpxAC0ikyyB3
DKi6ivh4Ax2edklYLAC2Or/FcRwQToYWoOsYV/nHLw6spS8TtrHt3HqrUOoFOHfq
vsUvhUbYxhfFni9pwNIYK7MyGN02Wi3gMuB2BWT192IqHDsg64IPN81QoDp83Ee7
ieAclLkqlKSL+S1SpPdTmCdLYUJqA2YfBExYgowBuHh4t9u1LKNCyLyz2BJL5hg8
E7zhP2XmhaKnY+lVx4takKo35iud0bd437AbXc3S1bpyMJ/M1Rq3JwkRCEhIReG0
OIYk5aJUB9RNGOw44wMGtV1v/WnpE6Jz99Jcjh1Uxy1JlfssIqSy0Sy/0NvGGMcV
g3iGF2r5hDpHxppanJIbyYUmomfvZan8HpK4un2iwuNCjxBAl0oCqfeZwnYpSyvJ
+eLr2mQUDCANJDRqX9E+hfWGjBTYP2mybl2sYV7vzW7fjupDiHjYHs4Y1LieG/6D
LFXbjY/wepbJpjgW4OUaZFNXi2rwFJ0sxei1pJHNedooTlZ3msxCaNxretyj42gj
Vqxtnz5U+Zhq7UktComI8IIzt4KxtfB4DeeaXDqbN9XSoMAO/2gTHSzx4I2NHMRY
RuMj489X7zkdT9nmNz/skGqFdF+ZuVuq13tUtyHbpoaj5mOJzYosfTkxHxXPzjCV
f1TVKDDCwB6vBMG76+cJLvu+lCVMX+aWpQp8LVUG00Uo1Esl0qA8Jvnn6961n/we
QuK0/P/GH7xfqSlOQVdkqHh7aRf2t7gNUIrFOnd3f8VypxQSUZFztYuXrjsGEfk5
CyPkYBsUhJE0MGC+Z0q0xl3SVcEdcR6AP9ygm0WfCbgaka8F2T9oXLb8Fak+7TOC
8ovyEUVhzsKoWo83I1SU2XR5N+tY4amZRv8Lmtg50dlov8D/K40JD1NzURfuVQvX
sIeeVryaYmHx8aHuS90Dht361ZYsf0p5wLaKfZGwVcdkkA923vDQ8qCkeyqfx0Qa
TH0XYpkoc1kCmivSxliwpP1Cf51LTTcGILvmuiT4XxBZqwDWXUSNhLNYPuoJXChc
U5596Wf99OORpsjXMTjDMEm8DOnjg3+UXBti9Nj66r6wo2Le18/CsbywvqlEudG+
OHYCjFEm4dUh1NO8o2U+4oZtqPnn92lL0BLvVPlRtNK5ZwsCD/BtrOE/+8r9mbD3
/ksQ9CN4heytmGTaOCAasxInHnHeV1xJ0xMs7PmtHWTZ+bF0o76rPQBtuDhoW8/w
2is2+Mxrr6c/a/ImhErDTHXOeNgfqmEILYUmvi7Wqmthtr4XZsFKQ1IsShFsO29U
1/X/ahTohzm2I9kvEAHWIBLuoDE8zdlb/tjx2e8D0m/+V147XHpBOXig4NmRwKeO
WuvndjFNSr16IRj7Mu5k6pCRZlre8gFGZEtxeTCsr2MJkkNFrKbB7kwc8FJ3u8NW
U2Zre6lZXh6lgTlpg7c//y6EwxwXP5ikh0X1uF0YGH66Xrt6xqqTfgTogHRfuHj6
adF3VoWekwvHfSQ1L3CGvmet4RxG2rDnqy0bqJZf2+R2ckE8y628nV1Rh9eF8n3g
xzERqMe0bXQSz6z1ysaGRq/a9KX4fWcVSFIlf6JlUTr2jSFDH3rLYDIfGyTX6lKq
+DRr0vvG1Pnqb+BPTPqGKwzFBAHF2teeOCdDYUPwrHCwomLLjhsSkq+WhPMd0QM0
/29mAQ12p7POAjoTp1HDNgEwaB6MYTmrNX3vDH5nVf3SlYc2Nwy3TtahiYcT0JIC
RiRr2JNsTu+uo661u4MPOtsI0GVhcDkJH4cz8cdOivbqs5toFlToG9dQsXGsK1AR
RUiCqin7BzH86xxg9JIZWttRMLWWWG8ThkGCnZ2NVUFkxuMBsO/OvipP17jlSIE0
MFVbuEGCm7M8vsH1Bgmz5udE1Fwvn60aIs6xW4H/TFnlMAz6agR9y7/lBGeXcwfG
n0GN6PjGIAZPtB+PJ9yyvRIJl+O+s0pEoC/LmvEPO4TDhqkremGeSDw1xYPq2gAT
7HJQXkWUyTrWBNDBBPJVNCTmPe6VbEHAZqTCm2IwDhe0zUi67sJ+fdSUYUdq3Ds1
mpZ9pZ9sUn7uSSLnOyZg1RNjxnpFFhRIAMycn76CbGk/k5vzR1RoFebihc/q0HrK
LzT/3iTHNveIRJ+oZDaswEt9sNglXvh9bhcdCdwub2504lQr/gG6HJEaHfKu10IF
2TKvBxRV3gq63OrFz9p9c3EQg8cxdk2HQ9hLSEeWegPPIvhm3YZOyDKVGfEuGop7
y/rZaGtOWTmkeH26wh42g9i29qvIGqYC94syLp2m4l3+tVeLcutotdeox/gYg7yH
bixkN3mWmjt3vdJnLUpV/yI48L7iQd5rRh1XHSAfXV69h8MYW43V1/xlRdcm3CIp
HtGBSmZhK505nWL96IX3TROE/8lxpaIcl4ifFIRVWN2gx2MREbPxBJdn+dtTpm8M
Z5bVqX3FsLzJKFg/PZ8fInvpqWgin122pOjTHyB5TykdZCca5MX5UrLH6kodechr
V18TMdLoYW7Y8ro3PoPaJ0OE4j/mm/c3znLF9V+d3hL7oCvD6RvToXGfa2WJqNB6
qvI5uQpJF9PUJBUUo5D30/f333OTJejghlDqSVkoKCd6o0hgOIGPGEd8zM7UrVDM
5aefnqFgtRtYS5QDZmhD7lXDgBJx+ZZS94KvFdJMJ9u7DOFJcKgeO7N6Sd30f2jQ
AIIgBMo5xGCMrc2ctMFMl+UdGwMUuIj2gflc6L81ZUj2CXorUqh6VD4SloAC5jei
9SOiWbpLrL9PhuJ6MNsHtiG3aJsjbrC5R0U1OIs2oT5CBq7NVLld841PnWvYcDkp
cZLsJ/EBRZCu1tyLNyat9P5r5AX5sgtTj1+ps77HwkAOFl7dfe1ws3boCDa8iODi
TJrGQ6HV6Al+nYKng2LDTKdq+kz+bdSJLxzS4E5qmK6otxvM+d3v14irOnYeGO/h
KMvD9Q1kfTQ7vVn+dBp4Tw855HO8lYXSVOCUNM/TIHgwt4ktmiCTVVuwI4l6IbiS
4/f1o9U8r7KCWxeLeh8QS0VncD43ceRa30c+fSyEaBZHCmMz2k+oQFxdtSfj6kh4
MN+2MX4hfnYFd1rzss5VtDEGUQhvaJsB6uIfnE8Jj58DbIAPiV1XSuQF3r24JvHg
aGZmJu+9nEW3csoN6RPV+eq94QQStPomNpxqyvHJ81xvRk+rShc1trvWIFpLffJA
InlQbAomeHTGASfIvrOKrfa+7uNbBEaWLq3pXAx6zTwynvndhZONKwxAbAOlHKy/
sxLabJ2b0fh9BuXDiS5nGWe8U3kgtOjMkQtRk/azK6ctAkOXybCeQHIioTCqwF6x
1V1XFcF26AFy+jGB+alSO9KdEwDp6VkimApEgPeg8nhOtQyrW6eI2xfH1fr+mOJi
Vderb7xoDf84JcYntNXa5Fmxjcd5pNQvtb45H+OIyfIAnHpyEIzWDouPwShAesL7
RbK47P6F/drIXdpgcbwkW8d7MYWh+53Us4dg0aL9SF7O8g7NCgOTFx0xE+603VDu
cRO6p4w7v55Wd6lzpj8444AX71NkqucDi8ReaQhSZdvwmUHJgaexmK6NcdtQInwl
qnLGKBoo70x9rg6CiTkMfhZDOlSD4P2qgmqvJvoI3dxBVXzDP8rC6/MftHIzMPQq
0hKSMl51Lf0zwj/idiqPkTgPx9SLfM8bziRyGGb2geeEAs7GQ0GOtFiT57lFuVqP
B5EBFb7kUZ6oZzRgzOx+D/WX8e6EFY4Bd+GGCXjKyiBlH33bVugnReRnKy/sFe/4
ObZUglew8bfFDnLz3AhGzcWom2qo2aRcE0oyAZjORfJkkElwLH8h/hgWhsSjq/R8
bF77BBAYU6ZcdVd1X6x2yqeU1laCKs2DC6+dX4xcJH0+svZ2pgLzBMMOCqZnz4tI
lZyHuyaQvjd+RXQeTUr+VQFza+wBjlVrVlji4KGZNyY/08+s8W6wkv4DFjW/wH6a
AKmg6nqac+SKw1TMhngTIXvO5PLrw7SH0IeMZ0vFe5wxJN3BQfdj9IYzhHk4B0Dn
vU7A7qDUQGAUdSJIjTJb15GXUbHsPrD42AJEnN6qLYMQnTtEOGM13F4B5Yrl9WPm
zdGZQ8Yo2c4SNOVMglXEv8TSqFrCzmSBI909hUu3J7CQVjlo1IKue7amodemno8p
BufGTaLu4VBPsrYnh4YHofJ64ZF55WKr7MFGUANQz91kxuUfHtBKi36ao+Molurs
rnJTblohARQMmFb1nHZpMYq03Lv1U2qV2PgJr5lKdiumGsuTP43T5E2QYwoM8n43
SVx7O8Dc1MtOtYryhZ94AK88QFU05bOpmjC5RTpJh86pIgSKpOAVEok//f72j0bu
qSXGPWaz+UKVTlWiPBuOuHpC8dISxTWtVB5r2DKLirapg73ba2dcTWT8SlotScFb
wxWluzJ8Bbzy0BHzkSudEc1zu3Zjm3tJrFgLuhFDYS3aIEFYJCWqjYmDz+x97klv
Bb703Jk/RqjN0U7wQUiLHtL7kmPRKTMef/B+S9y4XzuP/gf87LENCUoeOLTCb8tc
HHFLwxdhJTT3SbwO9p9mvA1oHPvirBxGWNed4vWdW5yDSuXupN6kjPjEIuc7/HQv
wc3+8rxpkgzfQ4LPtBRkYpSXqI2DZm6loySfQb866STq/PiWOrgl6IccGLkSv2Up
AWtsYxr9jaenGpdIN+C+1kOw+M8oESVp0imvbflveNybyi5L9OtBxS1rezkjtYC2
QBhyhaHCLWG/Gd/mD/LJbxcPwC6yy3uiAnjqMNUlmNq9Oi6tOjWZs08/225qvj/K
cZrXQdjRICzVJRQzcU8bi9tV005QFJPdNg4sWz63hiyDFzcS6goRngRQiFzuGSe0
vMcuiXnS6PgBVb7Kq3eFq68+x5DE8rUXFPLS90mWgjJKGAfZnzMso0JZija/cLQL
SFUl3P4wx3evhcPX/HLsReZiCEx8010Wf8rMIpHvK9dtzDfQnKWhh0L4K3hT99kc
gemU2QBcpPa6ibMDlEA3EAP4OXhZqD1pcHfR5E+oxIweMDFBh+6M9nC3jXFilLXb
JTCiMHQY72MxLyxXdQMNpMIzCJvybKdvfQAanPsi/WqXTx1XNlfWsUCo2REbj6bz
KrL8UQiaOrKoCNq4M4e0xNEW0fQxs5pzewMGuB21vBisorVuGyfMbPTpL72jvqGm
tv0AQoNUwvmUELj/eoeDAx25AatO7Wtg0JUODMt7bDa2F1SHdO4xprqbU7z3FAkK
+FxECUcRW+bis4f8rg60Pubw4hL20njPCe0y3UaavMANKP9KSY/uFu5hcPIMUnIw
YNpOiK5xIgiaSLYi2++6Nge8840W/AkkDWML5PSGxCANqfIGZYST/0tS9LPXR+xf
g6cG7X/P02TRPgJZTs3PJo5PaMrmvmIBgDZjY90oE7gpsDBe7OftOfHS4g15qsAP
MixrSdFxGTM17vyvxhyQD+1HWrAT50LqdzSNxZm4Q3Tg2UgrkwfGCJ3YpYejwuJZ
RWnf0EGfrFmhIAjlk8tpgKyBnoDjFYY+L2IDcPlXE1n6QvoVmOjQAwStsr/U9pMu
AWTXRd4R/93eF0+0TXSorAH0UVEqQKJOyfIYaKEH/oE02LmowQTKfcm5udh9UHMj
wCmxBzZ3+20fXUGWfmmw1vdDcuJMR4nryeNh/87cMLEWs8pQdURsUUyzxeXhXz6D
sg93AsG7nSTxXJTNaLFg15ecVO1SKR6ygD0E/4glU3tr6459Xrw8zXGsQb1bPxtk
J1zJSKk7Y2wxf6tIgjwvzbrMrnPxD/8e33xNP5aH0a9oR13qQfBLk2+mpRFerdMk
8Uo2ZZKijyUVENXNegK/5FJDWybM3nJToYjKvx8aX9MclDj9zYb33gSsYcEz7e1Q
4zx/I8DCcKu9y/Pb9tWUVMkyJ3vKl3VdvcTfjFLCW4OHdWnEQGMl0vPKeYYnLr8M
Fp4ycUVQ73IVULAbbA3McIdiO/ZXy8rXJL/2nrQ70JzONNC9x1k3hJAGHjXYvfUK
ryZ0ah9aMlh7mv46vYXyf9OPeDCUXk8H3hV1Hv5xlbJStw/SP6E2/mEAIBnXNv6C
P3Ujoc1E6narDd027uAxH6/gXaj45hlyMzlJrhsRS/0+MR8vHVQrg7h7kN7Q+MiX
VFkY/FD7e0NxQLWO0YJErRE3l7c6rdWaPeBO+CguPJOyp/pTfR2MzXimRzbFYH1b
wIQOMXLlpw+dJ8LY4UQCIfcEhjS76Pxq382pDW254oYgORsN3U13gceJKeRC1jBS
BB7B1kfnR+Rzv1Vf1CJ2LvqUS6DdA5F6Y229K7GiKTG6wKYhBktHua5p52bytkdz
BNdd1BlVbExOl6NdKbubIDK9/j4g7nko70BAw4CXo4dfjQTvIO5sj8y/0FtPoVVh
EQxT7yLpaWpouaMxEUTaH6Z4n2FFoBEJdSAAUgyNU4IBI8blI5+lbKEZjvltpN79
vMfR2fwXX+lfVhnf9VmL60Yyn2N4vjaCLAjxXMEhdlrdTZAjnVeK/XIxPfnFSbJ3
4nnUOAfwoctbfEDPJk9MvqFu21RqTyDJl6GJ1PmNEBZpRriUiFp+4ILTW9PR9f4C
IWmEfnL/ydmhOIdzOE0xMccLQ7wFD5mBCjxGuV+E3ewGYbb0b4En7/6Gryze6IAn
rgD1fJjPL3afNwz2TvNCCUU4jATvzvMiAdqju6f0SO83poJs3nn9ZoFOqEvIq4mQ
2Cnee+1XJToImm/AIzOreJJoqsxoe0X68xLAY0XKt6m3FHkkxRz7iJffg/jBFv07
7YXFc0u4cMAHcDEcsbl9YdEZ1MDhiOVvFLEv/xlWdpyaLGTo0JEZk+Hyp85Cmz7D
gdgXm13D3C//HJqv5pvWstKP9btOgYrxuCCgoJdlE56t87vvch8qFICGM1wMa6CA
tfBqhRuVr9sFLAXwI7rrhQPDXmY9U2e5XfCouxHM4lIhwcr6yBeJt4RGXjnvuS0g
tZPrvbaP9qRhsPwsB6PDximinULwJxhor5QxAqbHedOX9lkOIX0YPtIGQXTFvpM+
qWwcb6r1dJLI5r4WvyhnVBFp/EWcqvdROAxWojGvGJQAJVuY6A3UHoIEyKirej+a
z7YPZj5FR8UMRY2Xx5OUkadeafpEPW6NvlER7p0KVRzyxHyFaykQjmV4q9iDsBil
lLj1nhlHhisHSZGkc5StTsZTP11nbi2Uq400VsrrZuPalCm2pedSpPvS2zh7MJgF
Sr0WU0bxxFY/ELBq5Ki07xQYx7816sNZ/ujkMEKcnZXnw2t5TB/yp0qKHRRfL3qg
CB/3UnMKKQgmy1dXfMpzLoB6pGM8dQ/9zVoGNKOXzsJCVGS0Hl6OEPDbWyf5+mTd
g4ubKcACs9clCb7vM8Q9ac27FjiREe4yH+yAOuWsVDX1RiBLFta088N76OvNzbQV
NID3xEM3yici0HDifoPmyJQeT82EhM0xrev+yLIcxYKlfhyBiJedi4eeOqa+B8ZG
CuojIS8H3Vj3RyGY5eNBy634H/PzLeayZKbJ0LoXhynFrup7D0GeQFUzixYxp4F0
zEXLoC4LEnHhJdlel9CimqCG/YkSnDWA/T0td57Gp6sX0FWgmPQL9A9nkaUHLjIE
k+5/P7rg7ektNBvxGcFEUoHjifKBGp+bQJJaO1+vIdey7zJskWMEFJHVfEuYFbtx
YALV0xUGcvzVBAWdDIXtERoR4N/txMExGBjjZ+sJ+A7zhTF5hGOoD+8sVdi2VPWO
A9EFKN4wf+P/yEsEKuxWpX45MWn+lm+Bnbzna/25RAifcqKBdB+h9FDCrh843SHl
VDaTZ1511nMIMY7Qth/+C2enACHVby/H3KPiHTCYXvOSJitsBKaEpbCttk5gFw6N
y6X+MBExLBgAoCLFFtm4wX5jBa6dL51SwNi/EhDWiFf2h6oWR9EPvm/0+OdLmQD6
on6odA1dKYX7RhFM1zMWLW4qnfirx+xZ648Z4g1jWB0kRT1gDS76QL8CBlhjqw8u
tw+1giiOXXxHW9s4lhh1LTGl4p7Snrbrb5O1vqE9DRMm66rDNXQfOnnpY5Z6Fsbn
tp16tpIapIR1Yyd1Js051rdXJGFPBmYzyr5d/ftLG4P8u8Cc4vFMBTNq2IkckcMB
gL+CSBlupvunvEL2FK+k0OJdmU6eWPMOsxf0IiG5Nw19FDH6f706JJXZgx6nuEvl
Eh3Pce18bDQI9bE5i9GV60cFCsGdEiOr9gc/5ZoNPZKWww7chLN0eAZTbl3fCOvB
BHJ5s2yF1uNCNglFqW49sigK/Jcw0VtK2KaLLymFBI2CRzK3UjVMxuZVdvYWE4gl
bQAo7gBNqMzmKUhiuds9GvaA5TWIYtpfr0QAYD9LjekScaj23HsizxqNYFyOEZTY
+21ECSFRPLB1Lp6sBVteTSyR9ZVQ3nisqJ1Xe3AfXJS0TQHIZ50rtqEsDZ00fWfU
sETfLI33xsxwQoAY3QyMgs8+FNcpp/ySemd7rn8mXllSKi3KATfyLrPDzi4HWgl8
CAYfGRl0NmxmcnXtGnSaLXnT00eNsRSCB1TAOC6MR8XvOvlfRAo4Nw+XrVsTnghp
ng/9QtUV3AnY3mE+GwXp5In2Q7x2I9d92BGLj5vkWuFJ0+MHwxzE26yu2uSLfLN2
gMS4ip9UX44AL1SM1klhW9+AQaepZrv6Z/y4w75asTU4ErLN5eaTe7nI8pqHzVAs
IWeaMPjojso77vg/iDSL905gHP7qLFWXf3Ljtqphq4Y1ngWzJaE+3K6kTNDROfTx
c/7+LKw0TvrvRyhPvTRI0JNUj7u5gXm8kDDln0y9bvWjggy0wXCLriYAPqebJLPa
ZbCPLpQNPgxaOZBT3ix20qBSkAd4nmBf6iP5JzqkGrSAGtP/3cFSZxnYDnR9m8Iq
FhCF+h2/fBOfonQbFqjNG3dfa+wZhbKqDxS/p16Vwhpsl2VmMXN4uyroV2Lblm13
Div83gIrQOs3QSdP9D28wuHJfHOrSDwhjP4dJEVQpg6O/BRSO9Q4VCRCPBboOdOX
67ppUS5oSsKcCmRpXeUso2saicpxGGSPDF6B9ve1Qxaz2M2X1wHPvdeC3/LEBXkH
fLPh4Yhr1pJvcg6B+RG8CGvipWFb2Z42Iis+URRYIdaM0zpRnKP0VNKXSwXAIDBo
JXVhBLEC93hNFTdD6Vv/qfULm+Imypogz2MdtXr1KI1J+ptmkRNYuOlKB2gvcrvF
8/di24XUrmlNl8DQMgkuFapicwkeX+n8b9NjTEbCxzD+JZUHyCY/TOfJLWk1iTQB
hDJqJsTxNDopo1Q2OzRTcis8Vp8Tu4Q1dx3dZv3aaLaaf1ihs4xX3khtCdrjJDmJ
5nYRCPwWbWRB9ukb88D8/CI8AdA+L3S5dFSmipiyyyErr85YYGMvr9Of+ByBsquN
JMIdqoC//qrAUYhpCC8OLhQ9BaC6pPJiks0larJO+w/TBThzHZ5pYBYPrjPV9cHF
O6NyNenw8jNmg8KGI3FxpIZZEALSRnOKc0nitxsN3GJdfCJP67j+wOx0X+rp3Xnc
eDV4mczX9Gu1YEvO6XLlFEPu+DiJ7bo0ms6xMLmn/HJ9uN8ztZY1qkMoBVtnLrXS
liTtfJs9+MECKAs4YUbGHpE0MQDkOnk8D5McVm/r7KOfADrRZAs+EM1G0oP+7MAI
PFrzsZur55TNYAzKl+VU6XB6RTG6MtvUJmsXS56ZUq2Y1mxuAUlsrWIHwH7pnDAm
iTO155hlWz6DV9gu1Y1PBr6r0mKE0hq3CqLO3SiAlPPjx1HNbjOQAGN/5bBIkEPo
FEdP0rpTqzF/jakNDdelDll9Tce83rGKcDjtZy/5h3AX9tftqxqKvI83spNiNKLV
mmJNOHXUm/W4n7Z7U/DVergMSuq7PTsqul/Bn/f836CWpF5i7AIEkf6iFIUoNajF
FaVCZQN8eMIK/mbv1YQmOqW0BKyHoo4u7ZVMw7K25UDCSfNMP9Qt+9QVFK+d5SIU
Lk8PkB9l5A9ii1H90mT7ezxSGUvoSTOGwPQK92wKBSwp18182oXF56/Ueu8qNXVE
7acmjWXTOBIBIv2FZh2admgRWFXC+MMEENfuBSKY3+f4WZ+p3wSd7LFDskkrGiHD
02tx1AzW3iV8syCgBCfL1pT3jWVLRR9uLCpaLAx/ig7HEXQHsRkTI64ql2ZgsWb5
gJTIA5gf314alXgi/fU6Tt0xbwi5fIVkd7v/QAn/iusjWs+PLqMnzHtW9kaUdwVD
zz0y4xUU0G3jt3PLtCWAUnND8NeoJAfsXK8ABuX6cq2KeYIgzTEiSLkD4I+p6TdF
H7CsGlk5h2mB12r5RS/S49tX8IgWNOcGG7uSh2pTq4jYBEtd+6yVHMCajzB5Z3zw
GXW62nMYhMMZDLkn8zkKuq8WYCxKuGGLuzbiEBoMbQv8DZTTQ0su6SLQ/qbVwO8x
N/1y8+1lGghTG9Ucddxtg/EZMn3+7DT+tk/tkCZf+FIaORqbTA4ZraArVkSzO+Cg
t2C5MhyVcZiwgf13KEdt87vy9GezojQuQllHR91M4PRS9rKkZEUg7m73vli6tYwZ
gLRNESnx9NoXzS0PTJieZxFy4/Ke+CMp4hJZrdPVneF6UIPYARKCN/PdStQOdGTd
YuLnPSh/9lOkFXjqYGdSSsvrbRwBlsa0X9tmzdTdf3pDcFpQq8cOko4Ce1JDRxO2
vC+QRhMax19JS6yA+dMYPejQI0RAaoypGYQX84M2knRCb5Gsu4ZoWqlXNT4h3QjU
q+wVoWWk3xeuYbzpO1D1ktqEAKjDFFg2TZT26KDFyYELTYIyFqizyXYpa/Lb00OJ
4Nq8/Cilg9PSzvSX8Pq+67vskwF7g3pSgwS0jZTSYPeRrAgq1SYYUZD2NZOLm93c
axiwt78SdKd//2TA+WoprtWnkhiZBCN1yxqDBMcTOkcLHuX9icygjz8MAmc9xNN7
369PtOzn19PupXRKfYtUmEhSutO+wq4cezX5C4o/SyIqASjuMeGdb7wNeNYENaC4
hD+thydtRitTWWGaxc13lEcCp/vdQA57JJZ9REGo95BzMgEp/SgdnSXxsZsZZG91
/FKsCX83jpIul3RUb7X2doFCChRAQIqnpVFDb6gi0WzyLYxMX/cvB7VvJkbq77cI
Dc19TAPKLdG8x8dqi69RqK4M6xjfCA0xNdfS90IYBCuvnB1cDMjhe1DRYbzg1pTj
MqXw4RkYmtvcBW7H2/4h8XzOzcMCiOXvD1TuJW2seK/OoxwyEqBiYyxn0gF7Z+24
8QSOMGKERvY1HalaLGwV+SMLFtDRVLXYG0pmis+RUlZeNdRNr5N1MZC8lZhg2fPn
X3NXi4Y+QePus/j0957DwourV3i2h+xsOEkU2d6BwTJUcwKH7031UvZ0/LrjVDbH
gCIApXqnAzqZQqyCQj2doD+r9H0CwrgZMXJN8XqAMzlOtHYKLB0a34+3uiXsPV4o
nqoLPDPlbWKgk6ZgAN5IziNoRgArJY8E28f2R6/2AaoZNW9eSnKzZPhM1Gt+Namd
m6wNvwjYDJpJ5nuvW0FNwIdrubinWSxoDtm2G7+RZ1jv+FYi44wGwCRHtLKs+iYp
h/3sJveGitgCTwX+cww9xbPe1t5pY5bdz0E6/T8qkDoFJJ1qPdQw7qMu1ppQbIXz
iwNWwvlgCr4KxpmyoURB7o4I2zjG6WYuz0dxnwgkm9PKURACvTUD0kbIBSPg5vOW
Gn32PgVUnyy9+JpR1O61C8TUoP8J1QUIZoeflfRgwV/ab1n93xnFKUgYG0+Q31CI
CVSdYRPt4zRXzYUgbGJyW7k+M8zhcqYPce/mnOvqVcEw37d8mvzukpimjTAjKoNF
S2X3Pny/CSpf3Op1btOyiQKTpheSchnenPWbads85kaCu+c1i6FeghDwUOCvMLeP
ty3M+cS+C5/zfhcQwZk0m48FoJuRz5kDCkVgkSutv13omdZLFTZt2WUwSwWg5fzn
H/Mzn2BhRuRywUtU+d0Tjn/zjes2Yh5AHfglxbypt8Ise7P9GfjP9ux7z4L8Up1E
EZRAs6fDEjA40OgIsnA3kBqWIHIYHK7C+O1Db6txlLl0ufc2sUj7ZsOjjV648T+w
pNnDQdk0ya8JsnNHNFURFaXNgmF/YbSDxYCUoK37C2sC3TJN/lyy+2ZgkjmbheIf
zG7atoZ14PhGnmBAFHESIplSkEjj0DnOvdQZcIxuyAGkEowAcWpda6jtLS+SgRvS
oTsxExhwgIFIebuGSxbrLiauf7grI3x0HF05IH+Js/2nSg8bdDo3dSMMkXAjvI8/
yYTsNlBsvKt1C2w0GFaBbZ/FB03G00y/W8jR3nPqJOMk0+bL8C7UUK+ecgJl2VNL
xl3QBXpxFy45cJf4RY3DrVv4y5S+59RfoJoNa3G55JYSMCp+Xh7twzsjfSFh+HqS
ssnu7LaP2GXcyTVY29sJdcomk106qiw8NaSQGGflJl7exe0H16hACltl6ni2yzfl
A7ApomPnO83EDo6hK88HE+WGCeWXjKmslfnzzx4aVjeegiErp5MoctT4AEJItkzM
WTdIBr/WIvdTX6cGoz98lVkCH0JUH5ExWe6zHipOQoAa6R61Y8hOB1WMY1BbsV9c
wO16Kb+P2y39IIUUpb0To+0LHupaaQDhDigQbKk4T1Z0/e806xS6XhclCKB/cV7J
oHFWkKVtu/o+i0leaT6pdJZmZ0+MUMeioWx+W5LD1h+TwofV1MtfsE+CQ7O6QPI5
vPeK4Zq/C3q8UQyZmwxKyEqEZA7TegBSmhKFoPR2kDZRTRvWQ9R5C2d87/cXcuzP
fxXWvmM9Q0CDumh/D1tXiBDF48YOm6Lid+Dglaa1L7RlWvuHZxfp8BCWv1YQYn2M
RmPiGswSQwO/l2622BUYYtDEv7HjIMkmw5VQ8Fsw+Q6qnye3XehayvNBNPJnmEIb
Li+annxh+sfVEUoRpZqlmIqnEDNFpIF9I1T74IM3sPdVFSs3mNY4PnPhqX0sfvDU
OW/zOPCusoUxU7rKgv/dpxkAFAe3spXEQkEc/owH8duHEgBhTKJk31U6yMgkYXJ9
RKa3PbdyygaVOfUhOWHsk4Hd4r33KyyAUiAkTEZP+znJroomaXyxwhu5iS/QQGfV
H784ky6ZBOGJXFM4/zRZtHemFqkqMWqBG/vOkway+iaPjFV7UttaO56PfWvKdy+Q
PP+go4nZnRrEv8SadRYwUGN5VNlUMAk1IJ5epHScH0QUhp3yWkCKo2RXbRv3fsdA
7O0H6HKeTfOxqDtjz4bZ8+mxI9cUM9U+oDbvl+Gkpw2aeUU8fBhqU6qNYNal2JL9
RIOQCnTeOPlmM40HIrgcVj5CoAJPcZEs48f12RMoFaThBSzITcnVSyMRAEZHEnLw
gvAM6SAiQZR/NVcd5SnDGrHU8yoP7i+XaV0hFxGxNlB5OoHjkp/W/zwOXh7w2ZC2
cV5w5TbNgj5U7YmsD7mncZDGtPPlIN7lPv4GDgXSZYG/ZWArIetPcgE/RCZ3oYnQ
Xbjn+P1KNDBBjfkMPiu+z0afM0kHN99Xp7s13mn81J5lY49EcCiWTIKvey+LNNlt
fZEMQFpJFdkCAY51mGZmouT8cqvE5SmauHPOtwoHkkLx41DsQS/H4oi2cXuRyip9
TqFqE6Kl93kYMe8lP0LCgDg00/72u8NfQcMd/RI+UgPMsMiblhFetXbzUANRICIB
gK4hrxaVxIqIZFT/tNaDq6Ot+UWChO4Z/r5x3hyoRk7jJ6TIRkRCoEaQd5hVBeuF
n892xx5MMqF+x+xBGnaO83dCcL4tOy1NOv2b/EvAIg5ymNVx/b2X2pkGnwWHmR5t
yTXtQWpp5YhHX5agTbH/r+o5XNVCfLvpOCO4xtC8vWxQ4claqsH4063JKgP2+0CW
Z9/tz9lvwZSesJLkRsFstmz61M3YR9gcnjEvdizikWQqmN2kjnAQbQmUGyfL6iF/
z56kLj664kPdqbMONmCMAza99vAAC8PrRiozkmvwysLNFBpxgwtfk/eelyrGqQbn
lw+OnMZHkCMl86JVn7fFF1dYaY6qSwyapwpQNoGnMW/eS86WqAUcvoKPu0B7fx0U
qhVbKFgIzTA4kwpV6l7WVk9kSyItlXpV501+4wQbdMVg5+tIYcJPAd9g+wb5l73F
huuiaRMey8pS+VjR4m/+XNyZK8FQqPt0ZQSOlUvBkoPibGhVVLWlXlrB73P+K2rJ
pNED6BvUH1LgygPKUflOffsu0m2bSLSrJT38uFZIsJxaXfg7DBQKhD0m3YOoJ/AL
bMn0CE4aSUi16+ygx8qednZBJ3rX8ZnsH4+aN8HdWUiVCr4rDoe3HfBeT3kf707h
nkiHd/hVRGFODQd+7t3t/Cip/V7+F9f1cTveFgG/4eZbYG06aKzmi1mXtoe9u0ke
2D5FOvDbrc5ZMwcN2BkwiDsO2SvNAUHzfuK07en0DLEKSy+R2urk/VdFVuu0DO7b
r3rcDPkM7/rkLUhoqQ2qyZwgU0dyhnYqBXkG6seLOGnPrEl8Mj+aqEt4M0YHXpzA
iW+D+PdJVwaaJQPvmARtdgl16KD91vtLXp+geaCfpcVz/PVkaPuHGBOSRl334ul5
GpVEu35XC6RydxnY0iu4vz0ERqBxhqJ5G4UJ2S6A0Vh7Lj6EjbpS39YdoBnvZw9a
hxNVqdqRDLxDsWXDED82F4BxtRBNQqYbqeImw8cR29QeInFYkTepMvwSpZPfFKTj
OdXfwHr3HxvWahyGhobhrEBKeMonZ0QrNANwckKVHBzqsl7N9rlz1AcwaSEYZQUT
MLFJle1DQM+j5PwvjnVBJD5L4Xul4L1J7Q/70JV+lQmYIerOTBM8zoItihCil0Ls
Pa+9vvJCOhgVvB6KYr2ZHVxHvVWp+4rtoJRIjbGO9BY6W3V2LXvb09NEsiD8g/RJ
9pD0TfFvz8GhyaXdpTi65M5xWaZB79SbSByoHTG5t3yHeUM8cX4dw9R5EpJinwff
vIAhGl/OHhhV+SRhXMLWrJaX63+Hs3UQNAoQlwS65wv8q5Ts1rXsp9OjDbngM4aL
/wCGapxk8ptrEMb9MRqa+zMyW/6z6W8XlDqJkMt/vX1Hc5um2YAmfZffyXzvXOAf
Efoxaai+txxpO4naplV13zxOWWgyqMxHSThwvtuwWFMsS6TOWqB7uYodN+rKC/4D
BqnsNKfsw2IIV8376G3t+Zd217J6vrJW1w9yVCx89TGHoDctujhSOEcsA+L1/QaG
VO4IfzTiriv/A7K2WAUy6ue0YNRWRfW1bhDES8UUH8mre1tk4G6hAMe4ZJzCqg01
HZQO3d3jTaBQpW4PMuD95aCYhHKZnvpVq778LLsCPRX3y1cWwr/a0IGzBjaaFPSQ
ME+bXrEZ1hGsMzPmyzNuhSCu3warBPoCc2dEfEDSSaogU5Gfcc0wp3iRqZgXSytj
sdEdS7pxgmFL/wT4Y7356S3Qg1C3liwx9c7tI4ZMq5SqYeGfJb3/uqKJ3vfkqTeq
NQ44nTw0W941DglzpuHbbX3RPipyKo3HUveCxnO/xocPPA2g1drox0Yf5UeJ0DES
gF3isTE8a/3Hz6pBNUFwintPvJzGqLaXjJ3j3Yml4z+AKA7C8oALR20qgmmb694+
mhOa5NaHTSesRvOeqqokoczRd0jtn9NSyMTN6vZDJXk0u5WbiI8pEZQKdltRsima
/FVbsdawn3GwzsGqi7C/M0Z6vSH2lUWX6nBtHMrK9Y34Z26XxaYXxXcFIcbSoIdP
aOJkcU02U1XhVMN1XZaLCZ5I3ZTc6dckyctgFQgzXDJX6wuMiQf2zFXR0kmRpoNn
BVZC4vAdX2bU2m2Ztms4SAyQQjCgfJTqZ49UygxBjKVtsFhBBcv5r8vDdrq61PSY
u7DE6PmWDAi4wnF41nZ2iWgsKaonQUJhkkhPVP7zWhmU4o1DT4GX7J1eZsABC61+
pNENwLdwCKpjQoeBae5GRbA/Z8bTQzbDXau91V8mSwPPgvl2czIn4h4KRhFZr89q
aYGCAgk9YTVQgRx6VIjQMW/wOQPRhXqGF6ragWvfLuILjs0cljsNkpW26JX3Uxnf
5T0AuPf1dMkhtaeP66IGvfBTiH/o+7PTrlJbcOKNNPAm8q8AoT+1KgUqKuMUQgy6
PF9065ZkfvFl53z1NaXtuETzsVzmg/j9uQrFtslWfnIZ+0UTmrrRdNqhjYGKWAQS
cWSh7wI51qlCVp7COtOHc9l8wwp0RyDdv8awa0lEZcz3XdL18901QFzbmYZZKGkc
ATYX1VSJaB7c/7aR2E57RYefTAx2xEYt5EkO/+S/b1Uv/PB+wlKOZKKbswMZwVvv
vG2yCh8uLdpj+GzFHL7JGYUes82A01OzfyPDS6ZHoc2ZgToduS5uanevT/uPOey8
fxL84oSOprkT5Hy+QyJQsX47kYk06dfvvwI8Kxm/RxlioSNuvqvcFKW8jr04ah01
hhKQA3wdj41ur3Zr5GqLgzlqzLmanQOtbjdp0xfuPqqIyI1zHd7q3qri3z3q8YlM
qVT6/kHt9Czm3yrI4459mTw6Art+YHZ9Y0jcoNOpDLO5vAOgtydZQGEQo788vO1o
WiXiezJeH5G+FBzq3/vdiISiEGslTuMs+a31dK0nK8HhNw5/CjeDbgkNStKSgRC3
yr1wHCc/uDy23+nXWX3QqqHlehBSc8kSK5cD+sQ8ZQOyXCWER3F8vHkrAIIHnbUI
c/mWZCwvfOugqWWbhW2QnRBKBFAKBuL1MyZKaC2sY7x2U9QRILpJF/e+EwRjtbkF
C37xs59vOMDC/CQJxJpD4X8qam51VXgk6zYoVYNwhjN7dXwgFpYx5saJW9UZI0Va
bE7JRZ0zOZxO+4WiBbmbTOhINHOWSlRUssAIxQ51yFStROQmu3do9BbjNnuIZs4f
WLJyh+dlHcApS907UuSHkvmGmNmo8rUsE7dxQbk9OAYtnu77xdz/seQmw+hZ20gB
s2mtPNsW5jKC1okVmitdO1/kpopvDaMq6iPwjgDqSsJrWW7f3FUMA29zkKS3CofH
1y/yxFSXq/x6TsX0moN0R4v/hoDlEFWafxx0l91GmzLsY8dwUIKta8TY8mwtdzV9
gsSrBdR8qYi4tre5lU2Gxx+kGkGAsHTxSOWXFqchPC84LL0vDF+uIZ8OwcFYeez6
eGKmvW/52/mxMnPvYB56mlWO6/5fERgqm5MXj5wsWG3U0EN9ayIRuZh6fBXph3aQ
VGcddO3lwMgNtSxlngIUb0sma/qldstjL4FXyx1uwchF4TqIIr74Nx0mTVMBQBRS
Q9fJcow8mF2BFsLfb0Kvq8dIcMVTb6Vso6M69A6bIZ6IpNZ3iCzyl5LsKzMwxbOP
+swig56qCm7vjdiKzRw+jH9mUveq1lM9YC5oTGBhHqkk8YZa7JWR69+Pr0v8UCFm
XmyFqxuLPS+2xtrqcuVuNnqGdEogywJL8+sIv30Dn02az0kvJqR19v+ghhM+Mrgo
m+zG6u7eP+GQq1aERIQ7wBUdo1fW8JDPxFhZwfAQDQw1UBs+BFL04QrJ4RkBViPu
ziic/KHmESXOdXe2Gas2lTLRhVSP2nsUwlPik4DhyPCuOZEUNDZBP6ElpcaRL/Zk
meSBxvBFIh1ODUZJmEQu+DA2lWNxC7Wlcn1CVmHlPpcEhqqdqhGQSnvzFClv1Dts
Wkbz+E47MQ2SQCvdHhnTS+VwN+vB1ZIUpBIb0uCgLzRDRrhS4elg3b4Hi/b7uO60
GPnKCmobMBBg9g4c19D9hTljS/k3xlNS0RNd/wEcQRiAQbo9SwsM3rE9KHkpyn8X
OnKvYgUTDY/08z6TbdIScu01eDzayvBqkfKpwvlCqnjbC9rkZhY8kzQ71kfJhYUD
87H3i7GNCIe6P0sdnzOMiLue5S2n88JhZhho5Fj3nyRmB9IWtokOtKnillaJmn8M
ZaPZZI9/+O3m2kq7ZFeFJpQ/kZro9ikExG4dkfUXYeJtYXBxD+TO7Ce0u4GaxOCU
+5JMIbk8QdFy8jXxlCETolNZxOTtJ/7y/DMu52zViZ53mkzc48hvC3UOWRqA+dRe
z9mWTtDEZrECN8OUeuljn55XF38QThosB2fJtm2oEqj7d3o40+aO7hD3SKX9Q57b
WfXyU55FWes5O9S6iDGNUJEEhW5kTBuYijarZLMk63ikr2k4lCwwODKy3fN9JIdp
EGOS3UBTIsT3BB7w+UI5kKxdUFTiFhI1Z6GRZZXKVTD9jwkFJCm64V7mVDoZNP3l
tnQILTZWfk8l8qoy3N16VfnfS0IjuihFNBl287wK3tIstWSq2QTjoBAI8sQDHjTk
Ps2COQkpEUGKuLkhu5OOGqjn0YfAtCMbKMb6YEnrblAJcq6AWQWhwxlY8fT0FCfP
HSme0QxEdWamlV4K6cFDlwXbk7RITAOSz5VFoi0mSJAtR5wVbd0OiPgHPvWkcgtR
nrGI1E3czBBe3aBPhxg6VdlFltAjdhK7HPo4ys5BfzViRstnfK42Sdu80lvF+diG
Mr/CfVnzO7fITC+0/Mn+cKypXkaX1SaIWlMhBD8EyClOkjPhlcJ1h5fTdelJMqeR
P1ofYLBaqpSYHhdEzaf7h9MDURWV6ZNHhF2cmCnbtvdjRAVKQdVwAwqUkijaJHl3
AdyO8wXMIb87BEeXHjXYvkpA67WBBx9ghB/tt59uUpBg5tHJ02vwiiIRjda4a53J
VkWPJDt3r5IeRQodaFKfFHvJz0e6paGBfMrUiHhwr0mYGBnIJrCCqrSkKX6EE4AE
fzoNGa1EaufEFpWJjl1JihzhNnRKhKZl23v+ml7h5S0EaqdT1SK4LSf2FOfu3QjT
5T+3MR/N/C3FKLQaoScdLcBrAaDUHL74Lu/bquBOidYGC0OgQMEYEgRyYBS0DSNQ
aP9sreB37IBLjGy8gaMb7u14xqOyUIRviTwvEp2FtQIUZImJJgimUXGy63dt7tiE
ZlTsdCpJdCQQ+eOkvpvufUEVBRFJNdywijU35FbLj4fg5NxvwZZTWSM+5JHcOXMR
zWQgY7P7RPwmkoXl3fzxGsx8Qwjd5jfWbKf9YhCVGLphiL43HXifmFbR92c2v+fc
LaxuxFAJknouUY64lYNYr+rA17Jf5LZRxh4yS4ScyX9JD8fm1q9PkXdEnjBMjxGA
Ngm3hUrltpPnPsy2YDO99J388MhUlqLfWVIDc1u53G/byTFSTT41lcdZR0a81Xmj
PjNK2EKDghvVJbsrS2vV1HzNLXaYL8R40gAe6PUqVQAgbw2r+MOQA2xHMW8T9GUU
Xjlxo4smW9DHft4u2BMr8QL2rGRR6l1k6XfwyNJOM74d7WTyrv9bV+r8ZIJyZ4Hz
gjdPoKgK4P1CxyLmpnFImKVSaB9poAXgusvbGPsDp6o0mQO3Wny4o9vyD180whOv
MsJxkNpCSbhvV7huPU92UNQ/cbnkn8bWQA3ME9PR4f+el4AbLehuERKCKcSCX1dx
lzvjz168Oe+jFyuJk0O4sxn9D1+UKfJIGftRFOdmD7dUz/J8xf+ZCojeGqTktClK
8x5h9WFzE262AvJd2N0AnOENX2DBlUnTbg4yc5PF2DbSK9YC8HrgyOLc9Idqk6l+
Cq6BH64vPFP8EuuRE2soZvl8dGHFMKOLSOfHwvZOKF26mi8LZkP8eNewN3vrHdUW
Uqflqj0QKnPVyDksQwoi6wzkaSbJcWacJfILn6P8vU7YQQiVlB1RkCTrkf5iyN1O
mvAZ3Xaw4PzH4sAsvaB8NarABwt0d8GCEmydDYS6adszYofHQtqWEB1YzznvOf4g
x4kSfAXCeB8swCOFnN47sVub4UtO1Aq1frbrL5W9CMrB6o4k/qg8MuNa48Gk4Knd
azauef0rxXTyB43gzI6Ivi5yw3t9FIT1zB8+mWsy696FkcYcmSQss+Ky04XQtGwb
T6FAbymVaRCkvB0/CLdwUFcnTasglvFD9/mICYr7JIP4RTgB8MlPRb8a/t0PEydN
lLjWFI+XWGMHv5efNzV0QipGbzLTIbw3mXhTj5uB+hfRqg0/vCx9tbQolMt+NbGa
G0iJFnww5/L4bikjCOmAf9SreRAYLupKbHyCntstfFYFfbAaAbUQAoYyWTucwfZU
dZgUYzNO9teN+S2dFOdPdM/WaVwUSetjC+EHey0Y6h19N2aOjQid3FFk986tro/F
2Cz8eIXMkvnczADUs0mgGO8ZKpcTQGiNEV7DmB7UmA3STWZVIEBBHpJXErzoberg
m1LXwiZir5N5JLzGgOUrKuCRsHvDTItKIPS2hiE6xqQhkwB5Dqjf/F2HM4WRe4/k
l4QlAUViCfv4qYekgWbIDdUpE/zPd42VPTB3JMp5SWK032/iEe+e/JwjUHOt8PVl
MzNGkInucSiPwYZbvn0wCZmkJU9AeRtXtaw7VbCBV1eMY2vBFlLIcfhharUuYe7o
zUPXkkWV1nA431Tq6fvr+TutG35NN3e0QNzbhhzZEeXqZp36WjPE5X/XrZYV/W8j
K/n2HSlIDzQDMtubKlqqnVMsTDLCAtn68wweWvwIu8N/iAJWpOzJdhKjoCdLBb7+
uiQIgj86JX+8vtxKUqtT5c3WL8frKOSggmtROfA4NgE3ZmaO/cOwsBwBGjM+Hgpb
J1AaKs7Swj8+okpi5rwUJOrrICtaiW0A5PcKHKQBKr0EU+S6Xjn0hiIhWI8yMx74
gA31tFoviCSLft20GTr6FnohEQju2zysiAra+N9qEYlL3rwNehxOjxqQStrEikfs
BMD/xMiCMV3ck0FmDTneI1Jbjatpii2vERyrmFq5ikJcz/VYjXq1gpLGIlzFQ/5/
G9NW2NU9mG7VjUxDONl4H0dmTZWL4FhT08rEe2yKiVm6ByMOmmSW82dRAUuaQ6vp
ZiZTis7DqWi9qgsG7LECqFCeSw3otFtMCUT84VDnYnA9Yx5t2MqEHYGIoZnnjeYA
XwiEjm5CEt7X41WIR9rsWKib6b+PX54aGoQIh0Rx0J72q5TVQ6ySCtUun8AVmgyX
Bv64lVHkpdJBbv+STAjlAL7Oyu8KDlqDmPCeCXNihW2w4fxSpfLcJ5jVVQy8ZhK5
f9NfWbYRervdkqaOEc8IAXLH8JdsRNKNGudgbMc6mQsPz99XUUpsVWZOaeChis8R
pf/ezuLXhQ2rItxuzIHKyD+smSWTLCDHqgPyqfQHBGf7iJtNVSEQiWOhX1pJ1EzK
AO1GLFztqJk/vG/siKlndo9AcP6MMsOtU4A9heN+YHH+vv7W4IqnT4TaLFXmj2eW
dyNr76HezN2iPBK/kMBrChKgcOjaZLx97ppZt/7BtZDxEIr3fesjKIOt/2fC9Ije
XU7fjqpENclfQmm1aYmAfdGUl6yYA5v7a1wBKehTgZfBxNfoSdb2SpFvim6KB9+E
avzCp5qm8gfLKeVznq2hTgWF20IkgqAoPN+dOwelxvsRphfgu0TBKnwEkZRNXav/
FM6hiAb9GmRmx8SCrb1F2Fb16e6aUxKF090lCMrEyOCYydl7wmRsgvRk6m++pvT7
Glu+lGWWmKK2nv49eJLPneDgE2CNokmJTxpcvqC6hP5Ov9oa/qL0R2XbbYnyhx/K
FUwnVtvdK4pCKvGTgc5zCY19G6vzKj/T0jtG9OevDmu2KAuLBY2Ix4CVQzKcGUf7
5EdcaFvwE6rDGadSvjLDlsp9iw/BczaRy0MBfUDgXunVepXnxGTV0v6aJkAVToUJ
78BBxGpsVI415tkZrS8Ozfqp9SnNC57VSq4H5FbZgC+AsSaEmyD81AjNgUI4ck6v
V6UxhTr0sviOSNyM31eHvH1HJdMjELEgOIDTdQ0MWp9w8TLMSK/Dw4WHFhfVhM5V
tMHtHKlsiWXUNuVxieOdnTF7yECiQaCd5gif7KzRlyk5q+FbFj/p+5a64okNgl9V
SLXmqQ1WT5a25ygrIX1WTPKb2C+pOkB+UX6x1AE6pShVODFBbPmqt6qGXQ3AAkDF
evPQpMwW7tqtLm/6Fh5icRVthIPss9qLIo5ohqjPWZUBl6dQP/KmspJ654bK39cw
s4hXtoNR5Fj+MxxO562xJ0SNZSuwRkv9AdyaGB50u8BNjhzYPbLtD/FJnH5H4a2D
DoXTCZNjCWi2Ap72lUzQ+XJFygWjiJJckB2CcopLsQ2T0jb7m4tsokS0EAy1sf0/
8X52Qwtp70Eop5tiF7yiyM7wvqYcCRXmhNqio2uSU4JDssOz/hLJcBwf7umR/lQq
smVOY1Pg+4PSqEVGKk3H/LWvFzci3tnv5AqYu7B9Wzhui+BonFXdb9CF8+U2Pgh6
GlRNjhg5j9xusc8p0eFzVQZYY2uNtzAB1Zshb9ok514nmZjF48OaTxFwJnBnroGn
zVANeI7dgkO8FVxMeYt6NyUuShnylLe7XVIcLXRLNY1KnKWKqqXHQ9DKg4eEPtSl
ioNlJwLIBzFO5V4LFj7jmgGoDUyTAC602N6sGRG2jymgheZwNzZV5i9c44Q8XVuu
a48EKuP3Zr9sNfotFUahZ8FyhRATt9wgpIaAUZbomruxF1dEmWOV/kVJr5sgyWh7
KNZqSv0b/ZQCYCHf2HB7O4076danN6BtMQtMy20iXSrXWxlJMNflEh6n5eoIaCqI
DwfMcnp96L7x6xFf8q8uAYAIspDwouxIeVocpPt9vjb33SPjx2rr30AaqmNi+G1u
3UnxL5tbaGsVQFTfJ2DKpokj782LrCHQ/6oDi9lZ9aQhcxjuI6jpjPrND3qX/0ul
N4Hr/zYCGH14CK45d22uD+xpi7nG5KkxmY+5w5xrn/O3wAAGj853ltqWxpIEfR4o
AOa57bsRA1b4Zgwy95TL6NJqo87unaMb7myfP0ELR81Pbj4cz0RJoKTzNT3QReR/
+hIEhtEY1915zpEFfkfRigtBG/G/1C2rXwMTONtSxbc6LcdPdfQT0JMjsYRvaiCX
PeKQSnASYK0sl5yeVthuQoHE2qK+LGHtEy2FJEFUY8Do+dLO55QJJWBaL5eT1NeC
x8O/DVzsN4jfaXXdM1niaz2nvRCSdbExOFv/B4/9Wi/Xvuht5p+bvCxvOeztI+gm
Np8mAukrsTipx8bz8BP4XkHhsjpWhoQfW2rII6x9T9RNJL3SCYdKCyaR1DsRimng
9SKdXiyk6+9kGhCn9R6cdZqbHUALNTCIiGUGnRZcMbu2dQfASsZVGzGpITQYcnPg
HZxhLcatuzm2TLY+UndwuKLDhkkAVp3zbZzJ1xyK9hOFJc8i+i5vSY20rcQxW+sN
6U46FH+uCHY2P0OAAr2uXEME7gPMtz7uO+B52+UejUtVi+XPSqM+gxhfDYOMUZyw
KvX6eociEdAKTMXUNuZhUYE9y395hQ5x35UWjWy5Kx1y+ANLUVpfSKKS+Eq4a22c
c1/gtfuNT0/H3Jm+JY8gS+m16sKsMrLmtWJ3b4arl7KrBTPnxIjSVOoy+s5wKU56
kiv6ld2cK6EW5Cj9+259tvp5JRLaqARKjshNWeXgOZWGchg2Pn3zz5oimm49jmS3
U7nEr8TxwNeV1bzx2SScQxBIlSfwidmsLQZgGncqiADK5CHYtGD+VSBLaBmSzya6
d1dDJkkX1MsgGLlbLxup9DCE1uCMtykQ38t32BtMngb+oR0U6c7VAK2qumRX3FRf
XgNZrWeI2XyO9h2Zfkv/d1YjVcdkXraUHK3pUjXK0OQZ/n2rZvMfm8Ti2gou76dY
FNkYq7ox7EkQ/azJnk2dkTMSyQ8Ck0ZnEwQ0r6LiD+kus+djuJIh6hVHrW27Q6zD
T6m4wOTFftiOwkFDj1WAF0htklA2mrAL63YYj0LsvjruUoIs4Qe3OXxaJtHRoWC4
PsmKi+vYJH1uRmw+9LzqeQmioxaKvPZhrYNv8h0WcPUaNx6q7AjYIrPX+jnf0GDX
oddefn8lFeehYHKannfRRm39VQnMzKqwdJqil/BVPK8eYsf8oVDGddkjbU3QNC9J
m03TMustT7oUFwyzSesdb1yFoItvK6UMAPdl7rMAglguM+YHn+QXijR20Sk2xCBy
mAAe55RFkEYB5DRGtFmc2dH0K2EvYu0XqXy73rClgaMkMGAiUyBXzijoe7EakLkG
/Aq2KDAykQ2k1rbLGZcTTBNM+pnUqLF+V9jd3iFIChSCEI7o6exOynqtr6JhnPvf
UIZuyXQM7uORzGrmcgua5pyGrvIKxTHuGNDpI8u4JMkYRpjHeHbE+w941dYFUXCd
hNRLS7jqLT0PJIDlQfzwEZAA1+ijJZbRugi58FXFhq/GRDJZ17uHpDtj4QcS+x1N
obUsfN4sM3HrMztzQceU6yI6PmpBZc4dPiCAD2RsZr6EinhuW/5V2XINxct60K6O
+RIbEJqQ3Sp4l+SCtk3a0Y4j+yc98H4qXJKUTVCVJfzWFcTBQC4Aem9AKv/xmiZM
dFzIu3mmT4QNw7Xqhynmxpr6zPfPj4EEvUaYtRPpe2AWxqDk1F9+xJzTryLdqJlW
QhxTNi3jNZTpFThTIWFP9b8GLuhgC6hDd9CDYAyeHJ0VNp4fuaOE1HO+BWWWLabH
Iu4quGyFCQ0pQRROx2eAPcLhLKa74eM7gYHJMrvQQ1LAAG4hM0jng0ucJGJZeJ3A
9gSDnSJIPGTffn4cN70Gs9ZNTUgydT2/24lwEZfjIaX40q3p8lSSeiNiABZuiGzZ
cKgYbNLcP8y5ImoMQhSKs23STML3C0IrfMiC2y8Oze64nYByZ1vFWhilocm32qpr
2cxVJBApgwrR5Z7O66hMVadAMM0krqNAoyf92JWn33ReACFKUjHff4IcqeM5KvHp
01fAt3Ta6C2XiWMPogSt7LEmrFlCMzK1BiAfT7Z+UGeLZhYf3+YlJVEbaZZZRA57
UMJC8t43se6xMeOzmwn9wo+qEgzCkoKnKNro/Qdx1OCUG5+B0cwuls+FIgPf5CNf
uNNY2L7Lg/6yvVx8RITk0kkbIPioQ8CXZq8rL5uletZmuNVxJPPH6tYtTM+c0cCA
gwI1jQSO2QZMkAtauRah3+t9Ve8eOOtoaZg22SldmJZIDMu24k3vHPCp+KOqvjIh
joj6Sn85TPBBxElz4rDS0akjP4eUHAngMv/ndFeWZkEluCjJV5FWfEEbKoAprQOl
Q8r41eEQjw00kTHo98YzKS1llH9sm9wNREbyY3vnUXwmUTB5upiQvYvOhdk3b9Aa
++arP98YL3MwWg0AYdUFy+fAAlz+77/YgruFZR/PRs9uzYohMkkUqOTXk6WfbDol
YGo32KVIt3K5hE7sG9s0sF8k7Nh4tXUwMPJoJzfoo6YlsNgZzHy1L3RTyiZ1uUNt
haEJLvzXei28iPOFPNZtCO06EZv471mmhLApKFY/Pv0wgiC63HcbpoyZM6W4QvPC
49QkwEtT+02RGXnZB5sP1du50A73uAupyM8sJ3Oo7Qr7ipBmKvFPix7ZWQbS9t3p
svw32r6VqESqiM9DQ/NApozvqCLJuS0ZxRXywsTqca1yXok2yqV3KlTsVS1gc6Z6
b5VEfwnKJ3gL1SqZPgSYaQoYldhMizS+NzyDfveYhTlQZOfXdvhPzM+ZrWbinvnp
DJwJS+fFGEYQxnTw66lilNT62Or8baz3SIwtcpvLDNzlvnAejRpKGxl8h1dKM5tz
gTE2n6DxL3fazoK9uQx5O46HH2Z96qeoK71JHDobnwZNr+RHtrZoxT7N5QVjRjpS
pQl1afe65w0XQWGdMp3xbxki2Osaayh0eNP+pPWWEYeEPmTg3n9U8z6RkjyJZKzX
ToINQ6MBVWvhoMcOMb2C9vQA6CtjWOEEjNVA2S0kRxNaXbS6SZ28rBDVQsUgP2MO
pdjQNR4BuNloJhbEE02GJywx2X3rMvtFwLxi7bIaB9LBkzWeNqQ2DSBC5wFetRYV
A5XVeWTMPYvANgmo77BxnVphm0XvAoJEE+inEVeq5joFK3qUwWk8K5uXIO2yYyTb
1FN5iT+IPAmsjAnPcyZIAVMmwKiLNOrIsFMHF9rVUeRINeW5eLsCRj8RL1MY9j52
gMtn+ZelExnWumpwKO2gZTSIj5Iedbbo9t9gDgwX0gf41lsPzk4pDxQiK2kn1g9K
waTL2T5/a7HVTlk38Z7k71M7mIfw1BQk9Wt5tpZl5n7nRxqV2kiGpFSokndPhkga
rRSg4fXort/gxsfk4sDpSfl+dClb3H9YgCY0sPML9V0jD3ut6DQZlCn9dW3+rjJY
R/CXXLwg0hdi52WziYb0JYeJNNU2/ryK25oPO8jM/e4MxSzqIVn55nG49YK26Vsy
wEtSHN0LSuAxjCBxCDYMGMusATpnpSbly4xDpXty56ilEL5L/EI/2vJHJB5Uxi2d
/un2gct/AJrkiTchkTvRsnQrs6ezQiJaCVmO1Ri53c67AjBtQp+dVnkaclMHa9AB
j+eEa+SULWhYPJvQQwQqPX87hs6jyIzdZqhbWS+6zxsJktcu/9m8vHvymsy85S7U
wz6UtwlWypWUCbP+PLXtwo9WTqObpJ1waezcDhhTu89RJ6YAvGOOLUCIop+PLbBs
Pua2Ra5QSs08j6E4ZTRmb7/3g7zgRxjOvP+PWjYSHp+Rg0kZ2wStUcxhS7e7125f
dB6yXPAr8Bu7e9186qoN0a3ix1MoyUiXSpDMEGZhUbeTYoz7sHNNwE91rZSS52pW
xjtOyUu72B/1isvxqaQVFGqqvwYevysv/XXtzq5bkCaFJIIgebG8VOTT4wdhkidv
fxiXkd8M9zq2lwY9+pxMMFzFeBEciy3/MbF+WGumPQeFpBGojkwN0RFqBPUAcpZE
84ukVVWX7GIuHuPx7oICLN+2EKtzlsHdR3SYGgPX2hiB3uOzx5BKi4Du/T++eafa
/RHiMLmuem4pfL2nMppEer7xcsWqG6o+zJz3hB0KL1WZD3AuW9sI6m+lSnulEReu
mQT2bCsTDr5qrKB3pWIP4uCbLPJDz8pE0DRRamtdMw9LFoVHOqyZ19t13hoQMA4K
bBayKMYAodypUY+aiV9y1BEZqx/Tu0bWXWL56S/o+N6qPu2pCjBQewSfguQMqV8a
8ISkCsBJzxTvN08s6rum7+ym3tleJllg1i4dQs+i55Fz6WVbsMmL4PyAZf6vtCvU
P+xxK+uTbPOE1Zza834l+bKMURK8IA9D3nYHlq2LlyZPSdFhkDW1kMpF3wmCSJ8P
DsZpkWQOiW7GWR5yab0vYzA0c8NcOavOTRyux5s6M300Wd8yuDF+y6rjo+ej4Tny
Xv7BfITz9NhlgkxSUfdGyWkv8rbB8L1BkYz7n2tzVxNO3dT/3X7YIPhqwUfC42qW
t81uGH9F8zIXNxuzfi8m5vlx08Bj4CyTnFf3ilyK8efPzbid0OFENQ7LMGGvIc1v
muhAyw2Fqhwk95Y32P+aoXkJDpGsS2UowNY4sSufk6KOk0m1C1puHN3fI9f63kJt
L33HWLVaaUpzjP9AvPyCiwOKg7W0ZhTOE4w3ZosOsTRufZGJtsm+NYK5hS9BQLM1
WS4K6GNV0pAD1PK02bz68R7izw/7su9nwKTUIrxbeRRegx9nElBuoZwEcNyz3pXq
z/XBgcaVBEtK/lsFiYgne+/uu3i3RX2yJJ5oBUXS/vOjzIylMRaycZHJGgKJjXRB
iV+qEh1mWtxMTtg6cLUkRDk7gFtHz8XIdkA2M7drjtTl2dbErspM+saVmgzyFbRY
URCOUkpUhh7ANbAiW9P90qeVuavFj/qKX8soR4tvXLbNUFfsmX95fpyVfx/0MyOZ
KdQds1tlaQao0JhzhlzkT2Z6I7Er5G5221AlTqofp/IBztqzp3mcmL6zMs1bSUvM
P00Oh4FvHtbAIVqIMaKBOOBRoMkJxVVWYTVmC34t3v1EnR8Tz3o9nHPW/9Nq4Z9m
+JMGnn5910xamYODrVJ/X+1IGTN5yBdeZgXGrvp0XBEUa5yVpFdIneD2tkj+C4kC
1KVajXXF/x5nR8BpVBnf9ocQVyRkxQy6D6MwAYGdXdCwo7PPdXrdtrHndkdWa7pg
havEYPfSGNUsH+CfAWmk7CpqCNYxC4jzCwdp/m4oG5egR7LmquSXW9tx/T5D82E9
5k0xis5PVhWymknG+emINm37YYPQ80qoWohWHCzIr/9aSFEgPlSfb2dgOzx3CfwR
Nq1mUh7srX/GCC90sHPowwJQYbbN2SXKnXxOIPYV+Fi/ZaVM5Ayxj0E8pDC3IzsY
hkGdzLQwkpfkNFZuDve26zpjv1IJl8JIFF757HCd0ChRPX67LKGxbLNBXzBamLd/
2xCV8vVwwR8LVgeaAeVmfocywpLNad5sio0kvlNrwIZU9tiSOg7QLFR5YxuBFTVQ
YDMKBPE6iOcWSCb1E490mgaMr3PRMSRMrBNwnU+cYUQc8YGc3ZxaRYgp44AANttc
KwykdH7h7nY4DdPUIkk4YakuNHaOwUgIpBhdKqu4ndFRp86QvitPDIMOjgq2mh+g
yQWFQem8hgnDVfynxVGIDM5GT5609zIK9E5Z+rSrZFF1RZAUJfYtZqzOF3k/KEM5
whVqgNuZOqWxNJ9/JAPjsTgVY0i2f9zovM7rj4Pi82p4d2LPy1WNsyCKIUECVcCw
DuKn7y4KadEHbtABZBF0c0T4acco9Ij2o23tOd1nX/S9Zs542cu13dulDkml7nZb
aswOE2QtNLVaGvI1zHVU85PsU097WMzUtqvEnT5NiqxtRCoUUUhxZZWTTtC74tbQ
WzKeLtVh663mrDpGHa0I/Toy/PdGZ28jzZoJX1LxsTzKGsDWdVsXXyia391QZa8b
PuhHeYuBGVRTL9E7RR7hB1uHAZQy84To+B8njIez8vTf7gFDtkPgkeaGysC46QEN
aUVF5v4ALN/KvqtUsPbCl7CihXmvSjtjv9Q7BZ9yNMkLukAWT3VCyKpIuE+QDKWC
O7scB3Qh9SN47W+hYTiJlu0++JkTuiLj8gPN6ZpSE+bjNXPcm+I9diDi6dDo+RYj
y9xHyVc3ajEcnz+k/0QuPl6U0+PADoCGwrt5Aqj/XfeYAVsu6t0vO5Y75npuUCfw
92lgQz6nksEbctim2QhDLyxgWYesD0Mxvp88xM5I4DJ11lMiEa3eccHKIBgP8cUr
Q3SRoRbUro30Lvl3Cby4uLuotCYmgD60O7ejlNJUDNRY+FCqzXdKyvCNw/YZdFdN
f5hTTpEhUegalonHh6/LNQqZuqy/2CONzigOMbt8OUzm2l8FFjhyYZ0siyIaYo0O
5kX9c3bRtnoboH1s3x8Q2BAGFXhf54k70aS7KgjI8oznkFNXBFEiBFKIsUcUUzG9
/qzcs6TI4jrj6BfLDbo8BeVhUEJEOnaliFaITsDtZInuV5Ph+DdYL11WdUOqg4a3
t3cQ1U2OOaXO0QtndN8sYKaAgE2kqEzZ/6GTkYBqujeVRmB4xqvLI2dunXFltnJy
7GBnIThCE6JPvbsDrRXQZY8f5gREQSDX8GSpgaG9M5Ai+IMByYF75UUE3lsh045D
VkRLx6Fq3flIjWudwxq4FFF5sx6yTW8/YLYY8ZofbrS4wgneMlcSXmIjk/c6KaRE
YaGqX67cblZb2uv8tnDhVIp3H7+Ecn6YmzHLrKI6jxZU/T+VXKw9OTe7lkrDjNSH
pA7HO8Zjo15MbsDTH/r9VtzyHqr9LjVjdnmHKJTXf0Yn2bjV569LN8GIS7PpTHm1
L6jjMwFRXkSWXeukOtH4qgaRy2sw2DS1ocdutZYnHM/N5XRTlQfcLC7GOAf8YsV4
gAuc8STxJTMb1CtusFMC/SXzCutrh50jBwm2zlKBBj5TLs9MDDSR6dFy5d3Zl/JN
LO9bTrTY93brxuxB1TfKi46IsI2Y2nusCRqr5ZFPGzu+6g832tMbOD70DDYljCZp
qGR71Amk4hYe2IP2oKPIbfwdi1/VPIrjo4qQ3I/rziin72jLo3+qN9v58VFMqozf
AItZj4uUe7MhjCF+ennYnXBh7tl5XmeVJ9LsSgknxS5ygT4A5bEF6zsaHtxeLbeB
y2MDjhDNHZQHDKEPfSVHR1PEC/2mJCW0HWZL852QiEB5+0iNf63hI5s6CMT82UBM
nSV2wGHxMxCKHxppmnMmZg6+BhKo8NlQyew1X/SrTvXb4ZkLifae2UGJy/6kIkxo
EZ1haPEiCbu69ZXnNjl8RKopa1QpOezU+KiOBmcFSayTrggwUR+lqYHWOaQtDmvd
+VYIccrMhM3K+OQJfqCVDAwhS/bLzAXrD5qH1huznB+m9uqAgqMo6YqlH8QxhHVV
TCztauqD/cPYuToPim+NJh6ugPsWhuI3ZldlU1/UPI+4IbbsmpYejwrZxzdnO9lV
fXhrzzJPi/K/CRTY7rU1wBrft4TBCnbpUSXWQE8hkBeU5+wlz6+vHYd88at0Y0f7
UCWbN8rZCbCXmLTAgvZfNdFm+EEfmPSy5gaV5nPB/6aEyKheL9NxdFxbykTwE5D5
5+3z8I3/9dL+C8ux2NdSD4rxOBuoRuH003CqNYvB8uiKz0YQlpQRD8mA3sa6xl25
QApT8l6EA3NAAx+kNCqEliVvMsVx1szQoMsPkxRAKDFygZoTA8NwOTOzU/LKPWvs
QrCr8FIKQ1W05pxor1H+DIPF3JdmK9DnMusLsVbG/vWTeTbAuQfQ67odGE3DQaZR
PRgx0rLAfI05OSggZxEP92IfSkHQfgCYnQIbXq6iXDqcQm7kTb5Z87BnLb0cCfwf
6zTvBthLKnFUqV+/B5EF+AD4ss3ZCE2P6YU0DV1Tpiy7N+oQrByn3LkhbRLOId+S
t4j2CkY4bNoKWjGfvkUUAotVk+T+wYrSbhB2DQdHa7QRj4sCQkPuEaILTxWZe0lo
eUZ6/AWn3NE7Tyk8aVQK8Dz4nCav6lXng45AOxJHsSQuLCfuVa+ApjzFMu+HCeC/
n8Y8to0vC3dcm2ZmEORlH3XFBVvpHREb5w4Q/YHn5Kd7Gm7xPH8oH2ipS3l5XzQk
bY91QL15vUvwPfmdP0vtWYoXC9xcBwirbcqur6erzKWxnh/meL86m+AA+eQTcHBW
zsfYfF8DDwA5n0rF/tTVywgDNpGcjPFCkUiR5gSRUuumeiKLpexkN8MBYBbwGXMh
EZ8xjpWaTKfnUT0WMKH0WWwCRpbzhOYBbr5E2WJ6bSgF4PMg84IdbGS9ABK5GoOx
OiRxYPTAuxEUq0mCbMJbJuwIip6KbY9FiZheayWqgKc/aR1VlwokUL3rNqf9Z+8c
h3ZzlsBxPlDf26ht3op6AjUOQgV2WdDZe2Bk8QNoz1EYURVIufXdB1/OKB7oaf9l
4lpKd9yOTvFRDbVHs1QGjU5x1j4wMMKc0Hz/XA9bD4HBOc6WU2EBPeDZZ7lwlktc
e+AqTyyE++4LwDL9rxBctcjB3PIyzn54eoICL/5dGXxiwzbpHEL3mYZii2vA3EXV
SjLYfb4f2yrWEfEBZx+D10yo7pMAT5WCU36ASvjk+Ii6Vw2Qx6eoSDp8aAVbXD2r
X4NAKkBqe1zStn885KQGxVIfzzK/7cm26a+Fj90WkyYg67YY2vOAeVv0EKtfra8i
dq+iaepESBtc3q6Sk0YO2mlUu05ussKDUhw7pi28wohhIVIfM6rDaUSY89E1hBUZ
bf4AlRSp9Pb50O51YpoIvNW021L5q7x4Gj6E1sXIOxxsPNXeifePmSMlxMJrLbOk
RYgZ/bu4fc95OGAN8TO5748ySToH9SyMNEUEnDFLIqAm9wmZYgCRJrd/07+czqDJ
3x+0jRFNExCD0d24e377FMcU1mgkymGw1CUyfzk22JbDlw5jRKWWTIciBLX24p1l
9ep6tE2y7bz1SAmNND8qHPrzpLme93oo+UcRvMtkPhFd85ejgCA4874I9wxCFV+o
dkwD0rxHC9A+kmPwq1gQzsoi4r+ZBRNXhtPEWQPPe/UtYB+OIoKmSKMq+VWCdmTg
l0U5qnIp7r5HIEZgW2kZEOljjc3tcT1NMe/4xEQNfx7sXOsYoPB22ha+xrxPRRpY
0309m2fbKth/D1Wt91P4MHpRljke5Am5iM/d2zNG1QW4L6oJ6CuydpsSUN3AIpWV
SC5up9U3PWrkZw0106Fd4zl0k3WBfixNe0+hFm58tb07seHSGTNvo0o0bqSAPtq0
Hu5faUGmVwBlfqbNeujhCXC6Lfaa8eWXgjgEmBIbsW87pgXkWn0K651xlcFrBmEz
HrCv6zGM0TZrt7Pj5GOThBkAreAlr58jZP8iEiM3fv/FPJcfYoOco5VMxuk/VUfo
T7WkH/jq2nl0mLhwbGRJjWOqy2nXCx9zTUILZeRA5b1qogdXjkk00MET41zmeY28
x00ZT1sophqWb9xMVK2Aa/5djW51v3zgV1ljHn22F/0/8IG66NpvXK47AZPsmH0e
HWLAkcREp4C4XZhqQKX2/rFAGJbpmix4Vf+gZwN0QfOAtUjztDC7/mjYP5YLmSIv
vS/u0oIovyO99bkwooZ5/3bivFJ7kDWSMSz1ljlBId+T500Ie2b8uD9CfsiFxnvG
owudKZEHC89JH+qykxxEbu0P3/aYG6YgZaa45TmeXSsJibWWI3eQ7IqhiK1TlcyE
6mmFPZFSL+QYSrijNfAoBkhviHgEHSPCQEq9ohljiqtoPAbKmGDZaBpxRoy2GFk5
JSrBtN/b7A3qFfXr1IsEaYLkfbAa++ylXNJQj//4mFYCYeg8SwHOWNU5Aj7cn56H
l060zuRO6nrCQA5t2nUQunD/VDIeFPyFK0DwwvYq0pI6e8OS7Y+4i9HUAKTzN4RA
rJgbath28egOC4kO/txVi6DRpzAwYXpT6m55hMehMyrJkmSP0O9qNfb83e8Llyxl
ZRItA0s+iYg0KEPkfaNSKq6gPJg+GGc1p1kxxo9KoUjuYXCararLDKvYCwh1ZOsZ
ZrzWMGFfUBqUJENVoaOxGC3WgjTbBzHFKdOW+/HNhWAPhcGY9hzXtZhAif0WIqm0
FP7Ecv6B38CoOlKgIFQLgHwsItXie6zILAPbpVuqgx43cdf7fhxscamgmPZ4P4jA
DFIxKgVXZRTL9D7L8rKF9EbnoXKSoDdPnVRLwrKsMrKI3N4PJGphS1XX1SKQFlyr
YYPfJAeZaY/lSVp/F7xLjrKURb5jVocZP8R0BOE1PCHkY6skrD2XENSk9H2wXou8
vRUqqcLxC31Mmyo7anaLQ9BFrJB9+TYbg3M5Fo7lOy9exSjkM1z3dqPzC3UdENd4
otHAfZlboGHRsGOm8JVDGTozrFUXtJxl2NW0XsLMVvNah7KG5HrzJ1KcfUQlGog7
l/JhgmKP7HOVA4EHUC10/nTmlvY5mcGbl8xvgUS/C9Z1nsKeZbtqld+H4jFGJjsA
K0eAmjQ35VOKC7NtqziBE70vY2sRIG6YQGhOJNlkxPlP7RQpWTuSj6Ve6nX9MFug
cjO/r23Dprh1y32Cr56syoNnNv4UwfZZnCBPGTpVZBHr8BzRHXEIQYOEB//fU3r9
Tepacri33AhhcwMC6He3jZpmooOGLhUi/21IPBWZNppj20UYRiy5IGr9Gh2WdG3C
pHOZIPG2joRphcOVAsoCTnhmL1e+fek57skrzCK1bBCpMfoK7Oi8RrB+8ESqZbXo
AyPJsUFLQFHK+D7cgNvSaBfO4oFdi3YM9uJCGqI4hPrc6q/3eYrKitSVe9ULg+S6
WdsbcG1fF44C29sRbI+S2qzL7cm2ZwNrb1WYvNGfxnv4Yb8WykIvGbA/vl6vKJFC
/1rhzo5qeEdf1dD07nQ1vDNme0GQ4w5qHTmjBJ1doqJvnAKRREobcvmAhZs59NUR
hVi5dVMeRbLDoEraO+4yBuiROUYt23zszzo8ogCwJViKpUqy7/hYU/snS+585OfP
LFXIwVUE+0aZY70kK6ELUq+GujWjt2k+foinqJN7N4O31nYDJBA0rBNFwesJJOlR
Af+F1uIPEfqfwk0pGPKyuSIAiYlWWUj+hcFVvEkwUWy+8G8ez6CWNZYKUFUjI85t
n1U5iYEKb6SioGybuN7b7NecWtGWdqyqwVuxyVzA8VtuFTU6HmO3zpVr1fQQjrv8
SWd4+x2b3TN667icNEP8wSmuYJbEPNNf/aYGnCt4lXaA8IiO+n+S4DklREKb7tm6
zyxQ5Hemtr2N5fGGoTqqOoROpjCmXa82ebmDv077uHOMznuP0IMqq1xVpX1Ucgp9
1EW5L1M1VCGoXgANt+ZHzopVdfGtkezP657tVNR04Trhv9mszU7gem/LIa35nP3d
p/uUMqG1KE6NnPS2OpXC6JAdgVE1QATL61yh6vOZmtGSDLQqRHQAA/T/2hHHJhza
yVWObtB++kjX10znH7B9bu6jTcqE+hDla/s0/lVt74lIlTR8YvFhsnCU/L0O0x8p
GtxOAxvNT9KXKSe6etxzphhJQh12CJx2AVZVp59jgXM8dCVnSOQ/7n7FE1a+kidN
fDaPb9xBwebUqfBsROBa0DrGtLmX+QwcWSLhfU8GVNrmsggJBKdFfygT8P+FfDND
fxF+bHN8rOEPFk7nS10gH4o+dFiKKmJpt2fZWI4ZTUSxUi9mRxKlBoTcEtqACnfU
JFy1K/3Z1HZ4rPzP+4AAK811mIeJlbeIkl0/enEyYuAFX/PQxqqNP/vh0UyGUsQ2
rJ+KIpxtIgHEr0brjCZfE7F8Ry/aryRAoNUiLj1xgqCZg8onjBhrWs35n2mKOEYH
/32aER8J0h0L7Jt1fYoBmUir3H2sF7RYeYvd0HdmFCII4P1W54u6pNj2T9pVH7Qf
wvPn4Ye0YtNIdMEhZ80hGn0YQaW40Timc8wUE/etj36Ekc6wbfzi4MjVEaa0x08J
0DjVGHiHHUwa/KOaQCwg2P6EtQXPO4C3FGIx4+3q/ZFWkLAdW8Yb8+xOD/VZO1eR
35KAs5L1PPCcM+mM1o501APBjCH8QxSKLimmwjHCw1OH+T4pyl/92LL5a4flEeAb
lK7D4syNnf03X7j/3f57lB5AgYF5f+F7lmDC+vEb01jKWDQKAOMqKo2HADlT7mfN
3VnX0u0q75HPkB1Kv72aYQfiZ2cIsRxKQY90DjO9agdgzR3mu4MiJd5BaQfbqXU0
u3cUdrOCLe0Dx/fEyV2bK6CbtEIJUC+9t6ZfJvT/bcswZqazlqb4Qa74XXCeaPnP
DIpLRX3rwwJHSeBezoGG2WbkA7qATQnQvhHrLDjjlEfil1pqxOFovREA8y71MUU4
/iYgofanZO9B5wfJfL2pxGO/epDLujC4p9KNuxmkorjXTR/2fGyNeB5/av0OtBho
gjd8AqxymltmmWFyjAbnPGBiUpRtYtAnMDcVnhjQ9aAjzCc2gioPnUCnUsdhgNgl
GzInoKdio2OwFu5u91Hi5Rk00pHGpVzxj5/1E1jXSVAGRBTCelx5xTkoDlFLOmqI
n703g5a9Vw8gdU10DZb4soHykD9d34BTTfdnTDlpCwKJ/+ln+WGCCdbcOH+zHm4S
FNRTCx+tuRuhP3saNymlQk8/xnvFI/cskXvlQLfo2VNuILm/9Rb5UUymgNAwJszo
tjFGS//CaQRmLE/UQI+SRk5olsINv0PMH14+qTT9l1Xb608XHjffqkdtJwCx+jfK
LeGFgEPWt1y/SeLF/JtB8KLWRNXPCSamMMcmrb8a20ZbgoEr2qqUKKLXDnu1z6uz
Qj5AFX6tzU4mB8OlrvSCXNboktmNWfMgco91T5ujPtxOqhOQRiQHOYL0FkBfaUrB
OGsltPSXARnh9LepH96AqCzxyCG5+SQUbL0JeS0dX4GxEYXHG+E/HWH+EruGjr5Y
6rvPMC6saAaYSC7OP3jHeKXjiljJzfGu14AQ2htzq+MnksaFsosnShPB0obPUOg6
FvwqdCkzcCWQtfbMk6mMO0RnEClDwakp67LZGheWuAhq/9UOu3twRU8LZE291O09
EtUUT+6JrL6BX2hVEoLmfGT+ISGwDlSdVnQkIVhZ9msbc0Tx95VK8ix2rDpH0DND
Co3ghex9lN5Zz0nZsLVTrlvTucgX6ELpGDeBXXITsOMQHFzTXn1vxF7UWfiWZv/o
BLPBLOe1zhkNHY/eMwDo6yhkjHfJ1FaWbd73jU8tBHuBLd6EqvZEWRdE9Y9dLVrs
fXPGly6CKV8W9grUDjXoJGckadONw2ANa8rSU+ySCKUWXwSgX5sFGKwI4W5DpFhe
wapu6al/ZXpYx79KHBSzdf6h5urkPnC1Jod3pA5oKdDvXtXjMQNOFu8fnSvXuZAx
6clYexkHyo7HsD+BGvzGCFX3bW2a+UINPv4tzTDzWhDLwHgWr3ybVpuA8tNnH6Gj
roH3lO8qcmj0+4YCBCiSrWA4TyGferqUOs6FZ5EhLG4hD1NwQaV4E/yq7UO81Baa
S9Cvd96HLdlTJhrtRa8MXdzMSnvbBMXDtamFV7L3MfeGcdjFuJCSg9XyWrbuioI/
ohzxiYLjMAXhaJXg9pK6AFTZz2ZNJtz+mnWwUNjPeo8l4JQ1hgYe4THyvUAFDFQu
689fdZ1T/MdWlmXLstLJEevagZ+WUyzZ3sdf2pS8wbAVDl8W7zRceForBlI01UE/
Whe4SS97mQ4r1Eweagtnf5esN1LPnBYQwKKviNKwzCwBMNMPIwZWQhwuEDDhbXvZ
Qh9H33lrlvnTEjNj11edmuQLgnpD5GLAuGsDU+B2uul2cl6wT5u9oi2i6BDb+QMJ
Gh5luBDXGycqAgcyN+YGVio3U1UsBonW5r4ByravO/B2v/aALc0wXK7Mr4aZq4Kr
Ehf0AgS+ygFgqwKKNkFTJwBtv2o9rXR0sr+g7GepSzhb8excSXMTLXGJY8t9jKSO
cd9JRy6VxPlGl0WorcVp0DDKbO8u9kciwsgWsd3QDuMH9WpnxY3WUuaFHbOe4Kgx
2xkDraMkC1ZVrWeMMg5tWvxmro+IXjRQI04lbBC9nVmgV8ry4GMdH+oIWlIt2wHF
XOrFrmSsgJ9t0idUk9Noh6XfSdQwy1hvBDdfCaYCXCLXEJyPtO+cR1z/A8UikQk5
NqEc44iFwYK3gMG4l/eEPq0khL1Hc1ZuXtfciSa66BSyByYySFJ73l8Bptkte5nl
Ht6HOT/ON80cfdB2RSXXki65pQ96o78tJwuNKGFZWgKAYwTdboguMi2M9hAbN3gG
FKVTttyM0IeFLeHCZ8GSpH0Rk1CaixB7UDsr9YV66TLW3Iw/SRZwevTDX5cF7UnH
TwY2QMrR81BU5FG9vYJmJV92NVhnLt5gbMCsLg6Wou6gkntW5BGcMBMiF0zz4iAw
mrqVBUlGz5U7fEYxf9J+ILZUBAkP5gL5KWfL5URpMXwOLKlEeJa50V5UXMIz3ItP
rjeLJpn1JEoq6epUrrP5PQ4cDzhA5Hc2vOIeZYnnWX9uDvcQAWGQklkUBVxxhyEf
CEniD3ljzjkwFHjz/w//mtqbVsTh8EpdY5zOP4GKpgnExzA7oTHQwQv7+Dw1hxNp
BbA021aZAvoMf4vxyz6aQ3XqZIzJhYHL6eul5C6UxRDR8vqc/hoM/vnJiOFiviBy
hvYdV3Ga+neClUWSKn3tNcGA91vm7HMIKrAWoyvT0O0ovW1J9fQR/8W9GAjFg3Sy
R/MocvAruPdQp8wNG7IfDxjB9S/u/gcm7VnxuXhRQO+2dJJTtR5nxGGtRtYzet90
Kq/eGpmiEtIjvd+4mGZ2fGsYcdqtIUyWWhP6GtCT1ak1u8QNjhWyqUyGfsrizyLf
3Da/sAwcU4XUiE+3BocUhpI9YxMhg/IhbG+0L6IBE30217mKry5zVHjKFu8rEyDC
p/bqop1uLbkfjY5y8wQpS1LUCXECc3fuVp3t3MibSNjifvP+iHtR9VAOQXKvgC04
9YKRkCwbf9dAsctRwOn3vAweJy7QCznj+uar/b1TkqC0Bt89K2o/cPuj22ga3C93
GsmwnAhzza/oiTWvoBk0XkYgd0Ubv0K2a9RqY2FswGczjKhCIGIt1sHYZxm0wdRz
HZNlBKOF8+MiK+VlGtkDNebfT6cL1Sg9iZ6XGzQlMUJLSZ+Lf4WLryeav4pkr1BH
7VcfU2CivvDb7YXUEQJFivHzL4npxOrPai26SkiFAS5iYjy6kwSft5uXA+IZWRNn
4NaxDWnleoU04nR1PBuGoNLVpk+29xS17tRr2YiLtuWKbYDgxf9VqXQeBg/vwat8
y6Ad8vANJK4nkZ0XemkHgFt9aMDzCtryd7wswyCruDzIbdAOiegHZa7jSK9i2GvO
a/Pr5bCfND54k5TbmJw2FqoLEzk9vsuKz8uJfeeRDZyOjE2UjI308AmmhMxhqO0k
fysj8JpVerpuwcSWcuTPxxEdj2kKREe1oQfJMTKlZ8UeIc9v+GgZgsRQmI9jr8Ez
yIp29XWJqlGPvbNyEHxL/wfeSQulPd72o/0JoY78ihGPXihYXa9IIqYOThSMdjsz
uEFCFyR3eI4sXcHxu9K5u32eluPdpIKeCC4+S3k4sU7xTGRLibLIWb/1XrjNavrJ
NdwJfTT9igyK+WWaq24rLOgLrr4w7mAuHbArcGlLyXqJhkgwK38W367L0/po1JLi
XRnl7qMZX2xo5L9xQxHI7SggMdaBrAAUTyuPS5/Z/ljK7Zeu+kov20D/S9rYwuPI
CWT8B2Ip01xrC1H5yHoRv7cjkTEw/Z8/VO9WCkEhqgH2fKMqDNug0OCEDvWk01Ny
8RMfSS3SIDF5eh6CNnTYtweBu1CuM7cPO+J7JhoE4zHsDcHAIhvR8G0ehydTa5wG
ggzYPtGzsrW98c9aFBAyRL775JbZy6te7oJ0Ce20lSDHhFoefZ4ra+kWj5zUSWOC
yAW+hadsuYV5W6OqSImEUCRn4SNFO8AFKuuJi6NNN/RVvvaih6oPUCmvUoSt0/l+
WbEcrfy9Led4Q/7FsrEdkfhbssFs4RFo3U73p+5h4iJx44cuowA4pFRcHJLRtDQm
qMEFvSVaO2cPqbPdXrsOXZYdSCwu2R26K+qqL7lpHEs2i/goZOaSznxUaRWAh8kX
WMrdflY/OlZjrnbaQSH05O86QM+WFRdUED5Sbz4QopiTcf5hm0VBCcuv3n2WwT/n
uT6Q8y2KWg1mdxfVHnxYNEUC7W5W7/R+O3H6jQSz1Dr4tp4Pq6JQ/1pAPMp2Fm6M
/rhhrkLlwWaaNk6V6KjEf8X8Pdhy0NLaeZ34z9TRl7OBG6Eqy5lNKckY0ne7brtu
i5CBu8Px+AuQhDrogynwkp82W8bBx3ng+BRdWMcjbN9bMUarGK12AiTj2Hr9PQ0Z
yJES3PBHo66YGj0dfNpcbrquvzth6kcjfLuUG1vg4CyEjWystFy/ZKoly940YLhF
BKMBpk8Ip2BQu4da0idgYXP04Mj9N9Ny+vx9MWuQ09BfzVu8iEEgTPKp4MQ81SX3
n/GhjGiyWkz3ePNoaSLB03TkwdeISu4PBIiMgKBHgmHVw2NmZs+eY7tFMHeoUB/f
I5vCf4bIvyh/tAp0ZuC62Y37AWbZRcuQUzUYUXVRc4XvxKqWWuAjiqhOo39i7Omm
I0evCzOKKpi7slOSJjcx+BEJLXMKJuWBzp/+vAXlikjUMUH2Rim4KXSrEE02rVN9
McEyvMZoCA6S5QmjNzJlHIZguc90E5zy9qhORxNNK+jnzTKxXuEcuhGHoltNHNt6
ff8XqTOXetzJWCMrHM//RKSzBaeLCQqVQrKF3/cJVHVnNqkdHQMezslt2iAr+SGF
Zwt6HwvVvregSZPDjHwniTK3eJqFlfl8Fy6RhjiWSjMvQ4quGSHBUf9mRqzGR2s1
VsP4yN51oCChoxnj5qgLvS5eiss2VFgdnbtpPLpHiPITXco7g10qJ2y+jSfYDFBH
ufMWL8cJ20VTFvAlYx0DimBsFyHAHCdQwa5Ef/IRJSbn6iV/Wn90GCcDyohD36dZ
n4ZUIGpTtsjUJO0VG2VwdpfSZBXzMf7h6rHtqXXzBbG6EIKq25Bt19qN9v/fBos3
I5D01SpZICJqAiKwcOsPVukwU5ih7G1Y2rnAuTQfq2Qe7AzwrvJlHaXQEifMd1Rp
nI19fuKTLHLMPZuo3+dGqcHrS7OjyGFFGpCILFndUDZc9pmAJ7XcoeraNJZSR2zW
IxoZ3rqEAC7qPutcfchtCdiTqmkyL/pOxncYog1lwFwVxXunLcG3JzGz4ruEGJwm
I/CvbpZXumJkmlrLfvOH9KG3ndjgC6hV/CWuOr+2nv2t5kyUHkw7a+Wv6HU+X3Pq
Y+bSQbaVNS4NLCpMK2Zj/cdCzVsFEwc3osjYoB5Mrh0p/TeJweZk3K/DCwOFYpAs
8SHMRCWpOEK33AMH0dtbEK0cfxektk9ngo5SlTGaQd87yr/msmHO1+IBsUT9j7fv
EkFq8zXy3CCGLT/+GBWV3K83+aDV83+7QVuvVI3yTJ33hdK2jaRdEfZC5H0MvXjB
L0RajblzQoOC6mjQKhDgWfNKjFN/T0Pg50YwGeu2yNg5Ytei6Soth5s5/RRG+A/w
9WDRcDDIN9MzqP69uGXKwNO1HPpXnP8UUbMReRYBSpmXJ9C6OySMDbdAq6Xzj66a
ZSmja2BW7YNEGxsY/6wWqoaKVz8REt2FezXSoZF/Aceug7Gg34UVl66Fh9kQ84rK
k5VNzwgecwnFa77Zk8GAUhW6kyzaNewqnl8QTbVvf13vu/eQpR/4RubWM14TwbDd
Xjb0Od3sPYw9hFSDR/+Fn9jvVr1hQ+r7veXV5nBRBtwnP2UBlsWBBXXBJdQSaPDG
kdtrtDtQrbL+SHb0Okd2aMzw+58jPshe6scMnmtLF+z+FN7NastD28HZKHH8KcU0
6uGsw9vYKhGZG+PIuqbVlxRmuO4UWP9WaoD/L8NJd5erXxTqjnem23V+q+Aobt7G
sUMP4zw5KQujdi7pSmnKgBTYgN+/BO3WIBXmrhizhMtT1kD7t/hEUDN5E2gVg+yN
Fdkb8GeUDzuz4th84gZOtS56lp6eVk7Zex+6ZMURQS2iqOqcAPee9YLiHZVS81ny
U9p8AkEsWT4rtwpOLrHT0IxtyqfM0xUsCZNZrf1AUwNTFcTOHUob54Dk/VDnQoan
vyeq938leWt6g4rAEhSOrjYoCwDI+RKaxhbt4Wdh7NLqZgF84UCiDbQGDyOfHE7P
J+jWm3DGVAXWBRGPyUbBWNtj4/rH9uKpcVgBw4/aS0k3w+paKLwnnBAt1pAuYLs/
ONqb0hbtm04onepACLuHuSffHURyTCkx2kcTeBzDCJPz/j0vdSag/jYcxHTduHVr
rEw+7VagyXxK0/WGaTmbLGX0JGvV2IuHv5DgX3+8RXxlABkhqWqGsb5EWvBMPvsQ
JU2VQXZMfS35HiB+wqlZigbj/RitXb3t0Bh/Bb91OS7bFHiu1Mv/C7b+89PrepjL
yEXYJ81FUJuB47KxT4ADSTDQL8caKor5q4psKULb9J9rJOh5H6aj+9Y46sXXpLtS
PNEUrICeF+45l5soXQjXMeefuoUf54jw5gyJXIBI32IdWHLoswA3Xd2qxrQoMBm/
aLDQR5uxbKaIPK3mI8wLJU5whPJfCEaf7KeZvoC1+Rt0VnjCevR9HTePZb4VBzSO
F2mFeLtVtZXa36fbeZxeIDWqFoFA9e+G2nKSnGrQaBpC/SZiwR4RN2x3KvswaYcM
8d6nhVqG4qUMeVpdmET09DKcpFoSbkRgESalmUd5oRoD+VOf8F67JjIPGbDPpu4N
CUWHoMeIybs+qsRkqywr4taSGbRm1HOjFfDjbBrGsjOnWFvjHdysPkDmc2oN/VNn
lN2RrH47tK/4734UYzNvQhWjN1v+6kaKedgqcMD5UXmQHWHVLUf1q+rN1WQBPmfn
s+gzPQbTLdFX4ThLVWAmrT6Y9H5CBqWf7Y1jXbcGKI5doBzFSGER5Vt7zRzcnDKa
01lP+Jvq1S5ZhsNzG9ccVp5YE39/9oaDkxjnXfhRdy8sf6pKpUNnSqRfwgbazLgn
+YIdyQcJJdxWXGTKLlxIwbu7PYcISE36ieqK8bRc64sUHsKQRB4z/g/93aOUkMDj
d10Q55R/9tOps5mZyu9jkcDdIITW0UXEwQV7/uVQlM38qlLHa4FYK79l0ky8FRwy
wbQH8HKZ1iEIuG7oboPnaM4CQxQ0V6m8q9ze+CjxU914NeQYf8nEWt+u3cxZp+9W
RRIIH3xQpgz/3gk8VP24xUwt+yZdV7fGFd/hWu1XmTs8DXN+NQ+bmHMIiAz7p+N6
VYda1BtGc6B4SzoAgFtMjDZfeq4zSU+FxbinfsGnzGO4zHe0ZijuxzV6n1wougNV
B82aSllJLnUsbBtBuAm7yM6c8LZmUYuc38XOCASvB+1GE+cgrwWxpdX4PRxPimw9
Aw/3PC1Fse6V7oYImlqUnwemwK5DNyRDGfTsXe+11tzLkWpSckGtNQ3QFtHLw7bd
xvgjNxZiTPiv3J75dqPMzd/avQKEnaFum6CvJWyDQhzWHg5O6jMxoBOACxCdkPcU
YAJVEGIzL2trLNOXv2vmj1pId+ohv+cKrbcoRti8P6tpxOt39ODkYD1r7Nt6wSvh
M8KN1AnlyzNQIUxxPGP+Z7lOAzyM2N08pgu/i5zprfygXWWtG/fDiWFfopI6i/Zh
BxwIrQIj/lYWd1PyS8i6CO1ucjkLrO/9yC8l1MVMicCVhHf1vQY78oIKBVo5BHsV
WsI9LH/hjAqRA8rhKE0mS/jeCpwBzZPQJC1TAx1/jycnwHyaE3At/mcE2cWbHDCd
T6gntFNQ2/sFt7Bs/Lk46Q5t8UjS1AovNHJ3WKIME5VYsVP7Nr/eO4mVkR492nfZ
3hpxRayp5V5DXYtyRss0LzLr9/m02lv8B1pQ1ygeyWS4t9gulDHI52wN2VGRf0+1
+xn+VivWfurrzw4aQXc2XIEJRlnZu7J7Lg1tJPe3P3a+Jj2lp0tG7oHv/87ja3Kx
Q8n9iRRf4FRqlNuOAWTlTn2YDuHQXU2npcB0TQzcacDZhnUpldj1h3gBheFUseol
t1gAKmC6ZaQacNIkrb/hJkG5zpOmCL2vKdwKCW3jdN12r97hf+CpQUdRvupjOsr/
Rvl4vIHvJz/3Kczx6/G8/DIHfqYHSaQI3l5DdcF9l0IFnA3AijrmobyXIT7TFYA/
Cf3KMDqce4pyWWKFsTyC1NoChByPykG+D1PcdIW8u2YhPYzfCrE05oTYcsKI8D1s
9fIVjx5KwOrmZgMHYWC/F+FgqGqVwHP9Wx/aLODtYfp03kvNyl8IRKSYQzR/57M2
Qn/yheKDV27cUCRILNERNOni1ybbXUs0KlyXxE+ZdzJIp1D2UBg6B8ZTRm9QVWo4
ome5Upab0AiOtwl6TQbKHPK+Pl+SDdlUEaoB0lQGIa8uq2Rn4x8/9Cu/R908qGLg
hh4MRdvZQIv85Z4NaqFkeWZSgAy9TyAM4Dr9WxMpRJaU9Eqk1gHLjD5zzvgv/HkX
rvcoahP6fs0+UpyKFto+AQ0pQ3OJHA4QE1LlJMpqI4F/sLPF7xD1wBoxsIRPe/FH
rqXN/CA3AZpBmCZRbwMkffjg+gjWJ47y7q6oiT33iajcC5idy1edZ6dkNyKOkRnE
hdJThtHaO3nMQpT5F3Smdoal15GSRDPL4qK4DPFRQ7itly9sPjbOuKdav2sZcKFV
9xUbHsHoZzTgS0OEbL/OLrrNVDUrX9JsSL7Y1NlWi6neswjOL/Va2UEdrL8rTk4M
oAwSztZMQtjpaOdqVmBvQc2UMuwDW9yv1rW87SdID/gUZMmPzFrHYQA+I//VPXMz
v4LH4Cl2eqbF/pl4l1DpxCBkyi6Th1tpQEh1CbhansK3zajJ7kcnqgDTsWJopLe5
gQEYPuCcH/bugq8swz5f9oHZ8qOdvxNCPPb/E4gUQLVkn6E/ZkU52vTp0/B1ocnw
Zyw8fv+qK9V4URJmbK7MyEe4XyVnEL4V4GhWJ4VKgV3AA+ueip5k6KwptHcD3NsZ
G5BdAebs7aBnK3OJsIWbFNBU/+l8IDIwxAg+xQ2myIgbjK1JygMfD4iVOP68CMJ1
/PM4bOJ4ICxE5cxYM/wgWBoqDGQviaoyxTqIyxnXqDqVyuOh+3dsN5rspwsAiSQP
n2mok5OKL8MIow2dTYz6Xob4AmpQiv5nQ3MzMtCEik7cdG+bVGDBUrTiledUwiQp
lKpx+8Eqd3aR1uoMWU6shJbG8XHjbWJzltfkYkqDxlS0DE+mPs49N4BoHMEkdxme
4c58qI11hLGE/TKVUuFqVP8DMjXeHC5mtYqEQ22/jmh3iH6i+/AcyBtaLm/9Fskt
AxeqFIfwmUh3glCOFkVzJCoK1i47yXCOge3Suk3+JYmQPvrIbIQsCVop5Ikp6M+9
HupXSq2V6Hvdu0NKUdlEqX6ss3eFSmr3cF6tUb4qqa05qZvJqiucjyOtCvVg/D38
q9sxtGHDa71HK6qT/gK7Z7+meFgMLPEfc4N5SlHAWITyn2WcG7NnxrvEEYcr+PdU
nkSuFYR6dB43oBvDdq7YtB/AUUZUFoL7Fhs7AJvWW3rND0gfCsdjM57fMXT/NHXA
G6Pc3Ufl+JpVEPsKgDdFdCW0dlr/AbN7MZZdcCK2EbtmQpKoI54xSz8pWw2+XCRu
uI17vBTa1DZOII26JbxFR/PPpMcrVTc94LyhHZXQPzhefjR6DYwwPSW3pLUB9CRt
v+KIQXKYsM70xztxpV6Ly0KO4D8U1Ga9qA46osaA8TYYcpcZBLsP/FP7XCNqI8Yo
Hx61cbJSHN4DCgBo3YAWOGf5PSb8i7XbWnZXnWKLqYimXSIF5mvKKXEfs/bVMJmF
CjprrCArhNMf0OBfc73eiQ3OprCfK7OHtjhWzczwTTisAznlAHc4MpoAU7ablyQu
A9K1fAD7NqknBGoFAmB/O0QhRmULFaMxcyjmm8QSIGhsjP/aLhO7vYIssGTqGKDz
CNO+MiaGpPpsuzLnJuKRrzmBzurAcgcUCwQ4fQB3bFMucr6+mAjsQ/Q4EyNEQcTy
Cph0HzlMJlH76/lrfr0Sp4VTkl0uBhJmSVbm0q5lQUK2pSsTw6iNUOcRGvzxM+ED
wJ3coqjVe7YUYY2UXSGDs6EFI6ZaSgPuLGQZ3rVeLejHiHuURroaU7+gggZrs4Ny
pJs2NBDAc2FF40guP5DHULYdxgGydP8vRMmMBZsw7O7kIZlP+IaYVp50kypCkFUI
tQpcJgnkbC9rw9jeM+T891ImRPXHzpMjBV5TZSdb56kcXKzJa+3X7UKIVbRgNc3T
2uZzDSsXQen6RHbtn+whfvYI9SlK7I/GCUuynlCRoJDgWPhiCC3PbHhOfu8YQO4T
JXDBlrv9LRlGBS2IBBletlBgKelsmwiV/mlZgTCWnIILfqLZnu8iJFSh0xg3EF4C
2LxUS6Q5YRM6fIDZvy2zYo8a3VhuxjiYTS86PMYHI/3rD1mIMDUsVA9xIDs649K0
8qkejBerjGJy6JLnPf64Qccib+F7qEvUBJxYIICz+bJHLPfw84RtDZ0N7242KBT2
IeZg1nlbbAVSObbVZgPo2roLsN09Y9HnbbDHFlh8PnjTLE6D+RLf3Iu2X8icBGWu
bfVMvfZ9trNxZGPUvmb20ugVZaAF+E8XR+OtPHyBe1ay6/N6/3V5rTTJw3BoT0Ui
Ul2NouTbJKjvD3fSrdXoVLYU/7UOkBpZY2I67lGECRSFG4pegIigxF+cxwjde36Z
/cm5aKed8JLxVSYiDzTNMUW2B9i1X8C7gD/r0/YaDUHRH99kjeYx7XuSpNOtRhvS
s3vke9+Lz2wxGYT2hxOdDq4xpXhI2s6rgfb4042oaG9U4R5wqSP6bf7aQbIbQigK
yFuPiPZK976c0T3NILO1xdDJncYNybZwS18E3HHre5tSzZjlaJHUoMM8r8DXe7hZ
NG7M5cSpIcAJrncyU+TzOj9p3XsBmoFkahB8ME6NRvIA7R4yjvowwnCO+uG7MzC3
PBJFeE9Js4qjpO9WrekTuZEoZIkBqxPMM1TJFpvhV3H/ewHFUt+Uy4HnloHGuv1B
5rwyWTLJQ2zKzcGIORMwLD+VOYm1f9C2ZwnjnyjaAA+WzOEdpQmHs2CxlJLxW95x
2OwSW2pIjC5Y+gXmqhRtoYPgb5tfYV6WM++A2IPxnCyBkm4n+Uo1nltnBWx0nLy7
GVRHFldAzkbI+hDW3OvdxmcHeheadEm+fIYb4ud0YjjBAC48x/g8e/6EK71pd4Ef
c681+nN7+ft/2/cuMDiHVic9PpAJcHC4Eid+VXCemHxnkjjMBTiAsha6Ikzo20Jb
uGzdsbAzTXlhnUPknmeG50LALLS5ZAVpHKSFuRIPGaHAKir5by7GLp5cggKs45vi
FSAYJc9VyMV8v3B08vP0Db3QUMQc/U+aGLmjRpLDIEuiq4Zf9OwfvOVIBj5KXiOx
X7JmfP4IGsAjK4xqc/2RBMm4df1W4CG1vKTc9b7AiLsAi8pRZU7fR9kLx31QjmF7
0gZwNSuT1Kjn09StA5h8NTYyLIjy8C2ZlscCCgho/paQsjWXpddvbeSc1VZknkWU
wlNtcMuvT77GGmb8ljrHgBaFd9e66EA8nBSQzdHQc6xnBRM9ctazbfozGMkSIprp
Dm0d7vVX/PogLAgCYMvNr8X0OVoejgZhW771GV58AHn+AAx0yX9EOynmUrf3+N/b
EQNKkYLR00Fta033nSg0Qal2cHjUqXdFykocvLpR61OzlyyZQZQYHjRzGku1U/Jb
uJdM5lbl55K9kx0amiB4bu6x+f5oKepT2Ngxh8+ov+LqkEZwpfnjwazLtmNHgT7m
hHg1pchcKM7Zubx99oVhDlv62iXMAShD4JqZkAt2QxtvwxvB2Q9P1VJ7r/0PvzJs
7LVnOEbHryBSqcOztxPSG+hYGW41KtHxhwy7gLnMeoVzbkwkzUCtE/1RxZqtDIWE
CV7p5OS5uqsr6l5aB8BdLkWOzSB6VGcKroUYuWcL0Kfufz6krWem28d1z+Ju4OB1
4v+3qhCGw35COx13WuheF5k9AAtH+dXE2lq0FyMw3pR7jiIHUX9RFlX3lqls2mmi
K6JweI3VEaePKRa8yY6SaCLdacPrbpFDB1QmD9AHn09b8zIT3Uw1FFOcVO5h7hLP
2X9FqIXXuquzQWaRHNf1K+RzDF0F5VQBLdMuy5iXsCxFOWeO/S/S52/hq5FTllyy
ObgT1qjDQ8MyG7SM1c3s4oivkhfT9IN3BOaH2gmR48Llnb5fBH2/q5dbvN4plYTn
8yzLLhOxDo3uDmAU9+0C0iqreTEYKqusaXeJmNhtLVAyjvqnWG+BAdNy9ATy4pd/
xUUKf5xRqTtithmJZkYhrLetix5jd/OrgzMwQtmvBi0zDdLL/+l6CWcL3o9rmbc7
i3biZtD1ly6jjebaVtqGwwiTqnr5eVbWc8qlyO7MtqSPEYjPh7HhwO6BHXDJDodi
C1iRIcI+uslUkMEv6kQBLi8FHzYu9r80tVmqXd74MXzC5ClVK2MOkyfDzA/BFQCn
k6AJYFpP1qt1S6Wj+mdPxIqk41Syhi0RV/kru8oi9kJETRvF6LT5IOUipOOFIyvC
vDUblKf6evPlPujhjAwguFLbRLXC16LrXSzriAzdKLAwrgfPB6638BqkSAcDRChO
IF01XzJRnDFZoSNQtAE3sT/W9wRVyLMQQHzIOcyx8VAZ4HE0WqwzS0KWDdAEtzr7
bF+eOzaDdJD++NZz9JRBLgDb048mprWqtg6roCjiVssZjG1kqgT1elPQBs4YXMMu
yC4Up4BymGXdtK8DhAs/Y1LpqlQQU13et8fvR3VoFdcufF1qL8qa3Rxft7bwKVGK
bmES8WI5Q7NdOp0CCtYkswqh5rnFvOsQY8GTHUpjDGc6vVOefEPotx3LwWv8jBPy
VZwtzdi0Zmyhg01hICIs60CchjndxN+a2fBFuCXyZxAcIi7bqSO74vFdUJNoFyM0
uNrJC7d1X6DJZYpTUhYGRbQtXTZcocJ1ywTXmpqB0A2sbwZKsil901CD2ywHXfI6
jY3TOgQajtEGuXKMyiHjaAVa73/f0lk1heAtsy05wIirtaNHPTunVq+OYkAsYEmY
cSn3m58DIhlvevYtMZnahZNNzg7N8BQx8aEJntSgv1R7Sy1zlcSowJxdVXZX1M9Y
Zu+97V3YZV+1EF6mrSCFy7aTIdIZ14vBBFrs2JHgEDhrbqwU6S9YYk83gR/FBP9Y
VioWzAuwvz4a7ZeJ37AwtGEEsxmLPIF3FTfVPeuzdanjgraPJBnUwCa6ZdL6lF7Q
8OX3wn7LxusznRVN2AZfFxV7NRjbIFwl4/c2C4YSdPYtBJlowupE19PcB3bRvRfa
sq/Mcjha7KtfNdhu/gyZXOWiB02wxBMC1qdqjMBpRpBZqLiu38XoF4jtlqrzzTSi
XgvrbKXpbKcAUFKmUv7k77bdbkPF4h0RyevybOyxEpsrgE9DJTCwrhliCgXLVbsB
4Ye7Xv+hlDIEoKzo3JywVcQzeuZMsxWsSJb8PKgu75+dKx/uyNZPEYs00KdUw7yA
I939SCPPNAtgTG2wZEyx8njB7zrhp9pEzyZUQ8urn3aDp1rixCKfudwDu+PAKdSx
/i4eoFggWpzhhsDiNrRW2KRoAdYR3Vi7Qp2ABBmbOA0ayaSsWiNxa5/0uVhqkG7O
JU354OrPmPl9+lsSQUocoHCva5wW6bUESelnkB5wnuY2yJCqNz645fO/QWhCkFsE
z+rgsPRgPG6z/Rujvze6dokkoxg0COWpKbs90j7mbNQ2yaqSVlR06KUFU6tsmYFm
RGNYVq7h+O2L90l/8YrYmKa2UC0MpHBmlOHz0y+UMX0eMw8KJPjIIeXrcL4+GLo/
TzIpbpa/NbGmo0lFuoHOwrnznwBb/VpZN9I+KNuVKK66EbkfOBz1NWk+Nn/0OaVu
IMEehRQ9voKFxElSOqAND4zxn2NTIA48N4dyYyDSL2ixJNozGQEKYSIfJPMuhctC
oyYAhOnMYmMdKh/VHj2u+ow4SOprRl+TzAbYzgp2aRtmY45jHvkzrknS+dAphelc
8pxrG9L4Qs8OwH29wUUWTLxT7avkgNjc5Tr8p0as2xg0WBQ3eSTkCOMW4Ukf+FYF
ayuFfUedObxBhCh2Ry0ANmgGC7FoAluQUZiNXCYknkYlcqbrYFOJRRyIP+ITk4bd
6Oo679GTMwdz7ot7FBIp4vbjaLKcPnVkYK+TjaHz4UiOZlRyojKh6XmyAtSqgOEt
AgiSaOR/qL4EBtnPhy0IXnwEsgrqplB0slchkNnGaneVEPfijU3Fxr1VElOg0EYW
afNRTW1SELE2yevaF8K6ieCFHVI3f6mJTRTIGFGaAnVZ0bjJOILTFbCvahRzMJ5z
yM++081gF7IlRAy8QajZezoccIBUvvtlvbgf6mPRzrD2sHPoNaljJcW8lZQi+OJT
j0ie+uuf/Hno6GNLhxlay6Tw0oyCSlL8kMkCQMn2KvzBy1FINUZ4ci5FsBZ4PNZ2
2kqYliCOfNCXCVNfZE16DKypEsnsp8jRcpJPwJv/MMY0oaB14Xw2MbRa0RQ9ZFpq
4KUZgeqi379+rDpcBchnmwMWP7C9TRZPcU6/h2u8AowccCFFFmReuK6U+s82xsCw
cbzIQv6eNc6YlXMwRXYl7QzW40BzsBX7YblDchpdGoEQ8qnzwcrq+oG/JG27PWxK
5o7ymqB1kPyFEz8jyX9T2GuSLKtR/8syCnbqEpEJdXEkyHu+jEjiZP8vM9Y9Pxfc
RGjBnU56jaUP0LJ7HaJ2d004NPmqol0SkiSumSfsz+VlrqBt8GAeKWekvYbUqleO
yfHzegxEGzcZGgxjIpdzLCHUgLKa2XVP1baw7D2IRs1pcRTUkGXDwrIhWblPjmoa
X51/MSmG4iXDmncZkoGkE6Z8V8eZ27h6EWpVe0ryGm4K4o1Z/z3cUkWmDqiYtuVa
oM8l481MNuzfLDfte1402tuFpUxyEIEoQsd2Lt7itYGg3TE8jF4/z1beTsBW1EJc
hmnu6c98cP5aHxlR6wIYmv+RCarGnS1FirtYyTZj6ohPtg9QuBTUMbBUx7TznhkH
g9h5dyeIfGp9a6rgbH9hJb9gojsXzhR4WSgp/1/Uu8W9UWt6r3dI0fYxwnwv6clH
zJ6kyUz9TusyW7OW7TSC8YY9NpaitEFjXenmp2Q2FPKz+sk+b9HyvTsbZoShlRA1
70zhuPe13nA/J9cC0cGLEKFWraTrN7anq7WwMx088zjbVBmPwJNjqh48E79xZbF9
SN6Fk06uJXdpEgxhgbqcPdU+23xx57pAwIxuhvLYzQZKJZhCHIrlUucZ78oHleH4
aA+CtEp3NGEp3LbDuD/AHWDAJhYjxGsMGFWCthru3GLAoKOpHEAo8zvudZYlOECm
7TnXGyj2dJDxUjeGnGeMd72hpcdWgSvM2yOzhhDUIu0Vl89lqZgaLBxck51XIksw
iaJkuCHq6Yn5pVGqAWldTnFML1OvQJSnyqAyycYel841ZUX/x6QUKHLf/My8Sx9n
ytvdq9FB+jkLPfsFv5OZ7aitFM1yhhmFy9H8k//nfqyyCxQJ8PxO47yhj1MSmXp5
Fc2TZhQa8nJWH1zfJ3dTzxxQZkO2+ioFa92inAG6XM054qUBAGr8t4B4c8ZV81iP
+xTCJOVCUJpYL7e9o5Jo2FuwbZxn5OoxawYTuuR+AZOzejRKwf8QwZpq+sTs1W+R
xvkyloFAbHcDkL4nQWV1XABQZJ5mvU0HgMkUJh80aYwbdtvuN7vu8FTRoY35xAW5
l48moaRWuApOcE8rmaRtO9g12nFqwbxkkcMnTKQL2CQNOKX9u1X9cxRAIBCYGA2t
kJTSWhSVkv5j2QE+7jT0Ofl3k4kmkWD6jOTHk2UM/NmuI5htlKhiwsJqPPUvrXRG
/hKYjyLikGZXN6wnmgEazVkQXi5wl/SX+ltRwKPPcoJlzT235449p90EzJH/0RpC
Z6/YxfcbAx+AnHi3AD0KuVb4krmqz2aqk5+dJ3vc2mg5l2YI6nbeHFOarvrLBITr
57Xf++DmuoCGKm+7zyKs1SpyHUmMmsHs92LQdkhRUy3Q4rXsQghqtyiry1CcHcIC
jlG+6fR9cVFO0eR4ETXhJIL8NpO+wGNfhM/q12EaWYSne34vN8T7nHl3tfzE/0vb
3k8+Jn80k4Oqhg+lG1mkqQTaANp27KDuAuRBHoud3vuTTOoFNorkXl4umyAHmANG
S1nBYmX6pr0WlQ1Ii6Fds5cIqu5zSIzFSG4fZnI9rbNnjs+6aZNs0wMQzXGK9idX
ezM/JvlRSrQVXJwJUzAUKC1A3aXUEqo+MaGkOY9/YhuV6AtHD/W1o3MPBKj3RawS
u+IMtBa1z8gtvfsTbmx9jMn+Ay/mw28eyGAh46VqFMiCb5AQfQbOI3gvIs6gRahb
CTZsjuNK+an/UEWqmdAq3ca7uMVhuQDdHrSV8ImTIQh4xKslo8ROkFbw0zlLzvnw
5SkAX0HRfZzT9fwAeUf++btBX6RckeA5lf4+K8cMslWmRpTgjMFpxXi5vJROOCGW
8ys+1MlCS701kURenS01kx69TtzIeO/gd1a3BcVOYLQRPQ1C+EFhGXWJsR6qHhmm
MM1fyE9yvIgg4YkGQaRnRouDDoBlkhm23+glcVvdW606ak4Pp2/m8mHRvk0T9LLf
05bvGIma4tsHhkvleCpWMgGOM0M4MK9kDbsdfljZoQt8clFuYC5bvCUE4Q27+ANT
msKmhyJHYod4l2EY9s6smj6E0f+7s8TleMgx04cNYxachPe77yNhcJZ+DUNUfMmi
S1E7mVkbi6qhZaI0nofyGzzBINc8kLcDRjVqOHZVyXV3G64Upcj0KJ7rdNKzQKqx
k1Ov07/yZvnP/W3/pjFCrVdxsIaLzLnyrTG1IbA2wiVpYsO9sksgM1Y9JegY50vF
/FBGwnRC6YTRnE+S6gx2HmJoxgUJCZq7GAcrb9YgTwtHomp+Gcb1/6x2Z5nIe3yK
hCR739kN4omYtQkCFHyurjaQamevAklfftIkP3jZovSChctld2dr2CxdJihOsaHR
KdpI5LTBe7yaKab1j8QRtbYoGrqxAgSmMyp7GUN8deKN/kXSJeinFHspaboZH0il
rVk8I39J+WED4X7hp25SqTssPBEOob0HK0IawebR9enW8znjA53c7qWb/eqOUsx1
tzw19GT+Nd3owOx/9p0A03gE6OAmYBllWp0P6oLFav9Vz+h86gC0kI3sKLSXGOGl
O0pluf8+NWRlnx9Z09bV2xigOMTgx5SKau9lLYejCDsXmtKAewnWyplv+UC4HLII
ELsEVHxRR4/C9Cl+aq+4MjB6XvlRlcID7J/MtrLCC1Sopasy5SYkARahZ3R9J0Lk
Mv3MIlcULVWjwsrcGunOPpECTHGsdoiHFKJnye/cGMRA5mXTxrUPeI71v14aA73a
AGlQb1MeloCURtdHPAWTZ4sse239Gv2J/GaHX0IpQ//5ScywLF+RpqefOVChk4yV
BOPWak3C1joqicmxRMAGMnGrlJj2rG+W6zjtYzCqCctKKhEsifvN/xVMruPe+RKn
JI5/wxexuHTaDsZmcCKjkmgTdsaYXNAeCYwLGZpyxVA0hysTrQpIuLtJrdkDIJr9
a2LzP8aMRIwI7w1mol6vpIqwwDk6g9ptSKRSSYs/Piryn5aoowp9KWKvH7ktyFwz
wTznrLV2Z2I2l/65mMD96oYer3bI3DlWjBTjb+lEKo28unD1KuLoyWOdotgkqpGp
6UgOVSCPrsRwkJ4rx6fUWw//3yu7YY9OXAPmQdwvlQF0IiMWJt79m7cInOzp47K6
R86+ZnPxu1x3mbEyyCXHUNSwvyxIWSy4M2tycB0B0xsW0I7IuxU8c2YIAkQwTpkj
UQMP3rFqJkqex0hc3LrQqkIfMpU5SAWsPyH2DZ9nfH89/N40o0SCHrmsW+h5RteY
QnCCxNSzMkuJ5tzbFaCcVqz8t6iDuZgcBkd/pykWHNvgFJc4ekFTW8LNWshC66hP
dUIAmEv6OQUraUJOlN2jIQ2Xz+Vsq4KGllwvn2rhCU7LwDSx2moqDBYarcdrRg7c
hAMYhX6OErf4efmHvzNK7cmaN41g8ORhUCZK6A92yQ6DGgiYKGGTC6B9mSrHCz6f
RJt+ebseCrEl4a8huqA9qTvknj0vaFaFZm3FBptcFyfL+4HU69h/HqhIdB1XgHHU
FvnjvJp/xozTF0G2MrI4+Pn4bVIZ1cxLKg1/Cg7YaU26dFJUoYTvMgoOnEMKJWzv
0QlZ+XVbA2wrAIXVpFfc82eADz2rS5BNFudVpCp/YSaq2Eyrx6VkuZWpp3Rn9blT
oLzFnHM7U3aoVZLia+zXDf6/pJWW77UYvIJK9MDiA38XBvCqnLsA/hxsI4l/smml
ndUoCK6hw6MuqsLnPk429Ny5U9KOpHlq7CBbm6fyJ8X50qIfnnynsfIMGs0icpMV
dCRMP1Es1ii9ECd4dzMXRuEiHzHd+PYit+ff7H2X+enykH0nNVGm9VevocyUlxMf
lwLkDTIQ67dUiDZr79ajKBVIiIof92sNGk+WT/9nWGHsYuaSR0ID+OBaovozVYzi
BYQoHfcWWcdqtomJ/f1x/i9jMmLv/Va7FFhVxZS3vuV2xSWcqjvhHLkn1xXD2zON
lZx72/DVKrBiY13F7TUyFiQfISdLkIq/4dGlBRfkRLCMSXqTHtd630yYnOxg6tkL
qapfCL6DJrfbwu77zwWk46aQ4PW+BEmNiiJgtMCSqZW/B6rWH9oxVF/UYH3faDXw
Y8W4JzA0aag1qP4VuSiuT+r/deV7MYynL2HaWDUT0vA719SChnt8RToyVNAeRFV6
SDPqYowpkdbdfu4IArSFp7TFubmgv8yOWVtw5H8y8F7I0dwspd9IlqyHMpE5qig3
QwVknqpoEh4yUou0slke4VSlxtYt6+jURbl6EHxRBx8Lq7f6s1/AAB11CYhuHmR0
n7FRpgIEiXwrb6g/HkfVtn1IJGeTHVtR/1oJaIT9NTYf1Dlwbu2p9v2BmJvGOWT4
zjFT1T5cp520TNEvyZN/Q0jLMb4Zu+PAHGWIkAj3AkOefzcDogtaYb4EH7naR+G0
ovMZ8lr/vEp6P8eZWzLNdVNWVFcUB/S7scAF7EQr/fFnu5SEH0MwY3L5fiXPIYgN
hY2FvU46RykNZhLiYUMqoW7Btycn2ajINbmLUOPpgkprl5M3OhnEfqCPspZgbpPS
MF8TjLIUmNKUtQQZ4ifpdh6yKcXJP8dDj1uwn/ilFkUJkECQOLfYj2zFCSOkQZFJ
eBxbNQf9l8iCCeQgNJdDYXDrnkn8JoTJb1uAXNaU8x4AvHyVfa7bbUQ1taeMMIGP
8xoDyihhhKUHtpd6XQJLl2QHOzm/v3KKhYHf407dU1XamKqSlb6QuZTyI4Ggdzm/
K19+S9lzymYIhR0GQ7p4jDR9dIZn55pSqtewcxhJGzXqsykLX08R3XMkV7vsGser
npS4xBeJEZRbEInkCvElJ11jNFKmhT6pVsLPLOP9yfzqoGkdKo50SjW7/Z7gsJrq
9CCIVd/hMG7NGUK1s1zN+NTvSsNv8MdNHb7qGRvdYLU5Z+Ciyakby0fWlz51Z8cp
AovRsZFn6Mrn/wZiUItvVLePWu8UBek8SPVTjwYn6XtE7YjRC+d5cSMbKA3Cgmuy
i0xCS3C/Wo93cDwDY7O3KCEkZVRGM3NSfAOS1iBPX1shL9yO+s6RdzQde5Si9q9q
p0UJFjhVE24YMq4lLdkC5awx/Jc6cH7j+qNTZIPbyqSAQoiLCfF+nAsNdyTwfCHf
+SpJbynOqd3rBeAJlRuuHgqYBjNwOyfBpGYlDPcoz3f3jl4KZwNmd6hm6nBd+RCt
P8BNlYE6v091ofKYohotHPTQm+1+ysBI8OYlu1pW57qNYC2uiWTux2UjWRTk7s2M
XvtJ3/f2Aq/nf5P0sFnXMKkdv0INDyR0qyihTNt2hip+VnMbQiI1StEojZcU0TWg
pXFH5/dAq4UD+/8omchWOUz88H2vb0q0WybJL6Wq+F4bLjRiyH3gKhGiFB3w0gcI
lz8WJ+9WJGlXwCN3lwqLW/94gzrd/G1q4Ef7g0/zY6/mYzX2OHrZ4VTD8viqNBe6
ZgW8D4I2ZLNZT3gBCBuJeWd2zc1sIVO9zGGKxbH1MaF/e1PJdLFcFLC/e2uQAlne
Y83fZFot4fpOcOyYXo6HDpnH//5Nyd8DV2E6h4wdjv0yUF4TWTDSvQVEMq8CDF1w
qmjpIA19/0x0sOxTNNzQnNpeID67BjpRjEOSqS8SDuDNu3nyA/9nmno6Tp7sCyNB
Ds7v91iwz1p8DE+u6OrMYY+vMmbq0aFdE277YuESiFKzFEyAZY2xDtnjO1CfnYxn
uwZYiqABqpiXqrglZ83tnO9S4kv1O9+0p8IMzi6TKt/4+KsHrrCyDpT9yGe0uV+N
eUmB28lVdybj0uV7V6r+wJmsOo7gV1xRnflIxdg0ir8tpSkwvWWI0czAEOHIoUlj
clJzeLsQ1VHTVOpw8DBS6dukw1BWF3BQaUvw+DYsph6lpAN2jzaNe8hjQG4ajLRf
fO8cJgQdi150L4bsyJ/qTL6mTDWnTn8MIn/V5oDqYV/sUFEcmD83tLQ5JQG39cRC
X7LlIuPW6A50ldGtgAsP9LGCS6s5l4A6eWPVrhX7x9MoYxDh/6ModpQdIW04vfLt
v40wkfdOY8lFa/OYLtg15oHJ6GDFnVkaRTMlAO9xa09TjdwDHWATINi8375jkByM
fuQDFutLi+/4cHPJgx6YcbGgtau0voBgv6v7IR7nxg/ByjAAZeFxhxiORfXPEWUQ
0ifFHV1GNgTm0PJpfAk/SfM4fRhXxkt+pGUuza+vIEKX4H/m6WmzfaVMos3ynXgT
KqTZ9fcOZKyoh3ZuLnwmr2oRzaC6juOz/9wbrkAVnJov7Du8lVSa4KRG1OEZRdxd
0e1StdfdfY8Bo69BHvl+vTWC4py0/l3R0TC/Aupzp7EIdAr3bC/6SP2Z4O9y9xFU
HB9VV91so2Ej48Y3nnX7XTAYWGZoQWjrmWhptSsOilfXQxAkc9jkyHQSpPyZRTPi
Q5X/cgQgeUvnhHETSQtqqFhVhK+q/I49iw31x9oCgbJJF/PTc9KJfwDX6IxP4uE/
N3yCFU761F+hPYw5rnuXTj3fMLG8/46xLydDsExnm6Ch42tW5rqeZEauAjMCeSR+
JE+a5NgH4lUQsj9KwwOsP3cgBj07ZYHpOal0R71oXOPkGFcWCiBUVbbdMuZ4qT50
EmleGhi0VGfV3REQCZpXFEs2hHu733XTtsFsMWXQIjwHx1Pgwp6IgT/LZ8svIZgj
7K2hc+qBND04UAq9wBmeBJuyYzrQYMTQwLotdroawOraE6m7TuW1i62Adrfh7ZgQ
+ZX55sr4SU3Moh/oUOOA/dFundyQglYBH+BNEQp+UDi+FbFqo50eFPgSLtU1QU9R
NOZbIDJmf9P3FAfro52jYt2iWI3KMf3o5IO0KAQlu/hNB/ISv/snJK1ilOuCNXuB
AhQnWPyl1XWpJnGLjsdW+11P+mbYIpfv0kGshs28hAMYPgeqzkh5fDIzcmvzNv9+
JKl1CCVAG3Ba9bx4H6btI0/dT+vm6HA6NBxFI6WMTQrdaaZWzVV/YaEb9ZRGiwcf
UXbq2JaIdejooQrseOQVvoP2FIF/BXcMjHH1CmBaWBgkQ3BnsiKcdw7IrqtCol0l
CJJilfqKG06vFZt3fVYUpKD3fwrU5HAvlPKv48v5wj9h4dfg9ejp5se01fY5GCpJ
mmh/WTpDUsrraWRxZEOToDFFIXHhxG8vJDmO2fOSPpv34BaOXTs2xkAwLLnhQTK+
QuC22wbcXDTsi7g7CkzeOEop07XrPPQSpC8GAiX4itEEeEwzPEALvwpZtmM2uij7
r9Y2RYkZ/2kuVEWEp2mA9FMEyIn5dS/r+9WnMZhdKYYV7c344C9W79wS1QkrOoNC
kP6w3FBHguWevtn1pSfYrajUFDZqCmlu/XglD3fLxiKqXfNyRkZYPXQjkO8XlNC2
+KvnPAOLU0Wx4ZEI1M5bg7njdgVNZGRTwCFkvp+yP45q/5uvasUBlTyDXl+a5D6D
h/NSc0Ud20CKmd5ddfGFBk5/IM/O3VnY6FqosG8xFdiadJ/LfvTwWAIOm0EdwrjB
fEadGuYkuBVXS4Yw8kT9CZRlpfJGWsgu9DAD+zjUXBujbl85Nu0pvXicsGPOcgUC
9sHdaxljxiMTtk0GVXLXGt5sLGTwGkflQVRMcfEj2Tg4/+bkxmOiR7ZKHtRMxo4+
ZwupSCADCVAHJbWb8UrBSceOF3KXcM+za75ALRsNK0bSqDMPR+tHMa2IuPWp6Arg
J+7sHd8mKgIg5IKPHXeLe9GbG/Cm7fkBTZJINYZqlneZ6QlccVPopDcKu8DFYezC
pJLHPevnlhBEeLXKuHEn0o1fY3wOgNn4Fh/KG5LC3w0TGnPnXLLS/ZL5N7nkiyft
9oywM6gZReOMA76kwfGKjW11CpVMTURsL1MQ77YpNqMlKPJFYzMjyJe533yqIfkh
7fAcgFsiCYvdAn1Pjqyi0koUAcCUVletOdtieWDyNVQmCTcb/kO6hMHgM3mBLxoF
Iy2FR+MHzfmXizh8oyaXAh4q9g7XM/8d7rdGEapwAfRr9sQBXYGIHC6vMbZB6Pgs
p/CPy3QPOGt5XKwDngmmb/5k5OqPLnYvAarcC9ErjU7eeSKgRNNeV/OrbbGSNBz4
QK31e0EpJLJt11Uoyxa+tsRAATJyjlolpjm5QDtnqX7qNKLuz/Z+VnieRtgzfH7A
r8TVwNthAYDSPSoaWrQOWNRXujt85VPagpgLO/UZIr5qw1tS90kYlp1gy4XBbifu
mbZkLMsoPC35wXfVwQKA4S0Ew7ZXwvMD1piZfNtT6anEehdjr/E1VJgYSzsBGaAb
5bCJYzhZuxcOABar/hd8cpuiuWcDFn+Zh0Xwp/yN3IJMwd1Iob5RxjBFmVLLoX1u
W+6VrRgMe53xrCy9fOB4P3QrO+0SsKYawJg8/Vfm8Cqh4EDa851Jni0m4ZPbdSrK
9LZ9rtW7N+1ihHlmn7/CzQGQnp1mr0XKAIFbp/QWn+ZqMtZKlaoDckp6+VxluNJ3
kWlKi7FduCZyX1yX4rhgzGzaWyrDM07B4ys2llzmu+Txbdi2oFuUt+3p7gnJu9n+
TryZhkiRzKdUKhYdxKUzxyIKUYNX7ESA/seERvGlZHsp5IWTgb4v2l+m8QdVFIdk
UCkvbuECi+HkpGluMsWutVwBPKniDILqwMRA+sBTG+FJHVxxPC0Zqrd7FK3z+0nF
wXc9o+YGs1tRMcK4JUZoR4zIGO5e1Tq5ziBFtmLzYfMm0kueaO2XtLDzEwI4Tznw
osLWMIDZr2d48SacTXysPhUvLiTW/lP4B2vcSfoZMVQIKUNaYlwZSw1ujZn9rcAI
678WkdLeSfK480sStj88wKYr/PfpSEkt+TDdLK8MyEYBKZQFMWz6pWIYCA+bVt5o
y+yaji5jSXtK3QF4UAWLb8c6LbqTs+RH41x+4AxK7+H9UNrUtWKCsQgRlm+Wh6R/
3vRJ2fDGmCnhC+6wmQNPhIUOTubssCztLsgJ9FVTRUIJ+8/foEa7WBUMibD9fuYb
y5wCdbvL1Re2JNStxuHa7ULbVQFAjSPTpALeeITHVQk1EgCu1uCaW9JGEoBNQWu5
fcsl2U8V1Gofcp/MlfqKxcPmllxJpRqozsM6bDDTmd95FSxmkrI2L310BQXvcSZd
+tdlZqHFMiEoTAf9HlNdz6Mlpr+gJj3yE5u9Z6wYLpBkWEaik2xSIaqQSE25GiAJ
VAxAgHFFkVzx8UGZKo9XAyK0m+GOsKwZAovcpfTBK3zW6x7rxA5NNKWmqiXeCum9
GndjStA6q2Hj+/byzyJ51Uaq7jHYJuKGTRhlkcvPJ8E1IZAUxn/wPlSUzLW93hSd
Cr3XDKMl7HHRK8zGUl0iqbNjuEVmPaQjoe8g/b8GLaxxq49Th6DttFReTCMxES6r
aIbewhRssOlz0S2dmUVAXEyPV4VKMjPKhiLw9RkXHnUy0b/orI0eRIvwk4QLgZSs
OpExF+u1Ld3/rS5lc5Bp8daOXvygOovZZ7GV0Gl9feEDFbOPM4gNiOOq6v2RWV8R
hXnJAJAgSlx3Zb9B768PKu0KeOgtvZx6i7RqBzqItS+7nPKZF7eHMJ70QiXesrae
j5WzA8kRowiDBxnlsd5Qv7nF9Gz69znvJh3bU3NplEVEJTdX3ysekEMUA6xf0K0Z
QuHjRkmpvoN55/l54fN78FJbfrOm5Vv1RBySjrIR5kbraxYsnuVecCPKt7Qol2XR
OvbBOY/OZrCJ3taI2KShrLAiWfajk7uC6LnOnMPEmVX92RMXBmLHsnAwSalGmo6Z
fMZPcsUik5qFKflvMEy7ApD9pvcjKUOgoL/gwFuPHi9ilSs4Wwr0We2RNR3cUu+p
K4pslnux0Sy+prcvk37BzSksVZcWq4vQ7JD3jOckcYUcLsnObydWTHPkWh4n12Yx
By0SCyWGiYTBgqeSIjGWfsAC0z2cMTl6OHDDvKnZ/5XcFLtP2DzxLlSXNMKQAnVh
nPGGNmcywXMXUpDk8XQ+XwaniEv6+Y/0ixLsRVpliNKocCSDq4jYt1TxdEqPkRh+
78Irn4PjY9c1lzE0AvzwT7TM//LPYNZ4mTgkN43dyDMeYaXFoYIP3RWHJhORlqOj
3x462Wuwl/ulTBckr+ZR1G2Eu2dJ/GPOSzcmSTtgjq7aXbpn4PGbw5xbvvMilFOn
PxGqhlXt9BMhI9eBTrgLOXeXps7PvhDUfvAPgaB9Vn+1UD5ZwaoPlWZg4qzpKcC7
aFVPkpp4HDBNvu2bGJvHR4mVtW84N1ud+lDPkbnleE62EmWiIJwoHlUOmC3OpyuD
MTVBLGhB+9e5XORSjwzy8/cxWMfEr4nL+IDyvwDaA7WwA7B8P7VddOD1eSmQAt8m
9u+KdVhVaLeHDT6m+E+hoWGc9ZX1nZiGuFhtgtvr6+reKjrIa0fJOx/u5sACJYnD
J8eX0/l/Jgz0XfOsQviuPnakzNaURsVBdxJshTbPgkS4jGSit8BD7vLrmJBvKBeh
g389QF0pF+APV8GsJCxihFm2/U65QUEupopAc/v7dQ0Orkyp08Q3NSer1/vFZg7z
JCIgQS9auBaen1x1FbalAgqjW+uzZSx4WfeOeO90nngeryumP5sCMtzVh/ZdkrX1
hpPKX06WxWsyXO4ZfBJuWLXJ7JYIDy9+VeZp/8sRfAlnRVFXtIMu3ip89h9SFZrB
aNkV1tOabkeYhnJA5pjLGXt19m0jcC7YOhotsMgj8sZB+t/jMdl5ml7SzcNtqEac
Bd1U2wMxVtjg6xYXk/wjLpRL2T1JVZoMicxjmNUtRqbfOHrIxYLYBV/VZd3y4qPp
fNrGu8Ni9O8B7pC404Jcaemlhl8ZVz8hfYh+sfTc2VpyKVEuK5zcfX6/vbb8SIsl
ymOWiyBdO5e5LT856XfaEwYYR8cz8bNojbEaoNDxnCOaXcDqpq6TvDYueaWV13Kg
yTvwYKVf0Wn7tZnq9d8C9T4uJKP0HA9MhE2AYnfJuaqvJe/Lc77WUyl4zebROzYX
TwsMm150sHdbkNq9sFzhaBavfqZ7py/Tb7MZpdUjnzv8XYra8PpW8CKh0HbvPkr7
eKSMv07Nl5sV4EwSVSBJ+rGncD0VjO1BztixpwoPhJ154BQLtBnN+rWv9foqPwj0
oYnVaHYgAdyLFvWDt+pUubsorvnE1Cv5svHnrCGvL7EhDjijRl6bikQaoEeai44G
Nr2Tjr3ezD5L1adoLiS6EFIbDXZcUD6lpf0YDWcotskV90oOr5kFmk93LQ/ndcCi
KLfzga3QEWIesxgryqMGZbB43LrY3gzrkgvBu63RqzUtElCe0j5gFWrwkrQnZxS9
YUgDnbZ8Ur2WPpEx4HC1d3zA5ovnTOK9LBdC2zRlwTDH7sfWKZaeKtYugZcnRxO8
9WvXHk+7EyByVsZxOEUMskkO0hix/WD8krP/WpZ6SzDBbZA5M96MiJ6DvMb1LS74
1XwC0QwZ9mKz0XWtxtcPvtujgTwCLNFlMBIfedO0glBeiBErCnAUIcPhhqhc9FbC
OdDdfzHdhY41YkTet6DMV/iW5np9jftuhkH7m6LPzAkj4XkNscxBzFMq+C8wPbSZ
kJALGpneLjfXTRIXzRiueeUEZtseTLYafpa7W4EQT6hyPPmx3nPVjpaNLgbW8wCJ
kWNGCo1J70KDp4aG9GFnqn/Ei3MMvhytHBmaNhMTvfvaWQ+gEsdxGFSN3p+QTFAw
U3vrgIorWyDCVL3k97caX0kYyQHfGVL8NxVQ5RSixUkSsIrvqdaTRnSmubKkPqY2
gDUXgqAoXqcIMqGdBbWIG02Du+F2kwqI2hM/t7e9F2sWOqt5rr3N1iafO/rEbmuR
0JHVZ2uPXEqcSHvDnz9BrPyLJywqPDv/Ds1JSiSKEsVmp1hQhsmuPbwsBraiSBzU
3j2Vm04+v0Z6YalaphENp7cZtCU4wpW1Xf2Y7ARJryAkuLlglpQuT26IFVrvZLUo
sa/m+cQN2+ecmlMjUXuLK81tgUDlWLo7b896GwZ3s8h0ao6I0nBDV8c5xFYj8/Ba
0wAmZ99+2nGr6csNM8zPkX9YB3dNnqscoDQuK6WZ3FDvS/NBOuzoQFXRQoxznRW/
ZQSTmU7EAYZBtmCtvQ9BtbNJqEdD1Qf6tmzHPwqaK00Br9B8o5QKSdj4CIXDThuV
DEt1tSsHN4HxiyJ4AeYws2m/H1Lro2aI94RUgt+nYwRauGhyJOuZFTPczjZhee7b
6l9M7tyZoDawIWS6tQ5URrVXsZPKykktvamTT6i6tvbKecISLdcXjQA5+hV77Ikk
mpaW+3aPhJv9BxYTdsRwlFQZKYSAQOadn09xp96n8B9N9VA7Ido+VCVPOLrMIKwT
XV9ojiJevjoOL+kvOdU6U+svBbDnVjzgZdvB7dyICi3/yPG7RSIbRDrOCJ2IZzNc
Ojnjm4DChtT06aJR8liK7zRBnf4ht/AsuIqZWiKRBWa7wcdvx/eW4juJVs5Mb35E
PMPSFnkguP0iTWE6clcgw3OXnb7s2mNr/NreoZQ/8BpSq5loINVRZXRIFP+gUqh6
ndHsPkq8/WcmThzNzkxQPzy4SbyMKtMl75WuHXnY06pQuAJeNzAPEgAQtfv/Ixhf
RpXNAuBnorq0Psyw2e5lbRgwhCJPii3y8zLYr8FntJdS+4oUE5W3EQ36HokH80Oh
11ff8jfZsa1u9Wz5cMZavr16fGxONMsxFcJmXWnJoH9P634uBvgd3j1RwtP/Z4WP
JrAUuee59r/H89CRsmGb/hFlBIFoIUVB922S5immbou65uva4z243IjuOKCYxSGm
zKxdRvCX3QCzql2br7z5KxIiKfU8PZDNizzVKoCTWW8RHGp9P/pvuc1wBw0+SRCS
Mc4AsqCsRlaUV0JGzX5GSVD3hA3mlrVk/naUgXXiegruq2daMwRmccdLyf+iTtPx
paQCNiaHib1OkswBkqVQvGlhtcEfKhZXQc6u0FdpFLR/5lzDKHfpVXk7YxUxcpzk
QavfJ0ga4FaRgh3JVafAL0vzrY+QVxSjbpdS0VW45U5O9SvXVdr5ERAFqoW2R8Vv
pK9MY8mG4jTrlXuha62uVfHqw2GYgU7iz8gORYR7UavH8/1KMIwo4f7BfZUP5Qu1
xR2BVpxUuE25uBEL96hSHW1uAOn7GhnwEcQgHIwaGJLHFU8LnT10UKmbpB3aWPcT
4QosndCH7a93i/xKlp5eaxXbYpjAhT5pDjwg4lDxRmByr3eIhOsKEO0wMedj0ste
nRbEyqxhEXR3pSJEO/U24qz6MXJz2oR91FuCHeeTkGhM4YB1+hYvlBvJLfgqhTXM
kbAc212NGKd9QnTZ9yWRMM2+TobREDXnUOvum8nwiKM8syPU9NYh6aBvBjG8fVZt
M95M6fcMt6kk0abyWixwZhtUp8PPTEWCYlUXcYjKb5tzMH2CrXihrLXD+nGHBTIR
fliz74z+QrxcCseuWMvQji4yHa6YGuWEL1lpaD7kEUlbAQftjkBe3MUaCWlzX4Bd
Y9hwDY+2GRc/6jLbfDknBBmoTP/hpcnIIhk3Mj48aTj45hTAvCPR+5AIMwdtgU2E
mdKURsRHrSPU9FAlsyGAiYqkGNtxmaEq7dDTKuMfGmY3o4x3IBl5U+3kPBk/28xo
PGkpXxx428qiHohRtpHLSqn9iCjVwEVZZXC1RzVOdFiy/1+eGHLXHuluTWhABNF6
HSq5s+uObGbYJNsC7auB0i80rDZldWWm+GZu8njMJ/xLPCztPg1Sanfwp8JEdznr
qx30tAsVTT/9M1wdJd5AqJKhZfKzGoUKtkKg04o1m9gtQ2g724MkQFPYGCB/simx
Bx4amfDg0Bz8+CVOQe5HefCfrCTP2zM0lMuIOpEPXur3efkPp/eiXJZCuaoLuZAf
ftbqYzOcWH5JnfrCo7XNiLYwERRa4x1dF8YQ/DpOkyzMziMK50ZTBCeS3jaQLl0H
3kqCE+foICqey8iHODx5oOmAnMlxTTGESxGKvceFCGL0lBu1riq8luI/4hrLUfOq
TFlZyEuSQh2sN8LJeZc/BfGv3Q9ClnI5yokD/ga+RCgLn4Gnyl9sk4o2kUb94j6j
8qEEY42VZGIF1f4DT+jO1P/LxgunezeXWRVyL0nFJYz3ARu6S6lwaqGjWsuvGZYb
Ptg+8j3DOJWt8FJVdAnkyD0LzYbXSq4s7F8Ce1zvrwm7Zi8n7o8URhJkf9e9f2+J
LvxLNDkJbHDrIuFcLI7jpgZkuX8r/5eB7XKUFDcU3Z2Ad6FdWsK5cNEtjMt8ivvb
9mdd4TJjUKQO/19MokkaeSHyc5mEeo8wlYLx1Fwamyg99JmXgTY4mEBhOmS/BOfC
+OXPPJHimYd2+fHxjQSyIIlDDg9g1DBen4EPNJWuFoNh/eACY4S57Pr6sVo79+b1
ibsXdSGs/R9HLW1lwfEbA5HPBX1nM8S6/qXttf/MyK/IRiPZv9LnL7DJT6TWT3tf
NbQbn2Sjn64JuiG4bgt3SSFSRI+nsGaoeW9ML8XDi/o6PbgSKb3blFbTiHbW79Ie
pRAej52VO1YOe4sb3sidBsAayva7d+hsgVNX7VAncgD6D5eT+OpFUITLBjSZEdwc
Y/+zpkH6WM6kQVT1woCs/5Xc8iWarQpGK8a9M3QZRqNhiRCWbzcZvt5RKWvyt6hB
bDOVbrZqE/1gvYLWmJhx/D+tj7yKvTmSqH/wfVWGbz7w5FRL5LgRzkl3wWGMJYt+
CVthNbH3V9V3M/ZI1/cey7zNQWIwFZwczInOnReOJ03OPPuwxN0LY6moJY4Mfbr/
p5wAUUHvBjZHtR4Y/xs5VtXKBsPydRNwo4xYB+a1wgZV4zooFZkm931dlnydO8wp
AbuRAr6BOWLXkeslLmXIEsMqUCg4cD4UDC+pKOjuqIebbyh6hC5ttO7Udj3DKwDK
qBCFYs42VoPZHv/Di+N/e20nXCTf46rygyoBEsM7W+yzp/NhUZlZA31cXG1sMk38
wR2KiSfC46YN4IJsYBJRX89gaaPR43nJ0YzZi9n7xMUF/xjngUhsAtH+zTAJECpF
+5XUD0OfYEI1I9coFb7poa31g8uZ4svuYRhGUwku3E/lSD2MTuKkqbsEHqCwKodU
KQaOqb3/2oHVMMGjA8v2tsmw247vFZNlOkbp3EHuuJTjU2ZesZ4fGj9i8sh5weI1
dS+wSHoOT08325h7Vfmy0iP86REBP+Zj3I5q1UlUa5yuqmLZFmBAXnSqgX5waC54
FtgH0VVIK3s2l6WsWTi2FiitP2uSekE6y75jsH3VbmdVFJNFJlLcnfWB9YpgOnhS
3OQbkm8SCF/dWiK9jt8lRTA1n0PPBlfy7HK/aiHg2M7GIlt21K7Qj4z4a9TrYwGA
ZdyroDWhK+/Z/jA1rB9huHBltstjsuRZUxItK0guAh5yugyNR8Pjyt1VCvyyJe7u
vCr2Ea+3xi/uU17fj1p1tmVzWQGLy4if+EGqfoSTuiIhQADRs5kqLajgx7LP8VTL
KXKgCQyZGFMAY1WcKKP+cQH5Tf2xAxFb/fDsObICOi0z9OAShH7Fc6HRCPE+To9r
Fmbthh/g6ihyVCCbg05IEPD7FSte73KBaU9Nbutsj2HbCiDaGH9aq9E2kxRnawFq
pZ80X+H33OvuPcZStzJlESg9ab5kg1MeITWaRpo6dYC4vk4A5X6YSwJTklq7n6k0
A1GxEWoE6yVPHkPP8ZFEj5Xm4rRsgn4Q9diZknaK4m/AHYF7NYaioYsHDKcWBvp/
kC1vhcZ/pMJwinF7e9WZms3230LAXoBlxnQFndIwUtyIwPnOHSPkR/HbeLiaedNG
1TsC34oAJQiaXcUCNV1U5huAYmBWa+y/jljGpXWajyS208ZRXmI1S/Tav2mkyxbX
MZ61+ks9xLzKfMPTLIbRXJ8UKhsB4ZFTnRh306pjtDKCxuIf6usJ8XM2/rTPY3Yo
8FIKkOkLgcHl5wdCXdRQ6ouhKtfOpU5RLfFgf/oZlea0xmwHMNanNYsGkOXcq9jV
8XMyXQPzw3Ba8a2TE6589MxUJJWdIHGLzyaPYVtDBjC3BLjIfSWOQ4Uc8kS90ydv
gXUIUfFpaSeY/Br9Y++VM+hxOrRlN+P+4zq81O40fi67H+fmyhKs6cI2Db9uRt66
pbm/3/Dg/Wf+3DyuzPRt0rtrBZDB1lPHpU1huE98EJR6bIZ4dBnbvVrryJkDnvoj
qpped1s67U9Msk8VcwFdm3mUv1+TdmFFG2BpUQXNpYxKlXHDRS5pSmQdK+mKqLnt
p4rK1zX8lbvvJfks3Czr6uH+stwtJ5Awof7+EXBvw5aAErw1gHyC9xl8asJsT3I+
5kAqEBNt6N643BsNG5ELBQL1XuivlIxIFM4qnMT+MfYW9lt8g7vO2bylc1LVpR+C
6CTSww9JuRFT3DYjrqVhEp4OvR5den3F0DwkYPwUArSfCwe5klxGlOxHkYG5TqxE
tEjKY0usxfSyR+SrbusFHwm9plYWfcBdLKlubiOP3v9DoABZraMPENa08jSH/0gS
jO4SowN17a9NMj/a5wuuqfgC8tHlYHBo4CL/KuU7R+kQX94f5E5vBrK98VkRY1w5
GHs9EW36GPqDQO62qJb0Al+cRvEb2Vss+zb/HpLO1I8mphck89t/UDkGu4e39/y2
Py73Vxn68ktNFEbwa639LAqkgg2AjGsJGJSxFXw9vdMfhXyCzSc5xD5N6Se3QYZ/
ZHt2/OzVXaT5uR4t3BFYbSxrNDuSj6zkToCQ6jnSewbbdP2RszqNpBAb/UUygFsE
++j6I6/yMGaJTYpMae6DQwvH4wmiZnbye7qGZ1eW2vvh4xTMKIoKz/DLcG+BI91V
vD4b7zBjc5gn4wCICbZBW8BuKTG6n7hU944SIfyDRlpwfZHVv1KSJ0ewNrV5S9pA
hbXRUgF2r2f60LGPZTAmfCC7bhS8vonoELoqUum5b9cS/yYnaKcOlrXP376tg0nf
OpxfmbEaNBIXLZB6aHPUdmfkgkIDifuZ2Y+0d67sJf4Dm7pooUF8G55EsR4Cz9fz
gc5/e66rddcECDz5ovcTM7onPduulxdhNXItJ/EhhXFg9OwH3j+t+NZ+9CK9g1TA
ce847QS++HjPVUq0y7xBhnCHRyN7PbrIeGpB+nV6oDPhcsFvQ8MDAralLGJig8ze
9C1KDzBiaUeNx8/9tcE9kUgb/UFbdGKsxs1fK+UyeA85vr6D5G4PuzUB8Dqnn4g9
fKcn/NJbt9k75ezjSam8oKB0kyEPsZkuO35cdgJxHPbXPMi89mbNZ5JHfyaScbN6
UanddErtBU7zVpsrDsw3jU2d5bVCoLgC6zgpScV2Nl/KmOS1TCunjCxoZM1dHOsI
/eWDGbPAASjvUc3aXsbQfjBMY1XB5tMK9lxZKfoWA8Z3nXKWZ3CwymexX2ao2KTN
aT25DR4pC7rZBxxTEF4znnPFmZUYj4xVqIjdcQbm/J+21kZBJyXvdue0Z8s13zh1
NgY/xWh7d5+ypbzER4jRMXQbNVp03iSmd4TH/hEnLbP6bsoCySCiCJtKHYhinl78
OFSzg3NBUFiFd2vDTRDvtqxrGtJunX96kmNShq5q/Czxj8Wvd+ApVNJPQo+ZqwSb
kOMsJfh8lxMdeSkKFX36EYceblN+2GJxiAG2SNl62FZQJP0AaxP3dRSeVEypSnSQ
8cgIn1vjlWku/Bt3Lw/7gcH00SgI4FWixJsSisersW4WB6ZxYGhtOhypjjTFx5gb
wGhpEw/y40dFGPtJcBX5IgQoEi7camouOhb9SpxQeUatXzhdZXYijx7dUaSDYoxT
CJh7uQtx00ZbeOp48b/7iaafG19g+iYGWW4rKmx92fWKvtnVaiUcFDNLoYuYB6+U
NWnvSaTq1kScyUhDQvcOcKSsbe13ok7LIrPLsS0GPF/zYBJR7AimjbfMsFjsJGSx
22/y85gXTLIC0dsnQ3y4CClt+SZB03ELby4BJX1IxbrGgbVvRKi2/fEYphG2SHM1
SKuuYC0zbOMNRL3lGpK9AH6NvmkajcTktQvQ5+HOSnU8M2NcPTEmQr5ndcv0XRVL
sZVYYys/jfR24p5voJqzw/0awj3wpKZVbOhREo9PYSrwwq6dq34Dym99vnPsQrQR
+1JTXXc8MeQEFdeqONWIBg90QDe2ytnZ2XXmmByzMH45OxAXqiMLyYopUBLgvzgv
3YwLGqNICffZXqAM2gE5kYzTTl/5DUJOwUUWk1mTzUuSuYRaH6Qv+OvGKJypWJje
UuUVXatWBH9lLOLgjBHwszur2v3TWKDzB2Yh4qhQwsNlIVuFn71yer0VCRD1rIB2
/7mWqQSzIIUB30yXzqcsC8anpGFUIf6bTXggOwKiB6FBqFsCFHKpvWpulv3RGOM5
mgXPfmEjCesJ19gXEA2NlS6+bRsByOX0gXGl69YH5l9yoI9CHlZyZULpfeM9kZyH
GK/lvgkpB4Fk7bX8ct7EaaWUx7NYog+fFlDwOQsEDjtsiV4TRFtR1gxnVoWaGIx4
pNgDxBq8PHGEgXpfd47v9tLkWFllBSsWNidTPq/RPlOr/kGMl9oI9ojGM70vZC0Q
y5YcnTpd1cbCXVJnRt31dGucLgeJBKBV2m8MxytTH3xqgff0xZ4HHBRpy3Bsa+T8
qzxB8odDFNwp31HeP0ZACqNS7FQ+YXAYiZX/pVdeAkEd/g9eSALR6AIegsVgt7e7
8G4swnjFVw+rh3NA5TVd+7U0rgx8rNq127D2zqfmgJMEGr5gn47xHPjLPAZZbLJY
qPKBxCsaI2mRO1MdQ/ygHsE0MHWxR2RE6H1bzh3hYkBdraoBa5suI1pR5+vSFX45
HONP1c/YszMm2CrDPhcy5zP86uShReqzmt5AhMbPB9UKZhSl+fQEPKH7tDJ+lfqk
BlzlCzJOwPDrjIuFm/JE93vVWayzp2jPSirUX/FGKA7/FoyLne7zyBDdBnAvuqE2
lpTNXyMHN3jLaqZAs52+3alx7yJTxFfbTjDkYR3OOSwKoXiRHQ3l0d5qFjiXO694
BH94T4YqGC5MZZTril6Sla3UNqxQvZWj4YwARAnoZerDbrdxu3GJdfy7G0+xk7AN
M9S2in/vPbkGRNCpoU0LTUsEFEYT2PRz9Qn6RJXqyOBvu+GJHHC19/JcccHCjoFe
j2xnnm1rtsrTfeX4gcqpAGP9RQDb0P293OlIRN7+39FAWJeR6iQSwJn8Knr2XnYq
vNdkEZwpnzkUV3BFEDhmYui10N4BgsE+drPXubrnLH/NV/FEanSTmveT+4S3TBp8
C9CTgKjhsVk1SuTMAnn/4ggi1AnlkEnjKgjwmz4NMmPjZWiN04iKsuMYHtpokU39
Qb5IcJzQatHDZMkV4LcfRcYvSX5CyU7lKbNx4NpDrtRyGAuK4ZihXoBEuxx+EJUy
4cdVp1GO6tTy9XhI2/TB+K7cu8lGVw+s1AYbjmALpue6Swt8DTnIXQTBQvqeSrzM
2vd40ITCbZHl3tldnkYs+YvMM+r8wqrWjU6EJUTRPLxRzWKf8GyLM8tEDPmhan7g
mgb5qMtOXiRgvAQGa9KcRE3T3KxXM2cUha1b5dEzmSzpgEe/EnhLB1k/n4FmHJgS
zOUyxvP56QIjC+X8Zuw7LsrEa4AzqcRKbqwMWoh62YzvtOB1kkEBr7ruHQf+FKkk
B9AfQ78h7IKhX5iF856I/0IrGH5gdYfXWvLDu1EaVjEDADZWVIhxKLuMRpFKlHMd
MeFGomC+kYPHbksvbafoKdkGIdiRbUl6/cHkTcpo7eGId0P5bVNJoorNk1OXzI02
6dYyWljKj9nPtkRQ9zbkTP94IvlYmiTy6OXxJdqgnuC/x/uwknHpkt1svPfZ0OuP
sj4iGVrgw8y84COHoQKll8YtcCu0ajhT9NKgnK3RypGNH7PRXnIfc/j41+RLO2af
hJCub5Xd+2NxDYOpeSB0WKNuZaemVnFIhWJ71/uI6P7fpJy1ETghqYTE/joy0kxV
R46LAZ08d2C8fe1DIIaLPQEPSDH+DRhXIfMd/Ure82EJlRykRFZJsqBtHigM+De0
fhU7BJHzjRiB6QhEh5QbStoHxVbJIviPFCp0edANAnDEZtNS8N9ovpv7hdZbmo9G
RLyP9EFZ58Jpy+imTgB5pPZa8BZlQaL7OLvvyu0a4k2NkNTgmeHYmL6qSlPRdU97
siIwZzzmuYRKXJgc9lghpqk21WdAysSK6PQT1qRseaMprQ9mKxcimbRgp+BjTL1I
STs3sLYy4ug5U7wxA8FscbqVZ1PAdxdOnQHh+klV05GmCl0bsiBmfs3ctJ783rbM
++D+xkUECwud+y+oT+f6e+R0tzu/6H1KgDeDskNFMhluCQ7pPtO5eqkyuVAwAzXd
VxCiU/pvr2FrQpzfQ1PfsugfPYAD2rApiMtKiixPindqQh/apkPrjzeWwlPyn6lu
QmH6uDKI10Okr63FzMHzGD37xy0K1/brwrkA1fZBFjHaC1UjKWw5hYt9Ma8vJfZK
PyWR9NgVvHnzg7co70JXUAuSrQT5T1NrpYY19aVIfVxiYjc1Ds2KHcGgwHxefj1L
Tto3A47cMqTxurJEYzBnTp61nIpOyMb3T9MeiNuiToP8M/BKvxhZEvSDVBfc4Ii6
cm/TIkTDVdckjKs64G1nuRKGhxGHe2J37R1/e1JvoPSQ5Rvr5vDcwsKKNcEbS0oi
T9IwcWVKo3oghyMnzJLOn1dzeJyZAyjWgN8q51UtO2MC2dfshPXH3NW3vxoPjYdU
F/sSvr5FTEauyDB0NJedchE0/KXGBz4kw2lJhhz6WRITIXizgmZWOrIb/rWBAH5F
AEAT7DPFUB7+5DiCPLvePRl+0elFTxoJ72+NO4tPyeW5j2n9tDdBEomez2bSO6u2
znunCjn7DCO9mY3Gw6efBx9xPHHoTo3se/hSmEXK0JrEBKSPLOUz+HaC7Gy2BBW4
StiVyxpOqxxPreDVT080DppVBEBlu3XnRd191mw6yxvpTfPPr9On7dQ69lBSVT9c
1eOPsX53qovS/Vp1RYcotZW3eWpI5zyETjf84KLhWuuanqTZl7hSK9XX9fJRjZVT
Spx040UIQ0O7YxMGsuYE03idmw3hk+WbMjhipeXtmC0ltDSqgD6kgblkaVNEAoAi
k+/pmN5GgDdmA9nJzhH2UtmEOW5g8J7+RNBVA69DBLfoIdKwG76eh81mO1d0uZZW
NC0ZtbCP9Gecbop6UFBEu5nioXhhOwsnu5AR37NNGIeth0G972xdk4feSUjsZUhi
VrbHHXudicuR5QAWwye4a+PQ601RMn8UrF/p15uVQDCbs1ZmV4PImQ0D+1qMNozN
0zE845aQ3I52xyGH6raiEvfPgGBn+F/Nft+NwU124hzNoNgIs9noPx/TKadhvMd9
R98033LKx/AJw8+os5LQorr9CoSqzjv71Yo3c1dRyS5NI3VYRdxSEDcg9KM0F9iE
MVfZtTUMlIKecQgXVk536wgla0OdQb7KPppL6ktqYH73s5+d1YWj6PwDfeujwh7t
aG5tbW+c4WgJt1J/301XdCj2ao++nKdeq5Zj+6s7nOc2F4eNP13W2sMFnsIQd7RG
Zmq0ZP1eoIRie7n1//cJ0Og55LdhxQK4l/cieuDU5l59XN+f2pnb0vqhtgMST4G5
wrjq5NYnt9EsXTgiG6mPmAiEvUK3dbgNeNaTwitK31chaEiACdy/jX3MB8q3arMB
w6B5MKUdFtfa1QjXeF/98HUTOQQLi4YsJ2NcX0+ZKUHL09OEJNzDJA5IUdPtXs+P
soysBS38v+PolfVvpRBGiJzz4jQ7sJKmV1KB3EIvg0uUapx9jTWOr3/7PFURXScK
F8t5TqKV8TyQSfmdv4XRAHlzsC7u8ukje0AsGuFc6rML/EA2M6IanZHivCoVGTD3
IyEGXWfe2RiQN1wYEFLXZuJXdAelFnQ3CiFwgYppuqTg6HxFo9HZZRD1aOMLO3e3
QYo1sKkryflb1q4EaYFl1/s8E5daIlSov01mW6h5UrbwV/Esovt2T4/vVnVGKN40
xkpp4KRiosruvhZI3uhkT++q4QYJKOZDDb+Hh/W31Q5n71Ndnnu+T2f+vBPxoRgI
i8/YAOSw2D10S8D+3YpPJ1lAWWgeMW6WCh7nWe1rWMvkB4LMGSjbYmqrTJJWlBPI
LsLaIAMhdXHcv5Ae3gmlKjO81DocKMzD5n98SFPl1Byb4l4hOHeBDyqpvnlQi41Q
tlGKLV2yXeKq6NFJY9iYPagNUYwC+Z++yGmv+MOKebkNpBW8ntEqCEQ6VQsjpPpI
Y/wqdgdowbdVtp0lWnEtG3dK7lBVaUTQBg8C4Mfp1G3qSn489JUI2gmf6cHU1cJR
YTn2HxjfxNxLEPVrYWLq3cJn5BTqYL0v3dnm+BENQ12RfZ/pak+1GQxZUTMadkuy
6bcGKBbEvqYqcXs0jTQYChr/gkYDliRqQu2G/yoh25sKQUcaZ4tHQMwd6V56akMC
jhSGfmONpXQrB4ckXCeotHLeKHZXk06QPZwYJEdAY6TBTpaCdwC+yiFZoXo8risp
iAu2h1khzUqzliJsB+LcvymLC82dm+LTAFWBpANNEwuLE/2NXpE5X+xLQNh/3nxb
Ai5Nkj3TZyZnEBM8fc5Hs4/vNk9iTpu1Nz4MDfwt1nYeTE6V/wTRznmgMpBwUdTI
NbCOVIJWmP2sCKgI/8dREOG4xcU7v22pME2FJUafiYi31UIgYP0S+I8rzU24LaC4
kkBK31PSyVu3ER7uUKFsoSKzSkILTRY+U4rrNSJbiLarWMNNEPv/azuXnyf2OYAn
uciYze54B3rahuhNy63LZb4CDZkO1yWjf8lV5TYw1vCt7JT25cCXROYLVoTuAdOH
q9P1vBuXcLO+EQAzQt4XDOAoR4hBTRciNNM9HF2hRtsdqQewQJzV6p3JxPPZCZVr
+FMaSMHV9O1fKoee1wWJrNMTZuaXOZKOlYAqTl3T1WIK+Me6kjthRuWTEpW70x3/
UhE23bTrTLhFGjKWPZS1seIrcx1nbKlz2Wfd80/78NCkK+bwmsCcPFhInBvj12ed
HozYAhsRpn7jfeHCbhSaADx97SJkVQCCVOi0cJZwwIUwIflUb+Cz/sERqvNVsBan
nIdk+G5suBdqamrW1ffhnlGJpb0Qitb/ObBCz4YJ7YyKSo18W370FNstrupKLagw
+nIE4Y4Z6vfrt00hwwWrSTnlqY0FRpGtaEAd4aZtvhPF+SthrvR41EcwYMu5K+uw
F2AlJvCaQI52clF1K2t+BpRVlVBwl4x4B8ipmJpXPezvXVM8m5or8GmCLdLes95u
bUbLdqBS8RQFy8wEM2yQsW3sAH2Nd47XqmJzML9lqNr+pEIdb9NeZw8WL032zEsq
dPUkJfOwt6BhPMSpPEoveb1XP5svwP2680cY/rF+WhCj98rSXu0RwyZtEmhVyQPp
vRxpaTrzszi8l7nyRZUyTBgnlPEz+00ah6YzIlZmdYrRakjIyiyJTK1e067O+8ui
XGvWggvO7d/7EHulv+tGlN597RPwnk+b2d36HPlDS/sgNoQtLTVaZKib2cCRrynw
v9oKropSR4u7Z30dZrbrU95EJEEQ4ceFbNBufsbSh7SC59yWeyPSTK5T8LbOEIbD
L7GU+jDbmAysKWx9Y9UjCYa7jUb2ERyAOcUPqoFFZ1MvHYFUdYOQoWXVmb2Sd2fh
2XBKuNQMXDxfKbcow9h2XHlB5SCE3l3bp+VAwhhdrkT0XusQsRX3FdD8IeoQzuh0
jABag8E+1nCn0zqUEczPZv77+pHY4zRStP5Z2dEZb5LyHklNlqO2i2TI/C7gx0FT
lcYEQ6CPnDdxhfA26+RgwiZWIxSFxzzqJUc8vLPdckuxzIi5eyXaHapHxgV9e328
Z7S95ngfuITxK76DGnkns8MLva1+2CanYs+pESTRrT5hw9V7iDMgn1FjbUldsRm+
+OeJhdtpvJM8sHy3354EalIGmG9WRzzmHGTiBV23kn0RWrIzp84TdQoSfolRy/+O
/GoOgRL1/fCrQHx1ekDpXJPfcymSaiiLgtKObcnO0JB8dOh9m+0+qL3svNTsXK/2
3HCco/EKACd5mrNkLizGCB97AFUCgnfsHjULx2oYCFjQf604D0E42NmkOtGdUC3Z
Dl/bzNP+B8hDgBsWZSiDIEEI2J89gXeI6Ab/VEIaFAA05UrKspODCanRJ1332h7H
DbDq+abucgUSRjuHf8UagqPYogE8FA3jZLo7xWnpnSGWV+Br0chKwiTPq0ooIxih
TYI46FxnM/LoWKTKrzWAGwAkmupzlEEK3eXMn9GBoarRaXCT0EqpgvIrUExedGWr
PL47pIMbqLxBMxcBFbxqctW8f8BjUMtN5jAE9GzelL4yjcoPtENJdzluwrSAifw3
5WfbSyv81/yruquQZ5oyhoD1RcV0cMuGwp058FqBROw7trwgjOcPKSGdwdH+DHP7
XWqL4zfElqYNGtCGShPqx01BIkC5MJgBHwRaDMOAYr3HOy54B7AvmQSBo3RpV+5N
6NxgGQAvT1gQkke8S5qP5MZd3JaQPVXHEAlXnqKRLdGJx/sMbvCJaZzSgpzjyehd
ZIalxa4lA8lwxn2x3nhtGC+GRiifRC+VrAd3v+AsF1k7XCbjjPB35W5RkMRWbUEQ
Fo7Gz6QJ9dFQqea6y7o8I2CZJcitYG1o8TcosWhKWJW5f7ACCalcRDaLf2FHnyLv
4+fWKDzuH081B4gqh+fkUUNl8a7flT77O5qHAxEpEcZC/QHjJUZ5Zt/hImf0FcwK
Q/9oReHalnwihOfyYA0MyO0VkJk20dWv5QU9eWhMHmuofE1wzkjVRTfaJvyoo3uu
d+53cuGV1PnVDfgW7mpgjzYgCCJ5qYIacxxthbIjHErfEOHShG61N7Y+HIKRjE1p
oDJ/AI1+LZab+g2y73N27CmpxQ4Am8W+kloZmc1nLy94/vehUOBDkwvlfHbLsYAS
ecbxuO+vdbkX4vDjMF65sSR4/6TylinzNjuthIO+nddXFokccb4yxalrWLvw+6AF
MsY0v2JFAI5B6GyWFlIW9/AW31G/9UrVYUoyGNgm1/DbcEegHXxa03DQGxgdb/fg
O+1O76vULyXsFMsnXzHTUJDbd7R9fqdCT7dDsOGqIbJZL5I55XldghDRd08Mgx3w
40k4xHDw+hyvIbrQg7GO1yXojKKljp3lkr6Bp2EAbZ7b3JAmCTCEfSOAGNEYcjDm
6ewwXdnhnB5pr+l+PC7Mv7z8aRx/VQEjwgwGKBQMO0O6pQ3nlPqvUU4qHoEe9vI+
GiRmc7o5hbvyGKu/Fm2l8Eig7V7odsBiaJpkCW8Y73Z4lWA0psGUTLqGd3eBIe9o
ZlMrgd5PInM1fHbi5WBDhQ65pvpRcz19mFr8IL4hHK3QALJR0JPlu6s74jl3MOi9
Gs4wM0HhgeBsPOgdk6im4CcRIZvBSyyeAI2UH1K6U1wY3HLg6OPTPMrRspZKyyrd
G0pwJf6AbhXEpqofrqDRyKBwtUrQqM4Tlcj3dD2wmZQ6fPavoJpI1EJdUCKqKGbG
ezMZG/Nigwl2VWaN9xJsOvdsZ6fWZEVUcxSmXIxJMARH/o8yyMP9PYhjH60+7XQB
R0D7Re4GRcl6/MCaGmEKp4oa6/ZY1+ORnifjmarJblGLyUGJ8jPvNihC1gFvkNQk
Zro4YwetfZFy9CmrM5lHH6EJZJE4N3czkpJj3Ed629fGGairhhOgQT0EJjcd64cN
XJb42tpFj3e8VFFba9eBnuO7BPz0kXo/GReLUTy5sWkD+VsCVS7HhGhaeM5TbKPN
fh58Da9SbjWo49kV278z1GkFeWckaik9kaBxfMkC5cq4BW+7gnt5zctvHQBhYva2
2UvJgWt6AuCxwfbdVPTkhQd+SzyyJSk4R9gz9xkC3nncqQAw94FaCIxH9TnRFTOP
AFCBobRLlG5nRBwglJ2rUtSc7+3y1I3u9jNUnGFEzPZH/VbykxB7tEl/H1Gcohfr
khlNKRUYAgfdEpj8jzqxRg9e03K5djyFxsyqXhthz3GsoXififE6sqMcZgJXk8M0
QuC5y6giNNhck/KTBUi6Nd2nXfiJdH4DtDsR5vtzhJ+pdRp+RqhHkt2OVf/G7A4D
lu+uFkXi6kNhnnGWj8GQ2jUcozKo/nVPKz/yB8HvURr/hqpOEzK9XwuUkLQB6JJD
vswZdMDKlRsuLGbfbvbXH51CU2BjKCaUnkbYjB3+r12QGC4goxa5/ItXawkXIPM9
yYupjyCDtiTZsB8TZ0FqO+XeH7Y4EUMXooCqWRa2NbqAFNLRv5CJ19SRWBGqgOgx
qvzHm3svH+r39ohlHvgLV0wXM4B8Qi7SSl/7hffOd4NfKfDRO/m4+qrauqQllrBX
gDzbVqXGuEPqLrFX3Tfcu4tJoX2SupVcN/5Pv2dRhP8C8YejxP9bcjRvijG3/rZB
Glr/Xd/gg/XM2GwQ+Hc2/iTq13d6TEdW1xQwiwOjKRYmWB9OocZCpnQUJEycOkay
0ivoKm9ouVogveC1xZxO0PvBOFNZ5eG+LNWmUtxqnsjMWWGN2mWHJ0Pff775dafj
/+E3wuvRveZTTQAnDPVEIKcoIFf+R842XQdTz+sK9HgRIv7BXhf4xZnVXyy0Gw3N
9ye5n4Ec2ECUioMw5gys/UVVYSmN005OkvVwa80KKir5LtR7h2Hp6fFWw0KpGVoV
0jHD9vUkEMwdihIavw7jnQ91wa8XNU3yt/sem4tFICuWWAN2s0YMvRXgFfmfxgCf
cBDG3amNQb4w3/xOEb1fsKNFo3HTHxXc2FLuPnj7YGkU5mP/TsdMRU7YWG7paqYL
9LGAI1T9+POHWpwcPJh15Konf4zxBUIHJCmIsENeGt9+lU2A6b+76LxoF5yvKtqA
PBZ6SKhnfS9kyqN3+3cDBMCTkk9uWir8/JT69KH0Yl2OzSLrhOoP01Mc/sMeNnQL
iX7nTVuR0w+ZC+dj+I0z5NtXcX6y7eLoT98tj5/mj2xG6b398SgPx4mv5hCa8tUQ
AYQkykRdGgTSc+LprdxkHY+IOkfOEVcLTtBwvx1Jb5KsqzpaAupWKZ+mQvCLMY3V
Zu/rZLFLpX0IZOOwm6OyDuMi7Nb7cddUuh10hCpWXVyaSno1mgzeGyeFXz7Ii7MN
cUiAIuN+fBKEtpkOnaNkQ6AH8kPFkhFvAaoYoj7TIJ5Uu3WA0US6k5K6MedYP9Px
6umWkiX8XGhJEEEQ0/9HnZjLZQ0ZWgHVhclMNuHdHjxEX0z3M5SMwT7AXaZHeWJu
GkL7g3LrBdw2SWFH/o4FIq6B+V/qbpekPvzRmCVsTrQjDJ0U+GQ73MT5glQmg3tC
3d9hxNpZC+cqJyk6Fcbdv/LWqUmoxWtHRC5ew/YO5iXo962rAtbAZVmcYxfwxngK
XFYEGWFwz0d2oTiRHzIZ08nkL0sYBgOdre40W5HIpuh0NSWKbHa1MiwMUmC6ATrI
FLQHeaa6FwymxJxM6J8HlCvizwa6nyRFCQzXk3tRFekkbono6CpThdbNn1oRVWe5
IF0WzmuTmbhDnxHbtCMZ211cZBbHHjpGAD85m6inGrH9up0alrmndiuTI4aWMMhi
C9iUxt/B+HnT3/oo0BllLlKH6u/V94NNZJXn+DGeYpgDkf62vVHQ1U7XMZ1FsUAY
/+6HUmRhxt7KO9SzquqeaHnZexD7bxSvlHvGFFF75IY4BiRZ/93xeG6Iu4A2mXFr
K+dxK0Na04Zi/ciADgdNlbx7kQyuJ6psYKsRMaTIBtX7LITf2XyHj8RAgD2dfJqZ
nx8pgCLSJiupO2zpVGYjNF3l6m0BKaR26+E3ktwGbUZ4eEN7F+TSKl+UpUQ0kcpe
F0PHu9P8aLvSM8+96Cy6P0EBiNvzfX09SpBoLPXNuIcZaAg1kp+2xtHfgJtsEn7l
Y3a3LDuw7/YWtM0lUvISyQXL1zbj1IV1Bntw6SJDfxDnsUB2mRaHg0cTIm6GH7+j
AvZj3t6PeJXBf65tLPUHQv69XnJmWB8OPQUE7d1QlgQeA9YqfFFGuvtFGTYAYasw
aBlTEUWc5RO0OAjVTXDN7Y5FpJzNuApOcXJsrGPytY7jwxDNQInas1dLiyL2fFVr
r+9gVJYdA0g4krTw2Lxy0Uc/LuKhNv0TihoHkHKGzlHChOUliEF16h0fBvsP0gQ/
2Oedfcsvtd4iMzP7ley6osX1EnDYfZ7wBC9UEl7cWCtNkmHGiks0sv+4rFJMpAgf
1OjXgBceEf4yZM8nTmXlV9rA+tGJkSeCXLm6PNZ4LLz6b0zSkXQ8rBboL5ljaRKu
x20h1zDFQ0HymnKzVnz7BJ0cjk54X0dIxG4TbBuh+GQ6+GyKygaXicnx/BZxvmBc
Rz1cqEiyH7ENHTgxjgXY08wUJAvkEQ9++otIcGXHA4ji1FmzMMRRiz/+CVNxKxpO
yDIot9RfQarI3n+TtTvmjWeJsxDFXQ2TXUjcnPllczDzk48aNgVNeprKE9eSu1L/
Kzhj3ibCIpeVexX2joIcND68L15V9Ad0iJ+2y46yHFhBZJwWcvZftf98I4DduvKT
Vgk6KcrLGLANTYhEYdAoo8UV3qll8SOxcsRdCkPb6G/qAI6NMRPvaRzD0Bcj3RuK
pr5r76SOtOMdscT2sOLh5E9MyqHtBSwF90dHiSaU7tmQZ+x/TdrecWdJiuNpMKni
X5u4u8k70i7Gi+dx86wRDwvgIX7XJJJeoRCbqAbdK8Jh/wuuxgfhX0Y9NM48tPs7
/cxOJcXwRFRWHvfvjaVnrylc1qaEdBUnhFidkfRgdEnEMIdhmG/E5gMi2XA0AMDA
T5k7yPf6vmnHexf5LEq31nVcsF1MzVyyf3VpfRz0MZVTQsDbB/YXhnpzLZZbVjxP
Q5ksWjslKbj9jMt0/DtExmGFzjSQXLeaAx1P9nyoVi88eU36K/rKo2o8R0cS4zRg
vDnayQeWkfqLo/UPsUuiQMEudD+fDE/5+QJeJ2TL8TP6i/2uLeJTll/T0mlTz/Yp
++AmCVYua2oA4GvTfvpuj0PYMnUlssHKiyd+PX0kVsTnCUTGDIaP5awPv2Z99Iq5
SEykYubS7kRml/2oIM3mZ4OJki+hhdzAfnXaeyinLqv26dE/pn4zJVPu2oP6+31I
aJ57yufdFAZJWffEFAK9KlWM0zQDy9jyuEQJV5SX2Fs6zKf/JQsusNLWg+5azLd9
ReEQ8k2P9DclZVedbOthSH5eBMNUGJfDiPq172rYcxM00cjV3Urv7Q1J/U0EVbMz
QtyOLY3lqbhF5Ps7Omq9hMFT52pLllpI/jCzcToMM3XkzVTQO4EudS1tYjIFcaRc
d1YvnAoKXdrUcTSzjSjUAYgbOA4mtnY9Ekfmc39sQRDj2/BML5TaIfz8G4Kk3QdG
u6ZMxirFnOFm/LupPzFO3YasHVfBdLxDJzP7IsaAzCoIqldnzt7DHDz0eXJxD4ZY
FHuFl6k02rPZcyXLVdrI3JOG1phiq/Pz9x67ZYGlujj4QJHeXXWmTwW5xe5vIp8X
P9dP/Z9z4bLuzv/EmvGx4d02jA0bI3ygmarJqA9Wa2dzTCGmt8O/3nEpGjprEBig
nfQHk6xcBg/inkoTYt6SWFeLRlRIlwpB9iJ9kqz0WqNCkAnD9JHmGEhVhTpZZCDI
vHcHr2c+jUr1IP6KNbcDLaRhDIn5t4UMf2UqDGxL9JqKPoJd6e2FKcofTnTvbujv
382rXbYrC92vnUWo9wrS1/pAhRfo4fsO2JkNZwFWvfjAkPXXFZXVO9iGVSZu4616
cxcmdCniXQKspZQue8r184GZiiLNineC/b2gdknmEGT0qvQVLaEVR9eg4KWEdury
jcq+he4nBugRB6LK5OjDItQpwqFfAbFQv18YTuDDvODBAppAaE69sGf291nybt0G
EYntO+muUi1O7nMJSRXsm6U2c+uQdCOSJuhdKXhy52SlcOn0ILJmdnh6TMfBulqH
rDZh1vLGOxtUYDHprScRw0BV5w+tzGUQNk8urU1PLh/vQamERE/7X8gJQqJchLfL
3R2+VOsBr6C27Akf1CqitRSZJSmflkmPoILcVvEm9I/4oKA7YVs/gVAlRy7Xzvzy
yZeveIxLdFsLz1QA2yuf0xBXqXiV8dvdlZEmXaqrRgawt0w0+hO0pgHsUr0s+Zff
eA9sHxnxYS/KAu/kp0nJCXN3Jz2DUguXhap5Yhb7+eoMvDO2tVrf9hVu3kgMfvxT
UCrboPKW9aVb5jaNylR4ddMaNu5Wl4ZxXLPKvlAUAX/V6szG58jYfv9z6f+safqs
jUKbCahEN+z2nyDpNLo/v2uB80pjgrsqaTlNAJHbsF/0ukzOa0IoIF116yXSjtZx
eSvbDJFPojOJd39yAA1UsIqW6eNBCwNHBTagtCbTEUnbhi4KIRzirHMrcZWr0J8F
pB/LO+12hgJhVq133rjiFXaMid4voeVMCAExTcxSv55RgxFzHh+KouoFaqzsBwhT
xRSr3IJDJv/m4qbEFl2oIL6ztxLDRum7TF7+BdHSz0siYhlhGIgH8abaEhlSV4E/
WEJ/bt5gvZKg4C0C3T5thx5S8Zby7a4x2dvCIcNgwhP98B0UaIAQUhzs28wU5C7x
eZl2G9meWuFO84P/b7YqrTLH63tQJkN6Ln6rWTeZoWohd+aFFlCZ9OqtpAwWuzqp
5gA8pCOrpxM/wEyvn/MYxVyvcaJJZ1xN9qMeCVPLYGhNJ1Quy4wvQzJiX80T6h+G
ndE2FRmFlQeoTmysjtbuobPKKyCHvkz5ztvhJtBo60UsxNKPcPCkKQw2Uah//HZa
UCitFYDvJsImihQuEKYPKyQrXJi0QcTw7SHf/6I+qsYr3ffFTyDpYSBwRLwh+2uz
gJVcQB8PlmjC6NA2b9eDBHtYfpneLSDUswS6mXaFKmI+UdGH+EdbV/9XymrhZ/5w
glEYY9MfnYMt94ftI1pD0TFkz6KWJHZ6P7uFmeDsO7EprhWEu2nDIvT1fAdJZsEM
DNmEB4MgOCrbDTKlEVvntlV0MiR2XtDAbDW+X9DZ38RevxAyDsU66Xp3wPtTkgcz
qGMJXrHCMDYnxXfPXjSWDzUoaq+mnBEX/Bn8YKBEfisUZOgWc9saTiJC2fuLMfDl
HUeZpTyfVtB9IqeIwM9Xe9FVFZmqHq+ezDlDlOQ+kn2+mtcRSdCis+J/4Coo0QAH
91TeiIIZGzoEH9gyGgmuxL39DoyqL4o73rrGA9w14078nbzfgI13rkvsOeHaBILP
JwtyVVRjh4rjBKr4glpOLjGQ30QNmAB4GVWkELCN/Mb+GeHkrpw+sgd/b94gr3pm
UEkSOA4g5R1cjD338gA1Lz9v0RqX0DtD+QnC3T4z8QRiqEeZkdM6QiA4CEY5OgGA
TzLaqwbqNaj9zphIjcbgriABBzvZAcWbFkl88b4xe5PNj1mvCoYTfJXKYQSyStH9
WxITi/ELMujYpO5Vsv+4+ODDRZ6UHRQE/mBCgAIeUUGSHd/p+R93qkQ0ZTtUgzTN
/84toTcDx23zCHp090RQr34OB+02pfYcvMUxma8V5tVHH5sUyeCQCQW1XXvKJpki
38RXAlMTP7ylxiHamYSieCqrSFs9V8OR7tacLPVzmkLqmRM0FpahJkZXG6QnpseO
dR+bV6+kW5bdTETy5nUkZWlnjjep7czidCsHcS8cD1RTLcbWRBSulHzMCA53xvOT
T+5toO7yULrRsEX4vMAHDSa3IZubQ5/f244BCGZGxxZKrUZA7GRYQwAD7KsQ8ju3
BQAWriKhT1LWhpVNUPI2t11ITUywwutcyEMrjbbRYHTrETp54/B2EWGkyMjaYx8t
hFYy1326stF1eYR/veWAJrnfe8GDVGz8RjU4J46fO4cZ16tdbPNeRrWGUsma7BLY
XFkzMpiP5Xt31fY1m/60peQ+V2ycGpVqVY7i4VVehNOMTlMT4WVVTAVVkU8ruZKD
8PC+AWJO5v0OpmuuAm113fOXII8gb2BgyLtXmR2FkHjVjLw3qIM/yNSgZKYHWAj0
99F8KABDhPs5TClXp4yVZ5UwntCh+E/lx6ZpdFYcIyJVoJo3/obmYarh+H0lodNO
BpNjDD97OUQuMowdjFF7Uv3rPSkQuQ6KVI78fVGr6p6eVdVn5PsZl/tvlaN7km7W
YARS3g15vG+8oRhWYcyrjjNvDYeqRF5WzsfxIDQfOcXAn3y3lzs+wlsCZVFPfVMy
t3odYXphZszCX/H1eMgnB5hM6IEzPP6OQbMtn34BdYS5lVegywwJxtw/uit/3fvU
GW3gfBD0vG9XQcqdQvb3gmEmTVQuBBkdoxceT6Krrl78lVr+NsXMgEtdpTJMR1cY
adUNRErgI2q9fRi5y/Wix1825gBeE6xETWN1RVQ4iESHxdraYdPM58eH71KDqjf2
8tXOeMPdFAg/56kHgHn4eZ6SUAe5b8PXVHQur73PtlMYMEIn/CT4x9fpYvPppGdv
/L+8RGwhp5CfNf6cKnpUqCrexZc0urDLHoG7dc7W/zBf05m6RtMtEUF3RNYKGeDy
H1QljOXRKT8J5F8s6D1i0JXJ2FEPMXW04bGq3+mXcmQ8TdCZulbme0DVayKi6Inu
uAc41Z5v52SD93n2cvzfIN+RIpcZXFvjb5xZqAH/crM4NcBYUPYkJpbRQV/tZ6ZI
/pO42noKezaxARMH9jHsebUQihEpjeUo3C4fUaOm/Pyddsu28fgVqMXfp2qlj1Ny
qwG9hpSoZcvJIgFSUOZahISODHeFqe+NtI4SuKYEe5cZEQ0BvmpOIY+6RsrGnNyk
jEfri2DND68/TGvlxKReEvvopHsO5nrTHSB/W/XtnycADE/ysw7u+6bqgp+5uDxk
iy446tCVIXQaWcZX+AP1epe2Qb/P222gELzncyqxe5htijstigaiFvFSVmnvM/Dj
xc/wGj6HJgOWJAWDKKUmiH6M6sCdJE5uW9ROr9f5FAaTCEWDAJoU42tGDkr7BS4j
+jmGLYTtU320ZhS4f4OmY6YkgUcsJQhln5uif8CB7ef8zy1tkRQc+NRR39LXOVum
mRro4HJtSsRwjVkMeApZhjBtPdo9JTHeHwKEn4mj3I+gY63oufPm8qhvVrisk1rC
uV3JS8BCfIR5U4bIWqxYOegStOemLDZkyOEo8vR7O5cgp7ByoEcPOE+EeZ0JE+gB
WxZ+myomnhyJZ+I3Zj8JpEwkeOjZJJAGYXBu23JyCtKefYsRiBiQzI7l/SFOZWv+
LJlKIt+FvCpAxH2L81R/A+f5rA24Wbuwi1tgApvK+4PEfJj9g8XCGjpBxQYwjuNy
4num0Ya7xEFKXgBnLhvAl/J59MQwX1gXucciVtIM1Buh4lcFHJWynGdFQes3CPOW
2yZzF5nlYQdigUrB5jd6Una144eWng/Brmnv6gCsaNjC7o0rWfvGLRYvqw0E13e1
J22F8r325SPo0Qc3KnRrUUSIEM9LiAQ/xCBPmdv83RBphe5A+S+yDTbyMfr4oJ0O
/0Ra7w5JmKrswHgbuURB38HNkFJPHLIuhMXwxgeog/Vi/wn3cNtFWerDNc+dt6G4
nP2EZQ+w1gKJZzE8olFKb3W3LPXXSDNhojoaattvgY5+L+l11U6W+6tLdK/9JVzE
qF6tcMnTuDj11h3u5O8iEbIaAb7kyDP2RmgSQsW28hd1u8TAQbR8InD+mu4RsszY
vN0Q9OkDhrCxf6ZXFTPZeEB3hPkVl1b0vZbkC4kT7Jn5zKk17sbptLpe+w9BXrp0
pE4eSQ1cpH93k6FtJ1RwfZeno+VcSehI0E9xhpfl8nwgjz1zluod24E/R9ngrc9y
52BzA1IBLZjtZ40nD/+cVFc8nB/q0TnT5ATqfu4pd23vJaqzrfeGyrqLtcbeA0EZ
etXUCL3PqCh1Zb6Kc5M9OxrQwj0NMTiRcLK3CrMVF7NM+HmNe2eAAXJRydt5Bh9e
z9XsboRHNXIbfkYOGVWnRL+Vu08fBMPWGDtZuFXgIhq7xRDvM6eKgSae7wZZVoUy
uwFzyTfFugptVWfS9KJnyruVK2AbsyjB6KLpOErOsvQO3k6LkfIvB5XIsuDEvcL/
Vay/nphwfhQwFAPOJnnM1GOiA8TXLam1SpHg+MRdzof2oBpK5SoCoq71iAVENesv
ZA4/hhy6oanB5o9WOmqb0Nmpf1T55R3OmJFJZGfztKduMiiCvMf7OSvrfnj/FlOM
iyoDN5HD2MExTtG0Y9FwVqAw2OBUBPKV6TMiz+AUZ4YMbBH6wjNAi+SCTfZkQzt/
CqI1gjBD99nXcH+bCsx5+18Dh5J+zxpZ49DiW+eSnY0giE0RzZ7FUw0n8/xwIOC1
Lh3RUcco+5rsWdm4Z3MYAymKeinPREDpkaqeVbPuGB5p3yxvd/w89lY7t9wVDdrZ
++/ilYqV1cseVzA+MxVWYicyOZDHK2Uuxau4pol1ypqq9Byhb8uxfn5PhRTqjmM9
dFtLajPBpDmTIxR5AhHsRRVUZdYFDuaD1FwXqWxwLDY820t2Uhrz00DHu1H+8Y/D
mI0LNUw4LodGppuEkRyC/9LtHyPrUpuISq3Mmlm/AcAlNs0AdtewHF3chHDo+urb
++Z7Dq7mz4z/qytockfNJWiohpVsUomcD3+XJ212/mShaoQ3rpslFjZq/58iHFll
njHfzx+//1iVpo+OW1Z8y3iCwz/7+70FZV7/Gkn/VcxfspGDskTJdbHDpt8SA6/A
4GTHOLmmWVrXoYsWOnL7+tKMwdL0n6WkCo9ttDINGtCuJ51seZq5vH8yShcck5D+
lelclpYqhTHOr8ak1KKNGcHFXr1UHKVYjT1tVs1QCSSl34qe/58jR/YEkEwJZpa+
N8adVsYD2PrglWySDK19X2KfidAhTO+5QBU4ANshH39+DAGbXvHwdV/v+4sQHMtK
TsGpK7rGnA6DjGD7+wZeRSnQiEpSJ8pfzDYycQmqGlnT4Oa2d8mipXbzZ8DEuHZc
S9O6OoAylNDNA3/cQ5wgZw/ERDx1oI1KNb2ea4pZSHSMYnkM/kPWXnFIOHfNrbqH
vUDp+T2YbDvPBC83g4AmfRfz17306y8pwwHzW5MNla1ApSfGZoEtWtAtoACoQeq0
xv4iJlsI6TvTFgpkufyWyaY3ffE5MLmODd6RVkJkHuPgBhJ5d0RfGsVsH87OtEc0
N4o6vUHUwJ7iBQjWhGn3TI+bSzJyue/N5MS0mrNpsenrkMrSlCgDflIH/P+ml06Q
9YRvZ9WeBEjfTW5ribaPIpa3Xc3ba3lZP5JstTioFGO1GnxGoAQAFjQc6poXzYiB
mxYYWE6QZJuQbzoxw8RpKZgnszizgykwBwqnADd5qhDYdusmrnezEs0FdcdlGo5w
wGlvvZJnATNlHIH1d/Z9Ah4FO6sJr8vYty/2/WbsMvJhsRouQXXApaJ7fuJTawkv
aWrECwoDyxOorZKRXr+A9LSbTwp+NFuVhKt1tgJ1ENP0S4IlHA7VA9zPSgHIiZNU
yKxLWwUlvLV94MeSpMKqfCnJtS+y/KVSIC0kun9IU0G/qoKfyCpmbOR8Fl9phM64
barHcJcYH2b6kXCd0uETYu7mLZdsFYRAuWemtcOVz/WEyjOKShXLuJ9+nHiPP1Dg
mEskZ66+NH+WgDtORL0pFSozVNN4B/wtnF3ek1OFGS9HRoxO8Jjvd5xqtBbps2Og
WazCP60yWWqdxKQoKrOmlPylcy8eNE7IiOWZtclPuok72TIqPEgzWTjnbJNTr+tL
mzFDy1r0638KL5ivmivTSA6ru9qqPUIvNLELKYX0c+IQyibg1St9YfGXGSRQJJdL
ljSeOyCWT2Zn+7NBHTxlOo89dj6+4eCXuEQ7hVKXdxsdehOJB8PBcoMLjCVDs1CZ
ItfzSDix0iPaiMatNMJd9trCk/rX5aAK/L1NI9ayQjXMiUet7H3DCDbNa1GF9Txi
eGPAucZGn6i60aJMxWTOWVIIR6bI37xvE8NLqbNMhDHBddE16hwCZrboZt1B3Ni8
SX3cA+cOIE0o2bP35m3xZRLP+2Eb4e64MPDWkYnzCEfuHPLkVQR2aAR8pHt00/a0
oNqt6hbX4WjZQNg0nLJO8tfxEjKAN1zIGE7cbSSaGQfH3dOIz1BRmOhg/6G+OBtC
x1VHFU93GfCKJr59YMk/+uLSLo2lskRjBdPpkla4IixPklC0MdUFIDct0dxVVZ9t
hp/FlHLtMsDz+ATqMVkFds4JTdLjfEIH5p8hmOH/xIb294ri3mCrrQbQq7iQu097
/dadKnWbWnH1V5BUrSNcMkE2Igi8IYNHjkMRv5OHzrBTQV2W+HRFdVjjitp2boYF
wRLRbLBJ2D+QxQOoog80ulzdWwhOB4SqG2jtq2tmNFEytYBbt2K3tkqHnBLhXRGZ
sWIBFcAVw0OCMETEDu3f7AlQ+MHduV7VLz6nvgX0VqYH1g5oTp/OHXLlgG+cr5NI
823r8hduQU3ujshS/6NY6KVdZj2YIx1NDymvdND0dS4oLYYNbz9ZL9gvIuz5suG+
x/zgYIq71dpbfI0SM9f2w6+6qroF7wej6N3iyW9ucs6iCHdRTtQpJDFLWuruuyDS
K/yBb5UKrUTKobFDpZRa9TUqfkSMIcjen1qCKp8idFSkezFVspsgS0E62wYA14Jm
T8sDxxbjF/pYszktOAvWpg8Oiv8H07y2qGJNhJbG0+IpEbmbk13OaBZLOI1xwMeX
sPeJOKbYxXMGfnnhmaj2LBfYhSYX+ozYRPayBAsLLmNgbCdmw48u7bbkKVUnaGsS
HfCh23jAHfrgdiGZbWjQqOnGtPy3aeP/hE1IptLRKYLyi3PaTTzGq+WHcmHyYudd
SoWv4gHDo8RKqdI0GbpQtbxUbWedNpPT85CN7gUudPpo1Q5IGeS7wnc42JtbXnsL
FF8y5U7Jqc/H6T1tOZ4jaZQLugX46Bbfj9gPQmeYSezVcXn69cFAtGpIiH0z5E4+
QLX0FnHmKPrX+Q3mEtfDcDvBmTqrt6DDVqJTWHI/Q4NDT33chLw2iVA3VB4ILaed
SzKRRY1Rn+smy01I3ahCf821Xft6VY0PNDfwUjcop121ZQnFF0VcZ4cSi4xgvHpN
uJJqGl8WqRPBLVuaAfo0u0jvGFsgIAlxmsFcLagCy7LvllP0Sc9cVlxCQYgUDt0z
C5HxrD8xXeOH0Osr3bN09OmXV9gmQp1f9vQ6ANUoEIrwax86+oFMPQOslJC1K7Hh
sUXjwrTtSwaNPN0XY5or9cDNbnjnJZOmP1CmdJUqkZQS8vwUkd1B7MZbEPbGKA3z
+dmbCpR7n9Pg+ZehnDMR/xIcB+/eJ4dHNOlvfiRdaJPm/JsloOVuOgqArctHUKhi
45gK6BKRBY3LsGy7o4x9wK3l+n8fab2BVnMn/LBAMxCcIJcXbTJBzdSxCZQb04bf
fa4zCHgQFHeyQXhLYM0BMdKbhMKlzur3Sl0cvJHEgoE1bEzaWDteMtXknNXAYkD2
TaleDItFTEk6lQrjP5i5739vIvJIw9B/dsBM5G+Cj5nyd3HahK5NZp3+eCAuhN16
1KUpo1GLNPSJ8vXy+dKlPb9IPKHt7OOWSMez43ZUCP1WWURnnoz9TY0C1GLOe4pv
qOrkraU49remXTrmMCMgzOLuWinyoBh7TOJQGFRyFOygaQppR5Ednx6TibNVaHi9
luFp0O4OLdKffaeTEtAouMo37BmxwzC/Rbza3itkhpM1YfM+DA0BW2C6NDeI9IDK
S40/qgJBoI6YshIaOTsKAkg5aqvC9bKhGLWQTv1/gMmaw3a7Wz8w2UNO+/Raqd0+
nRYKTF3MWPdRHGT9w+c9/w3ISrt/ap0KjxcIBlq+8AUefwI2wPrwmq8ZA//uWasH
PR1jz2o+XTMdmVjGU3ARRoDVrhmGPJO6uDGxavzhD1DsxI8VWiFEdgKdYlnAo3XS
f5yw17C86hpss0RS4kNhBRBCNfVFTvMi+3SgOhVQBeMZFvaWoabHAwf6Yy9RS2Zv
YQ3eDMahD+2yCQcXyBNU2zqOnWN341qCgedGkNhx/8lIJf/BMnL2GQv4I3vG5p95
GRmbjIEn+j5agWRF5hpxMBM5iestf/soG3YOH/Kwyq3JOKz0FePXd/zkq5emFz0u
7rPA7nONXSsdbs33nYTbzwLSRs/bZe3BzUqtbCuxMD9OUi7h5/rGlJ7UXfGSS2Ay
ziLdBWCOKkuvl1pYs0AOiKHRTeQuGGvo+Iqy3UL313DD6LNLEh/TBlUZUs77ILPO
cinab3AHyBJBsBeIifAeOvC4wxl3cjjuVwbn54RcdW7Qrzhd7yy+LhbLpD0cAeun
4TGIebPUbl2XsHuhi5du43mbFZManQqokXx/w7E6YpdEevVay9H+lnxEkNNRBfh1
jdO7s/dq2u6Ad4dkdVp8MsjJ01ii3Ucgq6dFK4S0MRSj9cvOI5Tbcb6YmChfaROD
cSzF88i+2oXhpxLfgp+Adc2+y+BORwvInikJPbBOiiwwKkSpisYamHqGDfihni1u
/Lxzy+4FDE648mKn8uFkk6PMnV6TJn98NJ42MQxnypgWD+BKNkZLKgmiHV6l+EEr
QcQOtuv5YtEaIdj1VitPS793Lbk2Gf4WvikAG0sz6uE8vOpEINC3VGNcMnnAWnWJ
9xBUju2Bzs+k8gZLg2EM2ehzFWJs7qHTT2+r30PuZLXY0l/QNfz4LAVxOi02P1re
Os62Uwm/RRicwyiAgcwCy7QMMs8aZrDfpi0zR+gZ5Dmaben1LBgLFVfZvWXAQIRK
fx2/9vJYXkKAW9LTz9C/3e1mPi8905r2MPslnvegx7XyZS/l9Kg3qr/8PtlhC0iI
rOpuptF3ogM7psiGbdScX0HXF8RVdm1K1qByFvpFTklCOFN9RlRwRgxhu1tOQnxj
YBd0pG0a/YZ+2+alsVR/MzbBiF5LnGHz6TWsopuR4iG2U9z4UrY4fDoQ6QXwbqij
EmBKu2I6hCfvNIa2I2Ls3Ch+LzhPT3kAY5cJLCr4l39vJ3aNa2d47qX1/eWzsNNU
chfLE6g9kCOb/qkbhnDVG13jxpD0LDC8o8HSKBZ8yDbcnLpkqKNc1LL44ekH0Hle
aatgahkQJW7jVfVgZQiHcUCAPLDuC3UQdtO94iK+D3rUmVP1UF3hfNWWUxLph1W3
X1V6MAuZJJOOEH0R2vfP5QPAeu72/lGVXqrw6ZS/Uuyprtjam9SD6fgfJfG5iKzj
7NY/QFAZK7yiTDlgiLHfCpFo0zcdthS3d94Q3mqX/SnCRwEqzzS7PD1yzoFRv5Q8
Chpj8333BzuJOCXBjaFNfpleZhbP/e2pF3itMPafaHbrbiKawCxNUxO0Wi6J7aIX
HJIU8eq8KM6UcfZEloAG9isA+7TFqCugLmw/Qc2H16vPS25VefB7UfK8++ulnR5r
Qxgk3DTtL9Y3kUQMSpxIspgxwgD1z8V2f5QhdDnpiiGnLZHkcFh2u/4AUm+rr2cw
O8g/8Haofq36y4MeMAQzbYs6zIVjLf09QeExIp1tjASIZ4CT/cejVhFXrA1+K0sH
fqNTFqBjsVBj0Lt//14rTZgdnDVLaqC8U6XMU3nn4+WU1KwBA6k/9qvX+sjZPAoi
AkhBWeGwJF5XPJthpnVaoQ0DedOPWyZEWZB9WBJ6t8Tk0VPX/WOgiLbZ+UKZ/7En
HpKX4BXHixP+FhknCZICPnnVr+x88YQ60aY0nAZvgMD5ocknT7A1ZiPE5oCVs72A
/jaNWsxkAycmZNXOpa1F+v7WzzxA1jIHO1pJdCbKrf0YOtDVrcolVzzFun23yhg/
QuAwfw7ngoJYRhvuQ/7eI0p+CmVugwAXeVDvWXQFnvfeTjIbGG80xZKT7e8cDl5h
JglWfAFxrM+rF0DbqGA5OKzlLFBKWdpX0ukMRFtbEKs1RMvjVIpfBoWISjHj+ACU
tZ/6dkI9uxU4vRBi7QSkCZ/pbqM3mz8/KiF1/CNJiJHe95H6t/8yPpTq4n7Y0WTh
yy2B6d3WaW3ed1Sane6KT1s9nj3LUA66xltC5xPF2fOMKA5y960F3eBtUcreDy7X
tI0cFCWs/QQmmXHM03A5EexHro3hm6fWyelwIoQAY9e9iSYG10XD9akBZSaiMlor
a74hVf4rnyKaW6QEv3OY5KpIOfQoDvoiB/hOqJqBnChNZ86Rwc2yihnJ04t8CGNP
ZBGs7OZu66X3lxOl3x/J23tEoV1qbvWfdNziU5VV/X3HdCH7ayv4XmtKlTP0Kn18
lYGPbeUZGfsLCKrOOSNWSCRT7JseTeEiIT65wRDsRupu5eeVo9RR81eeyEg73crT
1qzXjfQAT0w6w0cjo4Np4gmtk4Q/PRB//i9hB+tr/swfQgDuawhvmXt5X6KuOMaX
NumNMpoz15FGjQOzur0b10gfmWfXJKjUMEEh1sMW+Z4IU5YOphIP+CvBHWChTu1J
Yzk60evjI+yxmKGqy104S+15ZW9u5PfQLgxlXYZALSfr1RKC0Prz2F0x4H0GFLRI
N2ql/cBCpjjsqb/UzSW9tSxXoEZwStsjVYQcPwNm2YPLyrBIvSdXQdq+vJdbAyTB
hH2EOmReS2fKyBvoSyswy8YZWBHYW1hA3PtndqnxZPda+dv0UxKGphZ8D9rxr/X9
vBi7LGcZCbamcZ3hYH/hZukcjPnaCvbtJ7ZG8lwztmRXl2n3ow4F3roMkWgNTuRf
dRWeKAKUss4gDuat3hGWktxGWGM5zKKT++OkgEVHmw0pMZP+tfxxX5RDZR3N1fR3
mNMYaqfUAT3dCriEubP2hzLfuKM2bJtR4UDplWEypDFQJdA6XxUMzsVbATrWSgvi
iSEFJYTnEX7oSzr43/wFG42fdZ442e2A72Pp0FbbwAKPlzpWSM+OylRKhyDa4LPA
40Nvw1C6pld7trvpdmVcB+VPlclcqWyZZm4TZuyxAgCX2o3GLlNEm328Q2qn6vB1
nlO8CCqpxBtpBr4klkuDb+VwUBNbSPoQeP0Ne5/4bqmeEdY2vru4pFQ9gvmJ3F4K
xoLfO8HVXjiWN1Rt3+8mTMLQcCbafIZdy07OQtUziMRB3rB4op7c/etlWrLaPtUj
gKaCapL8R7siTmzVGIlQfsze0iEfSxdjxkKPycQgk+bNVUpp1xeAxhncUB6R7e4B
7eifUr61luICihFWwcS6xzj8W6Au9JgcRMDWEBJeQaKSLrL2hefch7iP9W8j+S+m
8uvFZtpqT0ELvVoVvZzfTbWykxkx/rWtbYD/UzfLFEErDSv7n2BPhGdlNKhTQA2+
CIEoVKE66PnIShFu/QgD+GuzTuqum3Jb/aJiBfuC1zPGy55xXIkrL8zkyLsy5/tM
oCA6dG9rCJ24Fr+gVg03dWJLv1mZ0/zJTGW2h1UqAGd7bXjHk7H8liFHM+ieX1MA
RAR56jWPvNjUrbXXRXvQGzBjgAFddeelmZ+NL3XEtg8GHOKEHbwWnHwdSIVXIgDQ
OqayNMmCh5ADIf8SfvxpOIQbQjxccjYF9MtRprS7ccSjBqEjJi1byKWcNDYp8n8Z
kuyxZG11dt2eSpp50aS1fpnFieeIlLXLfeHeK+MZZvMoaVequrEGc0HQjGsUAUik
BqeJFzBTF8UbEUK9NN7SDv66dfZmuZ7X7ZjN+DM/G6gHlBHHfm+ewRyz3zScqbsl
Mped19rUZI2WSrk2qJSA6M77okf8QD31uY8qd9mhgtjcVGs2ZIMaa8jkwPAuStJr
vPGIkqTJDi9JN6Scl4MNDf0p/uFN/9b3CaxW92HpzCkTz3r5x7CAo3CRW6NmzYY7
9yDsu1LOeLI0gAnLmdLIrDCX3PHpQhEPI7Na+g4hKZU9dd6h8dnnbEiESudr7u6H
5ChIkB6BkIYvImCcFntskf4jM5MWXNM8YACoDbFpXlMEnUa/R7Uqga+UvUSr6MrQ
tcKEN54BS+OukKEAUwcUo4uSNydla9H0oDJiuStU24iYO8BRdkF7YIP8rFeB88KU
EFA3maq0QymKF/XHvox5+rE7zPvrD2Y2eC6UnNi8WGjOfvEtfog3eQuRBFPMhZev
0wxCQyz7ISvsFcwhnqGehzOQXbj3ZgdfLpyWPY7IqWozF0f2UHxFgmJHwEHcgQ6H
cihY6mwRvLsrtQxHEz/HWRsbb0M/H5RgnD2dkQoKi3Xk7p8WJcIAh5fk3kdcOFqf
fq29DQ8DTshBqCQ0iEqEiMfp/pIHuctWm1VVbH0+SSrgm7LHP7YpCz88e60usnlC
BuRYAZzkwL60Zw928Z+zijgNSbYs8KMYsgQ2Rr6/Vgn/AOBh/3RX9CPXNGh+Ij2A
4quU8/pJb5Cqu3Emu1xglPgLDY2VwRU5yFB9xNfdfr82usrLoMGjBnG51e635/zp
2ZRUBJ9IUOBC7pN7jTD+Sb05HFxf36cS4corBjTTgnG08ET3p6kt6QdlZ8bMLWKh
ltWAIq4UwqnXNFQUN5R0GohpC1ikiCviKKsbeWv6khEmtpFPfT5mEv2N9RSFuGtF
hTPN4eXJPpHYm/rwQ/F0fFhQB8EOHiQi1TNiP5fImws9XoByEMwHsYAKg4P+M+vm
0f/xFuhlFKhvKC5BrvHKkn9S+4+kCKnca5VCiJg3wLLsa+vQmNve8cbJXettqxD4
2xufGWxd537MjBDfo1CF9ztjEiEAt0kFbG+t4yegf8bSlVe8qEpZQ59LOvblP8EW
G0NFr92gLsr0jsZXRHXnwj8LKB4Sq88bu5VH7FO+RYTvfsgC1yHNgUCwjhLU10vV
FhBne4gseVMsLmeJqXOgGjgKZUnhXhuIXpVSChVUIUNRbi7FL+cAtwA/a7pTlyt4
ZJSlSLrrHKbJgj20E25LOvJeVUBcLtr+90SWMvvHctW+HyllRCaIXwXxMYyBv+o7
p+4kkvLAj5R2hZFJWhRhyKPOVs2MPWn0UfLyuERvQXqEBoyhxX7k3GAujhK6mZJG
E9ndKKDb+IS1xsWcYb9y6UNNYeV1YJGDYgWq1ufW1PeX411Yus9lphMlX/gg/ZSv
yV+i7wfJwON2GZf1CBEQ/pXhkE6FIQ7euJ4Hc2xoHiHa/Z5AVSFwbWZBuHBE5p8n
8758doC4XQCOVtwRR+h3QM1OnAUXbsJ25c2VVneJzDVchbRDKMme+eoMWQOsmhqP
AB41ECCSxPHHl0+J9N83uPnFTQOfCv6bererSufsjnmntsPI6LrMOb6tSSyAxkcS
OBDJ3zQRwNyRXOuMHEdXj+FOBYVTT+pCS4AuIWzLgIg0lr8vVDedxoidOKXy94xK
/6WVZ6HzxCG4eH9H5L/R6nArW2Om22Ttuqwn5zlh6Ehqd48jhaMpQ6CX/hGZLkVU
DhJMv/U3TUxrXM5B+eksXAfYkAdzgkbMjjQwz2qldMAxNXt/VvJNSr1d3F01iY3S
EVXbYuZ9uon27zGZ5Od6INUYmzR6Ygaouyp1cO9AE5O4PKnLCBWC03v+CVX0OJf1
G7CBIym1ExuydkYQee/Ui6Qrezv+WD6zPWU7ZJArW+6rpCz+Pi0TAcbAwpqVlKLa
OiLIVOCoeYor1MAlu0h0NVaNTmDtWD89Elc9upSq5bJJqtXPfPujTQA/IbXgn2P3
9xZb7KxWLnBGJ03KSbno6RbtbGJ0Jy8GHe0esbki0jEZxl2B75BvRTubS7RzLAIT
ZCNFh6WBETcaOPxbP/YPb0Rqi2BEdrl+pU4LntgPwpIfHz79xXdoRyChf0lwKYDF
eQ4R2V96Jtqsgam3aQqIkAgDeTzf/lMg0PM4YP889Wss3x8PzCpS9q4qr/yuzxY5
DinG/e5wyklDt9CkyRdFDG//sUDJVcSQ5p+GSgA3OLIOGB0eoaIrfgObSl18yL2h
ODIkg3GYR5+d/Z2Elg4KNG8KqaYguT60I74CT7juWQb4D2Za6nu4CjqRu0AajbjP
t0Z195LXCn+VkEII42g3+82RtuYS7LE6EphqR2f/q6+bhQRL++UeUYxv0mkTIqDU
ZzShx7ugqumjvWuTkj6on3Mdy0+/kTbqjt0WnR6NtPETC3GKuZMwpVBaYGgWe3Qz
yPftH8RmpQlfUi4XQhlWvd0WBBpySWdY1SQdaJU1ajP/Ka7bMvpWXIZ+bw91qfjI
ve4tXo+Y2RZHVphGmVtBzsIW/X67IbVCPuHu8xLKhljn2iWWblOnL6Gcgmv/7Q3l
T1VNTw2zkiFkM5YTlCcPZevB6VDkY/m5YprNXnpFjdkvnyTvc3BcPu/kfUn+q0rD
ATZFoNfC8ba+VpMLBmupLfzjwSOehK2YWlKrwvJH0TuiZGNa0uCKI7s8vQsP2Md9
DQMtoQXk7jxh45tYVNzz0viIcTzGLJEPgpcrE96834cQMiUAzMDO1fzcMj3OQDFx
2qCp7s9ydGqeh04RV8y35lnx0YQndPw/qOSRz3FecKXcaN5NPFJzMwhb9Hy9hlBx
Vju2BGl+u8Xs4RF5aZW5U/s/s4gkmR8bBXAIuGX4l8eskHweU5AUIkyMXYUttSbd
S716DueYDSYiC/MbfIO/KALm6lJ5REUHzPObRj+++qhHmlLNK2afYU1jiqAd+1LB
+g9q0+4indf/kKs/wvk4nKlUnb6QxJD1vMlJtEX18YQ0bq4XKhVU/XuSQGcBiAaF
f/aChK0wGKUJG0Gd2UGVryF1EeevEOH0T9kHTpdEV4Iwxb78nwZ4K3r57PUPTOq3
x1j7TawNvvGCYPMlDtrWbYi0eF4ljrBRdI9FpuB9dgNyOuMIxX7GTpo/EuneOmfk
4iKa9tsg4KddzIU19QXcKZ1qeOJy9caAbazBSffFe4KX91RUu04irb67ejCUPwMn
zM01VhG1uTSXPTyOEWVOXvBZUj9z5+mlakgf3KCBOJIuo3BZepF6gLlSTxxwdJQH
rSpaE6MG03riAxKdCUVFkYhe4OymBHYf3knAJAk6b4dmHePC4oKwl00f0M9bVfKl
BJxMdxKr3UKB7d6nE3hIXw4jI/vyk1nzOQQIJ3T1Xq+AYYNytac+x0xvALbir6G0
2rB4bckzMciwuYhpO+1lU4/T04zrtJyxyqL7/O2Pnupkd1mkq9gOGGgzWoOHE9Ct
nyk94ovL7WCFiPUBxvLSRGVU1W/NlfKtqYVPIWAX8eOQNq1WtD88MJtBNC05ZSr4
wsoeKKX4VptwxcM+eLArtXg0B7Bo5u11wwV9vUeQPudjYAAQ8AF27R2LuC9xFTiP
EboYsbCFzRgcBukq9l6pZ+o+qS6NFEQKsMkQkgE5iVAKJHsW8J8UjCMpoMr7GG27
DsAguwf1m5HN7g4Jdvd/CjkAJdH6YzJAZnNRmbufRvSRNkwSR0wuaP4v31xGT52B
EOp6eFZyYIB3viv00l3SazpdyPGB6oUeQw1w4GyFGe7MErw7KAKsDutp+LLtOoLM
yShshBeHr38/Ybn2P/pXnT2vt2l4LWSzyLrtNbo7qIAjzhfMi4ZiRGNiP+eLdz1v
G1GIafIffoT7A2O6UCxHbv5ryu9jPGpdDBTM9jSxbdpdH0UM1RgYKdlxoU1Se6k5
LNkRJsBC89EoFvlaLzHcAMl2kJYN3O1O4J5azopp6gF2UdYYF6JzaZ/hRJDSlN/k
14/ToGWlnHC6B7CU/nbfS3Ybr0YZdKz+pA2uivpRCiD4CSVYAoGKVZ6yw/PD1ax9
cexDcyDnZpFTQ7TdUsq7Hq2+4zXW1Wtel2YnxNl2QA7QOlWqZebkyTDuiV09nIcY
KykOLmHEIH2ZXVbbXLWr0fObdVkp6CyOwRSEDCLEy6zHd7hlXUVNU4YcDUHvHJN9
jTzjdlaGqOdE2t7BYcsP4Fo395htHZZADPWWb2DqU2oVWAcStJwqElahuge36/Dr
gmXUYK3fqpGWaa3zrGKc4v7/ufGwe0Xh4bw5/+9K89y7jHwLlDfmUKl/xPxViZ/R
WImStgqJT5GNyjXrzcvoo3vPy0kGY10/LIFgvNqPI3BuJ9R+X6K68wiw/l+75+jz
YsdYUkXlVbJ3YWNb5vazuFYgIINwI3pnxKO5mDq+faTU9YG9UgioCpG5bdw3ikca
I3vNBnLdXD+ZBo9fQblErxGVG9QGYU1aZKtxSqrya81uoIx+m/s1Q6lig+Gy3LSP
O4M3CC6htUX4hw/3bpKFJPuO6qmHiNi0xVMeBvIMiGua7UPjSLfmDoKKx6eEn6/F
EFwmdrR/Q+69M8DqLugRWJaB/vPr6O5Ffz9CuwV5q79sxfE5KH0b7Vra87QHVMPV
A3ZK3LhSyRce4z8VHzOGWfiSHRyd8nNdcsMckf63hqlnwDwkRRWQ5X9KchWRaIIj
Gb+SKyAboBP4qMVywTHoRlEoYUeQggl/0Hb+RUA1wwZUh86h2lTWDoVYwerCG1kC
5Wawx30fLmwo6nYxlUyXs8wnpDbqSa3aHQSCJj1AKv8TBmpbxO1/C+ABUHDmUtVF
4thGVGbPBzvrn90LrqNROt0nnTOmlxTMSc44qR1C2ageZCsWTi+KLdmICwb+MDLd
wT1Wz1+bn5vFZ3ftVHLlWST0qmsy2sUyEfv9LC4z31ex94Cp40/u16T3O/n8wUET
3Z3tfuhbhss0OFofErF2bS/ViO4TDmsvZ+53ks+1B5wyujH0un7EocD1uunmeSbN
rH9ygHvyoHyEIJcj1cWK6duxj5uJMMzfk5CoClAuzhP7tC6hYrdYdJAMGcbEbSMn
2087FJQ3itpPGkXLKyThE0dv0NkNi7NT6F0PuShjS2+f3z+K3O1akAx7lSnyluO7
N7sOI9GwmnFp2pFcWo1ROHS8Jzm6+7nxlUdgV8aAh0JPys1uh3gQ/qfRvboaQriY
RjUPYep3sqrU9g5wWEAgMj5kiMmWmmAbCu5M+WaOe7lpRIxxfT4yLtN/JqNagNEz
5yiqfekYbMd/s8fbPmiqi/cMe7cMMeeAb91GbrCBBFUaKttCI0K3kijZqhGInoVV
irK5w9bvgBO0SmV0lqmdFHqavTrdFb5F9g/7m+wqqcUXl+y5eatp04R243ULzJPa
D9V3k1AYpaQXjQ9qzJ3KvRgEt2yjIH5DhFKbHMaOzev6xLBi5uGdmip/tVqea736
+4bTV3r2qJfDR15TtpkK/FjoDqrfgQOrQqICIh0pSQgcCE209iWkHMsDkLEFSX4v
+AJ1KlF1rpEqiNQB/u3uwLBYXPj2WUWVfmlx8yUPC+55lMm5RTS/JgGtYH/7FO/3
vICp43F7FCzF98TbOaslO1RNdt55AySEVy11hd7mnc2AoVAH+gi563y8I+9NTrL7
8iPvSOYD9tnjNIu8yFrKOHdLADGbrwvIKi0mxLwH+h7Gil3BxWT1GpD7AV0Fw3/v
Fm5nUJ2Dv2tSKP/MGRg3WPQ9bu/PUPvyYdUOKm8DrGNlAzhFATcKbgl6GYG6fcRD
/UvbjYNSdH1XomtRyEjk3YKnkTTJq3k+3mqzlCkGTB5xPaD86NOatMT5EW0Hc+qq
nKX0tu5IBLPzB7Eh7+cyblv3J5+2TUHZfI5yMoaOGWlC7bOKI47Q6jj9QN9G+d0j
gsaLKKn6ItxUth+Q3uQoRer7Xbk1WMJ9URjIi+zz31eIiK3n0Xb429IUFHtHgmbc
eiwB4b4tu93m1KtDw9GLY3+VugJ0lxZc7ujqTW9iQlQrWqsiGKU9oTT9bKJ8VZWR
tWfAWcq5DfnBwCB0TFSl5eJTsXM5H/5WrD2KByDgDTFk3L0LoHCctaeXSX1QXADm
ScLj7xQg4TLEwXtOnL7zgWeLLgOFRXe0s9pVLHgssEKeqWMuVltjZYLvzygiFTTU
4+ZpHyVPsp2G92NYDguas0nQW9jD+h3BnB6hvjmSKgHzQSlLRDwTjRRxiynO1DFQ
reUug8kjGIJ/hwTOqOvWRgs43yMcO9F7bFNm1+D9LDBowvO5bN2m0hpw0YW9gGVG
sKKY60vnwbiiYnTjV3ewNt7hdGPMtdS2yQqy27WQEjW7+47xx3wxYPNj4v3svRyq
VGAet9pE6CfxxxxyPW2gIhrsbZgM82QQs753KjPe1pUZF707YmFT9sq0Vpw3zM9p
YJv24tjw0dPK4QG4KvyA5L1o1F4YV0818MMvLuOgXupk8N3/Js870JsZtUkmcPn5
ddOWzfEIlaNsxAdW+Q3DxbrPEvCt5A9wWu/dcVmPhs1udWfI3pslOQM7EAPaElhr
xPKv4mj9rF7tcWK5Db56qShTJjRRK+lvU+WjmRtjRvaXgUgg4rkZ0wy74i7cKW7b
K3Oz1NnARPSAzApcOU7P7FTkEt3JoFizM5W9MO0L3GwV5V4frRjD00LI5GCTuwA5
NacbP9G2bNDebu3fbPUtJeptQUy1REIaViKp7os0E6i9ccHaAbu6aIb4OSDfuMFH
0T+NoY8eP70YSFk78G2LP+AzNkG/WXbp0yqHFldXsAeyWlQFTTN7G9sznTeL+yCK
e0sDk2lDRMHFg8p/bNAmrnJpTAdZahvG954j8s8arDn3tDtvHQXi7OJbwWrYYoNB
tAkUrGD90momaHipn6OFRf4m/IRnn5HxmAlknnRyRAS1XyEffJS6lprV7ldJ9EeH
CPM3+ACoBQJzZGSN2u3fTF4IIoRh9RS3LAC6Eu05QrL4h96gbDo9s9WNbfHOvK+w
tI3qM1HIdQTVaexiqR3R2er2lkA1wk+eSNFcFM8RnJG/MPApUGPLBUHbLyiuB60z
xvGVYrpYZeuuLrnhv4xq1t6qNOHDiRmfGQoj5283Jjx6lmkvLAl3fpMOU1FhNrBO
/5ZKjnz+H8nzd0f9Y6NtuE8QHS4vgv5FYISrOCLTSKraXXoh+toaEW4Q6X0S687S
NMlEtHSjSDlfSCQYuceA6P7yke/ehJvNLXFv0iFiqxCoCm6pzp1K+Bc+G7/RSZvc
FqbPpB0+HUPqs9BCcANvp+FukDS4rtFAeLy1b8fQ6WcsStZ/cikinP0ViY7O046s
itoxmLb5vrv0bi1bFctmTYcMpH2Bm4NrkJRQyruzykiilH0/sTLoKJVb84WXdBnv
eF/mjaJkqCwkeJe4rIOnbPmTsqydOttZJFAwo0fcFMzjHLm7V7dGYk1xJPSBUjjJ
hVGj4iW4Cylp5v21s32hd264/HFOSQlG+tKc7rClToKhsaiMylKBF0R8iqbOXwSW
DEHTHW24FOTadKZBlMc/yqNP4Qu5IHER8Zq9B1fRi7wu/LnAy4mVF2U+SAd4bOd2
hufSGeFOJWIvW3/o95KdpYZNXtKPKgRfHt9Akr6dLkeQdlJGta9k9G52gUToWyqv
j+EFeS4avl06cFQyBKXzwngqcbIN3oo7jaYrtmzC2me35BFDbSXhrZJsDXa6MByR
1/G7l0X+XVkTSJwo5Vyo0sOgzk3g4hHMt4nqLkKjbJ6kJYYuI23vkuMPZ25FumL7
CWG5qM8Tqg+AOYQhkxH1lRsRDcP9derj7cWqR+n/uO8sIEXIu7yihVu4xZw+EuB1
qUY4zWqwgjVkZrog/o69kAmv0q3PkPWHqI31uvmTjGn6N+tpmwnE+rxcEglUMLrN
IeJNvS+92Q/H1u8WwakV2oxUmWN8PVC/q+CkwrbCB+7ACcN3r2BbThfzoUG8ZTo8
Ag+YU0ctNopsGZNtg3lgSlb1NvOr6t7HNkyuHWFKS2ISKzYgrtojT1pT9peg5CWq
lEhQJNRHc1hQhpy/hu7iH+kWGGkjMJ1MOO1WmNXcssk2pBC1F3PiERT/u04fnAqL
Pc2k679OJYgbRVTNgYuspxTkTAMH38gv5G1YA1wZb4+yNUrzVnBhXoovtpaW4nC2
ce8boplU8opdPEqK1OWmM+/pMkQ7sNvvBoTaI1lSfR5y97nAAr0yiQhrLfq/i5P0
3W74Fx9S3I8smYNAWKnPZ+N0iH+TDNJYnpzrWSUqG0o9yy1xiLE98oqCcMnQUfzx
6Y68F0zmPsCwk1s97FjoM3g3s7ycs5l3+czlNHpmL6ohXTiZ0R/495SQxtcSI3GG
LUj2QylYbas78gjuWON0DQoGDZC1032YC20eESWTK/wtyvT8SSMCkpSUyXMDNu2B
jWvX75wcJ3eEc8dUvHE95yGtbPhpd+47BEW3qLVr9KOt3aEvt06kOR+fD4WCYX6q
trwEcJJMWmzoSih3K68g3GvkusjoIPQqRkfWTgWO1wi10N9gy6vqqdZUUTwOZGrP
LSdHvktrTFSBlhEdU5xaLL1zie4aJjI63FiRHTTOhGdzlhFrI5Gso1AgTAqSjcYx
7H/F/pAWJpCYXRKw5K9X1VswMK8w5MHf0e87QAPV+I21GYloo8VFtbp7zAbsmz9Z
gsFbBfie6Iv6QG3iGsuQWkMw+aoI3bl5/+CsjFMeNEhy72ZINDZcA6f/P++0+LkL
J0GSN7TwY4LqH7MhwTK5ghtI7aoBndIWDEZzfVQKI5hG4D8P1JLkAfjyyQgPavCB
yZsqiYf4n72QiRGdraDfenzX+41jIvXogtL4q42WWKILeUvi7k70wJJP+/raN/6Q
QDcYgZaPiQnMDpC3O+Ln+LJIH1fghpZIC8zkvO412bbEX2cYIe3AZtpzuuDrbZQT
X9nwZezqVBJDXLSUECMdqKUCCZ6Y4kwvuwtOcPDkuJ65IxfT0YH29lP61H3pGSqI
AYV50bfj8tN1WpUefNXKH1+fYp8LkvjWstAtVaRD2lg1r9KXuHVlT27dZunt79/Z
t7Bmf+RCnPJWU/HeeNyhRiExtgHTqKl0IWDezRxpiPBXBWo14avrCzHo578heSnb
te1MIqzczpaWL2AJQ8MPEyEj0tZ8GY/HqlCOgho1lg3MBTszw/zp/9HJHr2zteDn
xfadET1EMv0Q704XkgpGVPWTsmCW86jX4B3tKGnVwlwcDUULDN18wI4qSJiDkjiR
yrQ1Z3DZnNQZb83lVZQFutJZogHdnKey2EzVK9kcg5qJaIB4dQ35mdiCFrPdskK7
9E0HbajsTxUOeDcDXgpPI2HmemCaevOMCux6PXyolD+Eh6xBlVKnHhUYcE/7NwLc
wtCGnwkAQ9UErrOXkDprSJ2E++4f3XwvldOHjvz0uVfsNLi4NTJHx3433nMc2NS/
n4bmFX0T9xQlnbVd8X2zjTT2J0TYRhtN/dYCZ1yjrqplVqa1phzaboIo41BTGeLb
mrep/WLKCn6kR2XIQAlrdqAjazMopYRlc3PlDd3b/n0GXfzoEVTi+9ab6bI0JfPP
yDeH6zl/Tbv2/fEAadhL63c/qOcHfQTSns2h7wZrKkaK8GtVE5VyLPEwRRxHOWFS
gf0jD4vVZr98+YiQYARRgPZOEYlMPmn/bL7RWORLppOrfZ/1v7dahbua4sGAqmXJ
B0bLXb1rp2sfh3e9uJ8W4H5BppGrrXTbXlrmrHl5/aYgftwlqUJ1ocrsyRA6AdpQ
2Ii7iWFxxhbIoOw2K7/gdee68vuX6XRoOLIwW77gYmGkP6B2Q9vag376A1im6rhv
szWtdWkC07paD39ebLttPGzvf6pU4grifikWPk9SH1p3MUvIDFGHVjBVC9QnOmsR
5MBzSFkxeBZ5hs2xLKMZGWxdBhlAn0S8vcUIbVNV/gaz5S/+ZNKJDIPOslXyIVcI
kOALv0ELu/aiBcmx9qQq9I4MoRp6180pwANsaB2lvxrNoV1mU5KmlqtoynYGtYsq
ZuB4qTIZwX/ZwT6F9ci27ECtvUsyd9xs9i9zWyt6vW5/ioftDpXjdm3bCPoX7/Yj
dWjWIi3okatfECxecyJdnPlr/8+94AHVth5LMUHRhx49xb+jTxVWZs+6xnYFJbch
Y93V/piK6c1fH17Rc9fbaAnfVfz1ygaaJUxmHwfGBpG1imvJKm7CvpJ1/RBMBBE8
WxW2sxL7II1yCtKmmdGG9MfezNzhxuNfpRahDNe25SX2o7Kipu/Ikc0AUaMP+s5P
kjEFa/QNDPdGfBjETpCwiHNBGLPmTTrg+oc8nSpXX77TRJLkMtHeZNRc4+rScUye
ZMX9f2tjNI6Na7lCl9/USrK4+OTegNnKCiG1BlQpM7JpzJJ9ZrFnfm+WQtUN/RcK
LN7dVW5Cd3PsY3L+nhX+N/kxBztCGR5E5elL1gXF8QN1Kc4iH94Qdm+FJuHfm53q
XY+GOdX2VlbqUXZWvmHL/rg+xuqKtle74h7ytlnml4A4Nxhuo0nOP5SWfGVGRYTw
eGQIJXPrWSG2dty8KoXxGrFPTKvyl2sjlpvb+u/OFH4g6OvH6Z+AdSQR3Y19J3ve
x3XhFSkVQGU9j0bSna/eRHIvfkrEMH2u2kM7DP+PuGxwfFCmdjVK751zp0RmDq2t
nmZYz4Tux+JgtaCjptwuN8oH1WVXBRMsfU2R/ISITAy2DVtYXU2/KI78uUh/md8s
XUQqpNWThYS57je78inVjB2E5587nNPBEqpIPopE/FKPEzJwHM5LVzBD8wr9k5JE
Pdd09lLZcytpdx/kbtbXfXfYHGpXnmKpXaD5ozVNKlbS4Dp9B87QJZcUFbnM+7AT
Cxfi2DPa/zu66CimEfvlJyiMY1TwtJHV/CXrnwtdAIhYL2Bjwv1CilQc24c6GilH
Tpq+lgcBpWrJdBJa1m7AASTKPWahQ4kLM813vtRKHmN0Wx+UIc2zMHnUuvBbjY8r
x3TrEKQvYSOYyvpql23GGVPSK8t3vH+1Vqwxksml6zzbz3CHBtmPRfy0raHazafC
PiCudiYpuqouJmfmT2jmWuiXkrurwlVT68n+Bl1ZjJsh7d5TLknKnunHHMA233eX
gNeHdh3Uz8J5uAr/igYP76l3p2ocvQElCdJTl9C3U1Pzmc1okGQGJMVH8J5F6QJA
QJlc9Ah0cIRMdjwvoknhERPPj1znS+HS/svlvCsrZ7JG7VaYVRC5Z/MytJyMT+kw
EEf1Unv59EM5Jr7QitRfES/CeIX14RUPj3+ZY+B5YqBzUuumDysm9WujEsqw+GsK
SZT5gxvyHrRINAYcMuoF9PAkE+Ny5HT/Sh1AJuwtANVVPOO9HOh6L/m10W5Le3iX
+dHdR8crfd8Ttq9WNpqV0A34sDlZ/4G3KYVk6Up+JQ8K+ttIOGvXZKuuYeHFG5VZ
iij4e4xUD9vLIXT9mUbLhNdVipGLopZ5qOYKMFjHwWRA/hRgPumIuNCqy8X3o4Ej
8soOxsMIHPiAMSBz9GL0q7/Tct17JuodQVXME44Zs3ivXummQr/9aC7X1JEukKbc
znF72MSyhBhokXTYJKmGmMiU5cGqALjRbIPYEG4OW7sYONJSjTQ7CGq9loUboVMo
HzldShf1RPBXzl9RXbNsGFsCr6GRpz+XL2Dv9MR3oUVJICXFwo3/wQtz1iVbxru9
VqNrUkZdUuj5khtRziRenQV1jHnzm0P4lNAryfFH9WGetivt3l2VxmdZDqV+3NHV
+qZPW81++6TYmxn31c8rTXWeHiByZ/7CoUZOQNPDEYYKKn2fjN0ghN3bAOYlEr1g
PsuZAzZuMX5Lw8gbEvKpsrZHSMUHje7J7JVSsWUwKOdlcs6SnBmKEsk82enAlyQj
486vHRucqHRTkq2ghmkgDOUToI8APb0TiuRUaN3KlAvWgfoGlEvDVvSN6ddJQ4BY
2OgFKlHNtTXMuPaC0JAQWQ+pYsE1qzly5w49AhG/CTVgu1YatDU+XvIletXW7iBA
CxoUuSS8tyvxCJvtBnIEqvwKGbcNC5rL2EsMQMCEHkEETHPSDKbdg8TPseAnPMug
sv3rVjxl8zBvMnrffukLDqUqO7TkvTMkewM4ApBYyhxscok/zNQWd4ibud9ZqJkF
1Y6QCyQcXilmt53nXuqS0BoakEAaGwUdrF+crjdUgP0ZFFFVX8heOpuZC5auoU/A
wwmipAK2+XpokBv0Ro6VxlAZNle4ZIraoxk7sMHRcLT0WvqgMhcWtb4JUZSjdagp
a6doBUUJE+X1tOnYps4QK75j0mdBXBeLEu+eHBFGV9ridNRrOveBPy2XN6GxunpO
o0X2KFAd0lo1FwES959zuFjnO4Tu30k5UA2zcwIDkpM7Z3Z0lRiGdaozU4mbvsHn
eY2SjFvsn/4B2qmtgsOAtEYzSwatHWrTBKZq4kwY6c4ABLAXZST7QWfcqgALhu/Z
ndjonWyKWjn2uSKe2tpQxuDOPpr21LUXcD2Y9TvGqxJRcN4bM1nktNAyxZsM9H1H
WNkFykqKRpfsEtnqwE0Zzii/8fIYl948K1WlHH5FrBsOckE4a34hvlTSPOqjKfFT
td7jjvlMUD3oelCLqeDAglLEL1X2UVIweQe+tKN51mJF0cD+QK1xB1vksmhkoEfe
Ng1mlKk3I3AP005qF/GAAw83KYiyfJ05bVBnB7d5ndh/06zxDkaV3y0TSq6R8JHs
bFFgIV99QnDS7mTKpyhiRzDO6gAXCQhyuo9YwaT2q0oMvwR+eFa++BR0IVCqtIBj
HWbDhGyrXhvir2t4PLel2HfR/OX4TWQEHw84TT/s6AhwQjHl0dvWZCscP3Gl065W
6WjbfmTGlAkqivzslPTM8f6gRUIr8+a51boMQiD+xish9s2PSVekyz5PsAXUE+8Y
s3NcTR/8ixhzg6jp06k2eWQL9ggJtCwIXo6pfytkmYWruiV4grv6ocXj13OtV4Ti
DGokhPHg2bafqmhJvMRiIyGosdGKJIXc5WAOyp2X4Dz6MGYDXVo/I4JwN69NsQtB
NruL9uXqWV+XIShFiGom8cKLNv7iFBL1lJq1yt4j+Bbtbfp9HbLglK2dsGSYahZ4
jcZE2OfxMRz6qWYFW6sdagROnDJgNHkGOP43aqGJELbJdZLE18Wt22qiEoJBVMRX
eUCxBvZw9Or1QLWWudZhhNAdKqkFUpAcnlvopQdpkmlZV41tsxwaIOBjuxpMQIC1
SzRFr002kWjw8UZWIYA4szGSxgYUfTDE0z09Ru/ve6eLXpJUhqyjHHYbxyE/puuk
+w9jfLgsD64cYHbGHnWmi7D6pbPIuxaVvWeO1Ph+rap3LxCM3pcm/ZxXm5qyHEoN
MjEcd+4F1kGVZ4GjipuW9patMkBUQObW1FhkbbYm5GNeyD5yiHcPjOjgeUXDQK4O
jIX7z8IcEoR+6RG5wtuqQ+4YOuEKwER6L+O4PD2OCr6Th4lfqU6NwEs38e/WfcQb
BBKpgRysFGTHGqh/H6UvvP/ccY5sD9gpi/yE6ffTSqaTokQJyqBJydY8oaD12bCr
3WA927kmLPbnMlRmx+WEQwyAej2tcHGMpIcHNx2onMiA+J2C+dBUBWHqe3uLSL+D
EwvMhrOTVXCpeMNLO3n0Aa1aPDzHeWLqRRVX0RbJkoanAaQPxuha+VgJ6xJrE7Dr
TMfyGYu2jVTWQTOOCQXxSzJ3KVCPCGqONft2bD0tsSCVrvZ0jBxPfJVXl0yDXn1u
BvN+qZtccpAkjmU2yqYcViDkzmtqX0cs5fa6/Dvwjz1ULxDJjEfcUXUWKJYeECBF
WpWHBntlXxjAcQxDQFMITDJVOyTPbWUvtaRzBhPftcB7vBR6cHfCbuJq5H5ahYrj
lemlXuks3QuFw1llsmhUTh3BFNRvp5pwkDSR8PBsp2+Ye/cKYgu6N+9fWCy9Ow7x
ynUfMhd7RpSlTsUlD2U0q863+T2YouTPEdL844z1ehdBgl3v/2YK0ZajdIhrPUj3
7a6mDARSmu4ls/Cif5W6RCBZQ42HRNk92F9nyy/6QCYZDpcdPIy4lmdOtcqafNqN
N9e1Nx37Bhwvtld8Gs0+qORmzCCj5Wg0z4jXU470nZ2x0EsNasgF49JCvD4cApqB
U2FaTfFZIsqyQG5lWZ7S3DuQUyZsJ0WbktxHpitapf8cpJKxIMAwygb97RM9xovt
PZLFYtMPsfpumFv5LmAWBCj8iJOWbk+mLN1eQQNwMDUu2cTtO/ynRjTquy3UFj8c
xcO60Disglcgoh2k5PmozPEMPnEeDMzJdTkkDimtPAHEuPZyBgTijFvqQOcdNHkB
AOzocDz2YQ9VjhSWdrdAJPPMVJSE3zZrJ0KwYz4x2bF4t/VwmcGjYaDDEEyD9nC4
ZT0iPgTsNWoNbvVbPN+SFaHkC3JJnYuDmOk/wEQ3ALzOzT2tIOQfy5H7DR6QMCHA
LVcYUwt4OQ+I6yU7FQVDc+1vxQ9F36kCWT0XoJy3trp+I9rbWVJR1LGHrTSydsES
7hD7hB3r/oBAAwDRRzPZiyIvkhmki7xttXP75t3p9H9LWBdISsCFG7hQia4DNpMp
NvtCS7Fxe3/SMv5Ok7A9BRMEc4zYuBvGfLtq26jyNagkeVhTi+0eCf8ghtOOM2Ru
dXfvQTV5k9pbwr4zhydAmKplGM+2hDigL9R5Dt9t5cWfONX5qhfJ4Gb2loVnbZ+B
5cg+GEecT7kHg3+tg7sBCBg1EaF0DGRgV8F0sqArLhy5Gs0xvF1mF5FbJhAB8Op7
rjV1Vw20IN4Bt+wjiUMnQKbTXQKHtAXbXEBLszSA+os2DR0HzNGBz5j3Jw1OFfbD
GIURCRQVQGo9N6fe2Rwwx/DzbsWFG7kN39pn0oT4JgZCJ4k85+D7NfgDA7tRa4Sw
0C66evK3O/FC7VK+wAacKc1TAJkT9r4qjqjw1JA4ID2YeS3WRZGePyw6iKbFHNvh
kDbWsC7LauUIGALd+Ybojz+Q8KCPr0/m8U5rwQprmlaRiVTxlgyiwEJZ4kZnuVJK
tJ3FXx6jPqAA3y3Ev+UvIMz6eNtwM78XPgI4qqYqDlrzA33R+9iyNRiSdJQvqLwC
U1y9LqUroRlRL6Sv3Orwd3yTvJCeNjJ9jvljVuA49TAXCLrrn33CwIoyCU3/QN92
BkfetdpYgmvy9RzJbhiaPc6a7KDFVuY7fv7eMD4uXKeM3CZmbYwVecnBTGyspzfI
3Iglb3RHYMzH6gxUK6ER9KcPbIVGz+c5rjBY1dD3wIMYCBuqnzEdFQXoep/J42KF
yIal3nZ/4fJtYa0reoAoFEvvqBv7z+AiO3vbyE5ogf6EoVvSS5Rvb3Lf1yjqAKCK
f5ysR1NbrIvg8ZC/fLHEhaaApB9CmRFtbMCd+JiZRrG5Ri1iGkEQA/9yXTur5H9Q
YJeU46Qc0bl1/jS84RM2yh+u5cCpbQrBkwafdG8wVgj0nfi/kFVa53pp/rrxsgbL
C79Y8dNZmIpfhVhuh5tRet65UU21WUq5cF8ELctDzUt+ZRMDinKkYN4SqCq8JQbL
PSurH/xvzVsII4RumAlPVUTLzzkyFbMPWA7rBlcw8Nh0SlrFWnmAE1ESWi/pVhDJ
aqZ3klcy2YgCJ89zenqMu3fwktdF+Nv49S+SpL/4Auz7wqPxml6blTSqp1GGv5Zf
Hrzd2EME0MnGB3E+6PA+eWLwCX8uq95Gaa2Gi5sAucam6BNfeUWWMQ42Lr7FoaXt
tEvm3RHCSsDCiysvkYmZ2c9Ash2ZJ5FQP3BiigCSE4fJoVOYLsHzPUcsOtLAm5+h
ANI4go1PlKkQOYDiMT68FeLaxq56KupkoMlm+h17AEj7eis8g1bWQ/mFHPotgU+P
+LbgQ27b+kVrD/Tua9ufPQ9BknF5z8BgUnjBwR1Ozlp1K3uW2bDWt/6pk+FD9MEW
u+TeuEDbjHxGpFb/AvT5UMi+uEPRs/RQFnrF7ErTi6X7WNgUz7Hwof167LhztPIS
TshImghK8T6VuAA6G42PPJBIhl6EKljRa75Lu/tU9WDaTZQpJJTiV5ae/LUHgn/l
2h3wuLHxaPLTWGZDQQIPwTsZVuSr+5qes4ooArBOkTu2oI/E7xLU/4A8udy7L4us
hUaA1fEwuP3TB+imKk8Uyq1hWN/UgedYQLYeG6esoPfazNxb8l2K8tACCSnJYW16
F5a/CR9lVgsMi7fg+t27NHlT7LPItyruW4F6Yxa4sHeygY7UnZcwpXXJE9XKjszg
mco8QdYcE/kJoGYqqgAODzlZ2gBakEeK6fFkg3fBKtw0gw26Aj/RCdGHxEP3YohR
1CwRolwF/TXzc18ASrQ/rCDNbxK0Yu+zkSMc5dFcY5OHuCUJ2qcnQgicQ9juVdvO
B/7yzCu/fiedpPAKNFC9d+onaqlBiV+nLoAP/z0kLssphtr+ldDw6Se0U+Cpj3hU
C1tzB7zzDoEwcLZHF2OyH9YTWjiRsQ9cyS4auiR0i3dfAH+blbSA2amQGB3o5GRq
FXRczIiSaibLbe4s/YhS6mS8j++NXJoAdmWvCiHXZ77Le1P7cydI/LSmcdLpy29D
E9S3z7KSe3UIlz8Qv6mq76ArVnQoPvNFV1UDwqO+LmxmgcusajbelLc8YQKrcjCq
csOS+mNVJ0+xOYs2iy5ZRkSR9qlIlCkTys6Kc+i/uDJb/Epd3CcfXL1vc5tH9z9J
u7p0AHUkJQD2UFSCIgS1iOCU7dR9lItlGzAzRTJNrhNXV6xkO4qoz9xk+Ts7Q6AJ
1dl51rgyj6b+wepqn8+XzyvoWtVnRm/1LxNcme900WqCRJE4eeR36h/RHuabyAFi
npxWd3k10EpMZOZTGvktT8Wg8GrUzptczzGr5MbHM9IJkPE4HJcI63Klzwd1ATVX
Wgk3gVbpwurcdrhEpYuW8s4IpdXsiOYH+roWoMeat4KfKtVyaoO0LX9WSsBbv1R3
RmVWsHzQ+IBgDkt30//a9QwNKPbqD0vbbylutUt9YsFGFF6+OQfX7DrDVfj+gNf+
T3N4UxQPRHOdTyYrE1AaLOSuSNjJtxVlTu8m0DNE5vzQ8a+hzoSPWC8JfgJgBf8u
BfFr2fwtfKHkoVc1e/IpXT4wykAD2p9nz22Tx1MGinaui6OOqcyAAEGyg8KI+Uvy
GkEu40SW2roCDP9PxQMbhIJgiEkD8UtnhKaGGFEDJm5YUrz9xUlgoIwEK/aIU4xv
IJ38eKiKHrJcKrDsljCtRTPSSxjwBna50sPaltoDcNudXZNbfUViAzPoCZqn0O7I
IrUlyQzHVVea9Hf+GByu3oJ8WdXrm019mAANyh6QQxaP13dveui0F9OrPzVRHAzt
JJcsPLGvZGh9kdYqlMGWhGwYoKwMwRktw9zkdE2xbY82xMm0NRYUNmC8kf3Kq7T9
Afsip1zymeIHXFhYspXPKiFOQfAWPDI02TYRg4wZD4+7fn9Io50i7MZZoZKsEJhN
3bQUDSAi6j8wUVapPYdiAqSF/BdzAE5zXZqlQhij4DGI8AYJVO2to3gmZNGrLUYW
cJ55EoITaJBawnIuACY8eC5a+xtHBV95zAAljIcr8MER8Zt2uSKdNv1GDW0EXTbd
dG7MoV883zPeaeT0dZkvBUddLnunPZNOsGqhIrihTzcs14IiJS3o2wf3kaHjILSq
0KL5HiULzzI128PgUH1aK9YyVUKLL+/EtHex6Fm9qj4Zim0Eso8Y/TVXX3srUOha
s6bxzWzym/E5TS+Swz0CqoEm7jkw7phr1uOMAwUZtkkvRBGROQaEk/UzY4bMh9ay
Ef7rottv2SxPZCRnXa9C47N7X0gb0fc+nWev4kQVdm3w2KWdpQcEbV0Dm0VTzny9
ELP9zbGXm3jjUsSgD6lWrYnAMrKGfJocYQAzYWN+m798mvS1D28lqnLwCPwdofft
y2QoKGkdWC34yZsuVgWgRObIVp1fpqsMaeWjJaHxWvYfB9RLuKFp/8SoU7N0LI0G
h3hwwEmBIXyv8Sool4r4mhApAl9t+KvNVw8cjJr0A9HRx6JIXjsBVxzz5BkM5QqJ
eE/MTjyULSBmRQVpkh/sEvzCj9Odsub8PO484iKlXGriKlAW3u9AHJjlSSSoaqcK
by5Mi2t4pcjcZpJ05B6saSbsxeeV/nH55WNSxs/A9aC7+LUuwdsvrEWiYROJr3C5
pZjgktay5eqvtabTsP4frc95jtTEipUvuymkaqI4VV2GFH88Q+kWf3Vd1K5x3OyM
J1EY+CdvP853aDyA8ueOmpbq/reUY3Cr7NK/+NrLI1BKcOJW4EkXmG0PGYaO6k5U
suZz3g5428SoJn1mzs80Je9SSwhDZFlEIUVpdTyGshswgV8TItZMON0I/ujMZn4u
2AnM0viT+DxV7Tk0LwJvzx+ebvlamWssV+xibqtj8C8FXaK55dbJTp4rCoBg/gZK
e7mwgTtxTkEQmXoYwMPe2WsP1uZZZONjLrbKH0o1RNxmX7rth0xseAyBdLJrO38R
Qz9rtal/sGD+t22PZ6ouOqk69QPATDtESRsTAOB47TH+9UB3kmrOmYPVFPzQXlgX
yyFb2IITIFTAGvVPYR/PGDQyznjkOGvUq2MC1BIXAWXtsuMRi36aA3mJKCvwAgLR
ihmJC7umMJVR3tbyotEKj2/IKLEoSvkaYcHcqNQM2AfY0qLhM+LW4IDPQ8UA6oYx
iUV9Oy/LXBaaBmJUfFz63M1I/JzltmZbcBTlmyt8eOmdgrm3RAK5EiosJXfIMEQ0
4WT3hrMlUVVOLso0ykcb9MAbhX+pR8W4ytnvdT+DgjNKxXdojzFDceHQa4Rhmp2D
NgT+oU1+0f521o1GTWscC6W53ZGf68lfP84nIvj+t6+8lJJPKfupd3CfNK8BfQcL
9MPSHBeJScWQ/g1LdCbjdLp90EWD7TYQ1kSlM0qNiFvMgtx25HMNN08aJE76ps44
TdaP0wOSskXepueMPh0cHIc21oY4J/giBP8Bx2LrYQOZlTbJPLq8SpRsNz4Cxzz8
AloHO2PtGH7t8jTHgXm+ceDm/KHclAF+D02VesAWsIcGFvuVD0e34oFgJdfYdv3r
aZHqYpCTth9gv50RmBYPvzss6HpzBws4Z+zCI7VrBa2Or/YSdZ6vwMbV4uY/k0F3
KL2EorCnATu/Ao1QnLs1JJFenl6Py6vmEvrB+iyZeS0NoLwc85bEuoBSIZnL5TDI
UdM1WncDzLPUyX4W6mC/Dr51l4BbL62jVCGALI0vtrLla6A/QOnuK0vYzDbRKx0R
EJMx3e9diY6GKOTOh04KHAtgNdi3hyl9Js96aZC3pGwWuaLq5glzntiuVLhpkRAD
VsSC3GcSvyCTAXkCBX/0b2SrH2KWcJv0UtEIjJ57294dcDDbh108bbF+OI9vPyKb
sQO0FlJdxq9VVkTzVM4qqWfND47I5IL75pZNyYNPyRVUG2MCJk4zkdeRTGNXSPwz
j8te2hgr6k4sDnYggAFnqFtwNHpaTc3CmXtBaxCPw39VxjM01BRvht2v7hlPalny
Z4BglduDdt0omFu0nSORcUrQbC7pKfF80duLiGrq+ktwTTZvdLRvXMrmbSI5NdK6
7FDcvuYIaNvJs9s4nvgt29Gd3XlptI5lZ7b3ELOklReQRuQFbOasaprePy1/SFaM
9MY32rukT9/A8bxOl7CuTKUyTqkNxBpE9IVLrJW1tHz3qpJBJVxLVJVeMUU4pBAQ
D8epRaNAtsdwhRm76RClM5nj8/9PFJRxknHujDVotzdl6d9CUYDXZg+AwGxFBvIf
nl4/AIPcaDJbGz81rj7JBo4BnJPnp/2HPEDdiGjkLL9QsRJPmNi5iH/2Yih9rWV4
F4qCgiF/1Z+JT2tAva6lRjoJlgdIJ6lJEmlkS9Ou/Z+HKNJXruuHTgRJ8DhOd9FA
Adbtyjjenb78RWboB/ftOHUCJC33z4c8H/+mhKhqZjJw0TP2mZtaw+AvSo9YBZw8
Hi5t/q9y4SyXccUqg0ZUPe2BO6KEz0FO3hVLY9ZAfsaA5jBKJrX7lQ3CQdQtDC1B
d6jG46tFVaovO6+7ah0A76bRf+kM3ZOSSZFnvrYfCmS1qtnZ9Nq322japmf3WMAz
cOdCh1XekQ2tS1awtaJyHo9v6tn60pkA6AKKAJ1iKArIlL6StV2jjCurIsEGDkj1
wkZSrf0CyVY28KeBSCzHZrvSnNJcj/7zzLLKznwYQR8/tSwBt7yHv23FdjajC89g
tdVUcQdUG+XTIrd+8lToGVCYfuBrLlXTmf/9Kd7H4duyFAjjat9xPU1DQjWW4uRq
A7J7w6u/cRuOFVOLzAlJPv6fnsYncZ0XWvtYYuQ8nHVOdRdPny9xgRmz0kD9vgpp
eZCyBvtxbBSRaN3gH38bYk18nof00LovEVDE/Ne/kwlbXrvI8lo0SELhbDI90nRd
kAs4YJylSnjLUC5GU/qLT+GWvZr7gl09pMeYFa6nA0RvJe7HlBaGdoL7IxoI4J5I
2HgGqPiNUE0LoNTpt3boGhJPnfAxPrU92WSIHzPpfnLYnFgXOBVevgGyquF1ZBRA
jyo2pJk/BLTgbZfqshl+yJbP1A6/lhN5vv2zHTDYEnwUKHdQhzGkwqcI11juxrC3
aE9Shgbxo15NWFUcxC2NPoRD8LqmAy6xZKztD+jzisIjRwtnXyR4sKwJWGXDvrPj
47U1vJ/lyLdjyTxP/FNGlAH7K5ZIOfHsV3M5CXZ4LvoJZO2Iu+VP5XFRnKS+LIEy
IfwCdAHpxSdYOkHoR2eYGzd55Qi+TvjI5eh5OSW/w3t/kygx/YOERMfNkiP27guq
PPjIIKEpG4X9EvUeeNsBzEgZd/aN+dLKYEZ5xeLXlRvA0z/vGKPpDto3xK6BfXgG
K7WM7n8TO2WBp2elpUd1IRbcKsLNlYbOQl+WqmT2I2GQ7/fE9iJxHwmDnE+sPMJB
C483dfhFl5rtmeSy5lkNc2Q2kCBvdGIO57XoKuuSgjLyZAOKaQUKYxaSFQVy7hWj
prxqoQnY9IB1bXm+vOwXe1f+XNPX8qgQZSUzQkxeD+CpkdfbiG709QPGi9EIu3HN
80S7QUt666jTj8amxv9tM6eMLXPRcyXIp+tT5CBnRn9Npk6AGfbwMnuAXqakGP2u
vZas8m5rooeRu//BwNyT8CsyTUMhi4j+0hnsKOfKUqraddO5WzmAz3WehwRZ0Fm/
NA0gXIWD0s6CZm4wHOQ9hmFr67b6UUtCAmK5qp/FxMO5Q5vLWkh/IlZgx22WgYYX
yhl0YulkFT8I0oNU4Mpjc+E6DHN3U3ze5zOR7B2bwlBryL7ochi3cIJqJ5o2L3Rr
T24Ufacz6TRpwmuAzK3rPxx9IguPzD0hppkpQm+w2fZ+sCyznYqjvfwVFRbUDHlN
XrmKnWjBvYCVxHWHF5ofrpvXSi7tfB87vUfo3x0uvSlK7wPUc68xcMDafVVNU26N
SZOamKT7lbV/2Sz908X72k/hM2bpIQKU3iUb+SRApgwa6e+5jQ7n8i28+07iWrC8
EY9lrcyFvHTsSPe3hoLeP4RaSyiJs6x60oB35JNsIIvcgCGNVv2KuIXK8rKTxM3D
v/u1JSHBpivdnqhLk5v71NAA5ritCs5nvA3jZQzUi3L/sD9e6GPenY3B/WQS51w4
XEg+AAFdpOFnyJdA4Tjex3Ye9y5p3QgUaJA7g78JM4P1Cg8S1mzFglqaari3jdj9
9cvVERTlota4tYSCf+KnTA6w7Z1YgqsGRF+CHSd2pDQ9a+KO2q9NZRo9+7hjlBse
WCjFgabSwdkiA40yyL5aXTqcb7R+7cdc5Zx5WZ6Bkk8bEFvqLd6QspLmE8WSQgDS
45IFYzBWbRiqMwX99wrwm+mVMNHpJWX7eSkFvW18h6690Rf1A6YFiEjHYccBCAB2
Kkvluw91HCSmQrsDbia8qMq5vMhadBnsw+oq97w56R7DFUIDeM9S9cakTbf3Q53z
qBXHWiXAoRig0IcjlV/4ddE+p4X1i4GLcFhYWxz8r4hR/pvdE5Dnf8ioa6Ut8S7O
vo/fFQZoYmv/sEi0/8lKrz8rZ4vwQvYB0rJHnvMI8Szw5Mn2HSTloQS4m7RHUmr0
u5KuYXIQGy/LL9Jv/zTqaJ2V+duEc/vjbBvJ5KUF4Gwf5ar0X6/jZX1wr+7fjhH4
ZmXov1kdi1RQmFIN5TrbI4r8wL1KRXJU/mLS2v8XFv/HuLskTVjBTjUD9deZiBv6
TFW2nnMsLC9+dHzD7iggpDolZw3yX4msB1BnXu+Em2gFn1dkjsYjFqpEHYODoiVy
XAzDERpZdfEpO33ZN2VbUfCmuf5icN4oDj9KbBmT9cpq5AqGmVNL4DRx1Ev2jjxF
K+H3xNR1phFUFDqOx3TuYiCw0wKwmFI0CewAqbgYtBFfkmabgjFG9C9UaERKeJZI
DOHFPWhg2VpIMqGUGJwQDpv1/k17+/c/lzkjdkpNs7h6UdDMeZ+UGHOp/PwioYpG
1chZTuxBmfebW+8bD4K1ZHbFWoksS6jGO9QZCvEO7R1Za2CwISWUO5rPhEzKD6z9
F2531mR4nF8BwjcHsE8VSpmnH8E3O1fTo5ycIkukKhvpP2u2I+WGzAw3I20KUKPV
03JkFMqqZimDqDFztZWOPi9Kf53uKcwXifsyxmV47DgwX5R2jf3rgEUrMrnUl3Pk
KSgVOPx561ZTFvkkzOiS1V1sBBTYpSTM19i9hpkNNmekXQwPr9hI77+SJgo5iEJL
WPdR3Ird9yVpQEiF5YXsnTCglwPp1mNIAGymZj3w+pYKQpAEjP63FZolE5+Emks6
MPysEc1zNqaF/qQP1eaKyVV31M3J0KGyC0hW9GZeia+rj4KXzgyJYlTGW/ig+XhF
zPHWUBGH/fm2HQJVipnF/pxl81cOFYqwQkLU2YIZR5SlsWCPb/ZxJ4mfRrZx5XL/
Jx1oZvilEmtFHO5yw2cyZZHQH8Z4UzRoWYqL1r+dKyP0me1AwDCc7x1sgkKfmyg6
F68FD4+QIP6B/PTp5VXBS++oks8Tcgu+UVmvfYoTa/cRhNmrhkULCBCiNEYRj8G8
CiYTNlfa61ASVHzGPnNemmLb3M4Qvl9hC8b5en/tcLoyrjaLHk7Gl8IsXMZDKEAk
gRAEMQ9fAk4OeaugSR+Fz0g/o3rLtsjB6iZeAdTYzYmJBwN17uTsqHZbJ4s3GQZ8
9nxABwswqmZKmbNnZD6ZJrn0HGYOX4Xr/elV9+nLfuLAVlBT5Bct6zC3iSZdqrri
go7Q7h0hmUmVauIPdl1li5SF5gvNFjQIPYqeoXBpZ40FykF+HUiBEG3MtGhegVfx
MMcMn6Z2hJU6J7FFXz4lGhOphzyKU9Vw9+17J5b9mvZYXUWLzqQ5xhXKB5ZWK9Ke
HD5PSv41ax6epkmpWg+fptL5k+Jdkl7h/iiBZfgTb/99o0Ke+WeeKcHuGiHzc58P
wt3ZsoiZU6O+v/GQMVt1cMYp69W/1G6QkEEWyxSiLyifJsyIXy4YLEAwNReS8JiU
Gv10xmzpap47kicOcG8JYg4sJYvVYFXjffT/JpmROg4NU0yRWv+NFVH/Q7wKSXyj
ljgNIY3WFVZ/Tw+AKPZe4pkpIDABWkbhuOPV95U64c6d7gAFlzo696fHZ4/7wV9b
NSUW2bAlpe4ejcNSCgr4/MUKdDmyothcmLIFh1Rs+yUBmHkdeVQon5UZvzACnK0l
pcWgqLu5fWdP2p+Q8pZZnoaJQBJnTBMsCPo+UMwfuE7PX/5Gw4KtNQ/pEwxkGoG3
exiIF/xI4k4iXzWEp7WJ4euykga5dcTqpI+lXaEF9NzDKg+PNbMekrHl50y1mVkq
SEhc8wAM220vrMKkPozM7kPXvSLRvQlCspjjOcNCGtTrNQVTCEgTj6Z+7kkPcU73
N6lGHNOqm7JGCxQrOuz4DyqELsMAdyTXn7CXWHZwNCGiZU8D8UaoU9CZax2/CTbI
osa93UsGCRy77+uKT5oe6XBqFfRFFSyAlFUFX0HMZRHDA3yOTuFVfWnbiWzw5kQz
ZzlahG+XZKhm/OuChDV1dYF1AONkCHY/M3T5guMOgIPmWmk7AUU9Kdiglomw1g35
3Z50ZYh4jnTOYlJmmvPEH1H/Pee7OgNC5OF5CNThM64WJ+Khi3Sc0YZe0sI7/v7Y
dW3nxtZRVFpZ1ODko2kgIIjjDURxXdW5OdFtDTZwqGn7x8jbJg22wBrov+vEbqtY
DPcIXNMjWvCIYOjLGKz3Eubf5wRSHrUq9hTHrltEcwkorf1kotXEAbn4bOHo0U3C
YjZBmDM6nIi7E5m5Wo+83WzC/QBLTp1A9uj40MtK5+osLmN6LVGoaA8huZSjhujK
KZOgH41gerlmLbWfz5gWxbLB+MKgt29ydZeimeiOe2QyHZpNOT6z4/0VobzZTtZ3
SDjI1PwhfKuNRjhV1TN5PG96tGSJZX0EhdeigQ94N5D2bzDYeIkxfOrcZLzp8Dxt
18l9EIMXRanrPYVy7i9RLjuI1wEzNtpvc3zN5tLRM6edrdZXX/pl5E9lLoQx6j9V
4byryH83pNMDfuMlpprmBxcCfHKrAN7SEUGQcrEiFp9eZb+IRN6a89foD3pRwMhl
PsO2jjP56v+tmPMVr18X5Ym13dhAEZzoA+g416G81GRyZnd293/8XNNtGqdy0xkE
DOlaIh6LpPmOZ+YWr40nNvNNIrerwmnGTk91Dz4K8z0Yx2DoCaqwWeDLxkybv0y6
TeQw7NRQiNPBtJNt07ooV2BvPvjTz5ipacZ1qyh+jZxQXUTGkZT2i3zlQwioxvRP
tkhFKxACgoH5QLmJS5PesUhHPRTkSIyNUeSlT4Mzjt9HGilrCTWIB2cwnb1IKv4v
iccRO3Oh+mRR4QkVEJhX5G0K/GlJECbqzhbyaPSlAI01zljY00tbcblEIPXYmyrO
yrBGKKmy3zj9p4kGcPYFXno4UV811DdsFt4OVRYGF3JJjMEWTdLs1MvIiV1oBLff
BEF6hfzVtqS1GdDFE6BwykQX34dbhKOCWIjXhKQUytdE5lVi4e6u4Hmq/z766d95
DcpPtYUvQexeKGtTVYmA+YjiwvHHTb7nAqqlKpLLuavIt9NnyofrSRy+AiixcTIj
rjIbJrwBgsC2yexJJwmkgXtN4yNqVEcbbHS6Tfl6QDxVthsClNIBxSTCUkPsVPm4
Vkx0X13ODKZ6J0oRllbSjSvMhxs3gp6KbDwfh2cRNlEeNUm0bzEbf72SMnmWXTiP
ai+A/w4wp8ouZEvDOHkDuVttlar7WQNq4bIEGh3mJqMMLNGhgCDQnXIwW/smk/5Q
2G3OBOsSeBtIsRB3fhHbEZh3S5xHQ0V1dJhiBQgolhvymjbBLL+3C/mXsJdlnmYH
YtuJ0of+osTQVNRowPxoLvXZ5fiFGkHTFSvJkE0C8qWSoJMeqp+xEkM47GIWIfuz
2g7phNf9+OuhdIYekJAeOmTJ8ivq2VkZBBTZTec5S1PcTpuewqN7fO5H+6MnIV9S
3LwIJx7Fy9zeIxOvMteFzOAqQCBQE3i1vWb+ID7iyBkboOdyI2URZ6wX9oSuxQcz
Mtawohac+lQXFMFRkTqseiFFl+o8fEtad5J1/0VyHbe9aLEqxRhBmrWiHuLLmsBU
UpvWmsb+lyJIEr1QFkjyuaVXo9YKo7sbzquAoZku6SvhRhtYE93ez5jmJSI4QjOp
BzXBQH176FYPGSszTHuDuSA7T6Y4a6uxWzjv+P2023UiwC8EkZWN15pSkXoC58NX
Chv43MrZEHXWdZ3TZ+i9NTWus6MFNmYi214QQAd1KKNwXk1vFOsRimszi2CnqBIo
UnBpSasa/XvwVS1stt/aWZyvVijAW46rG3HBbrrRZiQpq8W4g5TvCfZY2IJG+McF
IdjzksRv//qVbaVUpPnj7sFnumHlh8fK7gGljEkdcpt6QMxOL9LIbKF2v6TitcI8
n+lCrvbGJ11EtQyc2/si+B7GEL2R3Xzr/ve4CoJuRmsGSXUOZIfAuFcNbLLigsPL
v+H/F7SWnEa5yGLhOK+hwa3zY7uq4oHXKh1ebIBrAIJADBLPWVazTS3sdzO+32dQ
SseDnwSwdtuClJUDbPmRGVLxVaytHWNDSUlmHUgsHe/XTd+XACdKbxrLdXZBcigR
lLZHHO6rPQXFrp4j+5knMuN77u6fohSz+kPZzz6lEx+Os/FXPLUU8GwQCgMojedk
4zUxA1q5l/VI3BOoZ3WyR01IyzYmMKSHJmwaD+BnGyToOfNbDIUB1KfRGAU1izn2
sK3ijc0U5dpJY4q8hijkhIEorVMpk4ys99uQnnlHminU/h0I6wNYlGASy9XrTRVf
RBBIiUYvTz+hX/Udgecb/dK9HH/o0lKU6d7Eh3hn+oLdWLxFOmUtKEh4GG1LuvYi
H6ue57oRYG1OkFXoWwbOwHHeiafhXDzPFY77IzglYAL24qpRJhK0rpAzySyMyL/8
8cObM4X9q/W93tFWffJ8pH1czuxqbFsVXhStO8ftlijt40CWpmX0/eAvbsGbBn9W
xXuez6xInXM2hi3My6O6fGVHy2f5AadjG2um5vXkhPIqiB8mT4UROf8OAQ1oKEbm
hhjpTL+hm+UWHHgm8M5ETfdl7VOQV6hiQR5TQ9aotabX7FBJ8JJOsgEy5XBdYsCw
EPuEmkkkg4xA1uVhidnr3AykFiGK6Cjob6anQDY/LACeQAYKiQhVI2WZ8qEO5u4z
/1wphxZBJQRwR9LIaEENuxP5EkXX75GUXD6oYGWbDOVMwOKn1yLsNMe3ja8v7FT/
c6YmTuLubamRtBtDfTDVbH4X53bOL6jBJ1DV4rRSKNODBwHkoEvoXRVQZXVLp+uA
BCoJX5U0gQLIH/wS0SkairfEB636znWj06UZv5DgRYlaWJ1PObenj9A0ETLTvxYm
GUPvKDaXmBQrAJZFaeGopmWM3oIfoKvgqaX2ZcwOVws/iUcBxSenXscm3hDoyw6H
ZHGX3NgKN6hsOE8JnLlR4yx9COEvbmsUqcWplIPOpagkdDMo/vG98Tt8UTsQF+f/
QCudVxCyKCfSn+OB7+f94Iu6pvStC2m3z0JAm/mky9DAbrmrHcKetOP1A0V7JcT+
joFMLUaw/P5S5w05ZNeNK4ntTt+2ikD95z0x/+nNRq6LqoRHXcxJnyIz29bx4nFb
w10CNAughMgFbzubqsi31CwQS1HkT/Q4kY4U/8mufYOefbeNwPIJH7NGW9oC01zo
rkdoV0+4IE589QIoII3f33VNvTjrpy53qwpzw1aYgQHHKT8Dxhb6OcCxwXJLBoKP
nfNudSCQPhQTBgXskbOdxSqZ2FHdpjOBsPr490qT4X05FlJMYcgJVyDsqiMkUELG
Vuhr3KnL6FuS/h5GsfUDZCHiLn1hHKwt0Q9p4XgB+MGzI4JPHoTa/G2m2kzqYw3H
7skiKRGFwz4slwgyZ8N0Q3Qx3ApFO4gMWlEMXx/I9Naibe18PepkRKfszyyyAeIw
QZynLBCkKAcufK26CJmqfRjKtKSpxS/2tlJHKn1wqOb13ridrdZKJ+sUAjk+lkz+
8GbjzaMQF5LUIoz6z/yzjH4YrS9/GraU62RkD8PpRBhl6uHSRlCTRc+Y7CJ+PpMP
1veb+hOxzunUVbUmo8MykmeRw2rkeFFGyGmTfDhd59nhgALwYVTw3zd5CQDnhfC6
Uap7SB40wR3JGWZxgLU/tL49fjF7aimrnYRQED+c1gVjhBhAkM4Iu/3QOF20xaAA
ewZWLiFI0hk6J1nTWXJHhrNYQuiEi1HeMkdRhho7seEIZjapLTW8EfcZPgGKYg7d
bVuJqw9ZA1UbdtJDaGV9KjjuXKIkLmyeq3+f5OmTzWNnNLk0eZNZroz7Wivday0B
qUoOuUaTi6e1MdAwDorwzbAvrAtxKliOMTH6abvSCmyxEprK/XYUZxFXSyurwYqo
m+rsskgS4YNNiLJDlc1k89aZCXoe8cJxLNMaU9UVXJnjqEUlbC3L+q8jd048KVuG
Of/2BjGNwigR1QwyHBAznz0HJswFsp6lUMkjtP2TTQ+/4NJlkVhH+UPH37FzrH52
pfnF+5ckJvnV4UtEdtu0Z+YKUl5RFgQSR1iGj0HFemKIvTiiZlqqArNqLawoVW+o
1SAivLwDnJqRRDMgsK1fpgIf+0srUtGYv+CFeh6nPgP3U7fAsuDMCrmOfiYMUXeW
4IFTeuchVyz21KmT6THVno4+YZF85gYiQ5lEzxwD6gra33GCyCJ6qte2GHDruiIJ
J7UJlBXQI2D17ACidz4ZN26KHygl7yLtJLsHji1avBP0kTaWt5vacmHzkg0AuDlo
dlLeuCgG8Q8wK+flzg9JgsyFNxHEz/qbS5DxHY6CTFgRlp8vm5qiHHR1KbgMhEH1
91US567zEMGtl7wvL/RCYi8tWdFzZRC4oLFXQoeMcoRwm7Mcbjqa39N0Wlsg6+OQ
WBwFN0aWqEaTuJp2lYjn/Hm7PaJ7AGkBXvyILRzSZJ4K+4U5gAWY+clecHS+Zk0p
fZ+oeZvxhUbeIVCD6BrYbbhWmIJqGUjErWMaqhBja4iS6BJS8f/pf+MLTGNd+aDx
6hoD63T7tatA/JfmlFJm76EKnH4c6xmlClyvJxV0JsFGeAC9lbkvI1F8VZa56IwK
1Veeg6rVb7qF03FHfqJogtdxvDTFfhYEVWj9UhL7BvgNyRNIGLz2VTYKV/X9G+J1
3fW7gKe8Y3I+D+DlfvUyfnOCTRD313QnMMuK4ajXE+CAnqeiV6m33X4gSHOuZ8p4
09xU2x2cb3RkEqva1nwAWdrvgatudcheNMjimUzptdcYpWEVmuhFeT4Hh361/Mqa
a4fTEj0D31GOV2M6thORRvV4TdIna9rF3bd1EqFPoxXj9ZQ+XN4Z1RmxtMwQ0sxT
8FdbBG8ohaxil0l+BCn53qELy9x7FkkbHU53IlplqO1KCyiQFGwh9TuySg5f0ZFn
K7tiz4Xfe3xJ16cKKgI8ouPWyjApgUmM5mgG5uMMTaYkpSNej5gTUctwgUYlbSjx
8bfewuyh/7c7vGn+PSXXzUjCARFFYZoeVZyYH10/HpobS+hmEc2ol6hbfaxZHDus
7BYekvXIPwAO3YN0/hoZ22th4yntIrqvrM9Wyna42L6a06Cp3PzZxju7w7SK567F
Olaj/Ea3dGdJV6c1iApLXKCCcHlX8j2NmZMh81CMupkso9aWf6NYYqZxI/pHrD07
F6ljz/h9JNj2sxS8bvYRehm/ye+XLzCZEYj1Z+WhiWvf8bROv8576T35X2bO7QMU
Ke9ytWAIMWuPNH89HvgVCYz9BUpCw9iCO/wexjLVXFYLqUlQbRmiaiVy5DI+gLML
b2NZpvkQ7ikZ9Cw1VOoIbE1zscypBPtjOSPaVcaVzlbFjsLF67ZRRO2s8kJZaeK3
L6OANJp9fmzZuwCpQdCtRfXCXIdAKuftEinfQ/UvoHoRy2WPL6sf16uNhZ35E2qr
+pJ7vq4aqHNSkE4U5uHt4PBOj2Gmp8C7WwT5gy6OB0UkNhRMG+/CJyiPKJ/AFSzM
3Ax5Kzm2aQPJ3SkUNDtKETeJccz4rysl+2lTtcEhHhOxAHXkjUxxkIdk0G0ka/ky
bzBaX32qHOyqcZ6+mQrbhCyOuaJS1ZjYSbl11kUwW+3rNiYWX1W5LDZnv+oIvTBa
ULvpfb4ErDi7/GE7DrOC+ako73VAp+cgJLSI7h9YqY6KNctIhTsyesDh0tUBTM8w
yM+dEqUyEWdRSrUgKV0bN3SLLkqEfXsIU7dKzn+99DjRYaZklbVeAzi8G7xIFWIl
L5wD7WffdiFUnt9e5ui//eZGycHjd+qggu3X2MAPdMYW6DODWKgVCrs5GEl9n3GA
9U6jETXVyQbBNOxBBKkL2ejrzm4VbNOZAwDO9HdlvtOZbxJCfWgSQxjELXk4WEtw
FoFTNfrriLYqqxx782koJjjdKUbtJ45FY/Iy4Ou0bIh+/7kDueMslzN3M/0QrNRr
I0GgRizM6+Otqv+ZWAd2gIRPn9b+zcT7Ig3ZZBDSGmhJjFPFd9e1AOAgq7lgSi/v
4P2VVeZJQbd8Q7iyYs47WLd8yrdEYRhnzLQ7jhCTkazrWHRdriKi+/N77pZ04w4U
OFEO+MUi9K2IEHyxwzIetUOCJ7JCbNWdmhLIm49rrQ+6CLX3BKBNRXdY7glSFUC/
+0TBmMA8BETEkt+wRSq4h/au23lJ17P2KEhwcGmSzp97YVUAsXgXqQpPSzJy2YFl
0N0rmafdICANZFA3CzspLxNZG50dPV2pb9eSk3HDidEvGnfk/NuuWbe/B6eG5iDE
iv6FrmiPkvZJrKK72hvT/2cnT/FIU+HSXnOD933NSsMISBK75S9ht/PyZ/jFGtU+
VMPOY18GgJ6Bqhf2crk5Eq+9ZLk3vQbS2q6UshXdHgLqrSxrOK7VL6fg6ZMV/RiP
smPBMe3RbUF7BaUnEV1vomO5vIGfLU4hYXAKIX7w5KH8Teoiucvs8cMbgpkVkQ9U
Q+ojed+CdDnU9UTPAJdMjHP8cB2+fKhhnUquGkCVlLSkMSRIf1VG4LIHZ3ec0CDb
12eio8mvofotwcasGQiFtUBi9pvotAhhxGxbEywvKV6aKv6e6p+YUJ4cSrZXPVaS
4mp+oea2L8MyYBTeUgTV81hJQti7uP4cdWVs5QKkN091pH4Oa5ks5tAJkvtRCG6w
u14QX9FY1eRTYTy+/XPD3WfQ5vVVXK1EmmW4MR+vvKmpk3QNigjqQku2YweNIWmv
QOi/Ymm9gnbElQurn5Yu6CtdD0wMEy4oEBbMbFBO9qxa/ho9rLzYnrRt1+/HJ9J4
cc3UDsVJECKiESoO11RDkmOmtksMLAM7w0L+lNcTREQK/ZGdVUwjNa51Lp5ZBBVC
y2wsBFTliVRZA7ND5/Mwzr5tK3QuLmssJv9pw48BaSD8qsfEPdYggoBA2Yy9c5HR
K387qZ/qEOmOPRC//eGTZWOj2Q1r+DrkHwLELurnOEm4F8VLGbBlkNZqAmvfHSw2
cJu4Ly3NtLXKumZGtJ/Seb2YuQwil8YZgQUmqH8Io1vHWMPwDjhCZwQ5XKpVWwuf
gj6cuIDX1W3oAQmFlkdze0GrTSBiuUGDiUlYguq4v5g86hjuP43QJvwoVGsEX+oQ
D7DViWQ8NPyeUjVFHaa72H1pKeJ94DwfjLunEKTiWiByB9godahcutIf6j4NMAAM
YHfe0gvEyXfK4RyeA0jfjz/ONgw+t8e8Phpa9amBaK7LYkQ2RpLilsrBRlFGLVcE
iITWNfaHZbSPEAYa6MKTV3bZlPeFWC1d5gpRliBWnYcxc9c5Igy7GThx0HjkSHnB
vgu7ULPlr08+aVutFrsxSmsPgsj+s20Xiz390YuRSHiJ3nEGFckEvjWBKhyVRMjK
sHj+2vpCZ/E8Mcodm5Ov+QKVIPf0eT9/tlCYuCkIVGVMK5u3fjC7KM7m+xa3lrez
S0qfKxvblw63FYJXLz3KAZwf2E0X+tf2m3N2RmeaBVjWw7KjlteHWGoLAVgzYSqx
n0VEY9stuVa6ta9Cm1hHZH1bWLOOrUe2NYwoswE/7LDqIj98Gk5zRi9xQPYFcAj4
d4mDHTttsqu0ZoEAIi7sDlGivJAMUwsX2b8LBgSGU/ixmIKbJTY3m23Knv9GbYOA
b+PKCynOybUA63GdHIF0v2JRarmvw8r1yIFTibgnzihfISg0fI/MOp9rQhv5JVjb
Yl58ygx0Cn6ZDuyAiVcanLouW2e/9jGy3/C9n3oPoPIIgyUuY4ZBlNtuSC5NjKMQ
X8XnLQMfM26SrtQOptnE/l8sKJLkn8JP0I5TxXdBl46Sq+kSn9AJ7xgFF93c/w5N
/Wus5kwks9ASyXJjU2gRyLjM5wduyold7t7MCHT8s7ljQf21MiRoGVhkLgAtvXg/
alWH12r4hWb0Ydmmcf+OmrBnvzc9qTARPbeOs7EXOHM5X5/fa8qAeV1HaHAaV8UO
URzbbTMqMrjRomV4PxVszOk6XXqC1GEO371LGjsES4py4TzFLPAJN1R8mFdSfkK/
icJ4WPQbS8NM72HtvR/SwHLVRA9R6mBvCVmF6L0OPXBvvFsbP1LqQ+Awoue16Af+
qxjv0/vRJCFoIIzTG8S1gqnRVs4qL2w7QENtn/7B1rg0TPYDwQwFRJ/QspQtTb6K
oSBKoykCqjlNHTjUj07GCY1KanYbEhz2ysVN2jEUw2MSGdg71xFb9TgthqNosxuo
1LNH4TJS5lDm1D6kND5lMhjyuRKhg/EJHs0Vy15LAxjEpTEivkGCofwYiqSO4yFK
6wXaXh2lHlGz9ry5WmbBTrriJOOP9E9HncD0LgxUXzwi+zfh9DOytxtUv0eCKt3B
XlR5Lr3F5RPm8/BgdNyy8L0wZLnKyFrinCj/lNWkUNbyxWEfQZcvZyRFJdXAWKMK
CjPfbK9JddpS5OPVieRbfRPhl+za5Z55VDwx03iIBCjTpZN3nDWu8BzNLw5vq7TM
6O56kVr88IfRd1ghYT1aqTaqIaVvY1nPB3/INlDRCKK3kALecoiiRCwFPJK/TK+6
waVe7HJ9LU0K74sdtVIj162dyOlOdi/b84AnSw7PS/fhKJ/1VZWJhT4fylD9F3kU
P6buoMNCqQ0eLPBcC+8BiqIPs3UMvQz/RaVBec29+zSXY9cVL8vS7mpvXc2nPVbQ
wL/v46TB8pCoWkl5naoilF9+bDBoAFJBw0LLWAXqtauNgXsvPx8vxbSi6MQxR92B
SAc65pODH+HzeLX609ZdJGrFOLLbfFl4bkswc28UXd1RGPaxRCzQOVLOtNvBd+6p
riej+X56wcyFX3Nai9uF51GZ8cPJtPk1QCFQ+2q+XnQIDcQAXuyRUrP3632LPLuR
O96mO5PvYqfz8yYfLWEhv3ozzkniKRApkN54JLSF5k7zJyi03E2vGARk7HTd/Zc7
PyTNbmtUsOyTr8AVmV3YwXLfVBKxQ9deMGu72tSUNOavtBrCb9Ur7pZK2vFTLoMg
wwHhrWOizrlUoRJDX1s2QhhwFzZj1htaD6fepDSdn7dfLEBGjidPvwcYQ0bk/YAG
LwH/4/8Ov/Y2YKxJzIIc30LXQF6SBdbLvd/pB27wsy+XNGq5Lcth00Dbr3M9+KGH
+e4JcYswRrhK6ijpfpVJdutyE0JRXxIWAn9nd4IpMIOJQg1HMBaMh7AQUePJVNAX
q+HWrVYHsXMAOVtS1n0xe14a2RbOjdBMZU34L165kIjD9WfhScHWJRVY1hj3p75X
XEYJFcuhDk0CS+xj7ZAOyQ7VaQV8nOWGZMwUgnfLPueYtkzSnY3UvjuEaYOErq0I
hmj4V0yYbm/nFy9FLijWN76KjdywC4nPLtPaKC8K6DXC2iPr3+M09a0XezKCud4P
JvWxcHEjykpM8MUXK+/ku28uM9Zu8rh4QkLqEhnfT0nJC0fT8sgN9+2MDpj9hOKi
cgw5tTfjbd7COJ8GuehRVnFA9pb5/1S4SR3U+ABaRQZhHdKsTcV0gmfB3IIlJy1p
IzK9aTRTepIv0w4M8Rcf9/UzVaIC7eeTQi6LnER1nArm/JeXlmWRYPllOz+KlTQf
HFidjqG2E/eXDLT7j0mhxQ5HfpzTHD8Zp1BWqoD77mJTrfTWAeyHsxzh3HYsPN5G
k0Q0NRCL0KPQuyDRj7//22yKfcbcWyIT7z0KTDFAZSMETvmIAHf0bTjwA22okTkW
5VneAPBSqj/nGJAVun7YpFutfDFgmujIPFtgnatOUUR/jB/lD7Fnf4ph+aJzDWL6
vsvRUq5W/IFSz430sATmildNS9grWCznH9jUZOdCSqnonUj8hTaHQsmGI8Zrq3ch
JuLkrH1OHFv5KSmZfdERZoMjolhWPgk07LGyEcIpQiCvJLXzDZWLB+ArRfsKsUQ4
rpl7vtKXM7p6xhoYIXlFv+eit0Jy2Sj/oJzRA2lLsbkxB0mCQ0mYFYYUF9HSK9xY
qXEMamX9GUnh6f4T6YeYafT1bctu9osHoxypOa+3T8eVc3zkIS5IC53B9kFJCi+k
9iBEQlxehxffEgmcPe7lKAOJeIFq+Y2/uH+lZAZHyjht2DmKf1spIkv4JbLOA0sO
FbHaYzYEp8Wg38rugjl0YbDfQbnuBPh6Kvjo6zfOr+5YzdCgBDhmWj9aGMIhWyym
fK/Ygl0qOeZNDn/tHUvg0LXTpGPqeqW6U1qRHDeHwBGpHuF9FY6jerJRcU1kljs1
DAjvu9NxmXlMCGq3oddHADhYDHWA+ungLZCaJre9gnLYkc4fGv3b7jwHG9A/onuI
ZEfxJoVswB9Wo33tSbwTMhwWZAh9tiMzrbZPExWamtjUj7mSblbf9wm0or/g9f2o
Uo5ylc4+l/y2OAb/lRIcDsyu/2nj420ZyqU4Gh8AIYpHIh4XDm0yHKXxzG+JXGL/
70QXdNK0K5q9S1NQmNhfrTn5rJOTDVz720R5OfkikgIEceXFWXPTgKWamYCZljIN
GxYiW8x011wN+wExXpPaxj2AUgUgvxQYE0gfoN6bni561UWii11ozMxOt/SxmOoW
PL0lQbhXNTTJ54hrBaa+91yVa8L5LWTBoNCIQLlMGzcGUCbsPulhJZXgaUrhsHfx
VdU14acoaIYGcYsr0roe/YMWxy0A552NIGlHsqmShuGnM7FHdbR0uQSIz86fu6iG
xk06remgH+usuHp6Kam49G1heNBfl5351qzmwTn7RoMiTiKO+U4M2Z1sJ0Savnns
pT67Ln8vW0TSrbDoZhW89DX7isSE9VPCZl+oALehhDame8ANVxDwsiy6ektRGrOT
+myfazqXkw9zNX3FrR280WYm8IfqDInAlidkeoJl4V1OTskNrlvBy6LAqdUxX1so
72F+seqCVGindLpqdpKGbB56ve5U8W1T5aayIrWuj5o3Ujhfmy0QIOWxHMx6YEdP
rmhuw3R8TiolkWBwRWfyOatD44iVxQa8uDt3vTQGcEAPQ1mvctJKw/jI9u7ue+qx
I+eWnI+LsB+TJ+X+KBQSP4JinHVONS7UKsYCm5kOxPj1+uGxOjGAJxzjEfYslUoc
B/IytGTdSH1oChRhNWZToRXiclxTZHi76Y1/FiDvTvkHB9i4HiZlx7nctGwF9PMT
YVSnye0VdS62rFuSQlhg1FPdb4L7uOGIGAkgEZLIOZ7BV0FV6dJxOPxMSWgWqDpN
fPbO8CyT9j9/emyjsjnhN1gLXIIqNAuuIhBBaaKl8RESbtCvXJR3+53MBj+omv0K
D4ImgOb3E22+hc5IhvY94sYI0PSUl4oR8zNgtT59fIDVisb2KN3SJcxlasrRVGZm
7pMGxZx4gXuyHvPCNAV07dtXpS2wPO6gOHp4qsUGmBZvt7rg5yCKo0YhBUPwhVd6
LO3TtRGsHrnCXKsm8xRdzqwI3Y6nVqh4OLyMv0GmWYIfWq4dg7T8XSLz4GWRl34S
EnAJ1+l/jQLher0W+lD35xU0FfyP7ezfLfNZdZUn1YqdwK169RPxIpfDifp3+tHF
ZJxiQV7/xlPCAyODUhKIlCEioX1iG4gBuvokiVw5CCAfQk3yenEndNxR0ta6KIYS
RQ9lXk9ahCT6oyJtJawY3NXT2FSY4IKXiF4L5QbP5kM/optUIraqMrdJQZ3WthxG
bZvhH/xm4MbVXf1f9LWmAtUCj5IfozP/5vYPZmMto1SPfOAX0mdDW/9ssfU2i2ix
JEK0XYM0hMGcE6VdgjBk2fA4Di0PviyLxEDPZiTVZORic7OlF5/T0ydZfVvaeHUj
7pzqhONfpvNg7KZ3o8Kh4CU/JC2EvsjzeOwBm7f3jy58N1wDem/11lCgVWXv60pF
8xFa3LLGZFdtdSg/1M8n9kR3iXBPvqqaHTFSNWVvfp9XF0mlsJ7Tmf2q1XXmUVli
J48iCQ5aeG3qhe23Bgm/v/2K9Ksx1PKuCpVcfFCyYi3D/q8SQ7+xnPYt7pKATKcP
UuCBHzplJXm0oFcPrs7l2XlIwRfLzE+o1vkcVKg0k1TrH64R+c6dpuKRApJX6geP
qBo+yDofcIk9+3abNuLYQBcIYvnN+JYKMzjQanh+66LX/boWyCOGsAPMUx8m9a7f
geSuHTa7XcqTn6BL1uKxCWdEfg8PXaiY3GGjgG+soRpcwA0O3bFUuB5cfDcwryCP
23nF1FZ3pOS+kiWti37cl9Z8/KsmTAAXqDVNtIWbjMqSe1MlFWN6eh3uDcOA2aXC
+s65oh40Ja7igsxGPJC7p6qMbNKWXQrQG6nv2N8PfdMyYRHQWJvVizcTrzNwsw+p
5J57Z7d7vGOfD7EGbjsDXoO58FiwNZGQ1a49acIBg2LoTdZjOqQ+3aZetk2qxH75
MYXrFtiKl9VeUoHWQEnYXfszAU2nKa+FqpExsU/fBfU03z1Wi0zgo4BWilSaIQLz
wF6k76M4UCzu9eZys/q+WWHyOfEI6/NXmuzwvJhBFxeRKRZ0HOCB/VHbcAZU83B9
zuJcSxQpvocsJSDdQ2Wx61igrbFaY1yPBra12wzfeASqu2ovmf2+aDPCSXxvf8d7
Xbm4xYfgg05TJ8J2pUKKx7Uvxw3ScJ3IKsSvqZeUOo4D2IpkKnJgdNDmLhYEdLpm
RaiN4zQFyTOAFRO60W/hua/zYH1o3YoxxHGPOk38Dvo91M0Ykl8fc5K3DVbtCFYf
WuTRh4prcn5FnnGckK8c9FRzixjOHcNyqpBY899vXAPR1eBGeMf1fXxEvZ4h6G0w
bpTVtPunbBcRwYWQm/iSb0drSlAgcAtsteWxs7/WWN+V/c1mjmzH3GVTBEN1UBto
HwcDfN60aXhrruFKigI/D+guTvKt3RMwGnwC5rGflLRPIri9OUhJzI+m4AcU2vRa
Wm09xzzrTPTv86+TetOG89aEte5oQSA+AJ1lhbtZsvuZiSGFTSX/SwX4amZ8GBCJ
9v3wHsSJXgyNNutlTVs7S7YHQFbWheiKHywk9jV9zeVlknzFiCOhkavOx1orEhEf
JucRHbTePrJGEVERLVdyrEBMpSRBzs8tDVD78z9MWpJT3975LgF92ewO8jimOcx6
R9ybSGjWv4ACa24YRMVhAESOIHiH9Lu0IXRmwK0c1hn+3yuJMqFHVQlaHsAgIF5Y
L63QrbQsE8E8/wZLXwRjK5ma7w/I1jNYHv26ozz96NI4hd3QpeNIhQ1trUfHCM4Z
YH/jcPCNm/k2XgK69sMW3gbygxu0F7iWeadtp+7D/iDTaiCteMljjAyjapwNIEPG
vcVYqJXRnjKeur05//TeU/rKoWYp9XVR6A4a540FHt49gRGqBQ6/n3vZlv5t2qPb
skzdqbVMv0+M4guAXli2Y99rFPRohbQhmqsF4jFHmpH2x3s936tKIRkpPIoGk+Ta
Ryo/OzSCyTjb4zF7S/jw8zSSyFAZQ+EneoUqybJorEYpWRxbo1plWJbrnjkHdaaN
IeYOYkAvQ2BrijDJAx7JI2GXdBXSUbGlgTo2+42Ozi0b2Iwz8A8IpsA+dIIgFh6M
QfEu+gLAmBCX5ettkrg7W3m4uH1jwLJd5UpBOlNL7pvHH+g94QoRm2UcFcE/1U7L
ux2wpu7xzqg9K5tar871023pKhKq1R7LIeo7whb7c+7jVIV25HP8oZzCwpxVumoo
9nZHbMbfIKfMAsvx/KWZ7p3j2aXmuDMeO95zFnXHXfjt7QJH2dbW6o+ekReQ9w0s
P722SwkxDs6/FOYj3WCa3AWPzIqMmypPk9pn+ueX1offmkEgTAF2vMfDBxZwLBKm
/dzqbG++N9dRRWp5cC+aGHq0e2/Aw09QpPbP3VlqQLdGVawZnzhHT+8uT1V+A7So
7oxapVGdIRfB77k72G+umqXu7UA8hQPymxEV36nRy8zumvIf8zqMDY1xPBIPnzUy
m0MribO3lzCQIZXzEoX51gegPO/5VBWgp2kg8M/rCQw+G8iFEtNKPt4sClF4k8jX
QBxVuP6RM7TDjJk5J4guXJopVwFLLAAR10Lvk7NWv/9RWMhpfbCNp/YdWce5Oq8m
++W59G2+Mn8UUtZaZdcYbOCYO/CI9w/fJuG5vfcgrPUeayKTYTU2GhnmDobJuMAp
ZpsFAJ5aQ8mMorMnTqjb5bGkNY/NSZHZXmND6xZiGR9RZlCMnXqCUnFzMHrYpcJW
mwk20+q+rvylAu2GLwV9DDJxGdJ7axCtpcsSR6upXDuBEBAw81LDfSSkgHFyux6G
CPXzrz07TZosGQBQyTO1TOuc47DwYwRabcnvFEHs5hcJB8ug/dT34rYpwz8mKJh6
Cqi8DtkPBkQhRzPu97mcuafB5sAdt1aaTd5eXSAV4+VyCO1Di4w6OZlSMKrUyOTj
8uvju2DcD46FcNqPtJApoQUqT8sc0MmAWWWGDJumd8Nnk4b3YsFjl6rPUC6jQMqZ
4lb2UuAhn5EOmdlHflUS9Q4A5imbRr2wCvrNNICrjEDn8HqRQttlbz1VPjZJJ/1e
Rlq8VGDzNTg5EviXJby1TlyXPoyImHkyK7D1rHrG2GwpH0/UK8/JN/XgBx7xa22i
QpHNziF958Sutkxw/PL+vkt0dT1gZiNmqXjDiPunSHF0rYR9Qt4mtmehjhPOYp8H
K2tLFMUjF/pw0Ij5zFpeD/rJ2hBmXmyNZmnwu/cCxmQjS25tL0sy6pRXpfUELVtH
HkjNTf/ez08c2Z2hT/7skY4eT0ctnm4EFprnZTr1c5UFg6K6h2nPx32m/OAfdh1x
jHZs5dwG9PtCGz9fRAps2p0vFG75gBvP7gHckRKeBMfMQ8NNU3PtoVHYjsTLJUt4
GS2vSGLRxKeTauznVOT62hMAYnQ0kn054tQ+dkprm1RFn4Jtc2VaI0ve4W8qR4mc
YOV/TELTrxespsTkn6SyLXVhyYctmVq36rnyCq0oLizPFiixahlyykaaeQAQ6OqV
sxVjEKptM9gTVj5uqNrUJNCAiP5FcqgUtEOSoNf4U4ZzXOagUCDWe1EKhLrodFPd
1yLcoo+d+PHhiwHk0Qup5Gh/4PoOyeO785zGKLmciDoPA1X0+KRu6zu5ETQrcNSf
hYIm6uwGaQW7EiQG0qB7iGpycc/Q2MFvZeagvxr7IYwhm9lfhnScoD3DzFX7eD6f
iRW2tqr3ROT/lI7kV/6pbOqVVov9lwU1wjLjrufp9DPmVSEh8oHY20PfpSlVvGLy
WE3WBOAmyjO0dSBD3KT/GUaAEoj9JLufdL3SiFudGaBzA4lM+4jl/lO7aP3VBVrh
bP5ybyeSmBxR2bKwyclS1n8XRAUXZ1VAlVAbziezpBlSng99vj1LyJnUXr62GQ4B
GooXFGXx0xEvvaLCA+k8YokQ7r5t7KT1zfKKT/ijcvJK0HPgyBK5rx0FVcIc/ox5
XYpdjrKne5qNlrlrzkJjRyRHgKc5JOpZxUN8C9nlKKMWPfRfuLyRibRiw/zuMl1f
ooRhwUUa97ElFcaWd03JWRTNiXfTHKCd6sA7TdoNX/F1s6z5aWEeeDDQJeIkQJb4
T+w6aUGB32MZgdVyKbQdSk/59wBQXECO13IvG8rFqIPf3SalZCCNmzUFaHq5ZFyx
SvYkY3mpKR4/k3q2g7DDFRCrm/vSiAfulZexRjfbsOiIgPPuwksKOfQkUOEz/7aL
grwqT9Jzt86KXykbwQx+qsoZRBlFaJ8TRdh3ajdBbowpzXXo4H4ySYQQ2B6E0RoM
i5GbJLVXnpNOIswW85/suaHTEig7kjJvUu+jobWChyOUW3o+NqWN/AOnM3aXD6N+
8SASQKVAaQGeE8lx1P0RrmZg2/nTRuJ+cjG6pj95ae2/hIUJoDAZ3c/mdp3zJbBt
5yFphqeME3DKKIOZPxFY4vqO+KSoanwtY2oOI/oVeMvV2rGzgWJ9QdBpuu6FnlHp
q14pP8le5KtSGkJQV0cDGb5JSn03HAMnXRDh39c1ps3LprLs2W7Pat6zdoOId5ov
zdm1KpxPQ6hWocnQs4AAr0iz4N+Bi1Lhskh3cDDEiQW2iqWbyx4mIZyYuXahw/2f
W52ai/VQQrmQ/U6t45sCt/zdHAHkpms6DVYFOquGji4NdgA/aEmOMM2ctmQW8/m/
6D1RjgnloeXa4K2cLyCVKx8RznN4cJvQwbVmwB08SbE4duCduG751Th7Euihj/1A
YPNifKmUz2t/RhJMlrq3RmnfKYtSraTvVhYMRnd4+Wo2Ty/bbWobrmeQXicIH9w3
y7ixfLZ7xKrbi3m0wK743qX1f9pbYcXq6Si7aIQdBh3Kr5SnpMSRavndjVCoxspo
1mX8BM8JH6hd07fbEYxVfRGsl4gvCNutOOfVAt+nucl91QhpbC80t1Re54yNPWCC
GZRzOEy/BpUHaW3PFA67qePHeI+0DAmeJcuk80LkxaGpGbyCNttpPuOi1GRe0NY5
3yx//lvtI6c4E3T57gZAVNqvw3o7g364SXQ6zhMP5pYzbTjjG6KcGQrLTpXrf5aE
LLG6A5Pw5ZvJJfJvQ1KC0zNnxywgAcaxiJj2YhonKBKKDRALAfRzAAxejEeNeNY5
sOP/KEJb65jbggb5X+rtntMy3MzCX+TAPHPRRLp+Zswwt6P36B1MI1zNiBlkgfE8
EYHZWiWRKL+AyHZsK7+229KN37seKp5FqeQH7mGQ189nW55WRVIniG0cdJW8XnMU
Y2ghRslTCkkdaJyw9y6EzWJ/xok8gWfmqo2TTEvsDKuSsjRQ2bG6bq7xZilIrU2G
NKaEpUXymsSiYApI6RFVld5RFSCSz2bXvk1hFcL6+gB/swDxJ/FIQ9ApethSoLTx
U9VLWOm8C9ss+qlXOsFEFdMO5o2wor6fJhEoJYXV44+uGMtb21sKDqIAVscliY8j
vCL0JX4PWic6sr9MS+bR0J9GHjKobVLP+/+m13Le25ddFVwxM0++uwVWa0mkgLii
kM0HUZWr08Wk0hdEUQOWkhBzjRchSgBb2lWS3xdW9EMUTk3SaWVyoEuCS5rg9iyB
g4HjP5UzlS23jCkXetu/sVn/QG4JFyKyswFlYTlEOZ2CwGdjc3XnFfeHK0cw/h33
+lUybo8IfgjOPHZ1ltliyDFOrk3XDqt1ET5cvkBX65p/aHZ/2dRrp8B3SJ26uuXn
tpdFv/pIVObQUetONZpy5FJCrwUyLO2BAILBS8fKekKi/tYDYdhMHP2rENY+LXk9
yfSlr2QGPSohIpizeuhU3XVF5zLZwOF8ZyGTa8JSHZH+FQG7HFDT7mPvClG7FHKZ
yVkWOjW3Igcl0snpZi/d63QLq8oJlpQf9+DUtRp+aLJw6yUW2BzLDWagEsR4jiLZ
hq6bmRj93DtS/7COH1QlxuSsS0ge6/S7TmOlBtenR01mfD+GIjWMi0rUn5UDCFfi
PfRBOdC9Mb+iPBKO0fbyXeuNWbq87H0eIK4eMB8XV5FrYmoLYmyXdCT7TzrQxNJr
NZPWMPKgafivH/TVW/LZtxikkpHyTXUl18mc+wFD9XVHF8QRGO2dSaAb4icLA6YF
hG1xOu5LkfrzOLoEkECVtzlv+scujxlmbZR/O6SWlbDBHpzbAtDZ32ebMo2+AP4I
H3qZxCo9lCCGIUPYHu3wDn/4ymg1QGdEoGv037Ty18fFl7jS/WKMHHxbogffA7YW
ohfvRInV1I0A+DC0T74u0kVBDtRizAxItIXoKV/ddo8l4kliqzJp0jPWHOQF2478
8sogfwe2LTRph9yBHhSICy5ulj2yEO2lfdSWIe0epR4t7Mfgevk/iQd2/9hBwPqR
ThxWyrddCfpVpjl8rEJ5hD16SqEBHPGx1HQs1nhSPayeSkdhKb/xdTLfSqwvWMh/
3JVTsit3q/+6RNNaUsAvfQ+rkgfbL0l5RCErkrAxW4dftAZXkM8UzDpJ5a1Hv+JU
bq4LqwyLszXEaaVfNZY7AeLie5CklVsxSrDSsVnJw41vFiMXZ3uM0dedt0AvrWRG
W0K5HJzuMQjbiDYWBARXHNBFN9AyuGTUKeLF9wONJ8+9ymmyLsPeqEdj2xK+aSi0
i+SJlxvZFg68l8ktWB3rVKLUCHIXrUvgpQZkIdJk3VXD7tQ0W18cLXvPAVzMjjNU
uQEAevzC3bX/0cMPw6D+t7cWdVaaJ794yOlKhfWzvvtfvsR7QXOeLErLelf3JSPS
o6gQU71O6/PGZbPybALwMuGVwDamFRKDfynIwP1oXn6JW7gd0GRdSKaAxAQ+8r0a
/tFjSiBSlAA0PczA+K4wNfeIbBXfEQClPb0vTgYwv/CgeDFMGUytidVTOdHFwymi
s7sKBgGmDmQpGF2gTfyzVSoHDK5MY6oHtU/axjlFsHElbdyZ6j9XDbp3/S/rf7M/
p/qvN5HwHGZ0RJEPQFWJA9/mGJc96BxQbOKfO+toXhU2SHIyohM9wO+MDeK7fvDb
YOiM/EjaQu/m+1vPMvS/w3n5RGjKXfeWHUkOA5iU4h+m2nQCRbxYvqe2MO372X6X
YwObvbWCFtDQKmHbDKVECzr4UxSCVv1J+O7H39cm1lzVZj5TlaUn9rHT1mferfni
56pYOs5V53of7EuK2Kbk5/KFsvXODorUNZ+/IFNF+xafzTVpzRLu+AZhG/XXxCWP
mBlS+H1i1CUn9JUSvRvC+2jW0ytaPnVoc5CrBzE1WUyM88b/WKWrRvnkt9Gu/ZCC
42Iuxg5ebCWfeUuhm7toDHL6a55dsU5kWvJKHR0JgnizkMliOCmwRc7/n+TZFOoW
ESkg3k5Fhe1LuYqRUh0dh+YxpxGsa6j8905MFvZRvFItD/MMJMQtW7ukFcaoueFO
uCGA/Gm6USE42DhA6QDB6HRCjEZjxc2ZartsRPiCWpENPTLXfZm5OrkYsje65GV4
h3fE6JeXC/uTDFvnjLdlFEYghSoxowIy2rY+QrQiG5yMxTsIamwxNO2I0K4X4Y6V
UMULj2Bd+cThtfzShofEyZHgZ7+NWhAIsALuEcs8LS0tK1PWzPIl0k2CfWrF9Un1
DgAW8UrVYbvdWJT6g67DiR+BbdiL+3hgJ+StSZll5VZjqeRT57k1P+cI5KMsCVxg
2TiQQwbD4XM+UksfNU0gbA7VReibLEGwp1D1ETai3XNCQY5b2JR4Ev4Apvi7qs/P
zkTBED/ky6cBeWkIm+pviy3eRoE1wDYFlXrkzcFRRj/QNT+u4/3TfpUqjs49nJev
XwVQ0OofMewhu0KG3Q0WtTE2Lph5YzXfh4+ZLpH6uQ8swIjtXdAaVYaoJmhTS6uj
XdRPzE52UiYd7LvUQEyBO0a0CQBbI/+XgxGOWxWiKLU4gj915OersdcKW9jbZyP7
GzoROi+S/6+Sj45EbVCi3B9+uBIKh5Mrr4NqkM6zHL13Xa3h8C5C1BMuT1D+vEUT
+KkWmEcaSsXY+oHTHYiBw9cItuGgo0KpeAEgFVyFDlREld8HVOvCQXkD/9EOUjxZ
XWzN0kPZLHU9AyiCd0xjdxyj/BZPpb1eC+oPXzTpAN8cKCku1dB59V7U95eRngTP
HQJPiPuKqXLs8Rq6HFZu5GBLkvipUMHMtMPVSeIkFsRe45LHCs7JyZtOAS6ir5hE
yxqxjE3aYGCST/XIlJdIdA36cZ2Yx8IZWhKjq9E+41/SzixpdzNkrLJjrHOpYgNE
D9R0j34Iodry2iBcGX03uzYxe44LMLwworCTBsJ1oIRm4y+tcrEacweoAMTBtprk
C2MAh1a8I3RfIS6edyYAEQj92x1AifLTCUPUluIqofgeV5COX1iGER2nHOIaXzNP
fBAsiNqa5IkvqU1OSUHa25XVUx0UWCOaREu8kLvL+bAb+/8Ss/JTt0k/WTaVqstU
rpBVWeCsR05y+JnX8v76f9SCwmfjJHSnHaSBfSYKl8+srmT26cvH/pa+PP9hfokj
Oy5NnQQh92h/1OuZ1AphswqhOq9+HOMdb4uO9SzITwdnpzJahsC7Hzaik9U4f6pA
Fyf9M9TIbr+J1fP35H28+XDoV4QARsyIfrEEtyx9JUvIkj7LK+7NC9d7jiaXaZvZ
yix7Au+CyEQx/elafLk1kZU/21Rg6asTrz8E8Edgmf8VskydKxa/+7TQU9/z5tLn
awRsrGUqGEr2SDceXuYxEircBbZdx8/NfpmfyKgzIRsHOj+Ug00KkyRouUxsDMQQ
EPHigbgDimfsbkOfyMP0pOFsyObyvZKLCHx61tx/qrYS75M5KGfFK8XNHaSo1Zdm
D21suYvGBYEDZcyYHpPbkCpWTDP5KYyISRkAXe/9P1d3qLUpUVVURo0uFEg5IU/S
CWnSvDDimJMneAm0F04ygmakTEvUjGxdQ21pJeCfrfTXFV6VUwqLlqf3y9oOL/Ob
40yQ16hWAn7jgF8/374iK+IpYTlOgIN7A6fYn03ftQj3VwXdcFTAtsx/9tcb7Uxb
JgadQN95hHeOS7DxsNmxV1v9LbaZvfQKYEU+EGYFQ9ejkY+CypwCeNX/qNV/WNJx
FA/p92af/MdpgehIC628jfzpBrQHlnstk2GlBA+oxcmlupMswzTAH2ItLwldkQYt
Ov7FYqQHBNr/CzYyq2L60JpMKyk2P46ObCv/tUyNbnb6IAhF4pRumME0zjMkrlag
ATcRaJRZvm31K81Qb7zIBmLFyFKFmvnm/uQkRVJpuJL3FBXynuqhRMbv62Ns4OF9
d1qKDo7mFQLHFMMr1fao7aOzQdAMZzeoIcdAGKl+uVmHfPrZhwoAjL8BZeVCRlF8
tXbqz3RMy6TCs0RPlie7rPyNW+TWyKFTno59+EhPIDqOFrWJ1vb5Yxt8idfYqids
nvcTwcvN6FdGNSUn4/aATLbwAglGPji2nu6QPk/npKratKY2Mns2Vkhg8gt/BNlV
btVKxtS0Gq6KObml0qByqakEd4M6fQVWCCZd+i1Ha+KCPLcrXbLij3ddhZBlshgP
OZIhLVKD32DBlQSd/eGHWH8HuWj1s5h7cC9vMklwumpa35K+J1jlv26BJ3cvcFDw
Bgldu1mBB52Uk2IehOkamHUL2pMZLXwp0VLRVPxWIQHzLEpvQ5KjORh5TKxNH/aT
EoHHWJgiRBoK2Fwi8EZTTZRbEB3tFKLzYmYpRRYFKiNvVCudzV9rUfpzhqbEB5EV
wgMfD2m/vSettfF6YrwUSZN+ZTNn5ywRKI+FDv0kHg5TlUC3htUxYzEfxLdcqux5
xLRF/P6ddmzwzXnuGz93tZSDdYfthKzVt7rSPtXWHQR0mc0PrBWCXEA6aMaNERbF
8z1TIGcdQI6WXossLAVbi6CQMPjK7YyAe3FEydRUkMYfDkCktRLWBY91/Xolg0Sj
J+8CY3/gcRGet8alW8vFUx+R5yA4KMLNtAFJVHburtOoQYDsuV8NJpd0gW4UpFFq
FV2tb146+zyeipJvH18tKOnMwep/8iS33cmn/UnHi4uvF5J++mrP71OThQQVTy9B
SlJt/5ps6L7EZLArmhDqVs+wGsGUhifoTNopPGJ1Yvqv3weizp/4U4v0GT4N91gE
aAMaexfskQ/K3EjNJMkhXMz7zyUJLeLLEFAtZFQbPaa90O+Sqsp24hJ6UqVDbVhN
+mEQBv26CnKlxjQyGV+b7yOgJW413E0/qicNi9XTFFHWGTdWlRJu+aeUDN23Hpj5
2Fs02jKCY8XNSs/JiFKpyvrkzbbqIpcaThGfDbUhFf5caPKkwKejnG4AHCS+/N7/
vg/HN+56F6wyutZmL77YoLvf4Crym9ua06iCc0KcHH9VzdH/GKwZo7KrrglGWZ9V
o1HvMGeuUafoMJ5qJkKQ1zCjL1CylmeZmMBaa+kx/NViOkFjG1xeJtYgg0GfCclP
Z3wCyS0iwzeM36opad606GcMKMdsr/Mcj7w/F8J4gvsFg7nXHWVOg/0zUJ+GGc0H
bLBLHosAiFXGkUOAPQeJ/D6YcTbTL+JdhJ+x9B+Ib7hG+ETzAZG95OT/fsJfe/KI
G5eK+y2hOFmtZusE2vMI5PlaFGvc9PjzKqtxDwtunA0prFeMWtDi/sr/vkzSc2yH
Ko/+O+jweuP1op0i4GSZM8TSSuXa0EY3tHY3TdITkV/4KO1nODEk91ojrlaXGub8
suYu2c3ouBhj2eVuPlufBUBzCoyCIw8Uz6Of/XQwwajo/OK++rxk+1U+Yux0JHEj
jM1UHN0COdQnbjztZeYQHa25960njzvMfmkJBAEBLUEbVvm73y96vvGK+Htzvfq+
mp6ve6Kvl+aeIQykM1Rjtx4wRvlUh7fcJViF1iziQNp24VWLnKaLOFcHORHXJLUj
jy4lpnMow//t3S8/NC6Byz6nDeNjSKAVHnCXEF7Bao5K7lH+7gBs7IU8oA/gdqIN
gB7nVQVyQBvsXzyw052KdLRWdniNEMLWmBJuoM4wdOvSxLYMWP9g9U+bMTXpUKOQ
ahwIBvVoVQ7GKbA5bdSesyMJaT8WAV/ra3PNd0W2Tt4gboxmSB+EYpou9EpTW/jR
4ulSjsaFIRcM7A924GqdXa+T+M+MZd7M6Lz+9S2vY2JBa/Ebyz+AWENzmXRCJhmR
NcQsZllmb1oTSASmZ1CDdk8bxplJQpj/SHThP/hRudT10h1c8E0Va3IW6KZ8CiKV
jqFJCvWthIgoN0Iw+QXwuh+K229N3Pc9b6lCvafCwmry+34kqCExp87aOfFksKth
jKqcinGOaUge+sFo3sVzqQO88Lyoj2MH6oy8Z7IxTqIL0hwDROjTmuuh///j6fDo
cgxYiPeIt40U9V/FdoQ5+JSY88WhiResCSnI38ahACKFp1Q7uMUZjQVq6LM65vGG
40AzrNEH193SKfqBLVSUZOjZfOvmZ7wIycCV3+0sRaLTe662/1Q70GGnDNuux12u
9yC5nBHqzTpO2jTAnYhUkuTYX2s7mmFboEzp4zLtd0qa7AtP+8X24SmjCUhXHPZ0
fScNmBFFGkkOelsymk/KeC8SzW533bERN3suogqE7N3sozlsPwdwhxMDSIh0cnjV
8zEs4ZtMR1hJfVWGrIjxqeNpX23RSV0o6gQuM1NjvqEJmqdNsD6YYtJ7aZ8iZe/9
uVnwUcKj7u4WkGISON4J+MrLAcDnrPQ9FhP2qOYbDR+pPWU4pWoVJqsHb+Yvulz9
sT24P9BuMMbLODnjX3fYZKC0huT4520Guxfe0e4KHx8RtiJPnEQWMjYpkIyu6DyM
CPCPUxhnD8tX39l+gslh/SQHnf1p6IT4RZGkb+1IYQrAQuGmtcp7x3HuMOJiZhSg
6OBsd6bhGgOFZsZZ+gD/BB6hWWwZpqo8C7KJX0PMJq4gnVkb2Q/fEpBUgoJbrvN3
xf+2xnjZVD69VanjADzbLk8tNtJwnUBGCEr8yma1ZMJgUDjCdikoktVPScCYtaQ4
Vsib7Gakm2BmhU11Hua2SKAtqm2Qme0eKndM/Cjxpq26jAVAmeCZqUI6DKvRskyh
aiNvj5J/G8208yVcFQj+AZePcvIAXdKMYHQFa/EXfkGXx1XNVjveebE+hCxnBISV
XPJ6ErAw2ZqKk7tdTQyOGThFsJqzjwWH7QjG9/87+/Ji8RUZLtCKulkAUMb57ZpI
0BTTMH5uqi9mCZ6yCAlftNXlViJuPkjjCMy6kqCfrIX3+GKLqcGQkWIzKKpUqCKC
ZFFnUm2KhAy7UwH1NeVyUvkEwa8sN7snfxiNkcdkZ6HfW/wzlSloZSzw2U1f+I8S
QdmLXHx9FgUegYQKf1flZtqr7vxlGa2k8LPhu12OU0BXkHKuIxwEdPp2E0jqPFKe
gbW+W/QRAxFYpZmXYwf7UMiNWHzD2+ctjyltH6T+xn+F/m13eRdACEMdxW83tOgx
Rik/tDp/+n5eJN5PZNVMzDjM/5m8V6iL31O/hlutF7E56vdjW0TVgYaGdH7kpMjs
qa+eb1khTu9gj0z82VwZGgccbLc4zMX2O6/DtoE6sC1naDrhGozFbkAvuQfL0qyz
Pw+PI2m6+XCru2zMO1ZNycKJxdwA2+J7Paa/ThPyUyZLpHxNDPPO1SZ8sC4NmUhY
gwWq9bvt+1WiUCZkJzJBwlV8DPoKjLXsvUBtBhiCynafmH+elllCur2xQj9Zv/OH
Wz+tC6TvAD4mVcUXuZuGnhXUu9Zy2nhfJEeLXrqIe13GjLzGNvMIqXZqa4sOjER1
dM7iwfPope9jXADmUEU//XsvntxktfpWuwmnaaPUAGK4gbwcVCyVraXUk9h+ior4
l6JMa45lF+rG9kxwX3rq7NW/wEVx2XwtPNnIkcx+7jc0AvwIroolYQnJfBAqhTRm
6yPawOeeGWyqXWXhK6LK0syN0Ees631D+1xhpXl0t3c2VL/Cbj1QSQmwKdx1SPPE
TVTH1uUtQ6e3Mvw6LhlYP5U7EHaSfR3YRhAKcMPDklMDwN/ldwieVIbhztIqQYXG
ph2g7yq1Scn2gs2Nx6gqZqwbuf+HCLV1Q+NG8iGJ6kHNkbVcnr390BC9mUvDeOa2
PbzDbu3h3hcvQH6sANtbGkaxaMqasJJh2O37cKEcdRt5A4iqwcUGk+glTwo5E4e3
NvQjmFFiQMN7erSFip9Og2keOOtQ9zNILCwSq8pOAbAob6I4cCoHQgntW8inBWNX
k6v8zDA5DkrJg/wuBcWdYwpmd9v2ix5GgYcRpjj8SMj1mCt6g4hlyiKDgkvz9M1K
n2zgdPLVQCPg38lenpwlNSVjsdG9LeL3qvbgaPWP13wfY6lq5hMgdeMwdHNiLKbs
0n4aPTJt1a8/3O0EgQ9bouIG5bBrr8pfyz0NNX7KTQdqNnU26I12NwjMDmyElmM1
maY1Uf0YXSXJQf4jCQY+Rz5Q6NF4DBh6/Pyf2/lKLUjKRbT8NO4t8eWowrUwx+x+
2M95dyUaP2MhJpwdpyYb/q7pSTDnnBescv/atpQIau++ia1hRmcSzO1zsFZZvaG/
Vx25QcxJasPe3KuIZVLDqR81uGfpM8mY0VaqImTZjRaoHoIogOF50Cp976Rq6tpS
gykJZkEJ/POgRmiw/3QQRqnlvqAtypw4KzioZGkHLFEiCeYcusNp1y6tmpSakv6P
0Hgx6OrtF4BX77IDUEA1xloVkJEyBAMyR/pX7hq/epZdYpCGrzKNslx7iIw/RnSj
8tMqdVLV3oRvbuPgJxxjYopW+Nxu3kI/zc+LHUO65i9UTqxMomLLv4C2s2ZmnURU
S0xwM1rqlMavPyZS9L1jyOWuH2hGppgkeaQAyfHL+OInsMJg6E1jXdAJWuzxaNwd
HyvDKx5WZaaKU2kX8kF/6G+WzDYqzTT7lk6pHSjokWheYHLODjqR6RRaQA1fOtsL
vtq3+yUrYn6KuXfH8YpDW9ienK9VhUQut8zMGigfLVEm89C9dC6hT8px30IzoN+T
HSnzc6J95V2xDqCSrXF6fnIrgGt2TRBEfRSf+rfGkaA/bgOWKw661qcCyTxPZ2A+
Ka0FQDlTpamuPj6xZ/Rj5UHo9EYP/6aeGCuoHXOOX2D1QiZsax+Fz8db8bAdWJ7V
sGO4BWWvIQTAgg1DNVZ3GccSEmpfivCkfUrr11mQkMbc+b53wwO9reA7pSOT1DZd
ABXJd9S7tlBGHO4YBxxDYz2237/3ywQjEXHe+mrryBgp9+BME+eiloqDzykphQoc
ZUJTq31IV2fXsdAaAhyVzF69P3ZkxVmeD7G3Op1X0r0ZuVmsfKukTg1qPULW1akM
YPMYR/UoW6CKmYek5QmpX6UaaRNy08S5fNMEX4Fx7ZOYmZXEym5haGWvuy4jRahX
rrKpEf8FmPad28mUV0OUXOK+zVITtCTurR+05DVv6329BM1k+fwRtv1waZLa5AdC
q/fxFPyaJ6tGNMWe4YYl9VnwZOtNiHwsobEyWrIJNQQcCpVZu2EuO+sBq0Mv0DAd
mhXfCKE4i6uxAHhovzpv+X2swNQmz6mXH54WcXFyDr2wTiW4lnVl5YXPgR4lA9dV
2CzITH4ttAXVq7DdMOPTmcO4AUWw432Hjqr9QnHavU3s0fTO/MO33kgtHojeCKeT
5JTXPfaGZa1bfHJTEZBgA0V2MOxqUQ61llXE+owcu8EioqsM47Y+ienxCvpTZ9PZ
1bpnyFFcd3ja0ad78dnymafE8OPSIuOFTK/1bXd5YPrLbSZFZtiPlzoDfwQGJAwf
e70ReSV9UjtHhtQyUBSsQWsG2PzkDzgI9quj2+gL9TwFomMR+UVeCNdzdLGXS4qp
P2uI8MbICH0BkB6kDbr8av6+F4kd7/xUJLa8ivxtxBXhvAiQ3FTPOKhR79FMOByk
iAGLYtO6tQ4EliTR0KIH/Lt67yN30/YCvQpQ9i+U6gRE8voqaa+UMGUv7+e5Nh2c
BvkFzSsUawCp1pPXXShFP2vXO3Q/IwPZNllAuouj4UAvKCqMh2sAH8QPAaxpTBzL
nq9b5TAI+yhSC0XcuW4jqshSkVq86esZhUgoBPIbLbHIW0sS6dDMFszywX4b1KrJ
wmg2eGRS0UZ2IohQmlmMN62SkSnHIsx9TMRED42bZfDMnVewhsq9h42QkaJ9srWA
4Aw/eexFlqXdtdYjHx99Ru5Iv6u99rX2Ygv9XXvYBTMR08BO//oyVYg4hxiCO4zt
a/zBKHHJvpMRfIpccYKq/hEQ7ytzGUCeYRp5SP3HVQekbW5/+IFWEcIyXkwa7uXr
EXBFhl8v++IMhGMPI/ZFiyIy3gP1VBowxcZ3orOuHF4I4MNDfotsrGtHtwtkUQxb
rftNPbit3ft2B8h19IWPOCQaga1dAB2KRD6HQIifC24a9kH6mmd1zp0N8RaPTokc
iu8yGUEYuwglL2J0Jo/MoRxtiVThxop1DQCFVEUl/wukA2agBHD0a3D3DrM852X2
QCv8+UNUZw6cOEJvod+ctbaXa3f+OgXkGWUqYO5Ex+YA7j06a6twnmEnktVJ453n
KY+DS84uzW4puHtIp5MPbBjiwnkO3jjnLNUgHB39UrZNkULgsV8hFT4gIChQSFfG
ZduaFJf2zCXcDbYV3B8wDOQ2vnqhXimlGEPxJgkcdCqI0kOScnER8mKq6jJgwC9D
Sc26LwlsavqkLidHmdvRJYBwKw9EXnHFPg6bZU1uuwZfzqtQUYnz9d0NPPJYQa5y
wcz1kYQZXQAYrHu6brDYwiLqNGgqoVTjH9wYp1hUpABkyFUPvyQLiuQR+2TE1EcM
W312jkNqYm2hNsNN31xyvSMHNCrfXW6LGsPq0jw0EvPPk/O9MnIZMFyEcot+Tr9w
mARKYKxcFDswseLN0ic5NyBovzYsWL7K3B6i7d89JbKpfhxbbjbOfYHY1UQMP0nB
8BUaAVcYGYtBlTZWFdX0Ltcsc6cWrbYoFpXM15aiHfB1+YkAei7GZpS/Zds/KhXo
nQVzkC/H3kJnpq6QTSxfhtQTzHzBJKqEOl/l/4fcVqMHsEKS8If0uVul1irIhBNj
DVbdHa8vYcdjAz8VyOqaHXLYlW9b5PDaO0MALsCEWlfXVz0o0fui7/rfLXJrBWk3
VlAT5iPiCxUp+CO4ul3hqBVwicuoHzKdKfUSSUz8P8mgDkSfMll1pVYReJoBjJyw
P4V/yIKz83KcvWHgsxVjt4IF/i+RAlQr7hv8OIPX0jdf0pzq7Sk4ZL8EDEl17DeC
UCULb/oqZL10NHIXZxgeiUOChMwWIxMXBBBeRS6B7bSI1l4epKtPj5kYUVh3Nswz
U0bPlnmHUOLm4JlwNHbDLW9QoLJOff4jjbLRAmsUngbs1B/T2XmxgdsXMdJyGfh2
m7A0KYw00W/3fKUerHi6ilgC8u+Nk9klPJOUveBxzUNYoXb4fxQ5Nvf7yJO6lRLz
B8CzUujNMpL2v9cJO1IEKeaK/ULx8/aAH8x/GmApXsmyMBb18USYdE6yNWtbyeyb
IepbVQmHcE5ERSOmd0KucT/donsng5DaNAo/MpexYImnhliDQPK92Fq38ODCREDd
odXDnoJG3iyzPg5cFaBgJj6SJpKWgCyP2Bj93P6Y3Ew3CeBYV2rQHSfjlpRgSerd
CjVC6DDuDoeEoG049ICxPqeku29nSYloklZAJse5cuiXQlO3WbCi/e0NT/DMWfY8
gNdBz0n1z4ADytw3jAluLmzlm5F2OC0vwj8YSPWNezfNPCVZELTky5DJoBYoOot8
0hWQ0/2QBPTwnTbKJvuisaiWpHarEStAgw9/a8/C3IBirGUchmbB7VaF/ZvVft6b
7fZXtUhYYkIU51hVOsAqM43W7rj4Bd2pHfQMY/YitfSqygXCB6bGEMnVsxm+o1/K
5p3MLaRt/7jEyB/H5sZMoP624D3fHjI14lFgiHl2UBkhy2cbYIJ1WnedzdtaWvVm
MZHKEjJjRD9bbjNvzvmMBPsJCnPZiYt5mixlHwcud2xG/5xshFmw70Y2XG+0QbQi
NeKU06K5S/Q5hRHDU4x2MdyB0iv5vaZos+xjhJHNDpo0nMBa0AKh/4me2T87NMTz
lCkoUzo2UAwiEtFHjVwXA/3w3w5vrLfNx/HTC49xvQJsprYsxBZnFRpEWN7s+K9K
0oXVHCu3zywZ0pobulfdkcBa7iaULDrh6Gbf5pUlHPx9fC3RFBlancGsb/3wrkVP
rEEkDb/zXguE28jnwF4hx6rgkZoj1zBTSGG+SaTbYEA5LGmkiXvKWkFX3IrNrGTg
TvCs2Zxzo1YvvIcLIzZbry9/p1YhQWLmUjRuWdiRBnNG826dCVGSpw3ZyzHUOAKv
Xg0QL2BeSy5P93HeV+IVJ21M2sMrfPqvHQkXeR8oV2i4YV9FzUwkIQZjkssH7vWJ
KqO/NZhRY3KB7cGgsAnbWyCSXo+m4XdOQO3uASlfVzdfCVCJoaB+QW53MHl0yebV
epncJPFZjvYk3gTJk2YN3mDLlEGNtXMEpr8fQWDtJ63CL65W00NlEKnFqLKgZRh2
JbV03Ygj3CiybUlmasYINf3AqrQM1okzJa2u6DA+FaX6cCE1/TG8PDdx3UazGZIR
kMdWXVNR1OiETzN6I7K7FWyO34ZEiMB1n/6LWa0VbzjOxcYKP4nH88797Q9jJzCw
2FbDt5jLQ+5IEQbm+LnfS4m7yJXOoIpcM2/Q4POZvY+GGSy3XwAeR4/rjZM4Ng+n
DHvuizmGWMEZZforIEOIIaVYzci7L2LiU8suCvc875jQkwjLZCzFlTwD3NC6rrxH
I7e9cIcJr/+OQVVQD4Xs5hoS9XTv6OFeKpkmqkkOlpRSMt03L+B6gCUaj0sRa5AX
90dNEYE5byPyGkSRkSSshO0ckH9IV/QRcg6JrEPeNqhIGKS306SKTp7fN0a7s7g0
Zbem4If9FMZokX4EftNCDR4tZN0MwKX+jT4+rjVYaBX28dd0G89RS7gqTeuTRsQk
56ZMIoS291Xc9yJfsO9NxuR1xidGKXCJFEB7UcWlFOpJlD5JANgNsYNejSpf9IMj
+5DG+FVgmhB503/thP0t4S83Hj0x3qNxf9jnRG3GqtN4zlzoTUkjY2HwuG7cdWlh
/RmxE0M8qP6POhgq/3FUIE7R4jZWz4PnzXHmSCQHyQGFFVIvApeEAOzWyp4kFKRT
Hhn4QsLOb4riL0Oh1u2QsOMY91odzZxQAKu2oW7hdE2JOLICFBOG5EnQzPbZ2FQ3
lyJqdgufoNsfPGZTRVpzCD8hoeK2EsPPSjY85UpJQinbXyUQNTc5L3BGFxXpa+Zw
WW7kA2ZAKAUOeW3GPdnKUZ5N6tVy53xrDlvEJhHjI7zpXIoWYIt4yNWR9q5WMMW7
UiNT9I/idvIhhMNYqoIQMKFVZUDtNdBpjhMcOFIIlvnc3lU7UCw+bEZun4IgqhWK
JkiNAUXbpWTMcRv7ElyyUOIic32TA8V8JPw5ycbnNrTAEbeDUNDEl9WnqzlLQ/sk
W7JmU27xxWQ2xvB4VviOM+6+UkR1wP8rSo4asQekUDh87cCEeNvJJX0iWm6g7n/T
QbYZpX9wqmXA9wIysVV4tm8r3hGOKVmLTsRqe9QX5aweF4UNmSpHIGPOcqA3bKEY
lO+811I43kVo75Fjwst2p1e/CBfU59LyHeTUIT0BFxHblgAvBSJN3w9Sc/iLORx/
DFxDHcClA6iHN7hW9tYGnb9ec4BFVb21YbZ6Sk6+wl1MTT8kGKWGq6Pwy5MQkag9
aucwejUqNUJ5RGZdRogyWuiUa2opblw1eAGIssA034oRnj1EikrSpE++5xkq/Wez
sY9U5g328KPMZXsd+k4wwgTEo3+1O9BPQwMaXsfL3P3mEkGMRlflL9s0zrlIg6Ey
/ScpU+lZULygNZ/WgM3Vm145ti0jpDsJucI9UZ4q1oeq2+oKE/3EiGBjsxUwU8gw
GlqCD6I4kRieM6zXWok61AaACpCs7Sbjd9BMTHs0zZQJoe+WpijC1kHYfOwIf+rJ
00qfDrAYzRXtrKzy/15PAKajNZ44aEmtRLFw5ucA2w6yzqeJzysnhndNmQB1lqpu
B52OmOjP4e+DXkP2OCmZsH3Rs6yalQG+5zFK+MF+7Tvock34Ru3Vs1/hLbl3Wh6A
9curgnhCNRKP7ZMpjESTyyydJ5zFLGGFzLgN8bVk1SQt4zfMtl2qgkm/FmvuAO2n
+o+pAUCjfykRE8jaRhmtPERrDqaDdUgjF4GKGu3dJudXxjtHvpVZGEWjd4yJHtJq
C74akWb6moj3v8u0H9zNrY1NRPo0WWgIzBmvGY3GZm988cn3H3MWGhIqoK8/NPU+
PoR8//kJwruZ3wjDUK5fAiA3Bt0QjcKxzMcyVAjHwUMbwCUdHwW0b8UwWUl/P3iz
fvqjmvAX475bIpgBRfTJpYbA3YuPloPfUDh/+BdhxTpSQVnJbQzkmcxdBiS8w5By
Nyl6CjIRTG4NYw3M9v0dddmAnzWjnueBmGmvmQ8ePcQN7e8RaBQB/oRsKDAhJCfI
/mFQvdhbeWjj87wcLZWtjzRfkKfeFYt+fSzM0JS3KBLiyXhmsyUYeCsUhrgmX0UI
LuyQ+aLRl98N7aaqmJmrCqLWq4hQbS5qJSf9N3QWI6cK1xiJQsIYHv2iALWz9zdD
p3hQBG8Rpbv9RstTXzorv33NF3YFoQ22X14pme9elyA8zcO5rXk/HIpDDLAG+NqK
2QU3dXg1ZyQpj0Fvw6J9qr6kxMQl68Jp1HBSXSJGAAk/Mkyd4WhILoOnlx7yaKUj
yulA8bnhNauwTmeN0ph3EJ5u0A5MOYXh+hQzxuy7ICEkvdnbQ6xlCI7PVgFiIDNy
E66v8341qojDkxowpYsq5wnt/RTkNYClt4OxQbvmKIdTGviaWDOPhUNAKKS6lfiB
OfnCG/YoRP8VzYUREFhK8JFVTKiz4+tt878uKuamPylGxOYGaeQOVvOvy2BmjhfU
SOIWimPevGaGuF7RGXYpzco9mhEoxVXmfAYMwK3yTySg40LZrKg4hLL4up8+wCZL
LNN/IRbn58v4tkqjLYGf9n/flkca3TUF/jpl0hzWisjtH1a47phrSZs5/pQFb+38
r/0ZcVqtsFcR0EPe6LtkiiaU26fsSpzXA3Po7X/rsdC2wAAfjKmpBu9yAFkl8cgt
8k8RkE+hv0rI4WrP4Li8ojQa7LA/MpskQZ4G/8qAEOeL/7juweEI5kg9A+ORPJh9
H79osZZynb26eF/S44p7golQAXErTt0Z2jEhsYTkbI9xFgbVZSyK1k5PWa0Ey1Qm
mRbuJ8JV5eaxW117SyUIoJTcDq2rVmGiMVJwNATZk6HSClkCpLrAu+s9YHsDQbTU
CZZmRsaTyySq1+zM1iKmjlmqmO/+78yFNVPVCZkLY5U/zGATNj8dprfh8v8PUtTv
tJqT6+FcweUkib7iPeGyLEgbC/X+IgenUeVuOJ0mZBODhwcKf0z5Q85WVIPP8s9y
T5xmR918L2JWHgsVuCQELXctWJFzpxo2T7ULEBGCNipvDaCv0sEUZm01S78SS7o+
NLil4umh5Bxdm7B/inkOfTRypb8Vaw8tD9CZpmS6YHp3Qt72Hy7EwMYIGs4NKeOD
mt2LLZ9JjwB8w1HOz7fHh7WxXjFOygV4qoUL2mrs9xCFEnC5loIAjanRr9u5p43Z
Ipo9TwtWtmIEeiIYTPAO7f8JOAF9NR7ISdIdQxDJo5hjhid2NHq1L5M1do0UQB5e
Thyw87arBZOWWXrpOrX6EE+Uc9Pw/KTvpAPxNECFNK9v6Qby3Ng6va8uLzWR1MwB
j7tSTUM6Nhkehqu/hUDWJRXSHK80wPjNfnlXYNvgr+Op5J9zOqMofmYYOJmCfsf9
75kvVCn2YxgHyYvLO3hzThPBjGwv6xzPg4IUVAVPXPZhq1Jd4YakwCW1EXs27Sr4
HCkU54O647elYIZPd54hiu3eBaZbP2vorWEYJ0CKuEnpSpndH7wZNFs2LJlxEuiJ
z3VMN6XZZ+zCdmSqrl3n6E6PTLYjYYp82IBRrzZsafdOWwVKdA2NxtbfOXdTDUSV
NoHNrelkgkQyTBSeh95iavVbzUS96iVJn6m+Z7PTAUv+wymPysnkbPoozfgjpeH+
I86EmZz2ejGRsSCwvrECJzrvnL/+op1mtv8SUUWV/Mdj9TuKKRsBL6g3itdUEu55
teAYY2lPrLDVjwHhXyMv+p7XIpJTo9jiSqMAWwbsatUeWVrfX0WHVbzCdA30DvHn
I4JzgSijKTTXfF+UwF3g7VJYJ750Hg5Wza0X4N30PKIP3pFwJW1AflLMbrE45ERK
SmFR35AUyxFF6S578TCc7H0seorgQvIulLDOKD4CL47x+gT9BHd/eP7NUA08WDnZ
1THUVAVyKXDRCQ/apKJGSwiPv4XYTZUD+cfdggKC3pwIqgSpees1IXL4X71x4z7j
YSFfCognVE0spwOpJ9an5/Kg+apoIvD0wu91VhUt+xKZ57V3qWoklnbpO20Xm0Ot
mR/pk8WO0i2ttnLGvkuIkkJm0rPeOuy/Tv8LyvYh8KvffcGKEJwRXXwnhy93rRUS
A4DIwBVTcPky46ihZURMqT35mf/Y+usmWKeLSJ3qWxAwacxiELoq0DWUDR1v3tuk
S+4PPCK1HqsQtlRImvPBSjZKVAawgZBvj16HF23fek28vRZMud9tV5wflR8x6hHn
LMoQM1Cb2Tu6bX16UT5Itl8HvGG0Xb2/KKI8QngcRn2z8Dyfgd+xb3A5T4QjkmNB
xcoViPw8hHbsNlmv1OeEZ8uJicOKtMN6jXQzhLvj0j8hs0UqJi8mu8O+wVL3gTvP
zUVyk2dQGWz8mYdLk0h+hl2DXHmLNUrMBwJTXD/chrBzKsK7EuMdOE+RBLA+D7V8
f0vn/80cRQlx/5Snh73EB3gqjRJsHEUB8vCR4atxXAqGXwbFiN1laZx2RhFsyIu0
GuGm6Ne8wg3wkiewENOhUcE7lBWbXl1D/EkeoHewzFUXrnxmEw83DgtjV9GGv23R
Rs+nAB392GCic9ND/YoOV05mLMpVdGXSS52L33v66lhBJhIH/CWjvGjZ8FQa54Kb
tpGoJRU0SB8giRIyPF5XLOVIYBVN4DODQenT2Nj7qpGbyXHBLj+6tDkALxBlS0tU
cHKdU7RLZkSw10se/d/sR8BsQzQoU6EQ3fZDwGOWk+nFKZhHyBZo3V3UAfNvB964
iIu1xZuc3Br/+cTDSZslnYjnylZSSBiUvBY/UHzbAWsSL4Jj5oxkE1NKpTtJU9oP
jiYbiWB30N+pOr4IObRS3iqZ2CoC0KAxTbosaYSWYklV3vPb8aT9HWWiQGy+xlKR
qTP80TM4CysPHI7A6KGYGgmeGaik6Ep9kD+6WfyoVFxj9v1m1MCtfQl3AfhZj+Gh
ssEtNoxRxzhJyf6XKL/Ay+p3GNWRyQ5IdZpR5skGEV0uIxtQtLhQ5Eh5yeLwGX6K
sAyA8f4LG9YtvYzB2q1p71+US6NyoawAXuEqFGPKvOIje9sOuxD+/8oA4iomkHqN
hFgssrLqvOYMYMJPRtgQAW5b9Td+IwIIdECYUK27lvVX9V26xW97u3vjoxo7v2sJ
T0rW+7UHIGGJpHrVB132moV28NgtLIQ/RNJ24AbpDIuczT35DljFEgsrYuFVW5nh
smEgUm54K19MAqdn9RZ57HMzQml9oZyGH9yvUE3TPijKp+BchKNQjJOdUSzTXat0
iG/CQbZ8EWsQk1jjrAbghMnYCpxPB2zUg/5XRg96/GH94DOQKuU79ZVz0Wi45VIG
opmFwsj6cZ7b+WYiNFP6oNKc97xOg1XQ1EiHJRFK7dqgNrYWsvLw34FdDWx7CGMf
vsb/qoUUTbbabJztHGRlQLUfoc3s3zoMjV1xTHEH5X0x2jXyooUpIChAJAS0dUgX
vairjkgXkNMNavf5zcAqvACEZ5Dr9nvCAF1m7zF+8CYG7JR0cx5RVUNPt+rh+mpL
9DJo8cuuCQ6B5xYpKQF/CCrFPz4yfU0Ge+ApnkAa5poyl6qFGOVxwlodhRkjXuG5
rLkc2fzWJKdFzOETxvrt6Z076CkaHUmySEiu7plqrFaUjHu3sAlxhBTPRoi+HkXr
gpvSIAYLOs0aZZwu78F/KfRffcedGOAA9u2B1nr4IRFbGzoquDxLpCRllYl5sqH/
UFHFHEzrIu7njadzXeinEMVWXebS76sXtSGT/eMX2LGkw/lOfgb8OAX3PkXKYRZy
f9q6q2xczobNYhv600k85LUIXOaHAWTmCd3rRtZqRBztLhgJmFdntSLUYJc3zkTU
sFghoMP69p8o07NCnb/fC4KMMMm6vJ4SMG1J5Du4esBKr4M8NQEfrFbectfUPXqn
hTfJBgLo45vIBTBGUpXeE4IatLTq0AiomgLmRfjRIJSZFZlP28zIfeW0RB+/yVPf
2b6EAO30ocmeGbfLC9T2bcjTzhHPAp2VmjFSKiE1h+ZJY5P3Sp0LJFgSAKErLmJO
H9kwag5ecHEsBw8e8LzAqyzrELhOPur+vvXVd6GBWGYwNpjPdY1kpYcKxEM0wVY5
XKYQYjcb1/UEL/FZz4GWie2L393ZfUjhSW1yDlXqA2A/WIANHj19qagLIE6p2qQl
jyIUpxnorgKoakkOA+J8dcYzHExvMwv1H12elM654Wr+Tqj2MKm07nhg1zJrmwEM
PKQNXHFXbBnUjZkTtko1+lpVf7ywp7s+6w41gDUEqh0VArsek/cl8528GZTFYqi/
7Z2BxRNAo/2j1DK4D4W5Rla71Bnevyr98e7TbxD1CDojtIUr+do+SC9j1vYjQq1M
3rTcTcFgEiRKvIH/2p35OEt/whpDx7hltaMXzCuTRrabzIPpB+pf8aqVzmUfOBCr
hFjdtaBTvV2JsgGN99O/hV8iP8ZA0gKC85ISpRnvd+F7jppIwq2X69bWIXQE8obr
lrHbcNww/6jCqQwnIDKp9tHfeDqK0/g+9LudU81/iXSVsXgoAyQa0Dx8uE3WZBp/
6JVgVu4Jc1YAkRx8nrPrq0N8tWmz4w9rHG7Yjr1ueLIJn8vPIX0RmZ5KxzlbYzKy
/iq/uXYbzA8GHs+PuR57yq1ACajO53fILIsO9TIDDKFXdDJP/XuiMvWlIW0tGuYK
lIpfPdXO4Gi6tqfgIBlkVaDzdU9j1IzK4Jy5ChujtuM+/sBApZhfiG8EmlS3N71t
nIXaWCKISyB0WiUca/wFSAqe2a/fDrCjy0IMtPUEUUZaiBfJVXq1h9UxvIngiICn
IwnAGT56VqNpc1xKe8TBKsxK/wlp1hy3gt8/vU63qJce5aOF6F/I81o8drAHrTER
OSwEtPDhzvxKEptSjzgfh125XcW4XIWXmevDqVyaodxUjA1aj4gk78k0orICzsDb
PKsmiamqjCXMMRF1mMYRk6V39zQenGO5r9btJJinNVG/75Pzw7nHsS/rNXNAQEE9
jSC73ID+ChdaP9muJ8qHMSs8qz9pFXnkBBAkGUC5juuY4HXaf3ZurwbtV7lJ0qYF
PdJ4ib9lZtKzW4PW09Ju7kX4qf3FlHckEibZGD6cuCB8jesG2aONcYNcz4StiwjW
OFQk12NZC4XCHzlbpNZnmo29TitDBTh/LTk9sU6EasLkXvmepHhVNn9Lov3+lEvr
XN5Vrnb10RWBERN7QDFFJhRYjq07xXTFxcDFfvy+il+PDymr+qWPwjYAdIuHMOtK
jDbr9sKcsPwqZFAHAp2k3kvozaloA/NGmm8ECK5UaBB2lJtlvkU4pR4eWv0e+a3C
SPF+SQJ4/oCnC6yr6X0cttrBauM2+8qoZjUtqH7bI8QPFDzon8jj2rtDUkeKhZjM
NblzFCX9ActcVqPlaBzggvAvvAysRMN7m95gpjaTE/49moGLeRUMrbSaiqGUN/hq
PARui0q3tjVPMoVaJNQZQoq4VW0f78en6qNOknpRYOG8V1+9KLkfiU0OXgfKcj0q
Op1dj4mVuFm65MmrtBkUaTFcBwOIlXe+Sr7LKRej5SQgRvGPJxvUUBGkWftThEiR
Ia452QvL/YwhXRTjp7IpZxh5oyqJ47SBeWROhj4KHc1KfSUe5FRq6s9bPfsmmBFE
26bIqHc24GDOFsMisluGHucFFb12LwhCH0+ayy0RB48LoY54Ip44pk33O1Dh8nsw
4gPajTuYyrLeFBArHIon5HpMOpXw6MOLDbktFaTYXMPgy+y/Fg884Eb8OXi/eWie
DS0ilADsPGlk4sJ4JnAWGvrdzlXoPQsx/e6/EzjPZrUmaSUajqAYnQ4xZ3JSQl7e
pGUTXQog9rS/7L/pzwcxDy2l4wQa/tasYtVhOWia9lPyT39exnZn2eV9pZkePsCG
f7G9ehlGCRQlHcQ/q9fj3k8QWCP2nUY06XYQh7VdGut7youMLergYMkaOA0WH5tK
S738siK2jnZjJuuv/N3W0np4A1J0nO/cTkq1wu0QHBQKlUi8P4o4HV6rxY9MFz0D
7TEsdeYQHSaWvxbvMn0V3D6t8i/ywhbXWfBSAqR35qQ5VTRoPy61gx6EYqKKo/G/
vIHCc2/mBMcG2PL+Uvmig2OIpYNYbqJX4HCMjUlRoLSfb96kVpOZ5S6lv+3XYnW8
MACrmB3KL8HsIKFmD0PCWLA8nJrFaRVeYR0c+ygX0dswyTjLcajmpjpEZA+cQNad
vLDoP9G5n84rPMAjienqJU8XD+r9FIYkLqtvy2SXnIXFtSJg7JxBR/tQxzezeeK0
hnF5mlewe5obF9wf0ZLUCBt+UZJ6377BzY4a35JcUeChfUf0yMVXevaznD5zwA1v
PoJ9u0wxvH5BY6AbTt6IkstZnTxyPlCzlpvrbyur3P6dkjFxmHegIpqbj0CucH++
7YnK5mz0Num4mccnQIFanh7XVIGa7GtqGGxWQMvXzh4sdLYLDWyl4tT8NhBbkM/R
a8gQnQ2jnYr+ac+/nzDy02nVBZbWyGvrVEASYqAAXu8+UfjfC7Da20v6EeFFHxlQ
N4cMtSBTf6KZ21QrmJxHaQXuR1s7nHgw/bVNCWMbLeV8Lo17ekMPzC9s6o0DAtX3
BMcX60xK4j76dqKP9LdGzStFFKpEpwvBzX33/6ALvIKtU+xfG6YAfqqwWTu2sKqE
BH41LE4M5Rx+uCJq7hMxq02fDmhenmJc2bkcO6UIjQ5+iXRVSXlqmBVUFmK4GgkK
k6iPDCLBBBpdMwreRipwUernAradHKRFX6keOnML0N5nfODb2XiDa7t7UndYB5uB
xhnqhaInueO+S9rz31GsNpkZlLTz7cgG2xojENZx7zkl0gRgLzEMWkilCLX1yY7c
Sm9HDc/eRxZSB62zIHsvgnTDZxZZvex+UG0H+Zr689avVwGJOOPLZOkhgIF02Tzk
o5+yxkc2azyvXmMzgFGZKfhnzxeTf5j9kw+9uHaBGagterTs1tRJRxGtotIhJznm
R6uTeFUjr5VpFwN/Y5b3nVL5XZqBslCFa4QQ4QJs8+mZ1T0Z58SribMsxeYCBB7C
nD8RKfAgbh1cbL1/rH2LHnEZYFx9p3W+MB42xBs5DrBB0ZYtwVqecOz0N0wIFDXs
O+LimCkCD6Cc76Py+J63uf0NrAho08nicjEkMEWrMPvVwU9fyTq8WNg7YaipOFG+
FndS4QULOghs7hD7a2E6QNkExUctfs6Tz0tCEkGIcPjnbIGyCoITmZl+AFDUqlyK
mNmvocI/0arLmmgr7+12EsGRD9hxt+wh58G5bHKAhBXM7m1JloNZ2B1fUUvFhV2U
xeiZOby41f2ogyoD9YTk76eE7FLusSrFkzvWq0EwDbJ84Mu9FYa83SlezrPmOsss
TsQwwvFwRXxY1AB7KvH9aW2jnD3D3pjjFBrrGLVrpRjg9XOx4doTTF+/pvkXhs/S
d8qhx0ql881svVzNGlI0yuWs2ldPMDKsdbaUIJ48RrWq3zcgcjUHJdtM2aNUjeEl
d6g3mfJRbH5KfcWI6fWUWjNmjy4p8/eQ+bXxeq/0WAycPCjBEpxC3LJfR93o7IAg
Y/BcQe2NEpk02a/hb8pKTPTcPl4wBfM9/rNRUwRn1jrKikUz8IamErsOAQOn96sc
l0Hti77bFdqJ9VQacSAxpLxociRZ+uQ4zXEzlB4wbfz88bPfXFlHcPVH2/Dxydus
s/i4GiV4+ZhKGWG0kKGgoxpWmlwVXUJT78B/Lxi+73OI5TMhW7Ro0l3gLwIE5K82
FOQ14qBFf/f6HPdI/4rzqDAYM3WtyKmHMtp6Gcc/X4pf0A0xjIwaMDlX7lYfDDrI
+a/i1l1kpkPye4KfgFwRdSkpBFQM1X9MhWX2SpM/uz8B2ZZUKacS8LN5iG1v+m/a
euI9ZIfpLRQuiov1nu1L405nFPDMBYdMCKL4kM94Es0N/aq9w9JVl/vAYiUaM997
E4C2ySbXhVHPXMGzhYVx0Jfut7HdnwnjvgFqT6iMyrZODJAPrKMm66F5YYyQK7HJ
nxAvkToF1glGvHm4JUwIswFoTAFMtFpbpK1XIKJMEZdSEcQMwUefTGyI0PwXQjsZ
X7ivFVTyj+T4btIpPw46SEIHsEbUCStDZ64YXoy6SX1qBkPL7UQh76MX6V3FqX7Q
U7+D6y+rn53PsE4M4909oKarWCMr7rMvq0QjIdQIpbMcQuphu9Wot8/5hKDjlaXP
J+AFJwrpsjbRLT9+OdBv2KFnhdqoE9rQEfZCm/z//cpt9SwJp0F+198GYbuIuPgu
VOasrr6uheqoT+GUAqP5izh80W5K0MVWLFztaFCNIWvcFuk5g3N2bpTUu3bd0/hs
M7H2RNnU0WdYVdQZgGwBAubqRhqXXr+RreZvtn6AIu6cz+i/+JoQAQUmI/omk7C4
4bVfAXlTv3GLMenrHMhvyV4JpTbX2nyQI5MdUwh78HggIrNqkjrXh8AVGQwOQEqe
kF3gURjWqEHc1YOcYVCQeKyl44oH6tzPO4SprzVC2BGQ4K3rXkvi3UGpmVVJuw5+
vGf5PifYgyTQ35TheJNJiu1XDfa1Y62TRskFsOlAtuMM3yoVHo5dJwQLkdwHSgXt
ZH3r9j2JpSDMmbplGjF4t1iPh23FRlVhxh9DhS2MQQMN+vydhSOrHovDvywbZECE
+smzNxClxvz+BBRZcrtL5Flwk421CKp0mUM+iNCBuaFrDt0lAWoFb6ZlWtprpzf3
TH3qy3O9MNTLm8ihTqZxMZ9ZJJUDXbfFHZ708jyO3Mn51nKebvKbtSHImLhVGqgi
voBUGA2U1GckARk4M0/0GMAk2kubRvvcbvkam80JkZZcOHjcW/1NkAWtj82f7XEy
uDGzfechEn8rHw5ukuaB4WYi/x3RgQ+WuGFGpyzwwGA7nBTBUidS4n68jwYSNWNR
4QKNSkZmrWqEN6Je/0qlkntvILPVOap6ei5TmsKXDYRPalMOl0t/TlQ5l9c96nDY
r7iXGij2f39//mZNCyavKrpjXrdVAvYtROe/f6z/T1jyWQNfdfw4dVvHwOurs1AX
vnCxHDJkVrQDd4ZNpfw/BThZShG6bLBOfzFNNzH/EfB/jKZ18ykgCg8WUvGJ7XWP
rkxwzwTTBP6X+zD7plHZ/un4IyvX/ZfMyZBiYdvm1lUM2knxUXSnnUsmPlIh+YFq
mO4/BdRcjDuXTcvFfMLW539JTGCCBHL8gXQeVxyltHKWDZPCImQem6eeSaLS/Pvf
33dzJyOefdfV/O3WvKH1b3s7HYcCldCz2SeIC5eJcKJp6Vn5X0ohh3EL5CWaRzaI
G1OoF8QSAyLvDBhTBDZHNYeth7fsSiONhzd3XtO9ZFEwCfaZ/d9mfECtoKNNinbP
Cokg/ZF0iiVvWP+zkoQZmyUiGxnQzT9+VN6GdcAw1ITvx3oUU9o2ZK2vevYCuqi6
35Y4p/mhKhs6DoXU1KHxWIUxdecgHQDEe6lJdLWdVj++tPkWxCuvUJoqnbBhcg+E
ZyKwh85Po/VPJUYfBD13Jft5sJlOY8KWBLiOrDICVMvnOTeNGtC2fq/yyNACkGOc
r2QehcuqhLVnmzhI2YPLaR/E9z5kuVvXYvqAXlRTAfZAzEiQhynZ+/MgNSKQn+qz
+PHBqiVG1F+IYIOIchVRpKCxYpR21/igOp99+YWLytTL/t3L94HtqQ9PEOXFmvV7
4Pp7BJKOvGH6RuevQvBvpRwtfG/Q/8i36V6rSx9ClYC9qHh2/eN3P8zZ+d3E5qx/
D4wy7V9GNF11VJMZrVpVkOreqSiGCJaaQjCiLV304FqwsWBOY1p0c7qMdyVVPSD6
fWadMSG+8dvdAgp2BOn+VDN6MEmL7/5la4XoDgjowudoo9gwowey1CxGnzG9DqTF
8nCsmbIoeebhYWs2gFGabKkpJpwdYmF4p8GzzejniNg/HNlUA8+6awJId4zHEV1x
U0yyM/B8Z8FFTF4ufXtdjdFqNspPxZU4F2bCS2rPUHxYah19zj1MyLOHMlEMtRiI
wDdEJQwuhWZ4HKZ7bzOl4zzsiIsXFfzEV5ZPuEhGIhS78pOlj3fUNLIkN5iE57KA
6JjVPSjSbI/cZdEM2tD0lxSurIrQkI48+cI0E0Lp0Zj4K7nE+EYQqbL8cwV9N1xC
FAOd5OzJ32b3C6sj73wW8K6piwch7scocHEWZcUEBkz0SIBG+Btxz8hgWFbmt1EH
kL8Fkkr3jeYywOPXBcgz3/amxao5r7Uph3hHTRcdZxE4TBrAvckN5TkeNJYpRpya
G+ttqcEADFEObi2Y84utGnjHv9IcFKK9pvXXgUJspFCBWZJpB0DG40D9xIVFTj0Z
dDFzBq23RlIeF7vTa/4X+RWLXFLrIHefidSxTqGmBmXjja4HM9+Sih4NaSnwLhKB
/A+acwc0861WVVifakkKjMIY9HpLbmmi+UdOXdHV/J5k4ORLMAg4ptT093xjSekI
xZvnCgsV+n4VLcLmZrY8j3SBSIc3mub8jO/suPt69Zltll6aIdMnmjjk/bwdEFC+
ehJ5o3gzq71pNHywt86J//2ON1g8AHCqK8IR86sameQOzsh/Fz4fWvwOycPUVH9K
SD2/aQh2iJjC37wm6mhP6ZUuz9KNgANxrIVkC1RqGFYHreHWP9AQm3BNK4ovnhwh
EGZFoX5wl6di33949Vzj/s4AGSvhuE4JkIUpAf1+ZWmx30a8Sag2zSptdXKVxDTC
7apzUZXJ3SbpazD96Os7ubKcLlIognWuhdvyS0mtiZVnJ9Je0XxfWXTyelwiiAjD
uHHN2+9eX22CnbFe2uQnONKgiwi/NchMZ6LivXBp3f44d6YuMfP3PK9TNN0q0Hax
vMIGdcSvitmbPU9nuXsjYlceMCyGHzMs4cKFqcmOZ3HhPzXoNffZeoLaRxpN6a2t
M5RnkJUublnRN7sCG2x+sB45vpsIQUA6Xrh+elRZYcor8iOnT1IGMu9cO5Bf+kXA
oMBAXqMn6ZHxGQ7l3hkDs3Qt4/bk0DByvDItn6eJa5kONJ6HVdAgkOnDekBmejQP
JiU2VcMpGKh3GDn41VdpQlXXLa4ShUoL+zktRt1BSv10aR4BVKja4jUslJNe+K41
veEaBXT9wVSc4k58hW5taontsvPdv8ptAwy5mouQu5yK67atPvvcuLNX5Cw5Zpxo
cby6V9uvEwhoT3/Aq5iNpmxKCsE+f7ybxbt/+nloiDJLSlZvzz9AfwW8wzuQonlj
pDlQSRUnzfcda6LYLrJFikgmPh9+y8/oTQm2B9fl0L7BjAefMcaJE7NawwQym9Xf
h3919NFVUWl7XjzU+UiFNBsL1ZPBITHoeM6fxZnBVq1wLJ1Ey4v+vibz19WobKXA
N3Py1K2MZlz2CpfBOQ7c6p1S5tIFm3+h0YjarFoegRH9jm+ZuRub3o4EkeFUBj1H
c+YkFsVkid63Fyq6/3zDzJMQTI7Jmy+eryqE2Uu3pt/PRhzOPEvwHUol3zsb+MR/
qPm2JqAZzI8KUUJyeg8AMePagGyBqHnLaejY8Cyffgl1Qgl3akkkSQPws8C/TmO0
DhSUs3lUPNJ0zTPItN8x5jaAOQ+BhKfdHYAFlayoAVrHySZ9PdqVCzHTZRtq/oAX
aAHC7HXCwzoi1kbQW7AF9GbeMmNKOSXfIYmVsFhUbzmVF/j2YHfNPS+US35299k5
3AvdLViY7HOT6o9OUMWklsAHWIze48aQgCUHOsU/Gy6MCrngssF3AfNtBWKuM/xJ
L2XhUsGvX1VzmXeNAHbbCJkw7ehkeyn6p7e3EGMU3HiGib1r2vakfAGYiRyOxf2z
/WZo3gyaU/eKP69pjB2fpAfc2RWBmxm0T9lUv0XfRhU/OxsX0A18WMl3NshGjen8
6JWPkDrE0BzwNcD7dTeLHyNE/7Y7IeugrEWsknhmPz5v/qQsN6RWzrpyJn5WbVbS
kHvcBPQtfxRCdXwYDZ0TT5RObAZdovpKJJsWp8gPzOvI9bu55MHBPNSpPsd1aBJW
Z+Cosg9mjWRvl9yY50UWrmuPf8c3RUBShKWI8+5/Sn/sdMdYRB/sAWWury0GWxhj
8NQFKdQ4eWR5lpA+qm7ImTHD2+AVANdMSSK8fHIJykichNlN3J1dY011vVHJqj9x
Y1YpDXFg1+IUj2WHLOIlQkdd0ZlqwNLaX8uzGMTxU8xgmCypin9Js8t2WZIJYt1X
9Lfcmedxyh7AyNq9xO7nmekCEoesWO0RPTqhwA0abEJwLOnyZd+ZEDZEkMHKMiwi
0PqrZ6vKnb6TP9aFtBeC9Rgv+DdfQ/XkylFGsafsa8NGN2Sy8sKrKw2H/p3Q+1jK
E3fNYQRG2V+s8UGtLJiNu6Cj7PAcGUTPBAzMpfimLyMpCilMGUA4mSFAe+xGqGVy
T+LN56SmOCaSjq6MVGYx+KYfzDt0o3a/J3SN68AcvuC59SqbiGu2rklnSbuiD5h1
AGO8WB5xSXIkFK8zVbGxtW8HSiIUiwOKBTNYy9R9gt4DnGSNsYygzaLPs8k4Q87C
h0gkBiHjAKn9L8zJ/s17zrGqGkgJ+nT7yv1LIx298OBkPiY++WZmWfojscl2zUZ2
MaZcc96M22ahj8dhgOXm9DXwjtZdFqSYPoEGsNECZfe8oEcygn3/XEAVhSnMw9SO
g5+0VjYA0PpH4EZMdL5s9KyWk92cINzrawmtq0jEMPiokeGNSkG9eC+1xlKX7twU
9PH0uduRlpAywq1WhHcrlAX927mhzkeCLQTIZD3lMP77TTWbZPs64qBQWH4ILp8S
3M+d9kQx0KB94MtJCP+yEQJ+SKwfB/qscQjT5JeV7MvujygZpYkftPSdJwwCia+D
HbNHSd0VnCsTyYGJ71/xE++JPN7Aa7kIoaXi7tCUmZW7M/OVyZGpZ8D7RAQrFSBX
Lpl9/ac0U80jZpPotwJ2AvNT0w9YOg4ZpfeONcjs5C/3E+I5qRuaHq2igdVq2ctu
z0Ub/Q1Ujmb6GiIGsFYmO8oc38lNin3VR4AI7u2kN9XbdKV0ht1iHgf2C6FzGlF7
PwuBEn8UJlSgeez4u6S+1LhiFdannDATsPJr7NbP/w2PzCQe5cv/q7KDOwgtHo3W
gXYi7i9QmVdBPJgnEcH5N9JV70DTvRsQi/iGi5ozG1BGV8L0uPA7F6ahFWkqj5VC
DRUMQvUjrEPvqCztO4bfHAt4jRX9eSnCaW/H5YkSFyHrQlXmEMQTAny6loUhD4RH
xVRTycJIhWmcHm9gXqKMKAlI2VPB7YUh281GmTn7VnCBFY+7IyvpEIepX6Fun8TE
VwU7W0UQORAm5PKThrTODemlK5zalWWMDOtEiUbUwGDWknPGRoRTYRPDWbnhD/N9
vTe87j+cbId45MaeIQAKy6XnpSv6xIG4C72dV7gQYA8jnpJInN0H5r1FdRrgV3w8
OrnwYgOzb1t4qLcwEmpLcDMpoz8EHD52geitTAGXbTXLjWgtjQy21bOY8pHlcbj/
sXYt8voUtYidkHduY1i7V8c6dtg9DmRVF5FVgbM4EGcr72d4keffumgOzAhORweT
A89vZHPeG5bkhwJ7GpxGKBfkVFJgUoc6WggmbBNfttavstdrI0oRQvJGRT6LTcaz
VitM3BzZx05pninEjeYxHc1FibnGKI0ZO1YuiqEpmUSC+44K3/qWSpvaprUGje2L
Qvkepu5KH2lBIAu4qxLGdfLCXN5lyGEAsBmomWeTOfM11p8x3iyDry230yv83yI9
OnaGiemalUrf7nR2N+PH8f0lKb+XeiUcCFRFFopVN2oCQjWQUsr/nWIE+yWilMrI
FIsmui0tU+7FitEOWAAMJkNfQHULN/Py9+aNOJgujHpi/HMhR/pX8bFPD6mO81b3
DIc8BuVjk/h6sPDfiHhFPSaCsVwDwO7Q6WXWDpdwNmy0Le2FKqGrIJpOtky7F0Z/
N7infXpEFz6us4E+b++loiTt777BwCVx/N43jp6WsypXd26aw+9F0fvI2EtSqLQp
Y18emWkEou3m3KrNsN2+V5raTyDEvJzVLDs1f46H5da/5ZPNjEqLX0iac+Oc7gMc
HJNt20ilr2QSXkdeL58elFORpdWqhED5iRFYPzl3ULkADYn3CTqFrNiv38vqa+7A
1ecDCIi82flpULXbzI65Q8M2sT1srlXfWVWL8lFe3KTzAzQKfrdIjs+lpxyE5Vq7
jTlm+vH1me0p6nUJ19f3+V654pPvD/Yw4TRF2FYeOlxNIlhxnVOjxP9XTPp0l4ua
/VPDtHElwiUebIicqYrOuSpyWUQ60h5GOURZ6XdTM9UndL0FvkwzHwyHrBqvjmyd
QRrl04bZYFzY2gy+UeKRMaN0EY18T5ErE6I85Xl4tQe4srwNfCAGMb/LEUUhV+cU
O3keRPXIXBJ7nXJW1wGu2J8L4StNUb0W5dJ9lnxIXcOQHeu/0/2fCj/qmv87Ixj8
z+Q2TSbV8kr1lYHyA4XYsP/RaUffiqaydIC0qDmtykneuoe622QohuoikIQUhpEU
aHjsgnxKI6kXQIBPOSnHRuwdVvwU+9G/RWKoPJqtnOgel05+xRWAtVj12+1nJnjU
ACvN/gY/s9vIQwOZ1R0fSJrsr69iZU3H+NzMaV1374Ca2h4JMI++Op/aj4pWZAsl
WBdctuHPb91s2zULJ20u87DUFAFs/KHu674rF325UYrgFptClYbQ++gX/srypsP6
3bJh1WnksBQ6WikV22WPy4uSMUoEERqJUmQ9YWTvxC1dw26TDBD6BG2VfG6/INJ6
dOzHTyPIEWaa+fCKcsKmy/+jGmi5iHDppbxcJC6NDLmCBdET1UlxDaH6hZIxyprn
KN9vZ7JJ1Irt5TMOjIPSlkTopoubMcooxCL6WeZcYQ/JAxO8Wh21GDXgjpfIyfn9
csqfzwgJhs5L+5xyctpw1ep1Y3kneWMWke1Hoi+iyncLRgYDpDbgTlgwGKEPiehl
r+X+/BUTMcg5UxFOJNQ/kiKEJNS6W9DZpd+pQEIBY5Pm3YLssrPxTDfKTTw1VKqm
G4HoF02jOP+ERU5AALQWy3upILsGNYYsdhN2Px69DuCFgNJnqST4F/xrZnWdquIR
RHZLWnl0fMCR6vWdAMs8xlTKGWbXtJ0Sng7P3HYDhkFXSyue7sEAmlUAHPB9TlWE
uXUoxeRP3uwE+n7sNLsCyrwhn+GiBSfIM6X7aWu+H5nzopnbdiyXoC/kaPIwVRhs
3bEHjQ2hKXk/QJcPOUyHY0bGi3LtwFL/+EEjHe+6QNW1/gfxpQwx6IgfMufWlLdv
Dhpd5C7+29S5txiMdnQML8RZCSol8OYzjz9pCfUa8mLN8JHea8OwAig7YT7Ivhqz
SQ3Z/lqZSo7avTNMRt6cGL65Rt+GXdzqhE3rA+G7OUSpFk0D4bz3pVutLmq71Aip
gbBd8pfrT2Af9e4G3sca+3r0960vcVATqdC/O8HiuQ0QV6VE/4Fo59zo9Ef6hh9w
8VzKmZSOJBf6RTFOXzyR7xCgqq/DTyZMEfZO2hDjZQaW2+rW9e3bLtFUrvlauxls
22jTWtsBnAwiPnqHAJinL/iUjI941wxlRfyi+1RSYD0MwAT+3uwIdBj6dZFpOGsL
+csfCXGvOmM9UpQk8o5CdvAF0wTNFTLkQUNfDYxJvr5DC9pEbzYkLuQ6C0FtAF4y
IqFvcAMPH9cyD73AmdfRdZwELJTbYJILUa0erI6tX7EMwKrNshwG7wsuOGeDagkp
f1NfEAaqTU3Dv6i+YZ/WhUtTca6tSg2QvH3C+/7Zw1LlJ6W2QKUsiVE3YS1IYxmP
X2nSpYsigSz8ZQTot3tXhH6iWrAUw2L1sWAChI/t1zxGN4lKnNU8ZPoZzCTUCaU6
WT7b35i5M8uGn8wOLJwTE4f242EicqY71ISNTAtYtONm8J3Uy8tp+/AkJXBXKGbN
7rpNz5R1OpKPWM04coeemvTa4Sal/WCeyP7f4lQcmY0+VT7YJ+ZMNxPol7HMrXxh
o2JET80A09Ov5UOOeaE3ir38r6nh+w6/+J8PaKNM6ykOvPuoJvVbwLBM0CXKUL8s
XtZKUGP6jMtp0gcWzRBYyUQglXT5lxTpewujq5wCM3YbC4+wjrdyiKTTo5J2HGGQ
Dm7K8qDLjRHFava0oGTuoVkNRmBTesErNCw3iOCz0N0fL+F7OCY3uSO+GCmwZnMC
hgSC3LCOM3sR6wrslIV1+NYDKJjolu4Frh42RsEnasvfmwUEibpweDdrygcNJiqo
komlJW7mqu6fAAwsg5YHVa4ZB6ZH8JvGMMuG+a01I/txQ7OAiemhmNKjqhVBascT
lH4m8v8q1eCKqTy0rPY+lKHbihDPgN0DiRqVzZaNLJ1uAKNTr3sZwV1Cb9FO/0WG
OMCU/Pc5ra6Kii5H5Oaj+ZrnAu0MvjPZGRB4znkKlo2Qus8MZjVcV38TbE9O6ZHI
7525OzLkEduhAL/h/tRFsZpjSfK08WO6IUxsXr/1DoF4/4b9AsaMdzAy2i+W6vaH
2cA53nmpxaiWGx54xSISAGbDu7HFLWE355hQcq/TU47tB/Dr4pCwP3x9vpRQPeOu
oulEM7HGgTdB/Ax+MnAwwoAEV7hBksr8WV5zeKbJB6hN1/alfuT3OmFDgA7o+JAj
STCdOze9omqYER2Z3cjS4+O6yZR33xxxQf4hJzIL8/M3gRzEim4imEY70ZXaPL1M
X3YhUhLUNutwHg82BwMCYjEJDamNHdE2BvpE79av/kMG1BU6gmdLENoXNXiCZ2R5
LjAqZp9xBBo+ybqmgJBYD955Sb4kSPW6qmmmi7bKqNIZWKb2OwrKAbFIusrkvPMP
ztZiMiOITPq4NqjFd/u1eDluH3ZGCBircJMk1+VV9ppBHZl4NN3TfZ/BryIh2vsE
tasAgA/1Ho3irlFbR3SHAjJimugWKxHvHxI1kcecemG+PfpvGSsEo1a5f8W34uAA
tD5vyVXiYHl7Gf/ZQ3UlL2WuCKns2LKoBNZAolZ00GnXg+uYe7zqE69hIKkxIgI1
Cwl4jY6va1uVPGGd6MEieGI1yyte3b8pobEn6Jybpck4X8D2tU9jwVjItGJw3FQr
V0566pzMN+BhsY4/rBGmd8UwP2Njx0f62Dr3hZn1xTQLnvZGC2RUc4MK3e5LUpuv
POGlMNhuE4Aq/VX/KGbkQCniO3dwWhOstyyo9kyD5iJezF1DjDSp1Q6iB5qF0mi3
0RURjqKlxXtec+vYJzShpbsMU/XzkLyAsUOx0Hoa+wlJalgX/m7DhslDRsv/q57k
Z5aDVoBbLJwj9lRzZuG3QfP0tgagj5KRGdbLh9oNyVixFGGWdyLAcqQf4De/i9As
oV0bpteQxTF+wNe9BJymFGoLl4KHpc+3A8i9ukRf5+rv37w1xLnl9FsoVm/Aqcu1
wuJopZIBVrCvf4C+QshscUS/GmaDz0qZR8GcaMCQC5X2jc+ZUBTRBdwsl0uu2iSw
ntKRKDETyatoiT6AjOdK/+BTY1BvaJx6+3tgVcb8F4Xhqw/7pXrnJKu+nbUvXuWX
IfWHmPrMf/LRCIWEMpIzOKB3WMMTUlkZkS8GEVIaonr9B5Z+Rx/cFTN/EFDHILFx
NFukxgpz+Bkoe1g4F5pSK+M/iYg9p/TW5HBX5CRMc5Dku5WHfxzHoAF2E2IOciK9
xvS8/6/uweF0TMDBu/ILgSG4gj9EX+no45q61qDPKJqJpKZvXsfWldeDJHxXOhZc
L++m+Zj9RX2yJbVcdrpcTY01oPOht5ZUhd4nnDY1x490VEXn9AugtN9qopjrgG3r
QxIVDTxxgGvjaylR0v8x5jybRKY+OtTSeKAr7nuvqfBPYQ7qv91A08/8PBOx5mNk
5Le6iGvE6mSKTQEMTGYAA0swHDisAoBIos1gUyg5Xo4QEC/fNcWldYwtsZvvkh5M
sMKYvXoe76GoGi/vUF7Vu5auauiZTHs4Vu1oepKeypDOOORrw+QyIxezZB/USteH
6RuzOdSewIDy7J8DeeXBzU18BdgEAwhtx44Hvsnvm10NPDlfF2RD3DtY+0ARvi8x
8uyC21CYz/SfVGXVjMzMrhi8+KnDSmigP3I9v2cIXYt4Eb6kWSQMyrFm/OykYwi8
FFif7jrvBskjq7V3D8QiYSAeyWKx+awe4+LFs9XrYTV0LUwMhX7PozMzizR8pje/
gV/L/VYmjxEMQRuiPaHSqbSR7jGzFIFNtEEgp7SI25Oq0jHKvUe2JVOR1Ft8tu7K
cXlpMtptIX51t7oLDkOqfTD4ugOIKyQfq2l8gVycM+d0dxhzRRaSCw+wJTqRBEMb
EQIEN61KBSDMkvKgrI8d9xL/xPlcx0EfJL027B31np6FZJhK4lMUUcwPN+VEiVxE
4b5Kp+53eCpRt6rLeW0+wck88KbeBJye2CHUQAdSkrQlg7pe72rs/dZC8RE/DlJm
kfDm9yAKBuCGQSxBgLP7nrK/+3DZiO6bEF3oyXq50nMdsU+N4ANM/MABp72CUyja
mXMoLMfDhNiVzAwqtopyAFuRq1VMZQV3xYbcVcmYCHQ5YZbgAvDNcMEZmPvDS52J
POS3IgdMV5VnspzfAJlE1t3p/Fkq63RE9nuBEzeWCTOOfjnW1faGpm5eYhuVyZSd
g9ACRRPzOQ2y7152O6/cNfBdZGmCsBQEgMu0adHViuhtmEbuhzC/nwRa/kRzXL+j
AIZkfQownBX73uwM+7otCF/VWWFreCiuWoX6H+Jz0a35rjefLFdgxtTey/t2ybD6
0VxKo2Rxz7MUvioDsiH9MlaJPVQgaHIOPYuTiOFXeK1dVYj0wPK43eYEDoWRhGOv
yZ9HPjh2sCBAOwhzqCWGQxGFUD+58zv3wYkTH428M15xs4XbtijFpko0PsdmW0ZT
DojW50HfGjzXffHcXfN9NTOCA/nOGZBl4AaKZcnMuZ8JF4S4ca9upP4PpRSzPL10
zGYhd4XFLgrihHQ793ueDvzk4pZd26EXi5g5WIScgwQnFxlMCIqV/3IbHE93PMeB
QUgrFxGlVU3hC+lGkorxEhIgABXfSh/BPlmiKiI8cyFzmfnqzEfkxLHYvbwC8PK+
x4y0woC1o1hdlCbvqYDzyWDZYFCphHXO9edmsXqzso2+Bipp56GI0PS+Y+P6BQ1+
OifonE33ZhaXqpk3w9DBP+mrF8owmp98roR3OZRUY7l64KPHOvAxCrgQROpvJdwd
9B31JLnHJQnQvNZ2R1A15XxctCaNAOAQymiLzzAGG19IsbxJL8pultvnissStwsI
AUWMRLsOC+hYa6beN2bYAjrLwaI2CxYXiRH9KPQBsT8p/fBwDM3TEUIa5hL6/38h
Wh+WvmqF3RwAsokCv7M5yndlWNq9D7Mnns2Xn31WCE/0kNNAT9Wyx3S7dTTbxokL
b/ogMiW0IXknV+E8Yx30Sg+RVun7YEd4Yw/L+2vInobF0Fudop1vnlQEOMCfENgj
MaJV+SZzQxYfC6v0bSePQuc6P2iohdHQoOdLiRzDGYJFazLgpCeR42izNJXYvZVM
obXNsysL9aCCPXc9yVSR/KOO98iB808IUvqF6SataNFBQOgDrU1qgu9KazZerINO
THIuu2DuVBnfFrhuPnQVyRIgTBnKJWj34ANIpDpNkJxkRaPLhq/hJ5+IrGX74Ydd
Qn868LsU3WZTRwehNV6FZn0PWmAqDzfzEWUcEPZ/PPE4SO9FZOFeHUshUvXHYOuS
pVfV+biqwMRJkp97WzD+4THwT5Yu8P4zzOswfqnadNBfajTSDNKC9gePZoZ18zLa
Dp13N0VfLqYjySDrf5t2dLQiEm1LYBFlzJkDH5S3J47KG92I1hR5WuIAAbI5Ng5k
wNdAAOuqwC9+6DDiKHM3iwDOC9Ef5yx1qxT1AmFVnYWQxrXlrzPzPKfXpa8yLcaC
pwIlo4aYUpc+JpEU2hI1zcFHDSMbQzisgVzlSHUtslscN7OE92lpRaqXoICeWh3H
k5f9Bz+fPo5knNtKH92RWsShouERsRZLeN85VWvqJHywmZmUwjw8Q0AuVyYqDTgu
k3Jg/Tq7PUXD42a1+fVyEWLh/wRM4UbGs1ZFZNroztWeq5qN9K6HxUTIoOICGxLB
tFW5IreAkhU2lXbIjdc0SYJf2VzcwVvhySPbdOj+YAkQpicRapYVAmGzkqwJXvdo
5S/waOijdFK8vxDhCqabJqDnb+6p4iUwJB9Aat3nSNa4/6MF5IYPF3jIX1SA3eDV
sjwxMrvgWJDZLGehEzg1EcXznXsj5E9QMxle1R+U+fyhLrQwnWe6VbBnqt+By7zw
wfFuo+NUrMtx+bd7m2D22xaNDve8KVCpjEsxtCCW1j8BNnJQlF5UhFT0asgCsSxK
DhziZ9YHbnBNtZaN0UKG4NKUCsA4TC2jvb3b0MkS1hYt5qf8wvNbco08HedEi/6x
Rja3A5TpjmwvJVdMUTijVbXqroFVHB/fTELcGP1kF90Kkbanf+ja5c77MLsypTj8
YJykXI1WMTIKgvy3isVN37VWiflhIBuZcTGWJ73X7WI9VCXW3flx1c+1KFAACIpg
eIut/CU/A5C8BYDmJM5eRYHQoJococCshZMMPcjQwylG2NrU5ofT/W/NApcSmZn7
tVMxuyyfijVLY0OenOjzLmj72GdhLlAzzZ4KaXNARxRJ//9q9aSTPu3zzIaSsIYD
TGjcsEXSWge2ziPRJm8GF+WKuNKNaAi32fVd77G4O5Wl6LsvkzMoeisnk9+Z7vK2
j2h36CSadPsGeGdlq/N429Zn7clISViIW62f5MM13NopO9pX59coyEH2sEMjifEk
FErbZlMfr1kCG9EbRjqZcn9NZrhKn5wyMn/WWm9uAGWX745cgG1gFY3y6Mg+cNl5
oHWpPCjiTDL8ilUMHgwUgnifNqvLyZhkSrFrZVLtKrnmGuDG110khvwK7ActKG2D
zA3yULnBKX6GXmC/HvJ0w4uCZvUcJQmDyD5k7SadJeGwKPwQ6P/iqaBN5M3tTH0S
Ao4cCGplQKmDZ/YdIg7ZNYJNO5vabhSHq+x8H/LKNy4Ejtz/KV0NNZQt8BLL2xHU
gIzi9DOTecvmCqRJ2DM3JF1TlRkFse4B6HQw7zQbPfDx3LhYrb+i+ln4KYTMQhE6
mFUF3QCakk2PDYIHrExxJNxSF4JChUA/kXVasdy+4rD9uZser9sc/or4XsU63J/7
AFwPCFo3KZBWZVvoeoIEBedcHN2orCxeMpZ+s4Q1b8alZK9gcERFOnZzu9TAZbUV
J5jxga5OR1FrPTjL0x6t8c9JbmMAi72bzIii2xtjhoNS+be5tvRC9C+fhp5sKljV
5gzo+g/V+hM15i+vsjM3PZenD7eJ5mhuINCvWxI58wWetqHJKq2gL9hUzgnSI81C
gmfGfzwodNcfAVbXYSj5kAMNKhjJx6nZVRqmeApLSFblSehE6ASruh+0+TNWlF8K
c2zfgOBdVB4cFUaYFoEFmZh/TDEWFqkesBuzihz+sNamGo5GCKgSh0KA90w3vt1Q
B5Ph0yjZnGqTvGNXEzcNOTT7TBxgqgHBXvK8/gFfei4Tp1ztlL4W5wPp0JtqDejd
kDoyHLfztHtOTc5Xjravhy+Uel+p+88Fetm9UeHNvyaMBDNCoLxTPYJMWOS7WU6S
TiBTWgilDqEogxx15qaueD0t+dBt9DbxQ5/zx9BOBCLwdt/tH9/jMFq/+YycDMmY
2KuxMSUwz/n5FQB6i/8kK2Qd/0p4KHu1y5WDLPlMu2GCbhs+MtdRa2viaZPQFHiG
79pMUwwK7dtR9d6OWeGZ4z/OGqLqoIlmp1102iO4nkhv8d45iTw/HufMbeHm0TZo
1vzRVmaQFM06gzrB9XhiEPoD7gqW6daAxVapijPUodHMgh1a/pSQ4glWXFF1JjA7
ITZW3gHXO3XqZTuPKF0v8oslR6CDc8OHl8GIYiaJ1zLzjGkANmsSbudC9eBKH/V/
C+UXvqj+DC0yeVNWpOcnIwzmcMCE68YNVZgdicM6agJ0+Sch8v1oGueMN2slDHLH
Xn+UjnrufovP5cz2sftDFL75/MPbBjM8LQUY/5mdu0/fZHCG96EFrDVLeJJ4vczY
M5UR3qX7NFLvnY8m83mZS+/fttASIf/IBIJptjC7dXxJEN14NmUhMgn8c3UinOSt
pO27/NJnq0r+0pDh2UOocT3d4jDR5jNwXoHuK8n1+oK0f3CSIolUfLC+5by4Sk7o
hK3HVYi2S4hbngqW+eWbKnEPWgYghfcVFbh4Od+69CSfoUlRsML04GvAH00twolR
O5w8ZRTeGwE+zewcwhOiQksU6zvyTH/PVuOi0a9AWmPlaacr9py50yPX3xQwjzKe
3N2UjsOd8uTg+mnR8Pdxn3NrZJJ+nHMzVsXyz55zPUU3CM8g5ODGHpdGja/NQGEj
5gAktbFhGMYCRqKKfxwBs+lIdNo3i7tHoVeUoNmzQ3KiUKcv/0Afu7o43CFoT0Oe
HzQnNdGVs7V0ZmKAyAMMEZC6xlJ3ypMfhtiq+orPv9/n5+k38ZvQo+fpJzlq4+PJ
ygpGQZJt2EwUwaFP8FPq7k7GbHEeuKSo0DcCZ2771bgTyJLAbcuLVcYU2vMyXse0
1LCYtwdO4e1rEYqMw3+iLNV/Z36eQJXuTOKrU1UW5hN1WUkrZ6oVxtsEJW/eHRlF
bi3R/jNrMQvzPyc28Ub6gj4VaTshpZiDtJ1jccMX6KO+dng6MLryGHqCkoA1oBBd
bzBEuRi1otYdc28kWKjJXlm+N0UZPxQ+A4cQINJUqq3DSrUdYhL/Xc0r6nNSA/dK
mYbirmeyttpyfKLoGWmoY2uqKvW7zceTiHbzZTDooCTxqNdTEcofeGsj8UAoXSQX
D2eYFbf8BvCn0Tzbp90dn0r3kao9Mb9q2ISpOp91aYIpBzHIDMPoTprd2EvrugPi
eK9RxIqqe+ulQwJDddbEIpEQk8Al+hCiKVfH0Gin3+E2hQUqtn6hpUCBYRCM5TRb
Aqpb2825SQio9e8NUyHYHlIXQaXbmRCp8rAKbUidQ5pSPHvDbabfW9T4gHFYPXkc
8Se48IlcpQ9XXb6HT73kokK/qe7+c5CIIqr+T+d+EHCFBxGvYS0NzVcBxqGZ8ecY
6XuBbRjVDTitsLVfZMC4qBsjxqMdCqrcm+UscHoHu+LvYBXRqmxlrDtm9WeXK9Sm
1FcZF8ITI4RYiY5bKbmf9zJt6OliaqjU+nOnauQqGd2+tPE6M+hnAbMXiQ+Rhz47
zqpFS+HPjs1TK/QPD6DoL27bqc53YzGFN8j9lEGKxr9MYdG2xQhzlLXISM/b9vzY
hhcrqL7x7r5TcwP40YugoCFoJJfvCq0h+kRxV7rP7z40ijW7RfPt78xU/KM+Mojx
y/YXAJBo5BGfV6bMjlvXiV0xEji05fKfW4UxDXIPkhguzhyRTRZBE5bhoC5H4BPo
HmmnmedE2CmIvu+ozM9O9qm29vElfFmoMVKXqijncFh9rHjfvPUkGqnK1sOwplAy
m2J4p+cxqicmT8Pflk0GwY0Hy2s2CuJGUQ2v/Wu2QbFounnkq0IIAwwBwywc9SrY
OsEsV8x5qrrGjsKWJjvnXIwL9mkYj1vnhtr6J9xxLgBD05SQdnP+lxqCuuZNiw5S
tHOQaK35RvDihlxi7isY5fo8vsd0SWYkUea+srxmg60tOIIT0UqK6BqwLmVAXDmW
d15VcppFvSzl/1eZ5SwkcH4UzGLH7ZG6hk89D2Ig3ohcJCAEjlF7x2msMCPhV1Tl
3VlrURGpTT5X3R249XwJf7Em8pqkIgb02jwbcqzX5BqyVzQfjylwFWDj5XddLr+Q
jkjklt/HLJNBpcP5i5SxO/5paAgS3bWOgPKip8H/AB+xse/p4TaS1WPj2JxqSPsX
tap8Z0H++hD/nPbVCGpAU3ecCAplzGGYZC3+yiQJrjtS0vTwtx0rVCY0j1Z3wjCN
rdE1R4gahpJBIyOWamceucnYNtyr3/HEZPkdM+GjHHuzXwm1/XuLmLfyZ0mf83dj
cP4+uQ4yU+VY+yX11SRbSEYAkJxJhUThwIz0/Mc123RjiJsVPdwR5e8aRCaSqeC9
58bJzRaZZSGNFCf0bPOBc06gbkV6OUs4JKFZ7d+WtJBECDHGQmLMLpGBBMCpnbYe
wLndFb74E0QErqYC0Xl8iRpQeFaFE106lLDu1DzqUhxZ/1bGKvLcZJ8J0oyXZuSA
HG6zsJUghGALwPkgy4r1KX0ujUr/DAxYvuEIu2In7VpxOLpyuaOvF+mu5rYMEBX8
XwLb/q2CKlYzVXX67H5FoC+Ne+fsQDImjnMappshOpWRP4ZPQqKq0Ihmhk3VAleJ
9FIGnHeCycpYCDr+Tw8Uc84gKp+UrgeFJnvkYYrv42yeRbpcneU/OzXNfoX9HqxZ
yxgOac4Pr3wq33Au8kpRFXGyPSjx99nny87pcsr4hf29URzp0luRKYbX9qv4shqU
6zAd5Ix71JUctWd510zEPb0cV5wQ+WUsdkYXJKMrx5I+VmJTipFt6Vmvcje+Pzlr
i/x4u8giuUFcAbcJIFoR69erJi4y2WcXX4kXr5RiXUr0n8VTKD6dx9cCIRtEHt4c
Qk4dWOhta8h1jjNRqCXTGz4fc7fI/vZE7x+AGa3T8udIuj0znjvRHqieNEyHX4iy
dcGBUFabskKARduMPnpITnQ5FSZtJ2XBWL7SNYt7fe0p8PuZyUuxsm3eVW/4nAnw
izhXQDLNFRn5OJ/zOEYu3bKfkWx/bGaMXl6Ll8SS7nuWRdJ+GTjA3YOPrbsmjqod
8AAqeLqEtqdMZprGKA9R5FcbHjNnBXNf0FnmS0rHq9MxzsQk8UAJQjEuo+8DU10M
uOcF8cAIyJYqzBSZzNxJCAxIleKmPETulHhFPLhFV7gUdeF1+/4BNqO7IeDl2MqV
MnKkh2qncweO4oKOuIWwfUFwEZUryPOMHv1Q4NLmJEArt0033h+PIB/Wd1nsT0Q7
Rtkj3CML8hEybeW0KZNXNero3HQWTkHQcDytVi6XPmEKs9KSMkgE2MCBdzvHA1Ws
lUuURmbHlOK4lpzdlcZaf9gNfr+VVZWgWbG/UhqvO00RCt2NaLM3OKImmAZbZ6oM
Oj4E3yLB0aKJQuRHGHsI4HrEFLowNeL+D0XTC3U9Mcl/VzY5f+5ka0y5nXbRCvbs
eHosZeyPLHxRvCPYIbUECqXIcwxpgxXqCuERzo181W+UMHdgUWQ7uHhSumkJ/na4
AxoNtVVk+BMKO+bmJif18iL17EvU83G6Y7LXa9RUbookjputiipe4pbU/iqkdyJu
jpl4vzFcFjyj4xyl+1PiagFa6++4vUBM9dYzjPb/7DdoZ9isp9WiQ1y1Hj+xsthe
8/K1gCGzS/SuvYHr0BlA9EFk80gc2zUiBcnwEu7RjVUHI4EHPRrhFTpEu24YQbk3
VGvrpdeBWyGl4ypMilHIuYvm2mupLLaAIlkHQhWrGv2ub4hjUKm+yDdcewyiNQMt
uQFHiZkp+ZvURQ/ezDNF355BtB1zyr4BcYPf0MXGshAB3RVkyScdywYkx4wDun6X
t9gmyfSWLo/Rc4VTXJLjpB6ngNfzR1sQDQ9JmBEymEPJFRJbiOdH41cVRXOSPi4b
sb/W5+CY1JlO2W1ljmSev44fd1h0LSr+6jp5b7x3F/jCaW61Gpl6tYmcnUCukeSJ
uXXZ7nUtQwCZSgw5gqbz2ElFtwxOt//Zfs9x9yaL2KWFh7u4jdFx8W2LDUVVK6Qn
b00Wj8s0MKNx2HcEAuZUme3kLWZKxynzRM6wF01/FaAXvma43xnMMCG8Uh50ELnK
lSSX83ivG2Kj3bfkBAnviBmo6WfMeb1u8pU9ES1P0uqf9JP1dUKJm+O3rT2BwviP
uKP4Zh89MN/m5jSlnq0PI9YAyh4VDlcgCc1MwEjNT7UauAlqbUMWQqDMbL8W03ak
9l9GVVCfvqV/nrelLIG7vhIiv6tb6p+x5XReIRHMxtZTVEI6U4R8UA+mHv0L5mCg
8zW9YvAWzpMb3u2Relcmy+hXYyNoNGFcW/6/E9hejwotrCK4kveK4JxeyS0xn9zj
lx7DSy+QNYl/2bpoI3SF9MG8AblnMmHv/ghbBLe2zc6Y8IXwXslg0LdqcSrkYCDy
cVrv/0sJ9aH4kDXKsHGudWgVq/hvgrybuIdxq05LN7LOieK2zIsHGt6pnn9tYZzM
6Vi7+fVQdIhr0PAo255pvLUufbYP5hiZvgXsEWCxzAfRx+FipKoHh3l+mNNTTGFn
JR/HU8/NnrBFamDJWB5uhfTOJC/6Mbnqa9mXsU2CF++maiMTsSQn2AroRut7Crdc
kRl/1I3dVHhjHkeMzPISzlUaY9MpOM9/Uak9ff4A4hPiRo+OLVhXPwBuwgEQiW7D
n38EYDCBDGLDRn8l7yuU9akc0cTQLldzVawrUPWdTHwaDXGR4zqmJS/QPBt3BF2+
CMq65ffcsOBo6MwbXZ8SMX2Hvp9p/79NpF1mFAdBv8yly+pDcVpFTTXvcSh6ja+q
fcO2kgDOlShk8K/AVzGWcSf1Mhpjn4sICT7tJ7UTzC+FpYQK8WdWzThFqVEeOh42
ifE3pTczCOEqQNQ2RbW9GaNf8jYq+imTXYkrLApLQQJ6LQ/pD7fmdCGWbyIEOJ4s
PKzKDzvd7HemZEOlw4DI++l2k/wyXQUKp34q5nvfedVkc7cFZ1oE8AvayiLz2jMn
lCVdDh5Kop4AUQJmWJRQWcSzx3+fyGa5vb/1UVjaTPqUUvhOjuSsMPiWw8Zaanh7
r11bFDlKLMZ9YrDWMUpHTje05D5fw68eW+jboYNJWf0skoIoUs9LduS8uobIFwK8
urnS06T3TkeCgxYm2D5U0eWkCfazfReENChjAR/tfZBPZARupg3qwcR8hvOr7b7T
jypodL0o/5jtog8OTaFp4u1xCv6pwK5F770DR+2aNgVNV9ItQWdCN+Gzio6j2mKa
hNRBrMZwTVsnranjEiFWxA2mnIj7Tx2YfEdk4bd3Rzv+Q8uMo46vvaT3/yPCeWvP
xM0ARahOqmWhf7MIgLSlUDKOvMP2Mgvdi87vvoRAW3TDfjYc+jwXdEEDLjQ4KUWs
uGrHxojXl/L9ZZr0GlP8WskcJHOVdZNFyRW8WEj7FHXtTH0ZhEHN/IAY2SjWJo7t
R9xFg1iheYRgCnRSz6Ck6uUs8POUjW2SavCfjc6YVCzh9gwZo+60sqijprpAyUtv
0zGDcxzz1Rs9Q8XGgEqOkC5lEfVCUuKXGSEh+jKFSxvAWMe9zkEh9FMTk9K/CzBw
Oke3w1Hspe5EfDZ9M1TLo/mUdiwrSOgwWz1/AXi42VH/9ACYwQ0e/GeqFupjwkqX
be9kw6dz+HRhOvEzKw/fv4CpN/GVlFvNF6V6FkiYB8zszclXdIDYButDoZAaeJKc
BaVaM3HpbgLfC3tsihb1dZ8URCAwDcm53dx81e0nvBH161rKwdjrU5zu2NIb41+j
XJnMwLIWYnqA9cpNorjk6vQY7+GbQo04Q4OYKNnUogGpgbYccz1Js098fhffuj3c
ixpsxax38JiGOpn+ckUZxyXa8anD1H5im5k2+mju1xShknU/lQWiPPRP7XzRVZB/
pRACje1dS0GTnVXzANHbKw9jZkr1vo2/YChqkyDluev5IL5BKTPnFhwQKSwQm92j
fwp2dYmWcVtl1rZ2UO0SZd952XZP30t/qW8zWX5P4MBA8xC99AJdThfbvlNv8lyQ
JcoiOWstLGeipJh/NNjO0U7LEjwch4MXB0qSwTXijrpJqH1NQW2pU33QBNjMNiug
UrTQjW3mgLbwywNJJShapivxq/PhbV1tCyxk6y2egioGkrCriaeArEkP+kbucS9m
Tvz7cAZ/EAiHxpJDAl3RXn0/KpbbZiEwOQvLhpD+5d0VM8sCeNcqn4dH1uaOYhKF
WwmaejlXk6EEKJV0Q9Wa9X/svRpzXNuqcLMvch07DFv1LkBuFwwSq2rHBAul1rtl
Dwr9/9qFJLgXHAd8U2SbSgXcHW6v3ZpH3HQ1Zq1l3TdqlRJxf8ka+ZCS/LCcN2UN
EGGEMdC6sAq0b7NSmSObcHrlbrjdVaR2uY3DFJtwxbWXC21iWfJhcFY+KiqjJk/x
+BzIlnQuLQ7z7A1u/ay92pYh3hqyoIMjCJNvXYqxb0envg93rBTgTMnuhi2afIh9
5yFlz3gFa02Td80wtDwirz9uL5phcUhHBQu6KlN8mq3N19t9VSLBAA1x8URoiv7F
vGfeP0kHpqw2Y3v/q5Js/5VbLzXEKrKq6lL6VcBSedbg2LX2A7J/q6+3DfNqmHK9
FjPVco/JRxtGQs855DlWFcTBVcnZkxOcl8r77f07ec20FWw9qTDaDTuqmOUTySxn
PTVSlB06FGHBW6SHGalIn/LjUMRGEzzxxGsiNZqV2sI3dVuf0WcgJdTCICZa3gF7
At6bEm+Hdjr9UUItwI7pn9iwyEBi94XtmfEC1Q0xXUH6sb5x5deXCmRYnChbOqZB
S2nW++bZy5xxW85g99vSTSW1APu3A0rF7BgmrJFU34fQCmmpO4nC0K/Wqvz/HBc3
RjO2Rk3K+E/pnygPQexIuJEiOl+d7SN7/5TqRXOTche7iGtkaV1J3rC1lXQTiRYY
dkekrWc7vqa8E2kIS2EqrlmRWFsorrmryXPZoC8LboRECFdAXRmnsOifI90Fy4dp
WgOOT/BuulV49PSh/C3zJF/5q3mHPIvOLj0is9lTUeDVHAjW8jmJiFoi5zf2Hjpm
BfiQwyOO1TqIPUYkv50PF1IlpA2z13JhISTweQTPeYiowc/P/0DZiESV06K7gBzQ
2PMSwEfQ9D8kgwU53fl7cT6+89+P6u/GPf+/N/uSUAzd67exmr0i9Pel4YNOmuHS
yVXye96QXa6fd4Xv/6TpfOEsg3wzPehyuSFsl/bDZbqh1smGUY90P73o8f9zDE7A
pDxi4TMC5t2u2SXfB6ohg5vxxGy4TKoOJnPoS3yAVMUB6sWq6/XJWD4w5ySFljva
PpvMRYoWv4xvMAeVV2uhAClEUIgajqrVMDTyKi1ysVIt/BN8ojvaP4VJsZtwCB2s
sRqAZc4f8BFjkr8JnGjiVpwbUw4fXOxnfHVa8ReZoXQ2zQWVkJ8SDC3vKvg4UEOe
tHUOI07jNEnCHeXMuSBOqvONn46C5CFzbtiLapynEW2xn0ZPHP3241orXLCE+MTL
Et/uf//p6JiyDUXWvAXQc0KU1dkkUJgbcNHvPzCw6GhYQ9rk4QRBq6b0W1L0aTJe
JJTMFmyLyqOX/WIeNd28uyVSr959nDqVZWW8rfON0TkDd71iODjCCot22p5vy+HQ
D+ol+GHEHLILC/v833kdzFBDHK9zivPwwKVOGt1AKpQIHPSbcg2lYsHeHTH3Ijip
BbH2uHoPKVYe/wJCZpr2tWmFSoGnLLgXMJMauIkhaagdmCuTOGe6Ih6zEecTVVPi
ttUcEVCfSgfs0PUSugP89se8oSx+iSvpL1BzJvANtYhbI9hWD5dViSltqjcaQm0W
Vtxr8hd1wMcxBnycu7zCzJ9qyI6H5x3lTiD+McUStTD7vCvlj9gTem7FtrZD6t0T
eFDeusPfwhx4azyalW76/0STOnWRplJc4OeNNsU0cxwwLxT1Q1AkwJgyIAmayIq5
EisERqrEeA4517Y5wnKyQOh11kIcVJxV22j6Kce6w3BF5FI8SXLzrYRjweyEsdvF
Or32cu+AlBiQaP8HHt4SH4GZvKXG4rJvH/7bHjPavkzJokwHT0YXLjCLri25Vdt0
3btB3UqufXzZRY/rKmGhKNdli732ofR/Avc93wWkpPlfZDgx/0NHOkJYTrbSZRRT
0uAuk7I749SGva0DGVD/tWl1lfYDfWOVzO+W8JPBVDQ0IaFheMXowFhvNwV5eAyY
hYhwgYYDPpeAd/E16u7ABy6ZXKSVvXUdX1T7Zm0suv+hdyq/v8vJpMVjRenbz4Vm
nPyh4PNxSxJduGETJId9sJUo9wz3PZ6F1rG5BOOLMcpeRsMeOkiMZUgyDEsK6IxE
E6uzY3EbsIQ0XCPuVGCqjjEJId5GbcbBkRVQHToFUU4JkR5see9jWbglYJYShWKH
sIP8FWKLHM3sUSrqD4CGk6G/E3zQ8kktMMaOJv3YBBFzBscfL3G1LAQPpaxkk1fs
IW08K86kGKNwWchfa6ZoHQkYPjg6uQxpDZu+HsrRWGyOzrNFsLnuau8B7UKsCohf
FmbPPq6h5vA2kkoBqBJ4gX2wZ8sSpWi9Y6T2OGBttu4S87tgA9M6o7P/CGAHcL4+
ba6SapEvDgaTQBGOiYR86sASsy7Hih+zO0it7HnoNuwz6Aq3qHkpvRGmdjGpIoIF
UOS6tZYadGaNLxWhPZsTnsFYWoCBx9R5DF1l9GhHv4/5MH1vxgTl/SygXr/wQh6c
JTZn5ao+Ymk3Pl/78n+3V8TI24Vg2JyBzg/vMBqqWKyVzjKB4RbcOPxMhWtCjfnJ
3M+xduu+3ejO1omW/vWs+oY1ERP/4Itrjnbe94AsmwVqWzL3gjLnFXTrxfiPJPS+
4EmoEoCzh1TeTK5qV/3cGljOCdw2XPCmx7XX08oyw15cr3vQ9pFMIvae7uww91hj
KdJDJOE4T9nF+PDpkymDN2qmNUmReRN2RoC9g5Vs5YKtff3eZpEe54cQtS2yBz5f
bE+aj6EH4RrGpoky0uEvOMcansEIFKxny5QCHFOmvIPBiX/VKB3zQ2Gw5qSthL4F
65+tYJ2qKA63CPQM/tllLZmq0pZQtil3/88AuvXs5JUSuE6eIbppzdKlUEwQPFYc
jqgAZuwTuk1iXi9T7c3fCLL6fCABw/4D7XtLQORiub+vRyHFuF3MFmJ0F1zOnwtN
GAZakH/rtBOgnAd2LY4SE7jhDnkwAxnoucRy8E8AQrzSzLiaf9CXRV8axWI5cn0N
+cetT2dc7T3pUpzqACN7XCT/BFaLlDEdGREGDNXCl24qrDnxu4pI/vX5vlKOmXZV
oxxIw9TdvF34P9HrPWvvL9B1WQpZ7x4xns99qJ8qrTb/aFnXfbbHJmnlEah6Dwlm
aY2rfOn0IiysKZ1MkBVQ8xTsBrtwDdopYIaKjlJs5FIE5wnzVHBuzBzPpB3DPGYq
oXQVvmzUP0aS13Hz/Wy6Kiewk5qjCWU1MxThu6aSMDEhgImLB29MuhpWFDpT7cOS
MOjOkP6f9EhEO2iaYyXbqoYt/hLW6xSKQlV+jcok0BO+S1aYDjqeHTfIWhJN+jB7
nwiEuARMzB9LQcgiBqMrHFucund/DU/3/gBNcFU+iYnAxxBGuEYRYSFDPyshYDUR
fkqVZ/opp7NIDwoTQDhe3RjEKN67NrCiXQ8k91/U7/y2pB5lZIrc8AlK+PPvOudI
/gsY+VI080UbsHViKdGVafshhBPaaSexnNhif4mPLVnk1e7RDpYcJ3OTDFSvyeLn
LogUMjOUcXm35SGdKMKQ0VNnGJr+VCSs5NvLx+AYuEdttiJ36FAWxTOZF3AhDqgc
fsz/DcJhiUvEygxHgxUhPXsqkWMs8WoLEsIqkQPQHOarhUzYgboOMm+7GiG6O1vO
60UBSw8qFT8Zrk7WEhR3X8XKLCRV4vTWMSq100T5fA/wsjqThTKAvRroHP0ts+zg
qMokZWvrITm8ZBrFExVGY7hqRQ17miQlFOWNmP1WOuXi1JeQe3+QlyTz3/Es+hZM
waF6m9GIiWtgq9P3rY6ADZ6vLMrWGXcfqoTaxgYYpuAWzvWhYlL0HlgbFsCIWXmd
u0TDy/rJ+J/yvmXTUzxPPOvgaPaSt/4nX5xgO18GVRZy6KvKg5JwWnjdrOP0k74v
vDPmKRP3dYrhWgpdK+RmgfY+jCqT7CRonXSkoRoZFQCAgoQj5KIZTHRI7puHeEhS
4xdtQqlw5ePc7C5kazJMwcH3HOzb0Z7eeBLlsRZYH2VbFh38U293uxKYEED8Ciu+
VYrbviPFKZT9tPy2JRopcIMVeTOhv47cQgr7/GkuT84XT9fLeKeDejLR91B7SsV7
tm2B3zkBUF7qRrCXItvmBdld+Vv94H1roFYOKuGEwdNXRikTlHwtuOfGXnscAXAB
D7DcaF/MuV/oV/tPNg8yTnBMMLknYTfiRqWWL53uoH26cSldr2eRcvtx6UGnCttd
2kKGNU+ORVed21qG9uTxdJZq7YW+mQ6JUGzxNadkZcuDRUKVF1DpDcsWlhE97i2r
s+d1vxucsKbihOfyZes34MwbBypaootWCYrvyV9fOrlNRiJY/5IGhiLdhrLFZg7W
nzwkR2s0uOdbIXHnF3SAVejks3zEZmwlXb3K0T1OZ4JWukuydYbtq2EfJpbShXMy
LMPgEgN5GnIzHhekGd3oEwmPMQgFOCNUzKdYgdKgYnukJXmPLz0yht6zNGJcGK7e
KXjf2ujQBaLBYxO8eQb4Bz3IihndPoKFX/7xX2GJ5HSfxTz75cA+SrTGt+3M1fQN
ofZwxI1CHK5ByWKzfOsIfg+d87WN8Z1dwwJLUapPhVK+OBrgN2Su3/dglAc31oc4
JYmQgjYBvOU8OdsXOeKTh+AhjOElzVU/TORO+Ove0KRzfWG6lmGs7+5Jwz+h15As
WV0bLQYi22PjlEWqEXguAH9kdszfX5mYxCQ9LRIfWrk1+0n59G97PZd4COiGN35L
xArm+OWF1dS6AZdO7dCGRaLBVswR5YwGj5R2nisNRvX0g5cR4UxcWOXC/1yACcNE
GN8Xfm3tsj16u33DGSMjyiS9FZ42KK8tsQS4DPe16p9b7AdqC4fAls20B8+qiEVw
RUXKrtQQbROEPCQTgH+2vYwSwx/iB6EW6TsHfyUlW4K4twwiRINrXnCXBJOr11UQ
rTO5ZiaIDLEz155zwO0OdqVxJClDy/Ji28o8B4YxfCogWBx4t2tkR2MJVdeAewoc
Lsx0lt8wUF5l1xJg+tTL9fgR+O4Ht4Q8N1sB18SAJ6evsrL0jI04lsdN4zmhJF4i
DGkvEIG6a+O1q5dO6jsm8/zWJly95O71KTcbVmlYHI8fCbEt+fxAreNXHTQDg0UT
MOuPELO0OpvG0szJLt+MJ6Hv0gZWP1WP0pZkXKUXd6XsBzXGM1iVe2oT3Huvu+ke
2YTxcUFzdWq5Lm1veyNegDcheXGbWnoUDB+vwgk1Hv/ynndKcKEbmBFu9Oz9euEC
eWD03yOrA7KAdcoVSx77dcxAk2/o6ZljECG5zI0k2c9X9d52+kTAf3OledEGl2Ub
bMcZav7TqTR9c9BWAAIn9F7X9IWNtlnxnh/zbTTRj/IyeUQsOj7y/FirH8SKssFI
89/qEcePbft/TD8MPO47zI1RtZy4SFKpWGwlJlb6N72t80w3oVqJC3ildwBXohTs
lI5LagAB8f3H6GdJHqQFeey5CA4C2SGoVWZwOwWq33KUMUYc1qvk7jlX5xFLpPJb
a0BsrZJPgpYIFH3i8J7MoEdzm/2P3kD+wa6bWed8+9U8ol8LJd25uhJ7b8emGbqI
Nr7Lq63dmMQlHqR1f+v2yiVb6zkydPtn8X0IfBJKvnF5cors5TxPaWmFieo0sPsy
Zv9RKVWN2yLHtxPy82NjqKJJFgvqbN2EPcw+5tyqrKH18x82bbgMlINwqpXSHOmY
QSArmUpWWfNP1ovn/MINUdrvAXXKOpXA08O5FPKBw3nW7pgDaUozNGh/NJAWzAMd
xfWQ4yn35sC5RB04TKzbcglY/VdP21TeFGU2YWnCRlJ+bFFIDkRPhM9fydXF+2lJ
hXGNwNlyFvkv1IhYYwHqPnIRPoaTizT2PJ9ZSLCjipE1oMYXnqVd4Mz9RyGu5Oqw
ljr8LqUSB0WATbQNy61ZobEJ5VCamn7yaAO1DGxRFBvVIRK9RfugLwhqk4hiNGnk
+M/mVZ4sfnMtR/kQuc/FffArJKMUTE4kX1iNJ7qo2OJgC0DdOVdJgWof9rt6JvZh
wNdNHCj0bqDE7Q41xz4Z88sN4KaXYPzRLLV+XDR0gDzWACM/e3LTz14DwcOaBEd8
3Uhz4NegZXLBvOBB7s7C8snanQMKaD1ctHhzAEI7VQN+GdamyOJSOJiEaJCH//vs
LF5YDRJuD17WALZh1cEMdcOnks0Ztwpmzp1xY3fC2MrDeFgWI4woPL7epcKAtBqp
CBUjRTZDxAMlnjcZClc+J5wwjanifWCB5rxHkZut+CzkocgcJz8sYhleCyDnpgbS
deGfnz910kvCpWOi3PHEJUadLV93MdKn1sQaADEv4khI1BreBXh6tvsxqvSmE+z1
ha5/sDrIxMbHohdGIVzuXbAbyNoV6hzQvX5XwdXEaVBmQ9bsD7oAXtlDbwqCYB4R
YfG5i/mdRbomWJ0WE04Fdw2cZUTMQZBEM5xsOVoVe9D6GXQTrXNzLscG1HtrjZdt
COPxhaAEq9shebRgNR0dXWbE/GP3RiuNZL6EpLOlvxEvLx21/n9blJUu+LP5C6fp
gaayO4VG87czIWjkzidHlLqw7+4M+PuQsEmBNSd7Z2LrBeovp88FKYylNmkoFTC/
IshaDT5nNoefErDqUubEBc/JBPiOojdS1T0sWuRNLluXfAqf3+XNincdtJTUodVg
ATvQVK1yoSRI28ZTqA3opWaf4IqNTu84LihUzXjsJMjJQG8uamo2K9AJ167eA2UW
eyyQRmF7BEzHEsiVcCUg45jEYTkO4nuKar5cpX4sZHfRevU5Tzgm27j3WhkDrmzf
7OnovUFsrRdmeBhlPqKXEHpbnRMaHsH/+qSdQ+m3O5tSLh4Ys4NFAE8W4zyb1l6+
YW3Bh/ynI92x+fOx1mwLCZRBe7LIHignXwcaTo1WRY8mD+RTMMIAvvtpy+M3CTj6
M6czNDriAdFuiTeClLJM7Sgv7IaMkm8DKobV3S+w8TFFxgA0v8fLp+g1XMZ7LtVX
xziRBZreyY4hOyNcsiXUwFslDR18P40te+pYpgc+A5tZs9av275+eeq9kit6p1WB
0bi/5umjVBiGSPGgznTs1jc8josyHWqU6YNc2sph2I+NUlhVpFvLmCjLPs6Lgq2l
rOGXSW0K05fhg7SsfmRk8xu6r52MCYDdceTOFs7B198JDgdfnHFbrNFUQ83WiKBe
JbDzDG9epOuF54BkCTGIf3ZFOrYRWUqc4+AuwQGglbzVW+/kB3SguFDSdbeyhB+O
akuyALdPAAzQdaa5yoZfq24tVfQ1zSTZGAuBRqVhVNQlSkBD41psdUOwuC5cQsNO
gEsJq4qZwu4QTnkhhw+g1TVS7orKa6BKlyW/ZdroIYUoXmZnBcEaubdbMjtvm2cn
m3bLMOhTyDlPT+9hlEI5PsfR1l4AqS+PUYHZ5n7jDKAuUov7pYzgdl4izD6uZtaj
uYg/gkUXqjHBmqOEd6YyihIYKEVI4x8oLmVdo5cC/lrHM7GQ6oHi0ES73C1AqRuY
pKDv4QfxCmBtiQLlwy9VUTn7Mpqz/X0sIkDT+sT17pexpI0ILQsTVAOF3deNgDUe
v19w1zg2WbR5vFL/PWyDimwoyjuTSIHZc8BG3T4V182wL2J1Jhlv6+rloQRuRtZb
7JfC0DQkvUiUv0AK4yCCQnQWcClOrjse7MaplcATw6s7C6XcLgN7lXzl262mKGyW
kBOcOLX7TFvFlG02PLdZSDVtr9sezq2fIba6JKFTFFsC4exXasTYI4RQ2LDP/9nO
2HU24o/JePLFY7U/PBgpqGNLOsycsFR4IsMYpJZkZbMVyA6W/vbmL6lFI2SnzxmZ
0iUOpycvy4SoZdLCSCjFXdqQhn3gDcCCR/Ehgi/s0YGQffXoqxpjk7wQkQ+o7lzL
ld68MeBWH27GIvQhvwyyfEIvQfHK/hgfQBS2zcoJ4vv0IB0hxLz+7/NknbkKRFtc
jQKjRj9DQhiPeWS5PwcUBle/KS4DVwU/xG8r4n2P7tZz3DBl01mJ3Rctb5PQRlKC
OEsOterbq8f5KBSrGOJ3CHBdoIEFEAwKkU5m0nCTjOxh6FFn1N65oljMPUmwNtgi
OkR60/onTuwVvFt5zfmZe3i7cA8o7T3krQVnDuoQKHjfjsLa6JS3HEALewFUmiAq
TVWI5AtVZY/fQGHucQdEzbXhIGLB1smp24S1FMcO0UAp2vtxzYJR6wnLM2valt1P
ObylmVSbtRmDYTa3BaKWvoQoLpf/nVom8hCR9gXAoh/f95TXkFXQvo1VDAdY+Zo2
J16zI9Mv4R9aNfzIY/I45TO7tFo/MifjHex2ut9QIblJGf26bndbA0gMyG3ojIwh
0okyRhGQrY01aAwVtIpMsulgwhXOxDbVLIBf8xgChrCEicYFlyZcL6vz3hfTYUJj
4e7d33qxZQecaxaOlJgLIY3il0S4qTryRZVXCT+1bpzyKjhjIE4vD1TMXewM85fF
WCZBxehQaydAD0WnO1i+rTCcK4Sy7lug50YyRB6xQh4b2xl22mTjSlv12GmGQy/C
u4nqFCGcEumJpulboyJBKnF7x5+zOSLy8/LCCzPvG905WALnjGbQYBqeBl/GcuhY
fhlbXtjcywdX5DievslDPtuDjbk3g1lOHOTLK+WT/+czGrxlPoQSzqtXbUM+Ij12
M7SIN333hsrGJlSUdp89gli2DVF9cHzwmFZyJ7S1Gik/yOltQkUG2e+iAtFwbmQq
bBeM7pYCV5B5opR0QqbCvRcYThHG5kSwqU4YcBeVrvisEhClT6BrOsl440MsZGjW
WcPwZLAsQTSbB8sHs8pwl0JJLRLG1NwVBi3+gb4pQ25KGhYEVY07GtGNvirm6tSX
Oujb66txw1rzf9xZqWT5/Y74cfGcwnyG9Z5LMqzI47cUGF6qlFIFH2VoY9kenVSu
z1GBEvR3gt+qOY0CBem2K+zVkF60XMWO9CFeRm2RkxlV2njFR/UVIsqsB6rMpt9U
JKoEjMIMHoazyMqXvINxYvXYqetUHB6murmt4B8LfAlLUelOA+vytP3u4KRK+Ras
zvabnijar150Q1Pq3W9GIgsPbDfbzeE07Rm9lqq4YqJcvK072/8Fz5P2Kra8M9lg
omEiJTfLpVH73JgPIUqNk9AjKPUo6IFMNctc1PBqxriKCVm1+/vfrvRePLumV6gN
2RA2SZSMaQNhVBXIVvOl9hE0v2w6ItaZdzsJLHgMqg9jTiQu+DfL4Vy2hVdFBhM5
NInBXkXc7kf2QjhjgiQQRM5VYQ0tf2VvjIBNQOOLC315ux6kpc686kHwWEFtPt1n
4rr73E6WhaO5h9vHm9i+EvSjg1qUTvbtd7D9OvfMg5B4btud6o5MP6MSkSlyA/D4
AcUJNC3lJXdunCgx8NJ53MVgRblMzAwo7+xGUgL44OhaFDzuarZzs/YX4LrDkJux
NNCPpQOjt4ssSJLPI4e1zwjL/k5LcFR60sQ354gDQEx1Evp8F3fjiDvltLNIDEmz
lbpIfACQaCTAhfNRjzsPzFQH0q0JTj4csaqYP7sj6ylWvxmUhlaR+xMRqsmOfJvJ
vEVbgzYJ9oHSMO/IeeQ5n9VP7j4DC+emmIANmhzcQTXFxyFZFN3EfisRyayKnayy
d4OeAvuJrV53g3qVOXvP2xCRRe1hSKd2Og+oWx/oVI2oUt16VB9wy4GN/0wW/o0k
frJriFLJGM65875y5XgY9MZer7k1PMWBF0koaZCaG0t/ycxAsbAXgFsYFWuTo33t
wWOJXXulssB9XQ4X6MGopPEsLGd1AQD5NYhVNHdYw0bDYVhu1WjBDn1by/wNq/fJ
EWsOFuFRYww27yWiyV9rmuY6v/ivc3/cFxYVqEJXennqlLYH9uNbwPqX91ewlJCj
ouyPL0S9tpzYK7O/K8HYeWYhCgPd1QT55mD7bSZBlkktiWL5PEE6GiIt1fsRG2tS
BiLem7u8jO/EcVWo3NZcmBdV4LOeWUMb16woaGrP7ZdtFEWvglj0Vb5/whvm7hr0
yLrGIzKLMWfp5khx+GiM18Fqi3n8cn8tPC25asxwsCC/Qy12pPscL4t989FkfNcE
rrrvCNaE83b29B2yei0bbGWZOOg4iDQ4Dtj/qviBUGFqaK597R98HQfhZl7mbLkE
ar4g1kfk55PG2nA66HXFS4LG4AB8/WdTHt89jpwWC1oX7T9mAtcBN7ietlIiH/6Q
P7DueHZovy/Zjte34kbY0gjU4jDg94k2E/JfY98bbzM4v2B9EBf8Hj0PYoJy2uZ+
rbERBkwqqRkO3C8h2EG4+HZ1k3z2d84ReoUeZ97QbRxSggfOXNQYP4RIMVWv8n8V
xtk03ycBEN9+JCwfZEdQrA+6ONGdBd079ZIwTYb2ysqcSUqW38XYHn9WrKhNSKP3
Q7iCfdsiRvqjVllJFDbt69xkOMtpT551wF305wX1PKlkaJNAJhiSlGiZnYVo5gXI
27DL1rSyqrvZey1UAar4Pj8HZ6ycAJjmaWWfjfplCWIc6FlgML+Qi6Gau0LTlMge
YTXeUvurSR03wU2ZSmP8migdzmNvoIQIdAwWvowGHJ8/aboDGVE5RWc3nkW20+yl
KWNkdVA6gFDWUriLHxVG26AM8lFwZk7rP6aq1OYhzF5w/lRgICbwhlKPk3wuWvvv
oPI/5W2520F+sUQLTW1CXYsAc7SsTC2cz+bYjTh/RWJlfjLTUOvNuW/2f1tTQCDF
uucjS+d2AZ/8EHiOK10Gn9MMj3D6boiTzFxWXPA7afBsPnXUgvURDXUnpX6+9fQl
xY+xcEe74LcrdBs9+vbyizAnUsGWq0R8iTR3pQf/QHfqKSlv7vRovgnLZQZ61Ldm
DklMoR8lwsD5Did69cApYxrvtZatvKCtVR96tHUbXPtsOeV8AL7dHjYTg/gO/53j
XjzuTDr5oQSasDTDbWAsdpZiYyAshqkYXiQrsxCqA30+z/RQ1ANOLt12VZphMStq
MHD1HlNLFDU2rTPcjRwO/ogMUlsPLCNLgt7fr0oSqkzuktKO7Qu3Gc0t1NOJ+7CJ
gWsF+HOlCHfxjsdsvj1xEVfoBYcoEkHtDkvKNjBZvpUgG87XjERKWq7rwkmKPX4X
/VwexuEzVyYREQIqJJxCz710Hu04eiESSWnvtGLRCx6sAA3Nsj2CKhc/8PrH3GkV
UtC4Q4spUm3yu9xX8a9q9uXzSiuAbgqkvCZpXjgsgEP2oBdjV3Aq3b3QL9x5aJr1
6x9+XB+jK9wEQWlJeOjvAnXdgnM+wmkDfzuRaORc2Z+hmacNgPDaKOxehJ1oNcwQ
Y2Aie7wl8jYIzUmcD9Fz+bp715dSY2EoCdI1pc5SJpLd/aNbaZpVODsiDfoezxJq
sx3pMpWTsOqnoN/DsMkly+TSNM9b6Vpscn33Q0v0t7HzpkKl1wNtMhwmlnLeizML
rxp23+TSyzcxBTwbSr7FqlzUb9N3LLZCiHHRIRI20ooDKZ+660ecLAzd1eqM5mzh
rRQUNMATSOyLlionImzO0Pzj5G9eqtfXSz/xR8QYb9/D1fDKelO68eFwiJeWRG2D
9g0DNIbdbr8PyOrIoQl8x/xTxB/MKGITQgo4qbu63UvQHzssEJap+m3rKm+bO17e
jTsJZXd3H3AMs8OEdBkl/jMeKN4KOdQnfO2qOnchlJcjRFqPy8G/d3NTU6F7y/dd
BIPBAT3elrBxQTPsataML9J/cuItno/IkIwA6q5g2Q0LN0+/ObaILm6GrcStlEs8
0nVpWpdXu5/74Md/sOpxPKDpdlWl2TDWTxltB4k2gqL3kNRhvfivxZ2JizE2zn6H
3TvK1TcQXpfqAXDmCXH5Kpm8SyK7vMpAO/3ica0qwysXK46BfEtO9h4fZTj7Uhr/
+7dqNgk4Hfct69zMjaXrH7zDN0ndJ5ykXfvKIYusK9MSKePd0zHB3t/O0ZnuGzYs
5ZS0I4cu3D0e0t8aZPaZ0ZxLWqmicdaBc5IqTPUA3opyNFP18Z1G2tZzmsNltWwm
WiXlq5suVwmiNNbkuRhnP66mpDdeRkRxXR65pKCpcryeYmZLk/snvzhY20alWPcY
Ip/jmN5YLsHk/gc3TaDENUiaopxfUwyJGL4ftM+5LwmBQCp7m8K4eN352LTMYpE8
lyrnZZJg4YNi6mH8ckDpeIDG4TgWaLNEQGelecB3qEp9PlOdhwqdGfgJ1zZu4MyS
SZ2La4AW9Zn22P3Y3nWNBbKgZXroynpO9VTWRY6bz/o30srMsQOMO/WSmQszObrq
oBtijb8OP17wsrPJRhQDwF9AZKQeGIssosbWA+qUNG1bmF5jgnIdfp3lDfLi0ap3
WWirE/BayQD9Bt8dmsztbLN2BE8T2G/E83zFYL9PhzDgWHq5Dc7gOa/Grt8CoNTS
DppxlZgReC2Olu5JxXHo9oYICA4f3OpvdZvGoKptJSY/Cr9ajZn1h/AvClRHtaht
ueC6Z2YRcFM4QLAeUpSZcjOEHfZpmC/yHU46f8yCob+FZeMJzo5aTGoQUiGnBoL6
pj47oC3swPLlEWDJd1V8ofTUdSMZzohzYlhdUbQiXXJ+NEaATjFcoCTN3NpwjDti
IyJBuicj7GzGMduzjrAc4wTUooPBhId3OfYvTPThpI1fRfj+3HMdWSYPcrmQFXbe
vfy8FXz5IuR1BtZYKtJAnT2DlgivaaeoZzuxfalEJ0NLVltHT6H2tDEE6L63lTPw
SP3Knzc6OqTdOY2NuLLilBuUaM4t+AV6Htu4sDLssFu9rBbqgQrlBr5qWr1vkVa1
leCOJs0rJ2DwbC7a4cAKZWkz7skOAR+Rmui/1JfX+rsCPQB/gqHvJBbziXkB0AV+
h5d1bm4q6cKojQIkWc/D+ViMN63lJtEKxVKQo+a8jDL/O+sPkO54t+Zwe/WO+l2s
PXRF+EHsdvGTA/9fr3Be/PZI15mPexuqfNxO26VHveuro+qoTrnUhYviwrg7s15Q
IeH1v7WvhtA7xPLz5QqVIdOad00m+2QaZ7I8OMDf8GpsB7BR/JkictGvdwFxsic0
qaS+K590OyxfaeUNhI0TlZMHpMwyscqNxdcqUrWmqzgMgcPSRroptdArol8u0Ik6
M3Cq1/YMOt1o22aS9QERQyggjSkZy6ux2U6N0IdhmcBWU0Joecrt73h7oc4slFjG
kFvGvQR0aZkIlB+Ieox7Iv1cCLZdzviiVYHHTvIWdyvmx2PGmjLthncP3tc1b6gh
JSE5srVVKLWnGnZ/4dT4mPLfdlGgyYaaYEa29kjE2cKsVOaIKp29AlRc2TGEQtIh
V6UXpXGVH2X836rF7px+OIJX7uI0HsPcCs/WLWjyxk+V13MNc7LtN72X9gsmAZSE
9AP76FjUrgkY/IqT3GneUl4v3GYgReKSXqAPuqt6DdKIwPGVpNgmqhbHUI0KZXmu
LrRuWYnYDOjX1yG3gm1yduuZXcHRkx6wI000UR8tnHKXr85ZH/wuJ8eyjVI28b6X
fnKnR3PkMw0W+kmu2lvxdgwZSlMypnJT+zn7Lg9Gpk7BTecBlFVhzcCld3In1KNG
mFT50B2z+H70gaWef1kVx4iuaRizDUEXrbcdaHevjb6P4O5j5LtStLI0mHToif3D
9OFCZ755Opxs5oN0ey1yOAo2VLMI07/JfW4ihFPGnIZzolUd6PrySui4MVCPiRa/
lEI5V2ybzuOzhZaqA96NZGzns0Swsa0KJupBWGCvnlJDs7k/6v7/AGFq4pn1s3jP
dD6P/xZTHo24wdwQbM+r5ZtO/m8w0DsB7aIq7NMH95ttnBxmkMEKexpLOvSWEKHX
TVvmQcwOec4ePnpS6fIEBWJ53mT2WNZ2hGTqrkf4t9in5/oLg6M1SNSRU2xB7nXm
LGE+mASlSdQOwCATaTe/m1dld1uUlu/rrrg/rnj085NnBoNxsHX9S1+Fy24DBBD3
2fOIcQxZ4aJ/h/IEwGWCbRDgsjqie28jmq4FSdygYJ8jR+3uK7pX4tLLHHxtlnGO
swCcQl16WvWO12dgRahll97MKuaQwvvtoi2rOGlO6xqcpqODz9n28FKxNvZXAWK7
kQz2QoNzYQTgNo6QkQFUXnIn3t9HZjdmOOvYuEu7e60m7xLMTpkIk7+VhjNB4ADX
QybXqs8RpbWGW3UFmAxY13qordBjiZmvls0TZJmtMhFVvo+uYi8zYbLQ6r6tdGzB
8CWq3HZ2w7sjJMhst4gKyxnNHqaSOk/U+f58Ez7wsEuRVD5zcDuYWk4iVXTMMrJ8
orLmzN84Novhl6zrHe7LdZ6BQ/SaCCg7buZM6Wp9EeAW/D/TmS/enffBafiCWBsg
NmhScitEqQ6A3occ2xktMBk77cKFH9XZjbgdyeN2u1IutDWMrc78x9QTP/UEBgYE
eZsk7zzIzuowHH5SIZPBodS7ugkmkvDbbUEm6bbzJSqVtlgvFa6gzcMDEtp/FlHr
UwsI3AGQ+KpNhjqzAVu9N1SXvRh1XMKGL8iO2Xz1MAGkg3TcukevwEr3g4eCdBQt
x7QbXn1DaczRa3wLxH+OO0hQWaj3Kz/QBvhctW6uH+ZlXZtFRdPZCUxX9/3zgy/g
5Oi0uU77BN4ihOu8CQoCvR/bm4aTw5iKpvelQX2f+n+UsRdBIcGFvhd81IBPeQQu
y3ynQ8EiRhTrkOsZDSRIJMP0C4CZoG0fXOZztN7hXKuQnvniwFwPt4WG2DbLo2/C
1kEkE6KDjwWejf1CH/6ET6iB4LCmriF3f4AOTi/krp7k/q9saStFgXakFjkOgqKO
eKnw+hJIMnMCbfACY265VfQ27090I9ksHL2Frk7J0Gs1As+5OCX2+ezdvx8R9GG+
L87ecsml3KTAAXE5NEJeAMXVtjg/tRx3B9/taek5xPqAXyHXjpO2G86WT12sqvcd
viEHwPn/UZ1XVTVPt1xIViPZkJ40E/FMau+SMN1w2Sayz/s3IJ9n3NH8fj9zAlgd
FuhrnzrY8y/EkaHagLZIVLMRawIzx1j7qZFgXXOoSlqILPVc78lCua7xA1b98h6o
stRMf4p2O5/bF65eaMycSoeLT9hh1kusb22EWk9xudASdvcKSt0zv9mSrIy71dPO
BAH5/HHtAcNORqnkhCuBkQYHYWoNNsoFdvzraQwbTovNeArx9NR+qLkSQ6oydnhH
oFxPWKWfbOP6ZatTO3Pr/qxaM8bRVaddRpGRN7LeJcl4xsQibHQKMXwCnlIKyUg/
Pf4gooourjwyhPrgGbHDUI/PiPajy2/Fi79idVwFaGwUKJZgeYH+PxvJ2HLIvge4
XuH6iF4fZlNz3Hl1mbz38mmjwNVrKjr02EWOt4TkRcM27ei0MufLFeqMHJxnGvDn
RAaCfbs9isbpQHt7EqRGmlYg/v/zzzn0jonFTzpXTefNIARH/vnoY8nLrXD1c5Bh
T5GovZzRhMFKDbR58CFKkdFkBlULMoFo5nOF5D1kq/a5xgTdvUAuDaWfDXPC82qr
ikQQ1IJRgN7duDJ7j6l0FH5dND35SsFzRD6KzmEpIng7tXG0G8mx49CXd1t2u7Z0
/FHNPonaCCFMo2eYiu5bWL00owcZNnKIPSqPZQNGAW3d2LkNPF2M1WtzIuUJjX7A
ixOSiEpDf6ejQ9VdaFHygTE4yas1qA0Iz63OsupymgCyr9eUX/ro398yqNAjeqRu
adO2mX+SNO3ObVPdMZyDyzbUnzZRN8ppKMn5q3z0Qeyns1fPryRcfihCH8Qsr8T6
wrhb+s+fBv8aPd5OPvzJ2tl4+2DpEhFgZ91Muwtx13Mk6/3HEXtyhYNgRb2VzOuM
fdSvh6e1IIzFMxhumf3TtjYPfZVsl9xQg8wX0+NarODH9dqtEHJUFjEA5ZL3IRKF
jJGo+suSXNdHkqeoA885hlxMAXauMf26b1jXiQlFnK9sPtqeEv0PxoEOXFVnIp5Y
/MZzuLZZzIF+ioyWv+klT9ToeysDhLgdx72+g1hv4VYpljhxLT3kIt/Ae5zI5zVC
MajmHQCyYKz1YrhCleXaEsdxw53qLkTRkjZ8c2d1DlAc5sj21eqiH2UJXN+0mdnN
DUV05IuUs2f4+MfHr15ujdEj1Gi0CN+ocsYOVs5xfjEgueUIJ9TMU/u1Sya+mr1T
DIAc5uXePl1tiVacqVdTOGJdWYtvocOE/GH/46kTZRl5NbqOSuGeC+ABv9VIWMXM
5II13doimS21fMVjfaH74PYqZtNEeICHKyDbc6c4ZePLeCl+/URZuR8SyoasLcZO
O9OIMcZTeNpe6vw4yHAUUU39E0dOE00AEj7DNpHB/T1U1gHJDU3uM6quu5Vah8A/
NrhpEAOyfL0piAZobLp7PSZN3St/RCSmO7GFDCW067hIJ3CCGcoEO+LIBrX5SQxh
cEh0OZlNgIgXPtSv3RsBsPA5QGcDjIDNnejfava56lLxUxqWN2tfVeRnsb5/ZO4j
OzX+rLDoFF+/Cy5hKlQ7YqNG9yqnXz9Bs3dgcZqJ+YSL63eYe6FuHQtmrXuwY+t4
IVU54+YZNQ74c3XFxjiGLbj7+8sJHFOblUyIHEXWhiYDy+Dkh7D2awU8gZMKI/HK
5J0o/OqS3eEuQP8IOTCMNbs9Bo7eR5uiWq/hvme3Ew72r8pFzMJxcDQRDeHAqcZD
Z6Qfho8OPIT4wkpvptZv16RUnd4CF5zZ8Eq/InEK/WNOY8oaTS059MdNAflrM88M
I7Q5lrz+7nxrdJOjj/Odvx2HfsmokLefNSSxepTRptWAWO+iJzn+r7GM2dTSz31z
13tD3Y1W0sYESJ0hxmU8T9yU6LYCWclGBkg8iGer14Y9jlxNWBp87HERReIn5AtG
4/NSVYwTJIAZKQp/JiSwR/LfkR5MI4KrhnF8CYUziLZgWhKtq5lHfVzvow+useD6
f7j8GyJuJ+m0i4r/JMkW6SuDs+FxwMW6alUkkA8GISmRIJhqYRI86GPRJ6LIzuVo
QTOUxJEYlhD681fAwx9x1b/S4BVKR2edmUj6QwaQsA7lMv27pjuLTmoNP0wqncPD
zCAPhUQG4KnoORloWgmAiyk2hgFsQWyJIt+Ly6wNAA7Dsq7P6GJ/WHCIjcIN7yiC
sYULNtPE1ighBZ1mtHf9fevwhbOYyScXiyD+1jiEHRUJuNgkMbaQAq/E5n14FUrw
YQetdyS5FieJDBXZ+vPPKjyMcV7G5WHyS0yiren/5gyHeyImQMMy6W/zq+1amGqW
WAeI5IiI4Ntt+CgvKqsHAIKNkN1Qg8ClcCsa0OuMH+Lek8KAbcmGRLjuvqFVXeAy
fbsQzQb3kASqh57gWTV8qEXlmnS3P+lGSmxOC5a6kjuKZtLurSNp7ttDu6f3l3Nd
WRQ9Am7rkcKCh6eX1HwAc2pW4z8jUPqDujk8SAXkg1QCO+HHMWdD9BgL8yDSU6nQ
RIu5jsJcYV/HgTcBY0IaHNGNSV5lRkLrjAvLxNr/Afk/sJG1SqMyaMbuhjAVrt24
Vzqn8zptyqXBMpwRW2D5f1FcPVdde+F0yLG3ZlwsCMwb3wBcWEqZ/R8qYEfaim7g
R6aiKwyTi6r01KwwL90CRc64HYSUTvxrmGjvyTp+ipATFQ/AbVtHH+CEKc06Wpbo
H2iF33Dz+Z5n3dL8/sazQJOB/o2uxinbWp5dHDavSg/xpMlP1BbZKKQPAnCVKOAP
7+Wdz+1MhsTuA6zjwiL3L8XCtVRtiB4nkQsXdI7Bm4lGhqkpJOeKXT7KCEvkQ8gv
gt9su5/UGCfPFkJzJiyYk21S2xt8F0Z705v0+gDSvmjDaUSRaDo0Rk7t5BGr1TLM
U5dUC/hrnEEYbeLzFGrJa36hSD3vPWNz90Pp1dTq/aaB7fBQUrMPRXA1I3tdSEMM
ADWub0vQHgIgZz8U8odXNeurkcl0jZN0cr8e1kViyvK6H5DQzQviOJhSShXmuNoA
TUSL9gDxOOZFvOR7j+q8Ez21hpQpWV49Qz1XFRSMqT1Caehfr4C3LXGUITYyV0rt
nes5AahHV/DghoHc8eg+aZDFwGgMPxg3SVc3aVOMiMzl5/16CElQf/4CKxoAGl4Z
9KLhK6xHtBhh+KK0NiM2tlJshbKOCOgTO6rxrJP3VgUUpUmUuxgv91L5+epmgJYE
emZ5Bnbv+VoBFkV/VMIGJlIolWBn6MkxQIb90gNC7i9YGXW4u3av/G1GBLfQ/syn
ahepsm+E2jDHZv4J2BoS4eaQY7TQXK/Hktg5uwKE4CzXJ6Gn8w9c8mk1AwGW193P
+vMXRE11As0CPpygZXZXynvz1eAYcRJKKOUsfirDvIXOckSok3Pqy1HLszyqdH/w
oSKlQwjGfxuX+4ktpF9SCsnPvVP7T+duQg+OsO0TsVYRTgPGsiW6HQ+k44h3o+4q
gfrpgYOj4+cInMGD1UC5EtZ/0Tiejh/mjl3c2R4xrj7TegwF2gj1PG+gb7Lm5e9X
saFsbVj+vvdJEkCY+7n7JaWzHYSpmVytBXprt6g0G7MBEi73Xiiiui79XiorCAi2
cgJvSS87BvEZftjUFRpwd7So95YmSGUA3tRkeTC4vb5lYEbRLMCl4xuWsL87Vonz
IbopLLqk+cGUm6iYBbD3UBOvk4Df3DBAuBeBFQRHbXxVu4O74qV1/FHNeI4yxxMZ
km/iXR7R2hj+NBe6SmOanFOc72QoKeGooSdpRIt/uhYb34GCDDtVEq3ggEgfLPtx
C9jhRBr+yX76b4TSpZz5mhwXAK7ytn9/O46N+xAB1IWU6v/Ozdb/HWKC5QM+9hpp
kva99+hgz2wVAYu5TKiALGke4JfenaLj5WRyQ3D55bwp5p+a9427QijEnTO/oxP6
oIQCRySRHSUlOGp2TWwKdyelpffUhk7mlPH4++rbec4cjETbeBw9Ubkx1uBUNygw
oZYt8YrV8o4Ciqv0ROdLlJI5UJvrD7eEmy3AWmrxlC5P6wC8qUjJ8yj26aKNj1Xb
2+71A85Vy9WHDFwnSDBk3WbF6KLWDxsvp2M1lMEYKl19gIKt0hVKzhOxtG4Q8pnQ
OjyUotXZ14MREJB1/MPZPaJcsfIYkhQR4WTr7eHs4NoMTzvUXROf3NtAogPoSjXD
vRzZyniahCwqeaVn9ZIPVi4QIPtvrDVttkXl6kP8OhjroEG9tPUVd9mMAtN1kzEd
MS7zL3fsDA9gYoCPrq3lrCwpRVjmdYCY8FAIb6zxBVI4dXHiRPINclrIWHYN9WzY
WH2lMnT51/Rm1G37yTG7tsA+bdZko8HYyqMd2KeM/Ag7+AZ23GmvcpyJL7PKhFDw
jir5RAksYJ/HpK6y/dPi43uYmFbZkRVSLHVlAtGXknRvF+aOF1OXa19W5gvm4xzF
Vsw5tOyEmJXvh+60b7hlKRhc4GEMV1qViHQp+D2BohX1eeFdgrdm8JCw2I/ZPSl1
YLUQHSeovMV+63xMVlekeVtZEp90G5w5RW46F8LwDdgnhJVcyKmd98fCKJ/4EmeN
DzOYYxVuxsdFH+8fDpxQ5p/SnRNSjkw64UmGBFOBF4y0gp8OE4A2EawYQeQIcObt
Z7vIBZfesSkBnvilzPpeUxN3g5D4HkGY9AeY8eud7mjTvSyRcY3rMf4ZU2BECvhE
JRR+X5/zHJomsMa4tcJf68idKIhdYdJvRWGoBicJU4RmSrGXMZHjozwIklpFRCkA
80ZGLVImLg2c+aSnamyJ+AExejMCPlZAhO7F5Od1lF110+eXfm/uR0wk3QWitD9B
cf6vXhHn6lb36AWSyClMl9HOvwKN+Fc4+Gcm5vWLKvsrBdEX63qw6bsfr1+Rh4PN
U971nQgkXrT0jwMNfsbI9n0CRgGGO2rE8OblF2zaaTX05HssBo4IQzsvBvkzK2tB
hk/EJe+FxgCaN9TfAh72q7/0soluEKXw7hSOfetCsy7a5tl6+axnG5SwEbvnRp70
722b6MuDrM4FH38DL6mgohh3e4aVaEYC2fltTgv3xdckJBQz1sm+OynlThWaWaUk
8Dvo42nbxgkNgubPUiwyKL7xBIAhbm58Yrxq71xjXqxIQNHlZ61gTl4qKpIk6dfX
KkzVZn4+A6inKWLlUmvE9KjtrfUSQIHaR2qLN6ue/QB9towGKiIoY+Y/Ztx0Jlmr
TYiEfP4fqbx25lSNmQRcWT81CRBL1N9xQFzXRhlYJJoTJhWJEHUUMgjHXXbIb0Xn
7E10H4QxnGik1YVqRQma4sEMIGUiqgTyUOZ0zyz9pY+6I9KrpHGOAl/Bz/b/U0+3
bRGEO+wRNiAAcgNOt6qd9xpC1JdhNZfhyRGP3J2sR5CV1r9/SvKL087pSSSH891F
doI01eMAVsrd2Y9ezDDoKPjinEisZ/rWikMoZSqV5GaH4X4wWwPpIjM8sLligoj6
/RGca+6cPhIqsiiiRFebc2gfDScErbgvSGPjJ85PSkH9e4lPTDAvpi56ohGPul0D
KQ+bDu6LJsWN4NA51JKyDMTalZfM+GZy3OIeJgjMv23r09wQxwiqlZFjZ5ff26xs
DuEbKqXPYIsGeaTtlmLHuPeHKpvVSA2iU8tQ5nSZ8FesQh+xMj8j3Eyzf9gyu4I4
pGURHb48SC+wueTCjSMEGGF4vHKXEVkrNgPDRcNNuH3MuUSR9Y8fDgioiE8h0JSE
45+PqmOqfvJhJPbvGb//tXNIFFdQXpFNuXW3Ze0H2YIdTruD3jt9gz84MGvNPP7m
bH4tSL6TfuLB+9i/+tPjrgEA1jNd7iHv4h+TKMV/pzw5ZdZddJd3UO9MO4ybzAU4
j2WOKmBIgFWzNbqukfEyi7LOMv0ZKuW+rs6/VNISk5XTcF9Q0toEwU+6pF5QhKSW
2c79ETcE0+iwh4fEDO1Ik0qcMiO8fYIHUeUe2tYj+H0pAZORqp5OIaFi0I3Udo/B
3SD484kbnerNpNOcTo2AUK8PphhPSDQ3Yn3HdsaqzN06LpA3WUGwMeETePG7Oxiz
Gygjy+3Bhm0wvJJhGGgfDx0Qxt29U7r5KgK81f5En91GsyH9hG2EMELBDeq4sdz0
kIHFZbUor6jkCZBw4zPC7bqgmC9Gpm/2MPDsRTUg84rSk9h9OuMt3K2dE5Jw0zq4
uR4qUbKZkMClP/QqBmLQkdjuxILG9OMWxf0+/ZxxqSceDlM4MqmLv+sQ5caRoKVG
9o2Mt7NnWB84zoxfYvWtgCveGx5I9DycvJz0zsB0lsj0/nQGAYvnVsC/jqpSF17q
7pTLXnAP/BpOuI9fQ5PGXMn+WdDntbxzGSoBAJY7vJbDXHgKLkB2O9jdvoxNKtnK
jTC3mFAtZbW2wgicrFw/j/UyLAWuivwWy5mLIlVaczKop1GRYXc94MMxhpfGO8vI
7Ido72Yc9ABM66WkguSQumdUFcMF8BVyfjmtwPwGYk+IG0Y5soZ8CvXB1Ibip8Rc
FomQaGzCz4l55FYjXpt1sgRZ8wYL+jbLYv4bkgDk3Xp0tV5YK+Q6fZOm0nukFt1S
DPkahWDQ5KEXjzi8Snjsc1/hh75avQq2JLQ45jrX7W47VjDKih5+J7OOGqJuKsju
Vw1U7GtQPlLi7z5910i6KBrmk8cNjkwP9IkR8lNAozrVHzhyNxQhUsNs7+z/XD/h
sHmPPGkgtLOtP6GsOChrbZ1Afjjf6rNkATXe6yfuj6Vx3AH1R1b7Atvn+PE6ZUm8
rIZbcCsMzosWNx3X0IM6ieo92tekRRyj381eOJp0LOX4P+nc2rAqsJbhm4QZ2ZNO
fTYqSoaPqzbB5yvMlDml2gvI+jQzMccwsRsPEmdlBKht7yybpvlqXOYrTWR8Yi2Y
BWxHeh5uICsp187LxqkHoslOTjoNbF3lGPpkoo66yAXL7FNxA+a2zI9GuJLXy6l2
3THJv6vyo/2Z3zfVkEtvaZvzzqLYnAnaVIl66sNiZK/iGVTPvI7XX7K8G40zhdmc
oiMPh9DwvFnTFsruDZ2apV563iKBJGr3lEC8h/ZyqSlQ8JRH/RN3Lb1CxuBMZqDI
JA6f+9X1i303c3dsWZCp/+LGYYVBMcFd56VEvSM8ejtW6C+RD+6Ro31TJLtSI/Km
6aQOm9CqumLAL81uaKm94WXf9ngK0Xr9fHiACM3bBE3kSdqDrEYcRtBzIIelP45u
DwU7rC6TSfdfI3dOAfvokrzJ3rq0I/OWjc8Qm5gT+UypGeEZNzML8Me1cQ/1zkOD
mh2Xpunow9PmJNG+iqdPnPo4G8772kofllYiobOlhxyyaQCOJl3eCSsGqmPTpyOI
Rz0T2OlPAC1md0WZXWwNykIDfwd+X+na2yvFSYaV/Aciz3WRuodDJMv0ZWACA7hj
DU6DdGTZ8Y7oIRoHKFw39UN7ZJFRqIwPZxGBmw8uEZvsvyi3sBkOfx8tTKNhEiOs
u2xosj3HnJXGdhdJWVk713StnNkXeJkZUhGAadBc9CqFGWOq0SMaWnpLG3lF3H3t
fzZ+PLZrJprUETt2clAhzYHyzLFPzjkSG7Nk/2/F3+2JFqSJ28TTCE67Pisziq7W
LNc2hkvYej5I3gtCx8QCqlaFwh7fskRoiErfq1uS4UWGglCCdR9VuxoctGWVyVx+
1A9H3Ge3ymFK+Gzsavk68Fzo7lOeCySLrOxqC7miyEP3a7VCnqyWe3DjrB4FFrrR
WuAUQLpgMbioTlGpADXgi0As5tJQ7tpufNBF4ujXKsVv3BZzFhmObQy8xxIt5Ch2
QzHspOWHUbqo44ahZuanCqqv+7wa9/j89deKa23j24Grxj1/M8gyIKD6K9F1Am9N
oxIk43PcAh3c6YR3lugybl/oUJQQ4JgwF85bJUMsKT38C1cWN9hxksz6euTJjrxI
itu2I/tjYd+XmoxJ9GYBs3a45O0PqASOzWQFFBq3zgecMnjIcJ3Z/08G1ZGVzwP/
R0lNC4GrRuHuluOdiG4j9fvRTXFoA6A1efpJwOm2woiAGTqmmneKLSXACP50PhO9
E0aO6JprvXkwGayeWsG6Juqyf5oh92sS+ucvMYm3bHeCE6pVgTvnATa2a97MPZ3u
nHULWIAMFfbF6Miic7RZD/ftApqiPTStFePgSGnSNF21mwyTylRTc1mKIutMS8Mp
ICZbbpfuN5LaKh4QRm8rZTaPJUmRFwaZ5FQO/JcTn09hKjEE7806J8ofe2ZaBjEi
OJcgtnGwmWJyu0r4RUk9byST+GD4tv59JWCHGDvqkOLXdo4Y8GPOD6FBYfGqqCkN
13IE3mQeG8b/I4VvhgrwCUXK8sNKys4yiaejCO6bHu3dMhH8ZcnyKObAFgybUU7I
V28Ao9WfFvkzSg7l//97cp42g+cv4a6izGQjy5c7JE3D2lWqi0E0YrWXM+W0OvBu
GvakgPEMPluCmRfT7wrsWvVJSFdYdTGWbLWFRJVXik+YTjyuVVdXalmpTwLdUQz6
r9MM0Mv8AP/jhHcaZ1lCDq2sgrkhA/ruDzbUJ0JrroiwQXItx3e9thqI+yh+pBlW
FsXCBsPK3MDoDzZ15IXBEPfm/E6xco6TyQjx1U2VPXnhX39DsoGpjMwevuZLMkY4
ksf1Pv1YSMzgKzmNvaEIqRDc+zguPcrESd7QRzAIvRPR+ZtI+yfsASBYygWU449r
K4uo5+4Kn+b0TIdRn/6eZ0kkET8jgoMt5tavi7NeZ8KRzSgpIxzJzU4iF1Hqwswa
Q4MT6h/IlCwJLfLQ53A1tJCRf4WKWLQ1qhqnAQk1eAxybX0HFNgd7BuxeUBE6+92
uegTA72cAyJonzpOvdGUB9jHMcg2ob25wDI9aB8GS/M1wqn6Y3nyS9NbXAspRkiW
NqWAEuwIMRjOQBq/AmpVT7C7X9tS3EfBDLFNQSCSr8omGVI/187OWnKkQuy8BfOV
00vI5c4MJ+fRAc/E12LBeTZFE+tX/ZYbPrc7BIrT8X2rX5Sx1Ej/Pkg+FeL/yHW/
UfDQWihzZuXutWojqdftOQxmEVrZh6DOM7qDcbvomvQQ9P6HLmBJ70Tlt8Pp3U5z
PKAIsI49VpBOLzMxzHhjBhH9ztrPv9fUisNl5Q1dEy4V+VpzRltykCOrHgiiiQ9g
eOigq2pU6XSQRpmp9mcIsiSvVyRpsxYZbXNOm0f1gfETIpUpcDaWQrPefbA2ThcS
VH6Tov9cyAJnpVdgcGe2xklq7YmA8Eem2Rtnk0f92WZ6NrmGt5H9wdyVdurD5vs4
T6NZRDoiCGDJHvijbJChDA87RTd42bCLhYQ1oL1c5rx2vqFHcqKGMa6n6zWdz7j2
4DPFVJvG+Uhn0sooICzP4YxCV1AKT47bKDqY8s8tx00Q0kM1NRjt6Gb2qX0LCR1u
OScPMmO0aqOauOHAXwOT+fwjNCVuIwzMB+fzP8bPwHhIKnd8LNhiqMYLF8UZkEgh
pikz4aS1nybUgOFAAFMoPT9jBXtdCQYjMrYdKD3MxH1DYCPETRHDwXZ1YBHBGfr7
bNfr/pYw8DSvLO6kFY2EETgslXr0nfQaXAHeiOAhf5k0RlXGT+VMxprOhZUrRRqF
cWmyEEDfB2gqgla4TTLxgzvApZMB1aGdYhpuxtqjC99u3+fA/P9xBoylKReA/57j
RfqfypFPgHzvUwgx3ES8L1CyuzpcMsLv9qxkevAmrTGAcq9/O5p6pZmDlKgDdovo
R5H433PUX/TxJRodJQwmo/nepSqKUbFebMIzLDN7Gjq7IDA6GULQiOcqNyzuVJ1d
x1WdQqxIxzFEJdtm5kM9nETml8jm/bpNjt+YelIgy+sJA18PXHU9OsOPq/lQrSZO
cDI0ct4aCwIMCBiRzZFx3Ck1hZDSCwHBJKEQNLIdgavX6esi7/SuyjE6oSpK2mt6
XfziKFWoLH7x1Q7Rbj0AQN3dhDmlC2wOtLWmOf/RorXlRImhu4Uy2AeJCYFpMd7t
jOysSiwB5g0v5jqFd3O3/7osnQTV9vpz/h3XdcVUXyKxPLiVVC6JpZl6HJsqPDBH
TXT6STM28lVLxNZajj89uReAzbxvWdSSTjf2sJoJRzqpTcMWB5UDF0S4K+B1AIo5
u2zCsbjS95gmyjh0ZvS/YUZujknxIm5gpXRsPWT952avQEYMZV2TLVkmHluNqnQd
XdsdhY8prZWu5W0J1QCgyE5EzXQ0yXZcfgAOE1gB/ISI8NaLCZrimmW4BeMbpb0I
5ceCLMuxYIwwjkAHFrYrHV+Q1omaYlnpHurwOPa3Xqvcxytu8LsP3YfcB6K1MyVX
5D5oZMXKREH2ezISJPiaHkF4TB6QsAHHzA4w+3XlmXppNy/NyrkKjy7P9yyReC0d
k3L6lOm5dR+XztHTQjLo8HaEdQGo3gHlegMw/za0V5A3ld/qnMcJn0kCoDHHmKjo
iGSXGoWFk6tz86cQsvbASgKAfzYZROOXICO5F2N+MVD67w1gGgkym9VXlDZ7NNE7
IlSPOH0cJc3FxJdMq1GIPYayaT4m0nanaXwTg/0FK626z4C26iQtNvN+2nQLC6Ok
+4ewm9kI2BAW3xkxrW/ZputIBYjMCG03qM4LIh4egwvA9Qq4bB07KFzCHVrNRarb
G57WuJinzxaNdlphB5fUKklD5SOonanrVOX0mWtf/KmyyMiWY4EYB4KghQ3b24QO
lpNRflJzIqbxBvWcw3ls8AzGjnB5wa2neG+Usz17o9ZALZ5F/8z+1VRuPCXrEmI0
q5AgJwqeJMEl4JLTV6koxve7HnhSb5YPfR6TC7KFWo3AvUR+aEn0KYRr9h5TkXF8
Qk7xT/OiTAs+eWW4eVlSuc2zKUjXasRdQv51LWi+L+2ShM/W5jSI82cGPt+HdxBw
t7iCv5ZvyJxH5rRXdvMq7GhN/yXostuZYnnaHreejlXXkSsPD7ymIoIpk7qIShw8
cMnRZ15/H7foKFNIi5CO0sb6zzWXzZVtQjn+nWAfnmWlMabwDwzMmD/7tsn6OfMM
G1QC8A7qUkHxq6dzfSmeRqjr99nN33LYulQeaYyOlbeRWZaqIfm9WP9AyVPIVtHg
Qi7Xbr36C12HTPKYMn7etI+qnbvC0PyvrksFjoUDen2jrGEyw+tFUNm6stFrvGrq
jQWA2+tcMI6lfF6F8X+zQj2IxGzhC/tyPpIbBCDCGaKdSeLekgQ5NZUaav0AqfxG
HpC5EIQlg/Cprt3XpeziTKkPuXokx2C84yIW36iKkoa62lEUgDsrrEkba6IN8leD
m5dbDKUV+oqAOn9L2/BrRiIFz5l4S631Ez2/h775GC26WPkNl3MUZ/TDTOmlIVhe
DL5vrPMccNcLkBIua9ogt1Fr+TItGE2XfIXrCuamm/7Gcxi7l4FAh72L2SFgzsDn
VahXmiHrtKt3xaomwxnbXcMzPKjtt5xNaQiOoadZzRsd8ph1BtbOPHaDyUq60BSM
PuX9inKIPlZ03F2O2plIHTSmHed3hFZTu/FPPrdqny4ImiLI3LKKdQdvaFcNgUgf
vRXm2MR7uyzdXftU2beIFla7RXdl/5H324NCIChKM3a6JO1vzf/TKd1NaWCn2gZO
6Afgv5cdRqTjTFIZdCafVv2IsbSu/xmks1gwuPIpPNiaCtJAc/eyUWeYQzSLKuyc
J59+ZWYTUDw08nNpc144JPrJW2T9AyAaIwqWdo13V9b/srQ84NDZb2EP1zdzoy5W
iit4iGHJKDlv6J+iXyIqzkXF8G4TziLeMFFZXrulq7fdTLahZMXhd6zHIGkHKdI8
sTzki8xZV3dQXoJkYInGJlShLRbcSzmkMS/3TrZebx8+Ytfh6K2mpRWoauPI9dkx
9feI0uOHBFYotfNom5ebwnVTkkVVO6/YM93MXA6xPmscafoQ0wUMncLhDkyVsCOU
sUU+tYn03AE0+Jy0DJM4kMmBDkeIfJ6lxHNXIVla/5b3fcM7NO5C7pnF/mfL9sfp
Odk6wHpBISaDjK3qAmnRkSCPl5mj0caorHfW9duTNebhFKgC7sjFnCPIvLCxseul
N/rskKMYAh+feybCBIFlEDYyDhZLi2RlEJG7kLqy2c9J/rJ2hmtZOerUZZRWp3oU
dk49W09+hzDF54d4rYfc++onRU2ah9Fu6IViEridk2bLdFVeOk8V7nWI/B1HY3zm
KF0rUn6BWGuCAWmtgC0SOsFkv1HnPSTqUZ8IfNPu1i3OYtQ1pNZFGNbqK/ln8AIv
wSyPe9Q0NseZ9aLj3XrvxeBtuN0iP74Qii0Hbh6ls9iNPla2DfZyO4sv/JPRpZ+e
5pIvWV28oKuTwXnyCNEjEEslKBM0SyRAYc/07wayIMvCDjlaZSXBP9FvT7joRun9
vpVaVaN4io5QlXg3/MhWJijZF29CxODn3bUmfLW+j/ZH4grtqWFMPidxhZPSvmS0
bJIANuzna2CP5OoSFTsn9oN0flKhiy5nQ1rQIRF4JDtEwnLGdTai4pNtjudzZu0R
RdOxNutc4U1i9BQcJIVxSC+pfta4TPP20b20Tjj88TgJ4PEeFgJ9OTy3KZga9zHV
2IV0C8mIe6dwCdrk3v2QLNA1IKFJRTht9tKJu34owc/RPQ3qiAy6OEsKm/NTy3cN
6mOxzDE7DcsMUYiCvAU735ACoPadVhQkVMe86O8tLYBctV8dYuDSwkFfHAvTkasF
am9xMh4AadOlm0fhP7c8XHh5zs1AYHEn8FEq4ssrzBqvkmr7giWAhWXej+67zrvY
i5C6/LZ6kD4n1K+IqlOPIIp/7SFoqy3rbPEuuYYw5HZCcM0Cli8lgkpXJgyo2DC1
t4lw4Dpez+56W+lpRgcJddm1UO0VaSR6e24m6UCIvCKXTXu0IZudESQ1nWJEGAOB
TmFktzMo3JlaeewcXfKZ0rr5dxfkybGwmVlkf4Z4nhkGI2c09b3do8idtmdzmC2x
dS2vbZULDF+NwO+FHmmh0QMUk28RmblRq6DLnE0FEUqq4x87qzd39pguOZk0e6gB
GFb7CY4km+uDANeYD9xeUSMDGRGlU+ruhMlQjfM4z/39FtKO2hqyqNBNdob9TJ2R
hQGpjGyWSkp+e2fFBdkkug6fVLLESCSTuSlCqjK/dwiRc6l/aHUlemCvqhfX4CwF
lCJH+QBnTTYlEeblZoU7aMiRKl+d2+r8F2JXwyJ6mP2sIFXkzru77WESShQ0SI5p
3LQ1f7vZRj0LGiWOOoZ1dA2Y1ndLrQGmZlretxd+BIPLutXmVgqUXAflTkYKniSy
DBy1OLt3nqM2M+QUPGF+Y98BM2tVxl7sDVDMo255rdR/0vT/dlDoEgbX4MIE1TGu
EJjvkDHHsHCqEQP88NTSZ1JzR+9vVRowc3tL4Va/t/NDsFwHC9qeV5k2f9AK7rrp
oOWVGayR8VmHUQLVHbwRVm1xzQCGLUTxEsfXUMe3R0CBo8No5qlCi6x+VWlFneaC
JfG6b+RynnBN9CZ0gMYLGuSleJxGf2DrUCsS9//p3dQlifRMnUq0xECQjaEeHQSz
MttCep9ZZklEvC4nOkiuTyyWDsFLHNsfbgV1+5pmWIB/cfQwC93+a8vD4Xs0HFtA
BRO7S2fOG+rr32LeBjVuLsqgiBR+UxTYtNhf5oNNTTIjM1mXhbiWAglTL5LCUSoP
MlbYipm1jT8ftdh0fGtPOdYIMkbJZMO8dL7UOyVEtKRVNWWuisW8OCgyEbLfOfP6
7wFKo57H7bYbjeD+GErnQUDQ5rMPyV3GX94YH2B6oM8GAWJvG58rUWjgNLR44dad
vlYRj1TjENM1hhN9ZZwl/dVe8SGL+fV8dsFo6PRLF1YZeoaVsqx9EvwcSUFyQ7CT
Hy3Q3mkhgYMZ81r6HoAal5XjPW4qzfmLaR4+RaNvFZe1rreRgmKOAg8ahuKeVKWU
NSkSWJn7wWCH3HMS5KdB41dfpsnLE3KISmNDHkz1fpQq2NnAPaSmrXMuB6apUwHK
1Ty9rL34gvwWHU7tsY9NopbEJuUCjAfAMURRQi0wPzoU3Qrp8a0nSkZSw+QVBM5L
RPMqF9ESM0mrm/Tot5un0wkczv/mPmueLgw8je0wnCWiJ7anSIfYNesapGzPa384
Oyf/AAE3/XEyLmZeB4uIn6tLk/iyEYjiVWD3gjOFF0lRYJRq7XjyUwXYuX8WIf6D
qvRrim7biC7mrUUO4fJ2t19KUlHc5xJHefSuLD2ZCg7AuI3yb2rMDGhNHKWXu8Gk
VbbAYYl/d6nlEdnyFUtqFCzxsYlIhy+L4a8ZitYGJ7FJiUXVsuGjDMVKS5O5TQyL
PHNoYAdv/JqWwFSaaazOVEJMYNrBKs4ZSiuGObkKuwtv31w894okZmuu1dZrPpJB
qLnoxt6GzUsB2U/FFSLmr8Cht2FzYmxWJ7ffLF/wvU7Yq7rO3bq6/AU2nrLgeslu
Q4ujYlx2fXc/A6o1I7YvxwRcjGjWSsAmck536xagznsQKy/WoMaAtnQ4oHn0hqSy
akDLiVgzsF0T9yS5KUehgEPAyeoMXXvJ21ubGtwSI7c0g7vDaMO2p2mW7YTtReAQ
DI9xcrQRkl8qWUFOc95N21zReoUpoprGKUiGdZSpy6m17uMo4FbzkG/1cCmbBjRY
EmNylof/6BdwGexcyX3NCRn3afjxEX07RdK9bW0K+82D7rAkyRES3+9UaQ156/xr
Q51af6IJWtTvdMsnymkHv4chkXNVejIft8yliH1UfyTawAjrfWjR/+S4WYl2xO0N
Z1MDOeEals4cXWX1xlnq7JkO4KaolOxHCk5eNDCRGiZ2+b2pBEarCeqbnKI5p/10
lcxuQJOssw5X0n+4vZt7xypF1EX0LRSvkiWOG+vwRs7F1b7ZaQHmUoINQQXLroO9
ve8CkcKFfNuwm6qVf1XnFyUC0xUZFqAVhqxnGpSaTZnT2/m0jGx5AoC7zT3GMFg4
jwWCBxQkdqGu4po7viZ6khF6S56XG0/kwQI6Zjjpy1PkAv9BKunGiN/1BhGmo9ZM
UmJQRW+a3dGbAN8IPblS5f9geKl+jDLQLDE7EeD/3RqJfCa2QJY4gqAFQWdX8JsT
vy58RKVKE2FLD4svOIMUDmUDhz08M/dqnJnhJMU8r2Z9ONnaF7mNSDBaN31bUWZL
iBTeU5+0W1zLoSQFPgK5iKhV2UxZKi3yQqaDcp62nPBXwAcvcah6rcp6uetU9c8I
b6J6YQ8cZqB25ILNwsvAGxEIPeAPLM2b5MO56/EUlewsHYgSLVkV27Zw+EBMIzDc
DpNhrZRrCT4GGFOIpmusnzznmwuIM/9fhfpJMWjj7ZTkYDIXL6Ya2K7Ol5x7LByG
mo2KYyhL6Jqcwvd7MypVTdyLriVT+cDKbz2sK/jAbQuJ0iAOTGNPzdDnq/QW9Bfj
X48qdw7me1EV9+ZDCvE/DJcI5rVYN3IAN/UKkYFSUIAUi5jT3hd1NVbZpRSDphO2
43UmgYtsDU+GA+h3y7EEtefNFZj2YEN+SOPQ3LOqFzaZPGylS7HzwO8byDEMcWI8
1SZqnt8ddxU4BvvsWSAaDXorSmOr1Cfo8sr/lV90xA355163PXZUvtNlAsfGQXtj
xgx9WdX+nM8zaHVwpBqmjDf6XesAQMtNPC8UIiFpwJypAG8/RnNur7wruNqlKR0x
fr98XMSOmBKqkSLQgpCO0BJNAQpiEiDf7SgGVIcYaGkU9riDPh3de8K5TcaJQTal
WCR7IRLPqiJp/RxClY0M+zVD0WWDCy2ZZpRHT5xqPyCnbcCNvVVnOBGPqbHArZgM
fXe/Cx48qUD2G7RVo1b799ZMyhmqXlCsQToJYYqw0Bsrq0NCZ4+JbJI7FFEK6IBb
hswn4TVTRdNySaWK3bAKOd2Q4NUv+G5ya3ebYM2r55HH43gJ+nlVCtrUETl1UKMV
XnTCLrJuhjBdC7QRyN3OzH+wv8fAkvyXNx4gIcxE7ZpD727Ssfr9TQs9TLTFlWI+
Wgn3/uow7Z5qO9gj4Vp9IyzlfrSg57jIIgbNYJOE0uFpd8+wtzOTZbjbY+s7mIt0
Me26FvUqJSckF3Ymx1Iz+rPrbL8sYZWYZKVsYeZkl1zURoG6BwAPI4n0boMBZDu2
aI6PQEEGW8akgyMY6ssiWXJCv/YLW5KO3CWP0fY1/LGkMF8gkGd2JLeLzKfWF8OU
yWswHwNln7wUbM3WdQ05nNbGWE1x3It33kzf4+KeGKqEWovuA4TEa+ovYXLKXSyS
XGXUQ+PpEZ+6Gh0DYnv+Dk7DSfG4pi/a6NtlEF9Czgqje0C+cq+FSIPNmYwRlHEy
e8waVHJex1JQ6MW1+L9DRaPN8stxYTeFYa+zVbCSz8G0n6bZNWowOkQbPavZXdzL
x8XJE0Boo6cMC+/LLE1Oiv6uxkJkJKg+OrsCeOe8qDy8ZRP2RsyM33jrbNLiumXS
abYZSJ5ic8NWheDAaxrgVsGQeYfqm7zx5U4AiKkFYGKomsK+hqZH1VR8KqKCm759
RifM+Zn9SM5XogtK4oQzeXcC1Vd3vPpbhgcMBKfDz1T8OUCV35Cv5Onlrf7AxFzI
jIDxbB4026Eqg+2Wb2onPVAt9b9zI6tJ3tuPcFS7BJBu3mOwR0w6GucCGKczQRDy
DvbnmUumnLDIvnG13XXPRIA8HEeMn86zD5HMINx3iT47LRpu1jx4ETaIgERI6RBr
poLDgG/RRujJzQ7ASe5wRI6kKsHi/Yc5ESp+eZd4QVF8qq1sutl3VymI99dp/Ujr
hU6zx0hM3JPURHEIwd8bp9SlthjDsbn7cjx2bYQDahqQZH0dQ9aFN0AV1ZBW9aOb
m8Qc+ijFHXjAvfNarJo/L3HyVz27sVWynKKu9Y+00HJ612AzFQdnQvD/6y2NBmSb
B7s4NyMIqQkp43G78jRQr2Y/n6LNSDKkh1fsi0UAcdlXJPLNVfEOpZhJPiGYr13t
KaYWNljN+MVP5evQbc6RVyHCPC0BREA3fuH0sr7zuJ3il+rSpmLTQP0jN3eCmbAD
lQZ561iaK+mNd8UUbbbkqDWVrnxe9qDghH+W7+D2lHIZO6Zm+9NPzbNIqoDNV3Qg
q/sVd/HN+riV403BmcG+jKduSzKQZQqRMw1BRnx7kzKGf15pT3zAgMUXdrbOpXTO
8qBoWWewjGolEMPprTLHFMmSCVwgY04n0IBTT9xqNJLQ+VJbs5BXpRGOJCqzllda
xZwHFmTMwcZS4RAEbB9bIvZEWtskYFWCbfNQcuLdULmS+HqpBvtzeIZyLWFQ18tW
4WVQvpO0qjKmi9zgGr/rKdKEW5kBb/OeQjYdCiMwAy9eCkthA9SAMPYoF1vOXO8V
0fXxZO1hGXKvUuZDP5JfkIzSt17kcOEYRfPHsXvz2+LDwnYmNgz95kOCJshZsAv/
hpsNvqBg4HJsT33Z+WHE3P5CLozF9ofzPC64nNfCzsQq9B6D3K+qhMQRZL03i9n8
AoXYV5nhl3Lphc7k2N+QcbeANu0OlsLTFTVyLW8Bo6O57L2U4kA+MFIEY7SBGC+v
kI2kqobeSISSZnUoqX1nuXL1ZUWYNLIBtnwDdzjiO3kBMwbBFQ94Kbnt0hAINvr0
0zoCLvO4UEpBGqH1hSLma8zZzuIU0ifJjsDijzhbgqet5aE/c8+dboZzXaMgRYt6
joCcBp1pVpfKSm4hbi0A6LlvuVJTujWATyho+xuk4EjLc9W01zEirJX1IE3ir2pq
8kaG7R4jPMkYo/IOBN1Tod3WC8L0lUb0dQxGBiuzbBtofghIC3B1Qav8BPboeVIQ
55mjM+kXpNE5G1Rmn+Ekfa3NDYsY3iDgeis9QJW+v/nYNBNRiAXafQFGZkV0Mnhr
hRfWOt2LYXtzLtC6FmnOAQ1NIRNn7c75sOj6THxEcqXNe6qmLSGtl8J+oRl78leZ
V19SCCdnrlKV5Ww0GoXmn4105ufG2jX01sU56FJba5YJQqMWspb2bjsdFRLjMcAl
0mzzcyrvhGiMkEe54D7QZxsjCqJofeZFSvbjzf62gMYrpS+/qkAg8h5i8qt9/roW
pGBr1ottVIsaIkNIXccEMVn/J/2Z7VgFgUtnQLWp0E+UBOaZgUt4NgfvWnYQISYr
9g/bIOmBOlxWDaEf75+WrbUufwCPfBDePYte2OYFSidGKPX5vVoPvPGRpl3Ym/jM
i7/KpWFg0/3Nce65IVmb/Eb5bXMaRbYwbSbZ69Z55ibW4ImPTLWTBqNtC2VoYPuU
siOXtbQcKmNC5N3JNJNcY//JntkaXKHfzAhoqWxgdP+5cr43umqcjvQlZIRRLV8T
O8GBpWE0yXs5Hgh/DcEhAsekACX2fgBdjPlAbSh7a4zxsXgYloQyNnCtkjxb/g3t
Bs00MLHNT2FCk4dePC5OQ6M9caRosOwM6jibY8GBd6ehD8mTgosq171d+QFZ/Gie
lrpQXRxqBeiNQ34eaI1QH48q3OJs1gw4PiehTx/lRn64BxG5RrmU7FhxBbVo3/bG
4V1b+RBitFaUWJ5+IU38G0dX/4OOUQMP+7ozNscBb9J07nunG1ilB1bhjo2RrO+q
qbKiFBpqnziC73pm/QXzZRqClMaYfbW3JHJq/oz+gpHyqOxeFTlB4FD8JYkL7vNl
IGCCjt2b2v+De7ilF9lGlonbII1lSvMdFZ2PbxLfOo1DGe36lNouEzZeX9d3Uj8W
yekBNlLCh1GPYTgQdhdAsKGUnvq+gCctU1VYG0rk6q7tbPTeT5LRGrtcntDXheFx
otluWvMATHv3jFof997v3OaJaZVAv/OeONQfrCjINLf0vwBmieFdkOFmPuQh2Pzr
GfLljue3hZPh0XjBRvG7jrF8bsoT09PrAkWexVcZpgca32gNnl+ypEcSW7eX/9kD
s+VlzferxpfOTTkE6fY4I1h/Q084asruLXkSB1gMNh/1nYM+XDvJh+++8DgdVCDl
8XJ3Kgbzgsmc0NbZrufevAKegDJ1uepH1z5gyaPNsEK+ZLZXY/21MBfJHJrTLc6Z
9hz+dzLkKV9rrO8VgLwskw6PSijdODyuDKZ1srhcA4q0vzRbhWpqrJD+1Z381was
XRDJsypYhRZCeXlw8m/o4xzcfrHpD6YmBT58NzgQnUfraFczI3bSEV4SkD1W/jBy
ycXihyjJVQ12QqOx51X58elLRxxLBEcIxG5+srszyXWkA3rx4AP59GiSyDDhnb6b
RRQ+xDdJTazRb1kgY06JsiSMkE3++fdypsFYdctFCcfw1U6mdr0Tj6o4CijbKmYv
s6KKOTLo50cSuppgz1QEd7sxmAeseeVa46wRRux1OQMX9PJujUQBCVElesJSbbfi
Em8Pgl4bLcORtPPanieHdR6Q+6XRHjJu7FCGgc7flipCMs7HYsItwwJirUebY/Oi
0B/aSAGUsnZUlFHYZHxJT35N2cbubfvu1Dl+ShFwWGbEmQvaoqOnaLOMJWIFBp9P
bwh7yaWJNPUgY0r1kSXXS2+qhtEqN3FszCK1uflBVU/phw+2148/Lii9nJ794yL1
hjKEAiJmwozcx9etRcadvsW95uixO+5DcoitWqu0B+3X5vk0OpsE5PIW+Y60n1xd
a7NGsgvwLCioov5iFLa+ON2coOo0jnzFG24Agg/T1un9myxsVRp5x+SGuAIYBZ9E
tVuCdSRahg6tQFnXOqIB/0LJVDSwqdov+fvGXQqGOGAQbDWdhRMA1rUrW9LThkL0
M/w7xRmkEeerBJNgLonaCQRUvT2h7KF/YwCga53VFVyYJoHfGphWZr8h/vS/2OuQ
otQTugP3gYBpKTLFg7Tq1BEzpygztoWDcYLTEheXXSvLwvIyy7idWCyx9W42PXV6
x24hU1y0nmc7DX9mQ5BjpyqYP/PDEK3vwOPJiaxwGf7ZkqNjDejwVUojEGQLxZvn
BOk9pPKr0ZzA/IT5gBiIcy+CMdMaUjEfLvadzNhVwuXz6QMRbQ2meDazSsCT8dh4
nKXL6KlqAs6FGZdvcisYT9VdNVKnVtlDbW+6Ja9KXgCmak20VsxP22qAoK/pb/3s
BXQp6AS5bTwEsmTh7swqsjZkZXcoZ48o8Gt05oYxRYdBt6BBeGPT0iJJiwTcldo5
XytEQ8sjaIZfS9vWLCJ8rp/Mkd5iS93SpYqFfqNW46PsXrZto0d4HwhIx/RgZhTx
yJC1pjuHGzFbW/OgYYujz7eovKhlkjA/pKK2dSX3tRk3qH7/EECW3ObvqjYfoGt9
clEW79V+dBNrzVr2JKOxLDnjPhcgYSLKVcDS45ZDs+7rOYwTxgCMFlleiNsTSGGS
TUCyAN2p2pak88DPdldIi0uyHQWVkdMOT1qtCGPvLKLNLce3Bj23KEzbvnAXF/72
xtk2J2A2/X/kRbD68iTjkGnycG62U1oFxPj1+k3dDESsxYtk2l844QZdAOy4YMuG
X8DKa6fGuBA2+hPHIIf08HQTifAY/jmkkMOjRiRaEaIjomNvsBrqA6+FdAMz3j5Z
x1NR5Ka14xOnnwCX5AvVwTjqa9NIO1xDFze9BsapBT1FsCE6l3LXDj82joT9oibv
DdJI+ooJuQ0YjEeyUZuB+z+kwghy6DexPMl5dQNwUesBZDQ4HL6EvZ0EJ3QYc3Ew
VslmJFS+sPVa5JUiYx4GnGsz4h3BUvth5/Rmh5my4DDCo/VkRg+qk/P+DAWa3nc5
n6h1cyyLrozxc1RG2F/871rIte4bKoKYYRx8uqG8TK6iFPZUSwNPJNVSZErOallj
OXZFy35qMIXlucl3R+zg2oRbKoUqaEcP5Xii0C/0fhQ1VV+DVbAGxL5IsO5DUB6V
33Su2QOAcMLYHiB5s8WP5RHbTXb5zGzFrgF+wzVVTOsLnohiWcEnQDWnltM4TpGG
3enHPcVvADe8Njpe6Ar8tIF4+tc3gLTI4ZDP2PwATmcwv8ll7V9ggYYetcLWjHGc
++UWw9Fk44zr+HajT0uybw46gbjebD1JfbbVJGKy65KnETxJpnD6VYUbwmEM6iqU
HW4GOEMQCteEdYg8bnUXpcMU2O71hoj1FI+mzPkaKUjDh6XY0kkCIfT8h3+GWoEY
h1NqxADZL7r8rz97OdVsLiLhKVZydgYNJLB2W8GEItMpt1CXDGOXj6ezTbcr5DPD
bhgkqozOwpl43Qqf160f666iu38KBApDPbIIq4Pbj63NbbiEEwIyh5Wjbpq4Fnmi
xJlkGdOdCope+qH5AOppj58Y7Q9gHd4Z2oHqeiy1pNB/OtRCqJ10tCrOWeREFYlp
wTA7QJV16Y1m2FtZVXsau7c+/L8uxMSYfk0a96y2GIzZOqsRiZF+GdAmbHpQTLHL
cOw6tcLp6LC2+VnlQ1tTVZVGtM4nCXYUwiEjAEHmpkEcUaEfazpEn5tuKFpQ8AYD
EyLGS8l/I3s9zRhjRaisSmQlp2jhohJz9UjQmP49tPh1/uC3i11FYpZZIfEFGfMU
34xgnjXQvGhJfpuuZeeDkfCCGBWMz1jr55avwiE4ReCNrunvCIcf8Au6+rsZVQ9c
eIDFmvuxWeki6X4uWb7ddxGHtQeleN2fVjezBm3qHm40xHQwSbIoJcDLVabs9SOI
SE9lnLOXg9Faz5yvSYEr66Uw0SQB9Cm8wOE+ecgHylIkh3ZlWmEnTFDSavi5fjj7
zRe/7A1y7nXWYa4KgX9uF+nopEFcrG1Ol94gNrO5kuzPG3hAz6tfI0JO5KRiW6yo
4PtXjuPaMFd3gI19VrQIQa5wPfB1R1T+KTDrQBAPXkIOoNeM9ZVmO6ryZUg00kBy
CGqPsOc0/qcikQpEb010m/ZW+amErc6nDkLWc1kp0/YhJxYXP+RNHCj9Ofj2MjZD
vhLirq09UU8w/o+xZcHbzckVnIzqFLFFQzC/N5TWZo6tfOg2H3z6mvALaV9dPZGs
C/CcOZ1aLPHyltVC6WTH3O+esMsJhxpIj0IXwhlp0kDMDyDkInSjm6NF+rOJZVxU
iA8jA2cfsJfVcE4nO1iueOX8NTlLQHIwHtorBzdf/vlTBN6E2Q2KtVCymszkh0fu
1GzgeDQBLkstxDb+ymd29nULr0D96jSDiKLefOFwTzrphN1WWJTAE3lDwEuor0Q7
eyts4BxxU94KgyKU/00ztl0oDhTqsqDsFWiE8dz1YJJPn412Ho9CIK0+NOLyRyXl
3WfWLWX/Ca0mnHwzKVhoW0pOn5e4E9B4lQJFcBt3c1wS4yPAO7XBzc51RGLDBJDE
KK2IWdfiNS+Tj9WKTJI4Mwob6zSsQ2WnRUKXWLQycEQ0+8nSIUwzFwWJ9JnNZlKZ
SxVFhLevf/2DJHZW+G1mJgP23ywqIuksNF5eHDD/JJ79aK/xlUY962019AWn2jCB
muWnXJgxxYYLcGO9/52JTZZvXJPr9HyYkwIAekAi7xOAWB31HgbbYoMRuGKBNVvK
0yVj1aTA6OK2I32BdT0N7c0XxbeUsQO4H8IMiZzPA/RGAKS2WiCQ8JHte2wVbokv
tvjzFSc0ABbiaf2ab9Ve3mYl/Pzd33Fo0aoqZcgGEmyuaT3fZhL7aH88YlaVRKSZ
+vvJioF9dVr2egaM+nUEvesPxID7CGWuGXVZP6lKulOl+iMjLfhNpGbytGMe/BN8
RAJpv/USs6f/8V6mihY9jRT02N/pGuPePkHzdY4k0prnTIFfIk1WFBtWl2mZss7M
P63Oeo+xyJskyBafOOzGarP7eILBtuMX1EdlP2Y8SNwLz158EWCeVs0NHsIWWhY3
PhINK2TtMDY2HMXCLWrd6tgffyzuoXRlSDSa268fTRYNcq5Hd7XBXX/hjIXYMnQl
k4mhI7DQAQoYfhqiePuOCczHqNsLLEbORRjbutnOMgPdrU1Yvw+70Q/VHutLQr4n
O5NVbsJFbLbMsofjpyO+rThJJZ7LlCImCFSRajyGLPDCXqnQQbFq9K/mypHZcnqC
rPrxFoyZAL4lC3YU6yNzguZ95/anQmZxzcn7tJqbDySWbG2/YPTg/NAAmas47tMh
9EZH71csyAe2eNprS8Nv9OWr069/TxW/ab23+oF575uez6+bl/p8HhlEhTGqGDzr
XnKDSAoVOjmoun5AUQAxpoKIy3aHFWneb65bmM0FpKKhBqDLf6hY41nXefQTZjXY
oe/OYw08qoBCt5JZRABejCgUg78RA1CmwylEFZzSdd5oyl2ZsNlw53WD0NlwMmiU
PMpv5JEPCRuuANLaVb7EUe2ys2bFlVOiOSVY38OSg1Cvu5Nr5fIeuxaG/1U+6IXf
vTiDyc8RaMDcNuuAQh8nN42wutV1M51VpaZVmVWKAp6QtPh44QiR+DUF8A5cEspp
U/mWiWwxHI9wQzzPcGsNIlvOEum4Kqdt0ZRqlxif5CqFYj70+sDzwYt378pn6M3G
n5TbSVTJD3O+7OO5/qEohw5DspfwOfT84RGj2dVyLF9PMQmBHiz1h8mD5BpTOSK8
IfJEGG6Yxbdte0EcKrc0ftLwPgmcVDOjIgpkaW0YI2NmfWHsF89NyW7lSUCE1tgs
1+GTavzDHMwyNeP57ZSKrF1oUAIG+P/0QQ1A29UsbTiUR7K3L8bp+tYvyhyAuIyV
hyCkItvQUe3Y939VWMDGBYIjwC0NvKuEKoSPyZexzLFaeycrdeS4W5frHp/w9CTc
C2Mghb2ef637ftgv42b7bUsx0cmw1K7ICW3lLJNd04FqF9u4lRl+dRrYYrFeGe7p
SIeG29zGBBWz4la/XSkin1ZAOGf47j/PCdPcdvvdclHvlPE7rNMAWhQGQLKFccmj
3E8jgUlliQVx1LTbdMd+d1xMcpakwNkFCihwexhF0/K2I0n5mDoB/9eoc3sQnRa7
kBKeDAATV9FYh7q/wiXfZ1anuG3lL8DWp97aoGCxfol0viEPjBYKB2RkoOPmW9yp
kcWeHII1Xg7HrAAC14sesLRswIKEK02/jnQf073SpXkexOSoD9tEkdPWRAl54IdS
arbdDc32IvCjdH/E2uOwR1UppfrDFCNsRkliumzIQDs9Alc6SfF58/WroFfGNXNf
AcXt87i7dP7f6PqefH5p8dY2WRZyd8N13xLmZZqM23Ahw/Oafb2rFBdtjMSA2E7t
Cti2PllVFdTz3u8SXptBXYhIwsiRS8D6CZL5ZIkdcoFEvEPPO7amnmxENz+HAhNB
aHEQXvCB4j4Nf0q9/4UGGR3LjwagRkHRN0jbM6CPP1iyaa7pXvap96pY0XBI1943
RgQYCylxyLBNessqx3cjD8S0yMjfd0/U9lQXw4AEkNQyvv/29KUqpPqrnyn9pnt9
S3lXmotfIvnhX4SAWa8gIqagr2kfkhObKNr5uRGme4G7kVgyjk8/BJ5+iw3IamhX
YQ1bav0srSJsZPiPaP8rtSl0Bm+5jOscJBJFFSlKyKet6YS1Dxy75iZ4/KWLqkFs
pMNGtnsJyqpEpmOp67GWPYOgihDSlyb9STN0LXqK4GFp1v+Ev4y/gAOu9qUNZFyp
q0F3nGhpJtgCn32Q9IZ7sF6j8NUs1/GOvVrmJbvQfojWRjK1v0Jqnpd+K01AFuse
VIQx+t9dXj9WKtEc17Zb87qXRC1RlIXHPLzHxnfxmCTlmTVUJfnbVb9L7DD03BT3
X7wWobkQA5E2hZ5kIsyyIc9Jliq/fAZzxG9vW+t4hr+9Hl52AlE7xwHlXSTZu6yQ
c58U+jQD6ToEHPFG2WADibwEKbzcoDl4dTzcXkzDDa1tKUU9hXdaOJI7uOIwKCw+
m8/Jj3lOUuhf9ykPliHF+kEzX/wVn+zfWvDmfiBQ2T6gKZT7GuhpVRDV9IDmzSoj
5V0EGCHzAS2XSG8jEmpuyZH0x3fcjjyQlbrNsm1osYQNNtElnIkD+GSafY4QXGwc
ImW7ZvHNKjJXK0uGUMNJJwsmOKe5DGftf0DgQy9BvBdEc7x7s2096BCA314FShZK
EiR3WJFCmkR5uqzm8qXruliqI6cIBAF70ZDbCCsFKxlrx2cbZgWnUdRxldoJwxew
iV1ugLai/AlE7Efa40U7yiBQyICCqmQ+klkUMt4zkspq0v74QPdNzqmK2IiH5C3B
GCedU8CqnH4gxgxobSfPmlHwo087Ry5CovSV18lUYOHczNCUNyzRcGgCVIHcTYkg
NPI76xTg/vf2YXXMmt+rbtsuRiNoAptqwBpFh4dqYt9UIY7GHO8oKz7F9YLP6eyt
xAbeKpLFaWolvKmgaEJ/sG101FXEb9R/meIdo8pb+9kjIP3hZCS7fvHgfedmyV6x
ttXuHJwCrD0fgoftKYIjPqn6v6svSpKAY/0jQt1YvCaTYI9dH6UE13Zg3zUG632R
39ur2duQLrjD64d0y4h0QW7Sutnfw71fybsyzRx5VL2v5gUw49MGwV/bjv2eETWS
BF8GPgmi4qmXzBdmRfexvWj95oUXWqa0USrtxzVKpriTCh8L3SQsEsvAB/x8wAeO
LBllSn6KDUnmQiMkaJM6HABFdeJjANNJYY9l41RtiRDfPeTj3MDS7Ekbcs+oAa0p
md2SvDhqqBJLNsbdKr5CulPhzP5HiquHMFiU+xYCw4iCgC9j++dV0EXLlqiqtHK0
gXo3VSpGQuuArgP1TlidcWEcj9G9F7gdeJp38MoWbL2Yz7rVhwsCYjZZhEoYXKRI
i3JmxFhMhEde8MLCyAi62THYbMTwSj57x/psvQVRNt0wFmy13Izk1zoHEpSICq1T
M8R5Fn4ZgVrPbbSIYAmlfFMWTBzNold7HQ8gPR3UFXXRUTTqLRwWnJSbxnBeePj2
rdNGZ2yLJx6XY/vdFjvTX3Ud7k3UCavlwzOhJcvZdToYjIOUi7qfCT9yn2rG6FZc
GEwS+z8UZieoj6jz9bOrWPjYeAoV3WS+cprQzugE1E+M9qWFNOAAr4A1I4CnFwtD
KOhJ9iCJ7NQNyLYrFTjgsvxKyP1cQi86QHabXKP5wnFHDP+Aq7wMZfMAW1s2o9jx
oKDkmnABD7zaUuwii9x1eP0m3CRslhfpgWtFhhz/EWOGdd1WBNGopJUtA61rRaVO
yeJNWO2aq6teWnzrWnTQeDEJpwRy+d74Tcskd07q9XIgLKnE7MFJ38GUzLRzJs1d
GZ+B3A8G0Tmc/XH3hxvF2ruBNERmSuEZjl44KTm3gdrB5e5OmcNErClksEoUtmil
Iuux58ohLoswShZr7vlLgJAnHErYMoq3h4k9HTDuie068l4Tj+0G2pSKfXQQ/8xs
nVRz4hIW81+EQCSCy/u9aggMNyI5ETdjXTmmnvFGGmggYEyiw1XgzBBFJFqOS+RV
Vmm8b+oYrlReRtLBQEYlSfpuBne8d/oonXOMRcWPB68RDsLM0BAkgRpi21wGlbDv
9whDWkCzbbbC7gUqSY1DzA949ab7fNRmfeJjIOcqUvY3ULYPGRx3IRrcHJ33EQNv
nv+hvApcvzs7tTq3O6ILJwUB0meDWScFkwHtga4v6zviKvv2dY8yrFsjg/5ZqHzt
GhsRGGDyZyMpLBs3Rd6TByoqvqJ0JAjdiAj16TPAvtrUMEVmq8sPhLUE9jw5x5Ad
LRWPiTqPejHuCnVHN97ME22nHMu3dTEfZKeLET8JYw63+F4u/MW60VJAFZ8vYDqF
p41vQHW8OpzIRUth8R1eix3addT7dhRcWpBjP/nSO8UHRQtmrCfOHRnuSDvJd86C
7nBVGsCi8WDE1FljbH+HJ4PUezzQb9J73Q9nlqGGg4acFWArQY82w44wCJyR15FJ
JehoZ2pqlluFwOTyVTI8ug6cGh+AEqH4xd6iE96bQErvzKzmQqt0bITtb5YkkAE8
vwnNSqoXYFtWXlPH0Xmqu6yKXACHp8eSz9Jk4pMH3mCfeyghgRE6POCmsZSkFiah
KiMK54jDXHayoKYVa6sY4XhF666tgg2/L66XPtSWGRtsu09cq+L285syafSnZNfK
tntFwEHKKSLrGB1rGq6zpUK5WtDaaNbC5Psbw0vN2l+IbA4+4j3Yg33D1VqWeVHh
BMxBcAnoISpWgVH7hSm6hVSyjipd4Ouhfw9Wb1ohKx6a0nuwaKc45b0F6cI+D39F
343th5XVu4qIuY80UV/4zN6STjVWBCrqMUf+8/lMA5giWU8z629dOIxO2C9RJuLJ
ShNdCPpA6fmouBY8CJky6tpD0GGFNanUOraB/mMTxFln9R7+Ev7HdH7GoxCaVJWL
SCK22Kz+6KYhPzm9XDpXcbX+kEGKqTV4BpnkfYlzKiLE32aRfmxaFS6g3WyOSs/Y
QJZKeh9AQ6JpwB4GkHSpY4gVqqX1mIZHmBGRyEVQ7F4BU2q3jHZx0Hwk9oGIQF5p
CtbMl0KOR0eo7OdvyTBy1phRcJWnvBVTARBA41CWauzFQzXdbEolvgsCoNpvXnvN
pRKfYrudiq7c7hhr0sV3RSSubAMU3m44pJ4+9+qECreaQV460UQ3uGF8SRWwcWqD
hVvLFToVW8QqxU1LV8F/gtfAA796R2zmFj88D64T/u75saqOGVQvk/CfvTWxs92W
4BnDLmK4CqlatovqubZlOld/Gcehr/ovV1pl0XBVpgbvgMMXlP7K30kWnd7gZSgG
bTpFEHHDi/x8nJ5DZ4Dxj5bP0GiBm3i02M9ky6K3YNCvDnjLYRZniNz1iUYWgGtV
Q4T40juvycmKq78DDay9rM8IV3aZiII6uolGDz/s8yRdH3X+qm5FGNDlrETjw6yG
CsX5O7sGnoU1qFPxOK06XLSxSoP1fnEarSJwXjQ68QDN/ZpsUZxLCLXEt7TwSQue
T8dnp8QxjtaG097oTdU+da5gXBjEUWRUEduPTEzdh4wz8MECY7olzmsV0nyLDfo5
rIvJhMD6QRfgQ0hdV1seq5T3H1jc635WIfJSkly48rEGNRQ69tXJSjXfg6NIFA42
V4bOIrFts2V35cL118INOEWOq2GBatFvXTMCe3BDqWpW8X58Ra2r15XlIHmUzG9M
zsQn5t0LCEoFshwdCnYrrOzxFHSQqnmyTxipI4mU7DZ/xKsmbys757teZHR2hb6c
6QKyiASPPMq5FGmlKX3paQcXPLf6VVsQUPwkhphGxFVEoGoHt5JnjDL6ppi98Jgd
LF3t1sLBrDOByXhq8srAzMCX7FWY8S96KvQ7zcGFY1sybBNO2BWm1G5XSmJ/UZGa
W1ampw8sdaxYwV6H4r3opnb4l4drX04z6IzzJpLJpInFT26BBogYck4+5sNmF3uk
EmjPAbhJ9c5nKoHhAQvnKtCHrL73cba4ltKiKI1r+nrgPFo1jFvm6bZfbrIT86of
lYC2cwuqh0XmfN3U3sggi5t2GuKhqB/gWhOl+zg3VijRdMOJhJGOLZ7r26lYYMMv
vtag9y62Mh06ig6rcEPzAzrIDxRZMlsfOoz6wiLiHqKUDi+FpQ7mau7KpFGJ+Fe1
AJ6fudARqOKN9STPaWXERBVljDLJXEnIyA4ATP5JNI8jL03VUDaFKQXtSPojd+En
VwjCb41y5k2T2XPT5dzjlPttd8i7PcZwC7i423kZheUmdtrvWMkSREIa5TUP4SRC
fvF210OMcT1SSyyfMdRbSb4y+7PD87VOcsjK+90k9Wf4yFxZINq5D60EEHXpVONM
dE2EH1cju5Y6D8LMORqqOi0tNFqvcd+datMtnw9Ft5sDFHFWckulaLanwZNtLz6+
adR5sqt4w/bebFNcv74UraPp5gSAHoLMrC6QYE0yP5YvvOS6kIkZs1kp6cVSTG+u
ok6dPtVHUm5npOuDJdoGXar2dLylwEp4tGn2bi3XKbTNRVQOd9K8IXjX2vvSDSQI
raO/S3iwhWfWudp4O2KzWUVt/PjtgAlu+9DmcLlq/3YUPjLNDZG+tCoNqe9bRHHU
rN7JryhScHAT4EDkD4dNGHweMQYUAtM5semSqJj53Rx7RxJiJYGXl+4oRNr0MMA9
qDIDfrLouhNwP8YJPu6XWSdUraV7bnJAtrrbV/qWYor2SOQXn+8dR6rv35ui8R3y
+gmL8cfkTdCDMIcmvfAGBDwUs6Sxj5ED+SlVia4irY6TLBUBiJZVsHIiIt03KWba
n//WUUuMJAFSj0IVDPtubaPF8e1MhL5ToTjGsiWs5sUI9Csw4BmFV1RH7Pf3y4I9
rdFJhxaWOownH7RX0DNyCibuwfuBrdIh8pkIx/ywibme/51GKl7QeAdd8cyTGJtw
ShNEalkGnC7XrF8cAJktMlrosA/FyTucMRDDgSAwc1gI96pkLhBFHBFF5oXL4lcf
QAB7Mhe/02CZlWZ6HzlRXLzMIcnD+Zjanhd5rDps2sJ+mij81zDjCDDRTnf06uBe
FUhj/bRfeRvNtOl8caSgw4A/7NjGZp2k0zAwVzB8DTim2FDawF0DTuxXc7HntqRk
6UEDJ/Gb5nHEBF8AT6jJVhSsqtII4AL8UHRo9cxkr5o0ugfafA02LZK4TF57gfkR
Ed1oLunCFohitmKmRIp+66CzIhUs0UszKBmvAnWgAWWic00ajbvXJpO9QRBut02p
xkbWJwzQGodrfs4VqRZmYKnGHRl2nLEeUFmHJU+ILuPoNQZTsQLrybeQKFKIu7NU
4r5r7BSG+eESwKjEN42RUVadMmGGfyl2/rdiUKgl/tvYx1KV5eWNq3NQFkPsp3mr
KDMRk9LFrlcKoNyqtpD+1xeiUEUP9ZMFVj5EsoQZNmru7gWLGrRr1tmtHhfKj+Cb
Z6cyjqGAifo4yaEmEDBfQwejSeuEj6sshZTOUVBvyvTRyJ5/xPr6HKtqU0ZRjLpO
AmSv6gDd+MR7pUW3zJ2iILnv2bnvZOc4pT+dONSx1Qe+45a9G8iMLqb3DCOKC0Y2
W0r8+1jNsLqW3GQZxXQjO3ms2NKgbBQXyMcjrnHFmNDWymRgJlPchNMVjStrczJd
+YYSYMb4hNTshIzb84pyLgzTMaqP/WGC4Gp9JzSHXjLIcb3j2YXeh6VBJ6rZXZII
ct7HVt07BGtYl2cN/+yUXxTe83upfSJXPoiM9uzDvYGtInpxAT6NQesmGASaYiDX
gKKsah/ZhukHc7zizpqVJfKxykGBw79YjhMczJ6lFyZ+gNoia7+cZbtJ2KLGQqFq
1kOsJ8a7zS0xhxD+nCVdsvgEa5xZFcrHty7wEE+YcDpUOdx4CpwdsNqrFBwbqMPS
wQXZtt6m9NXehLBsxgknjoC8+Kl/3H+Fmkno4a//d19uKB7uJ5v7DpZ0Pm+FyRBh
GvCEXg4igd3gXv5rjOf9vb/YcQ1Kc5SNRQL679FaUz7twaW6RbxlC6SUzPNvCpU0
N3B8e5X5w2al4GgnJNb++EcBj/qeEEoY5v/Ac7SMb4XyENF83J584ugV6hlp1M3Z
vSwVQDKHWwnodplW+BAJ0pOBh5bdHmo60Muvsvj3wjYNV7IdNwsevYV9Iup87IBy
XLNcQKXfjlClHJxhutmJS+rOBbxWrrqXvesumQHDd8iF1PuVClQWR/acW6m3r/kx
QFbTWV8OGwjEm4RM51OvBjUhOVxY3wfIsvwbs9voS9JXutSdDzOgXTBmWgY8XZZG
awgDFeZZhEo1pDm6wogcuRIKkPHpmdF8uXtkzJVkPHQAveFlxIh9OgyGecd/2AwV
3ew9qr8ZJcIz0Xb0xIVynaP1zbsSH7Mm61I6/h6GhuPyr7uRzZTbPeWFL9rivvCX
k/uyfLZF7okGZT7aOnEifT055XM/yfO/+FHLOxwDfe9lYzACbZC6vjzLvOEIXYDc
/m3W9issfPcc40+dBjcsIARXb4gh8kiBbPu8/JUWUc8+vfTuYg3XL417d/9h9nP9
rcBNlzD10KxNpT1iYAH7UQonY0eZHUxiXnHn3K0jTY7ZI5JAML4QDYEsU7quLBsn
2oQWeVIRg+XYqeiit0ab2alsamyo7JXtp16wCRpYZwlORH0gkJvcXDRxWr6ZosRC
G1l5lTMD7BhImY/5N/bO+iRt8GRT8bPFVrslukkcsXxIrmuKiyBJFHSAuYuWwk5Q
DpteUDl10qw1Ig3YCUIPdmWCYMKXioyFNWRbSUohzK7o7BQGFRgDzNW3uL5PjbRQ
oQIa2LT3XiuQrfG6xJ9y0p7tTm31yh2YOz/BtPj8fA5X3HuMaLtHHtpM2UVUpsg0
OzyoN7SrPsN+7KhCPFxMbmNQRhz96TKNWEN9o4vYsJbUn2wOq+7if85iioMdqZqw
R1oyPVekaPkSwtA6Wu5df7TjF8KqGl776tLFciJ8eo8M4YLHs5Bq3l8PFjUpIrY2
wA57nNXXPDB1NMz0vfWCU6pc945VKCl8UDeD7C32HHvsHZrIOIdyievfGCDguj15
Skc4hwis0HU5eIPaXUyUGsPqORMKYso7NM/iW4mNZcY3ZRu2W23T45vD7ASTdRWN
LGIXSnL1EP3WGJMh1g0yfyGShNQb9ioVxGen1Ux5H6QPIqOVc0hL/+lOpU36xKm+
LXIjpjQpVceWeXY0YvB4yCTbaDB+001hklEsJOUnyfHHIJHTwdjRLypcLkVqGpXc
0UbIF6r+Jw7aVgAif+bswbY6tLLSlnsqWbNkbFZ4JVtwmiBiDtbjExEdLVZNsQ3e
TboMAytXz0eqOaZYh4H0aO9kZFgLv3+crJFpC+FrDF1D+Beenb6j/4b7Z8xzKGT5
vWmYO+pYrLPVEiZjOU4NbecBiiQLNquXGoMeh9+p6o5kx5WNlZAwr+mroOa/nE7Y
BJqx33ifoymqJFC9/kCKYJ/GSHskieSnDIlFtq/Arkje/89uFHLFJNDwpaU0RgaZ
gNv8HIKTgAL6UM1Vn5O7NHhe4Lgz/4y++j7/omZzeeSQiVIy2DjI6lucWX/FsxUC
xkmyIb4uZKOItP1MdH8ldYXk0s99WSY8mQTNHy8AZNnyCkNzUgNwciQcwqa8Ocky
/Cr3Wt+bvTCai+w/dM0ITWMq7y0VLI9dx6szvv/BUeCEg1iANVUB/8PTO89oGe9A
DOGARsczvqMNsTyWTJyx87wVTduOI4lqiISU7pb9sO4m1DjflGge9jkWyM8YdQex
TeWQ6ztAFC5C3ioFQNc6UT9z2k4Nt0s51uShVBzaQ/eMJnBheoC4lP5CIqGZTiEO
LjXN5/lZjC9pbagTyxDnPVkxCHnprPtEDWwU1YNQthej6Ko/KQtoye+u8kAO0cR0
KXsC5vVzVgTvjIEAewakulNUn+urC2TFwAwyBL7gQ4BfRNF3zHftsnHRiJq7utNR
SV7FUnErtQI3YS5anmIiQopsYaI5Tf0Om391mC/lcEr1jBXZvG0xEdqGbhG4wnR2
IKws+BeVClF3p5VyyuS55ixbJOB//n8E685SbLun+qPobvL8XdLLygmF1aFroGFI
cWhgEIUtDArKSPuyVxc9ShKaE2lDVf8DS7al5AymC85+Zh5MW0ddenqICDjE9xOI
/VN9AxGRYJEZfCyjGrHP9j8zbBORzGgDBcGIcoa4kSOq/AKv7VWytdJWjy3YeB7g
D+1bxRYABdXgWGdqhKtvZ4BKWb5XYeZg2eehM0+2RJ5Bf7bhIZZjTVeU3mg0ZS3l
/aTeYmhiJb9AWmzzi0lbi1y9b3dur//NuFleG2N0LsLP5O7CAr/5JGW7wYFg9qTe
6OV7srA/IjzY4vWuYNbu9jOORMW6dmzhr+sAOp6WI6L8DW2JNSxDfue9NNFgdc65
lAIG5uFLMiqgiaFBdTD+lY5hn8TYIwXx7nfGJHrWH4p9X7CCgUJ0U8rejAc2ndFL
FVRZX8egkHT1EE2dy34WV6WR9LzSU+QfcWi7SfywwHkXbHSLKbuaOxW7xTaBgga3
ofDsurn3RdYxMmzrrMJ+7gtDC6cajr5OwoqnYzpHX2vBhvkNukUQGDtQU1dE4KhS
wzG69xC97a0P6/t/KGN53CCJVTmzyIsUlfHOBxcoimWmkfYVO7ErvJh9aGBnbrQI
EuVNtmkQacfoGLPVCpzCcQrpXKfYe/JnNdip5dfPRfs/uosYfmCKTXOz8S3A3kxG
C8jt9RCWwGtQOf/PcxR5w44DOiEDVLROP9Ww0F9EVEaw4DixZy6uO6hcDWzukDBG
58vXToVRGErxFVEvuR1SPAWGwSZxXpQVjuPANXFTeWBV/T8t+Xegn1Lg8C37fvmx
bUlE4LxGeaTIUWL1bo7oGkosWh++StY4RVoy+KJSKaNXRmB/c03nZEPToyn61aUo
aH2ABbCnWKUfZwd3u6y34yySnaSsDN/K9e9b/E8eGDalq4zRxDuB2z7B/diVOJtx
BX/E3HrZwmYaIKn29MtLMc3OyEayxX+r2yIfIdex3wBpczgrHsPuaYBlU/4rBqpy
y3fr9XkAk6DXhILBFn6hAAPKAxTobwSJ/gVqmh3N21G24NxbbWo2icSNywDvpXWR
Y2Gk4NXoixFed3dJdi6zIknYT3zs9mqqVyFldsqssPIXejP46L55ZZM8ZYbQ5lFZ
l4pfYAJVndA+UamIiYhuTb/0Kbv6qKzHne+l3vQ9KpM201s8xR4HuwSn0nq2COa6
ggv+7Yb1+KTyOAla/DmoRuQSUrjp0FuUeWcvaadyxcsdIaA4HV4yE0BHpi1uod47
PRQ38zSzkaAXAgguGrCxLX8KfN7qGF9uiElfaj45H48MQBXAPClO9ck/NFej7T1L
0W0yI0XtcdhDDvJz1udma3+lpZVUV1yqm+70pR4RZ78PBbfoqgPC6v6lx0WEdR7H
9pNY9i89y8oHEoAHl53ICkbfkbcP5KYrBVmkbORcnOWdSKQvJzAN0q0nmfiYyikh
12ySeuEU1yRRuDlphdp8KuvFcmuHRRvsed7lo5+TzuZMyqBxz005hnN7lIP++SMw
5qRTkBcNonLXEPFVlp2OmOSNJEumR2rWPTjTloXrryyivqPPvSW85FIcLbPhvgN9
1hmFke3HRkHWEnIbHS6G2jjh4hyYgirr7R/Wo6KLJ/8OgKVXbvhMBvnvxQjw+m2F
/4H5BduumMrZG6UAsIMdWrYorcOgC+U1Y4kAn0fJtRaBCWmIGodwZX7w5zKAK2RN
sODQ7ohPwBylgAkNd9dQI0CuYZAbH8MYfhQuEJns4sx2ZCzZl7HESMQ1CPov3du1
QB86zIcPfl2tdt0CvwLWIeRYc45cJdAzKomcbRWOIFwV5GwY92KeM7uhApJCrZom
2R9N3m5ecnCSugUpTHoknEemuSmMEFvVQQiwXoh6yJ0dcSwFgADSDIYii1hVby+9
bTwdo5yryIZxDiw9xVaJf+c60kXXPSKPzhDBzuWX5NcVj8sYxwJmBB71HVnt8IH9
rDDCXO9jPeJhKa5V1PnxyB7I5AGYGBTPWWeLNuWLEHLzeNjbzBbM3QxRcVLTlFpR
llQdRDK2w8v69J2xM4Pz1TKcnFU44SmjsgU2Jil18cEtpFqG3Q4QBVdV54D1hpzy
hwUUg6fWqjOLf9cp5+KehWJNOmGXTHW5gmsP2hCOgNTg1749SdTIxz6+lD/1FP4R
mV6WFD4YU8Abw5Jswlnr3ERgTh3AhIQ3pv51RsmI2RHlfeZ+hmTGOCVlwc6C5b7L
5rj7JZ0l51V9Cn5uZ3oM4yiG66LHNxD8p6ZQnAwu9RB7+NCLfQNHorcol9zNBlKp
W+9/x6ws8kgCz8rAh5Rv1NqrByfpoSRE9iEWsz07hGKnQ+scE5omkYuHFI5tGeOJ
e6sKp9C3kYfRbE3E650Ou9I4gz0ngNAh+9E6aBacGUsnm71f9rLjb/XCnOyC3mOA
xbXXmIU6zkN2ek8WSCABdYFLK5TRDn6645Em8J5/gLM5aB/a34HbnMeZpivq7ll0
jSD+VaXysPTjTKpi7PltfvwQlMx99Z5bmWWiiIbt5SbUtHDrcozHwZzshXQj5G8V
EZPjbFv03urt0gUtTGIDF8VV48PPqqDY9EjlKKDg0S+foCbBUbQzVYcGMDRMNDet
70c0gxt4xPjWlfu82FfJA6fktPveK7AGUh0XLKWmst+21rZiGG9nsoOuOFCaJuRs
J6oybt1yHw7Q0a40h7qGCekRqkXZak856b1NMLWfuhAfYDnjGhk4rDVaGGug+OTz
aMWpHYLDhMqGuWYzO1PYNgQ0PS/faQps9SxDO+STFkwoZEAhpG5mGm8/do97m0+S
IULa9EeMvdxsFGHK+jMeuT9/U4MJyXocm4nW4JTd3cSwibH8QSRj3Ejf7etNmBa9
p7QbP3mQQrvQFeuaMqcCQSzLMckjxkHKtGl4yI0uzNk+YpEIf5/a6060fFiQDwJG
p5bVgbch0V1grhL0FKHoBcFvxyLRD4IPqWd8f09cpnd84wSfh3ODrLycDEaqMtrv
1J02Mdj7Iw5RQb6SlqYWtLEN5quiaHj3U+2v3KjMbFeH0lgpp5qPUOyRBajpkGfj
zK0Y3W5TPxUbxRlcJp85BP1B8eg7e83scw62c8WxkPR5c5JQQxdBpC6g1XRQ/49I
LGXDCKvJrubGfzsrfUifairDYTp3W5UiVW9UOiHq1c5Cw1OkYOir565Iq188Pqho
BNmfV4Npq6gVbC/0cpPXmS05iOT4QSdy6j6kvQnEYmuyE27Mui4+2iEhVJLMr4gj
IlXhp7qxd0CKKfbnE+lVrvF1w3br8HR0KbFvoSs/l363eLOd8uZRuI29MRPUO1LL
Cc26TimVqnED4oCDccorGEt4zbqgMkJ1rX3AO+C/lpURdJi0A1SHWcRrmnvTgkbP
FboJyDI0EC4XPUlLBja/3aTXTb2BDDIx+8kDiuROKLfxmB0J4fKBELCDh7fIQKyd
TaXoa5vCbvATZydP5RpG2UDnmbl5NOWMTYf6W3OWZ8S2+KpEcgBE0NVcpftQzRvT
qN14HAq/f3dka/TEAdhI1nfuFDA8mXxgLHHSb3UxBPpcnRvCSbBavTmn0l0YJlST
ZKht0e292lrYln8Kxl7B8nPmnLwQwVIZND8PZcl3gcxvHQQFR7Uk/tBdfND+svA9
PsQLWgxGyf6nsVUOgxw64HrTb3NM+g3ps54zK6EFWcR0x2d0pDix4ms2agaO3JvU
FwMnq537pBPnIngr71U0q5qalpYEceyOr2EUpbEnnp5UYJB8738hIle43DEC+5SN
Y2gamYLRbaGqcCJ0aERliRXOA/XbTOgMc9pkBhbYjdzZgrLPkJX7ERc4bXH/w6kp
qOrGbgmjscbMtPZdcHz+atDbbIplAgbpvOrrNi6HEyKIXMB6rqnLY0LMJcf9qNLj
7lKOdYD+bxx78B7KrqQY7bmCdMZBvsh90nlnskMSarzplloMcXhOjtfWHzzQFb0Q
608YMtUQ/yknxpsZ7erm25/ZEH8I1Oh2jr4WXaztzxoxEEsChkg2WDnEocnRdht8
syByXC9U5VPvHCE+X+z/GljYviqOE/gLE2r/sIcku0WFh6CdK9Y6J1A4OOAn1PU5
0ib+7NdEVkdwjRQpBbHCOE82Z+j51b/bhmXf2DFpApE/6cdzAA35I/tACHH0CMBH
M+h6krlIwb04XD6w94BMFQntIQY686Ga2PNqxXRBcg9V0W+ryMLpG6cJm3LCCKv2
ce4xoPEtyUCJ52DakvwCpw18q6bWZTsbSz9bemPPKQWiYOgzZqPh8bY7ufIweTBU
LGlE+ZRloYZfuajlmajlFMmPBIdH5KJnVKvDoZ5JiOcK2XcJrD341fJCafji0ARy
fvtTd8p33UCDVXF/bxhUmOymSosKIQduWFGToXMmTovJg7iIeVUE5NCugJFWUZTo
AVAtawC2FGiV/JDqvaLlUafNnoGvhGm0y77ZAjY95Y0qnK5QIM7OnQlljT1AFCeQ
24heoge3Yab9KJSDkCCcrkQPVRiEzLypWWPCwb1pz+qC0v36h+ZsD2AQHxe3VnlQ
47T/WKnSvAlWTxPH87nncGdXyAl/MzMceYB02Vfn2bj9Qgi8lGXGeH9h9lt5SqZt
NSl2yjLBhx+541jwY2OihrmqzZ3zSiO+rnKix0vWwDG/x/6l4uiRM6J75IdxJsIm
Fv/ubiE/cRb8PgS6quJIBgs2KP5Wf5r8DbItwDQF70HjCku9YJ3+w2u1phAQLjxT
06k3UNtz/M/L0le6TiJEI4wD0xcP2DYZd3QyqNem3AqAiBf79K8jbL/ZCDYm0dBg
WYfS+z1Z1zRPTRKYj1chgMs4GbcC6UmbL1R1HBfNBYrf34liVvSanTsSwlhhDiPF
v2Avvm74jlbzBZ+qj0FbCGXHYkLL9NItElxLlUsYclXv2tIbL3a6zGtfMUSHqsx7
49DB+OO4orXqVTLEijuZ8eBTzPKBI4++rTycSTsAJ5fWCwNqqvpx8gRR4hMkgPdS
p9N+/QgoqpwZaunePgUeTeqnrQvBj3A3FRTj00McatTv3xbdqo17QbWGfH6QX5E2
M93qcr5mtO1v8xiMPOIurkqbjelUakF/0t5Sd4B9HTlYuWBqt+fzWDVR6Eig4ehh
NNS2aeQTEylUwlIZbOKQHJTS2Dgd2fGYvCS4/QqxXyb//UnuCr9EGbQJUXS+3+CZ
fPeO+7AuOlvyJZjMVdEBA5nECXaSfdDfxboU5IFOUjHX7TSQY7WF5Zf2tL3Kk7w2
sfjXAd/z3WQKh4c2UEYwfiYUYa5CyQw1ZK/Q2JQDBPu5XZDoah3IS+KqmmRtG3Av
aHwnqUpthLeO9Q3gRdoyCTAYbRDqr1CTr8MwidePYDHY1Q2HyUNTbQaGdgjTCp5Y
oqBd4+0bjkXCl2lWRBrTkwH3mnRBpJ22CpTo4NV7ZFprJGeuGcI1WFwoEuokNxQv
kfMAp9jVcojD2JZfLqcKmlPd8CC6Vk/wJ9qF/rGcmSfylvuCPeUqY3z2jhBU6mxI
j8YUJ2pkDG/L/P2ZfbGdmA/U3vIGeE2lG31ArI2SrlywoJOeGDgGavUrb5TksU83
MN0LSpS6+iiu/5IpbohEO38cJ9rH7YRkevro0cMn/XFUBtZU9psMI4ifkZXX3H5u
auUaHieeRq6QhBHpuYE7Q/3JlwJWmLhO1cvcLzyxGSX5SWvNcdKOmzatmg8rNKf4
R02YMkGPdQB1HA9jfnOaBZQdZWa87lkjP4aokSiVnF7XmtLSdYjVTyWurz2cKH9Y
m3XW33Zp/4ZeA/ylWu6s5JyAt5+Vlg2CF77M26dQvHoR5OzZM8vUEwv3JgTBlWZS
cpSUgBwl4ACeTtARuk/lEl8M/mKPiBB+FLrwQGgE8ymtNsFG2qHh9qdcx+To3sdt
xZnVilQKSnRC4k97+mQyW4gao9npFJQc1JCW9LQko+yPPRye3mdxTr+L4aXX5Hbn
8ifej88y9eheWvbuwRXrI8tQGeN9/s5Cy3PkgUVZjURDbtl/GuJ5OrDGSHx2/RE+
1G9R1MUBV8owO4GO4Fd8qJ+nya2Q5+5CiIDmkJnz1scw8cxIvYwF2mBfEAUy+i4S
ZwNM6Egy4b81kcyGrjNzqObNlLWc8KzJP01Yb/r1QWJTdV4lZMjlqA0Q4rUceLfk
IMcXwVXyF7Bd0pyrA2/4yUYRRuplu/nifIAkhf5H5ELSKDUZYIIRbNjIuRAa0C9x
H9MLabTVPKEP5Yii06SElcDikQIdh6tJX4ng8FdUzUDobcHdDQEOSadntzVSBU47
lg1+9uENH3AyOtjmwO6+/KID3jegdC09TwR+zXP11+++6Cfc6jBVi7iMJ88IKQ77
YnpdpBi8duFigS5sDWawRTBnd3IE+57akhQ28fqrlghkwWWlsDwrRh6iuq4fICa1
1K/jnekNjDVQaREIXtGZZmTW4zUlxCWlmJuxxm6rWRRhr67YIS27CTbwEWRUxoqT
wdjwgoR9SpFLuKuQN1CQihx0atO/IyeAdxhukEj99RSPEBC94XfMf+742NNGlYW/
j5QexPM2qoOzn19haE6/IGGi22n3X5k9EJFqr1b0dd9ZjaxNeGJE2UlREqmZAZTQ
DXQtCPbRGEBk824YV/XJs57he/aGUheWSdH8UV05cAKDDoZXBmlMV6eItJR9LfOb
7JlMftZ71lDLAj4XqZc61M7kkLxBVisAAb9R27ZNtu30Wb8hTsIk7NEw0elKj8Q4
MSSl1N7VLnHjUXTKNO5kt4TsXPeTri41p2Rod5qyZtUbY2F1GuwbwE57G25zgljx
L8K0zOH3yJDn6wx3MkxBPqKJF2mu2wZ+envIpaa/n3hU5acFUcPtPOJxuUXopMNe
Mn5mGk8FnETNohAiOjO9FIJ827Zq4qVXqpM2Y6fd1GTO9dctKnO+llnp1RrQUR6S
G+wyiTUpiPdOuNZ+dZGloSCy6U/biXm9gAPF02xyu+Xdarxr+4p1OeIT9NGVcBfs
i9mFqMfoxFL8Z0On5X+XzkB65Wr8hI8VRDA4OpXgyhVeo4SuwhGWfp+kQijfWU2z
rKl3J6rGydCVc+OzBYYf84edcvvV1SEDx0CK7bV43xpJZ8DM0VmVES4OtumkiUXy
yUYj1n2cY1c2MgshzNj7IF3qS1p2PwLoCxUBDScBc9436i3HAMZwFaKCKetCe9q/
+qEs2j2zLGAEabCRngnIz/Jcap+n9GfYlSFdOXkHHlkWbdS7NWiqrBij8wrD6RGp
ZY7aNeGzbW0Z2biP5CSluADiMTyeSNSObryxqkEXDl1sUFoTafGFWhPw8gL6aG4Y
YVx9QTjOo8inhwo6gb4YnqCL5NgWghiUAg/MQUOVJay8lZg83tSHkZ6ay2MXnnBV
myRi6MzlK9aZ5/ki5CnqFC8+1sweUEnrK8kryifTCKrGmxX0mBJoL70pkRqRZ7XB
S+YjMQP0Mq9VRr6ckl9miWYTbLwFFnWnqN99u1cxb/F+DB9dkDXdpWeADGeHvV4T
LLzEBTKovBO5PQcBfUPnNwjls5ObPv7vFEfCh1y4ktJshQgcaF2LTasXnvtNiluk
7uml6+muMUeLTfb1A1U0Wt7sEuaC4OG/qAPrVynIENOmMqIijFj94ArFgGjgQyCv
SOS6RFY1Nu8nw4IhGTv1SvEkPL7XxAFdyUlwKU3pYMHIjGR0J7rUAReDWhMU1jLw
PEj8cHSbiKCUD5MORFED/Re1xIJd6iX6UYYbkH3WJigPCBczEvc88njZhv6xdTWn
gKEiGDAObYcriQdEEExaFLCuQyZkFcF3NLylVZh7sJX1Tgg4T5AGrTiNnzg7LOrf
i3Or8nWhCJS9+zsrGpxrOMSkcF6cL7gH2iqLyZMwxUG/XYTpjCKesm7emYAQTRL/
64F1JuwTSkYkTepUozhSple4tAf+EQGWCE9u+WjaXSEFoE0KH/Nwa+48Hg+CelD/
TaGhdfkzYEEf9tdKxiSIbjVy8kCtXpqKDFawMFudWCqWTDNRK+/mMp3oWWzWS/NY
jOZf0WzgUeM+hNTk23HbCsM3NKdubqgEKV/V3d8YHrLjjpy9rnrAyPt9bGjfJj/d
i4dSDus4LREJoQdnacjhbgql3oZt2wUh+AH3n9MWIXsdQrmzQJfJ55tx9CAb8bxg
YsSs1U2OHpjep1nxjcOiTXeOUYbDzWKSdjYVpnFU2974EisG0ccgppLHX/auHeAK
h3vtU2WPcx1D+Jwmd5CtJ1kjXDnSP0IX9KeWOSdYrt19We612C+442PTLoN9aByV
o0zHWWM/B0BmyfzYqlElXZbVIiZW/u577jUoH82A0ET4cpA7N6Q26It0Ch7MLPPc
QTGNrWIungzeu5E19wUQPmKZO8TalHzUWsuc3/c/zDcSFyVUNW/PkP9f6Tm0VYQr
o+MGIz4Fb0x/dtMW9UDNd9kYGkTKe0BrgxtxgG3Bl+inBQUeU/A1XZ7BrF1l+Yx5
s2usct24n30vRMQ9LpOHNA+O1zZgjDWp1/HNdfMnC93hvxPYmHpIEcci3mGX8n0t
rybKHf+jQzfEo9Hq97MOkEK2clKkNkKsnQwvv6lZE9KsK5jowLRL8ZPfWibn74MX
wqKcwgHn7H3eUbfd4/RDJZ2iRiXPAF4xlvcRCWBDhf2c5hKugYOBqdtL0MWe0XPq
3fhPd/uJIHf7Whs1nbjKWUPCx+ZhYVZfUBa7x4fgiV75RvFPUk/kfe95y6rEVr18
s7sZooRihS4Ls5vIua4RAMxqUavQpvw70C73eMzU7ra3e484x1SbWdetDcMXbq2i
nTbaa25vcIQxnV7HbNZL6cScPnAVkLWO4cNLMCvMhWNbBwPj7WfRyrsQL2ELD5ZV
ZhcqUCnmVbLW4OEhHmOkFPJMKhS0gqcMDeeiBlN6si4zLJ8PdRB+QS+VPBi0OOOK
okZlknZqNkuDwFSX1GT7eR578QicQuPG+GkGHARyJB2abrc931RoTHCWEKtFb6xw
XADt9IgzXHfTnSxyvC2YZzNqSsYoyZp6YjmKUwGhM8mMUIWFXJsiqBqKWWKHmWos
MjXqjzuGpWvdOAyi7+VPu9HYeZkyXYleT69gnofwpimnDwb2Kfqp5pXDunTLrIwg
aPCw2m8GiRioyLWvJgt9W/jCW+GvRMAHFlekrrxqAPCYVD0i/n94CcZoDXsQfvni
EJzuRKCgipe1bhskB8qrkngmV36RjpH3RzI/tbfAkENhrHxeGgs9Fu8jqTi7fTzL
+rhOKcO7Fc70qiEGuMmw82CKd+8YME6tdWgtjMRcF+aViKUJTI5lJwF58K5hSHKt
4jLfVJ6nMhBYk2db7XOiCXEtBqJ8ubNrpdO7TM22Z9MkmbbCdVi4vpC1FE55f7WK
8BDVvb1wURfgDWEM5RTokHsrY2irqs4SzSDcvZmTP+DLtyb+91BSjLePbGH2TZPz
idpWisjQngHkLX5sdlUeGlx70gjh2HbanYH1/ngNG5Q9Oxw4QAXYyh1+SEhCvKre
jAiGyKANth2ShgYKPqhEeAU1OUz5wKkFSsMISCpgNAsfV238LeSNxCQ+dPhV/axW
UJmfpNJib6dnyt+HLbfLzJU6R/AKmug1ZIMCT1j2gYkYpzujMK9tFYkAijynvZOD
LrAXqeHpO36BO6lswvfaC1PnnmbrPEfiO1UUuGng3h3xOHjgDqMlh8QANWk8a8Al
RY1xX/oRL7TsuZSuiu7NwAOa6OEJvzv5BUbFWzSwE4Ex2kOhMHgKHNiOV4o/21zH
0729Meo0dzhFdYxmyTszuYldIlvYKYGHa76BEi+SJwu4b8GhOPYwVfxrOYy0oLTf
HQQa/yd0Dxzvyr2Dn/+FAI23yP+VYD0RT+tD73duMj3HUuySXomZSXQJcM8IvM1Z
RPWP36n6K2wWPnT3v/DeFtPisF9hHlnpeVcEV8YXLi71EgsYG187/iyMNwTd4y7V
OEUfqHWc2lK3zifpZtWK0kK0cC0s3uMs0knKhyW9FpOhuVIvuY3diIXVnUnROtDs
HUIvxJT2leTEQrBm/QfBLmlJcCuVJMU8c2qvyxxT0sdGydUtEXchN2gMZmyJ+pHS
Sch1v+d9ZgRw6p3MGbm7KPUlwlLGBCnxi+QuBB2nyW8SUgSK/0CZKKOUlvJMtlgr
CPktwbZ6DINoE2g+bDeovIypKr54VxznNfMJElFeOddvzVCRokfk0qw60MXeYWZ9
4/BqDB11EYsb80s3KzlitJqnAbeIQKCwdEIPBw7IsWV5mppRfjy/8YFumyFGWFPy
Um4n/pwzB6AX18nh+98cDbbFHPXUndHhP+MN4+G/CMM8rAg6A56cmdVm+fOrRihb
HJwJhIEmwRoJh0DiklPsxb88A9HAXIBNfwZr+jloZocw2+SxE3bBnxfhbsN2Mx39
VUB0BD9aDRuMfvn0In/bnlm8Abhs9ErptmEP2qQdzuW8HvcoG8YetTlO77ZqBdfp
5dGaEFf8fQT3WcFxVr3rozf3N4/sD9jgH3m47JHgyZKNR1S59BYqiaJ6k0zvHnvM
GtyfnLzTf//5LQAH5tNpuM05ZyWMoGtRvT91qj+gc/PSw30IFy+y0yiFApeoGIAn
YwuzomuAbPqAZn8Ljjj18xFK/5QktCTyzmJiu56Q+cFO33WrutJ+lNle2hleFI7I
/tm+otMf5n4wCJ/Y2AjBd9wxXauqnWAPMylLsavK6e2qMYfA2PccU2fL5LSt1eJT
MHCXDsh6R7kqZmYuFshrLHwgBk9jHR7490rccdx5vvzFPj8CFH+g74xaMszzGSav
usS8aMJNhYLKwhQMK205sdnBWwaCEakqKSQ3mJ8GQTlbpHFSD2Wik69PhM7xeujg
hV+4ud74MGfAa1EEJk9jPDWoQZDugKyT/QOQfvtKZjll1nEPTHx1qg5GkCwLxevF
EEtAVY0UKjXkHLkiznzdVQgOIkhvsQLyluGwhOVz07232h02adzlVfhu7F71cYVL
+2ufqW7t9qnbB4XrlWJZO/WYLkdi4Rj95DixlhFdoLyGyECwhwv23oTi7JXL9wLS
aAlqFM8jdKUiLIBprtO5lKrWsXYjbzsWUU/MHX8RXaKs+yZQsNKGPtUWLVQWClk+
e1PTFph4pBu3q0PGrxK5/sKiC5tuWQIUQs/loWjM1c4TF8VMdVe3Glkm0mCvIrvw
FdDi3jJxo5x02CmP4HXkemrTh1I+J39fjyi++Ie7HKVLmnTFJK4yCTQx+ivx9VM6
05C99aFjz+wXF1FV12cSCLrHu99cUC/vGk8j0y2qS7dph0r3rkYg2iytfw16Dny1
WJLFnNIp/Sj+jx/eYKZoTKo9M9bMEQJNCp/ARCkngb7U2D/2myn6FO16+dq/SphD
jE0ZBhLEwJ5Bq36ma+A+GeILibcsy9Z77JXNLeAbyirPRZh+ws46gFtav9tObNrr
JySA8AyzNps6FpygIkrLnhZ7LbRrF9E+HBh0BAApKkTzMsfcruk5mucFCJc0FW9W
mFu8oEt3q3YBFb4kpXTJvWJ/B7a2WZxvmmdl3wC4ai/DS04EzZvfxyuMJpjOeHfl
B/1NZ2FCuQXCZM2d0w71TDpQKrXm/hd295oNU05K2Z6bH0SdOIGFqe5JPpYE1FcH
mIANNEcEDsVOTo0DDhR3Hs+YNDp5ogUFqXYaLo43TOYbPkssF40TSjJmnOSYkmxR
Xcyd3TWSIOpF2N1HJElE/sQB18m3GIltXXiXCxeRaPExiX5LxRR5VwPNkqI7biQL
45sQqFZPg8Ot9QECv5OJuLvnVj4WXy1Lcs6c7gl28ji8OSJmhRxu+GgtuYooUgsO
pckO/sXy59Ly+W0gGQJdVRB30jF+Oc3gbHCKlhmhBy45GWspePgdpK2mbSJOS5TX
Jg28GjH1MfVMMlwwzCXAtzUqF/apHX4bjO348fhJDYnRLUehmNh43yMhbnV7nm4t
rZzGIdPtz5E3csgOr3FNWxc8hRXmU4zEGYv9Sn3jz40iqWtvLb50Aj3rDKpFpaVb
VZy67Gg+mg2PWwdE82y+UV5OL4rrPx46j1R60G7C7WnIYb14hSSx+an2sBTlrzjO
LsuMkRMpZMsgZ0HYF0b0zXXjcJDIL5alXafWi8Ssr6nzYAtj612YGqqc9b07AZiU
T0y0NqllYLMV0Buv852PbmGmAIN9NwfzmpgCtjI3uU+hH/ZprEVrWtp0IH75Mq8F
JpDKFym+TJ6E1YfqjxprJj8rTo7MHgcoEiatBNX0KLlDswozMv2eiT7jtS5V+Vi+
yLD13KXw4+675G7sSRXdRi1TtIg80A3KX47K2pCFtI0A9q7V6vnqW91nE7sXK/7k
1gmusaWz8SEsdm4x6WCn3sjhdh5L+r6xf7ArnWzhTOMyHSIKPs1Bn91WJwbKqiGm
Ie+Uir3WU1aDztppVhDDmDeh5RoLUR6motbyvte2BGwb4CTFQHVlkLzsyKbqzRUR
wMOWvxsf4/wP6shMQg+EW8I0od08o2CT+A9Y0/KumP8n/NurY/YceDc5S0vJ+GlI
Z3ykeQZUgeLKyWTOARHV5fQih0x+eBDgWlscbX6OmPL7ALS1A3AZAbx/7Vg7niAA
4yXqB12LedXtR6joAQ9KoQECA18IYBtFII1SvrQ9dbt3L/L8wfDTQokQcaPsNvQR
g4l7XmhrPXBPmFIPrGdHinmsDiLjwjABTh/o+S6ZggEyJ/rygq7lvld6nvIeNjQm
JN/8WYlch3vWVqIHP5dJOlyRfc7Ohbk+V6fBFB4ZSGboz/cD/NbRsBFDHOtsEG+H
P2YAV1Di4F1qSi3t7N5RBm99bm1VfUXwrYMMuaO7wy00PkK/sD4n6VGdBbkjraZ3
IrC302QSX+zK/4ctzCnLstpSeIpMQRWamzL7sjyEZt1zn74A/V3plhyBUiKx6Eu2
ez+9B8hlzDpF+3ZbBop5qxdzwwkKLPALgP6vceTkfEXBER0J912SkNl1d1x2zZWz
iDeeNsJ82xSEK4N9kJ1nRasZ7v0ynhBME+lgBf/67yPfpq0uMGbe/GJjfLC6/3DW
uF2HBzg5j7ISZBLFptmSrNaJi/Ujhppu0heA47FM8YLbQy6lBZ4pWpZr/cFVnGuG
YTKVbEuWGEqWKqGrXxzBQOtn+hgZlBr1/Q8rk8FWYEpygKqb+D7I1UjqiE8CpDpH
QCqoBnxthMO5SVufJZQeQ6uDmDYntQzI9uAsPdJHd1Tdf51dvzncVePnYSLSAtah
4QRfNdrFyzcIwEGOIvuNMvJAcZHXP51V0PawljTaFzJJdibxc0CSA/k6FP2J7PuE
UdIn7qu1aeiCJmfHIvHBiooOgGQ1U+UNMi6rMpU+gXZJhp/YAJ2quDF+d3PWIlhq
B4KGPb+nJiqBFAZmhCBGGmMVR4C3KjSeFvSC22jpQjYm6nZ2djFLgoDUbpcB5QOq
5keDtGzhMsk7UMpZhOyqClJBDYyDDIRYX8ENHSXtKSSnlTk0sE1EtDRzQKCtqicV
sxWVwrIBUNnRIuqVajHD6X3crUoNK7WGtP5aBgMgiJpXfnU+xmlCupufOoqw36Qb
WQuVMuvay9RMZy1Tp1HgoMtQtUIik21yIsI2UI8HdXt+gozCfJLD47I6+aNiaN1d
kN0znVKo6xAn/uN9+gGBPGmLVFE9Axy4I/9jqfiFrusXT5KLbDIuWb96xIrdmTug
p5LNOnpwI68xbWzyDiv/GEzagz5yIhbG0caoLGybKn7Zw9MHcS5i82YHTHDQevzS
1fHgn0qYJgpqm17KAZb18mWXViRx1S3Y1qVSX1ynXd2YoKQZxwEnG+aCexl2tncY
wKICUS3f9yd5oYZ261MAN9xNge2zaTICFNig+iHkY/1RkGn7GgxFNR0u/jLRuIF7
C/wdTjHVZ9QwkC5djvqsGzJl4qIS66C5GcXGZuiNRp7Utvsy9QE8ZKOt4IgseFSb
ltmJc1l99vcw6TxQ4cdkC1XVgQ+grfi1lBi9NRpANEQdOBYLtA7gRbiAMbCG9jNn
o6rzOOIpPjCFTkHlLks0IbB6QMBKOSrVu7EaTFWRxbbZnH+cMomh/meKEfrRckn2
cDgYhCs8wTiR5vOgXiC/r8Uj+q1spbK8PjgcND1goz2e6dtzaUHFXwvfZlBItXZ1
trburERblxFvX4E/LYm5Z+cx5EMvNm8KUCiFWzOnPz6R7WYe0w2Q85HUNZQvNFRB
4FBgMpDoY8I8ptc6zWmKAnoiGmgOSSJ7MCg73dnuktsOAg8AT1BMswVgciZNHNXO
lIOVFnxxU9+92yOC6PTulALaxpNwJ6Omrg9/gRpU4COIufgh9ARGPq86L00SEKJD
5DeMhj40UKPzaGLASJwd9xsOibrxLFvWHvd1sPWVfncD74fHbtmWsmxV04RQrgk6
X78TSXNbb4M2gwogKoktQCTLeCODGsLTeIV88psBPBS9H5p9lGwflYjNC1OJQ+Y/
ucbdOxI9dAi25uOCyIw3kFyY8GZ3LuJRUO6xlg8/Jdll7SEo6vttAVNj6I3RCIso
qqE3Dz4ige3Nyuq1I/Y7t5mLlHh5r/oaRKOq179Ef0WYNwBT14mAZJtYSWJgbZhs
z3DcPc53aq8X9Vks6hxKaI8SQhuqMMaykpiQTHIDTODHfKl+SyVjNg1vJnxfM9sW
n7oALRZiuCeNhxn5uEOKrtyWR+65tXka1AgCirTlG6MwVM5ixbE511HG+gMheKPi
EN/5p5KPj+0by3/xkgbQs1L2JYJEzZvd6a81AxTQRbUaYtK/+gS59LMCYt8Ioemq
VgyZjId8NmH5sUZ8HhE7lsYuRkKPRpGZAFpsuAvdyyT38R5CpzSNS4L4ToqmvnW0
XQ7xkDeSv0vOKlQFxU8OTaQzAge2MFCqk1CmFc/OLrsSHRrCQgeks9iSQxwCe3z4
s46V81QwKUobwrpcx3TYTREcF6vqVi0qF9ijJz/uI8ZFejqM5BiSxFhvU/6hknrs
FRnL6qLm7KuWHysZgKwr4v8VlW8gArKkMZRuf7BAby8FjMHPCrh3xgjC5mDjACa+
H+lbQP2eyTzNk/SRkGeInyEWzgufOdFnA3rBbPDsLB09zCQBCgTui3asYjowPwOB
8qzSAbqt74Al3FUi7CQyvv9FNkAQLj34YZVF6KICwJO6Kio3PBpeShYgy53nJsjh
sog36mP2C+zsjuEcrI4BYr7bA+mkcIvB/EEUaxlbqXGdLU+lQQeDJp93e2RXJRtT
rvQplpp8ESjFcTC2ZHQnN3wwvqYjiGFbFKlHUZErQh7FZXqBEusRbUGe4GHGAr32
f23kmI3gF+0sltgwkqRQXmP9yc4nsxDdus0vwS8lKMsgNPSJreCSiiFjJjJZqyxp
e+u7c1eIXpL2WDwgYCrk2/K489F4wNvyGUNL4MDT5XrESGA3GoBJKuYbTFWLcj1K
BfCsJqeIvdA/uUwinWbd6e0Rf3UDQf4mcKJ5qKi5QxknbsnKtAJWYeHEWp5PYpnU
NW5lNRCapLWXYesDmffB/FD0NFjF1ya1hC6ld/6ziUHjU+Ni0sBMW/56l13DG3xQ
O325hJAzibWgYk4P+N0MO57dTZZiYgDfJZJWcgNJjjjtlKNv0sPzq1ajdJ3JdhSU
CCEWd4JRs0r7gosGVDsNAmAOC/3Dci7Afr/Jn9DQdXL1Ai7t71P8XGx2e7ybRKbF
0qGobHkEWGJatVsSjlsrVBjs7rgbyyD1zNAuvg3zeLbbljgo2GreCESpnhhIPFN8
DBflR60rYJlt87XPaOo8J0OAWJjD5BxutVIR0MCqd+c1bfM1ZsvPV2Ht01PTKVbI
EPyLIsBj//TRl9IyXbXKT+8aRw5p9kjK0uEP9QW1Y9nZUy3yqiI+JQ7fBer1DiTH
cDhQiz81cscq9osE0SG6K1PoFaZnxx3SgZmc7/cjOfouW9UZ7N3fUIjjeHhwjqY/
smr8UIwKc/4dxBpO2I4zjc++jdop534RCctsvoY4lAoQpqytfDF1ajOdcwkQKKKZ
xuHghIyOT2Au9KrBXGv2D63qHP5+UNvH8ffd1GxLGziY1uUsYxMX7XkZ8bSQz27l
rlnqeatwRVv2mmV56SD4UU4vJ/9pQg3atYVr+CEjrfqcu1LELV+984aayr5ZQZPK
mcXNgmv1ogK1lMKu8dlgmX2yESGnb16AwGRSQr8xaZWFqL0E/aeSx0lWWfr84FAN
hGj9+4xlAgoJd0E8qxGlbCO6k+P4duZlqG80sdJkHUlSlxiyg2QK9VUy1LcwkyP2
1SB34Z7y3HCode0OcnbByGezJAMEdDXbFt8qCIkU96l4M9OdGIKn/ZmUuH6R1tbK
EVTPKdMYa9O3dr13uFPngNqvIfH+nJE+ZaO39TiXg4du4zfT6xJpSqXAJKTjC4Bf
TnLIKsuv6b/4YLfC0NHRA7gND1rzaJ9MYvSfUFpFg9W5R/0nFQuJqxOQ6aTNvLN7
RzCASlgf8rSjqvkOF96TY2jMZPGS49xDnFTCB8pMz8BSKvZZ6/taXV+qjoX54PS/
xdyVLBQc+Z+XqTziXSCGYqD9627iPu7KcmXjO6wg0gFCYpO4Ln7v1l8qbnmz+GYT
7XrbkGRGvsVLm/3NVKnDIPbQa0tTRMGqsE/0ed3rdsJl5lgHvSV5g8hRn8j6vfuw
NZsCADgJu1eAKTjMa1woB3u84bvQ7YWL6ITF+lncrSo3f1VPSI6giLmWMhr3CSmZ
7MNgAjFxIFMwL7/vLedGWnqBWQW/cWnOIdXUZE5GBhxBRGdO3wMw3qskZq8qfQBz
62kAvv0NBJy9VDAXfzjkM27UMSmsoPppuul3qufnbkhbhluC45Y6cAkDadgdYpys
dQ/CLmYPg1QY3j0w6dZlXjt9CHU9C+drPSVVCjgUKZLYRhqYl8Qg0nuduIDXzmW5
JEjt2ahrFOaC1xAiiEOMXiE1uLyefDyT3lBGvmD5lhW3M4TaEH7THw2FNZEqujIa
VJFdN9fDLWEWkjh6mv+3wFt4LuehnaTTggVcZyMaIAZQL86ZCQt+CpEeVSLI4Hmp
Cc6vH6g10HwySl+I9rnK3ZAf2aI+cDJNZhVttnfBRO5KMAHmw0SpNnJwryeE0xCX
Ov147Y2U0U+uKcc7feMWIydLOudNm0qFFbeT/+DPYe+1zYhkNBlOA8kRvdZiHsV/
lb7SvXgKFMzdkXUCCSnNpMU+3t0gq8F0i52ppBzuA2/UgWEE2NQwfXx8olbK9dLR
6ltxJZWf0bWkQueFCb6wbfGtws2MAC994GJhiS8eBWCxMWBZzcrR7s2Y8QnkkW1U
PRuIwZSSbQWvr8sHv77QoVkNuwQ8LqTlEwg7NUaCgDXJCPcMR6jufHl9eEQTrsaC
LUG/JL9QrCtVEt471ndTXDpdoX3vWJX2jOVorQE5LRyjoh8D2qlyUMruxYBQ6KUX
xU0JilPe31B3ZT3f8CfyeJ+BTNfcz1alCMjkKx5axd0i2Dywkb74VbX3SXCwKcTl
rBIdqQgiOnPRSjvHDksRpNIsi0uYjlgQ+XbfNs76Dk2WZ43GC+1uLNYWEgXciJ/f
lNdYQiFxMr51Fwbt+ILzIBdek/z5BDAmK2YMWRoGE4oOz7XTc/w4GNTdRK12hKxI
63GVLIOrHzBVsto+cJD3wrteEK2YNTncaA+oLH+9RbAKpBlph9txKEXmXwoU8WKt
hZUslQeu9cBjO5TMWQBtZIE6jAPVZxupItf6M7Td0ODIQM4d5q5DDOeRWIhalnb/
+Q4822Y/B22YbvvaAuUcjwtS+T7CugSGmk1rPKJj6JalYb+Iv71HqScLn5bzXdPr
fN5dIvUMfsOGgCHe0Y0A+IedGJPJ++yqJRopudfG9MeHG/h0v0lSI28UJNZ0ImTy
wGt9mZXCfa458uiI6z45AJK/WQ4vup1qeHIiLC83nyq0I1CdQMZTjs9skj0MHxpN
rXknVIv8xmCWWBuYrF+mappnU587c8njbX3P9BC9qevFWZXgVx/up6cG1PHYntsP
3uAIgEm29SCkCQ1RXSmGAYfsJizYfiYtx1c6DbCrjMm4IptMME2aq9u/dyboIlq0
RDHd7b3H0qaaBx6lAntlTLXY1UjCfZWOWFkCKfVDIXA8+LlIk9u4EM5rSseASYXT
5Oelg4tfOOEIXilKQU3PdinhST9ZvmPPjixkuwcyaY2ySwIf+px9WD0nSc6+JrAi
aGAijd5ZQnyMLP0FhOQ4c4X9GXxjgqmU3dPnYrS8jg64+UQuTKU8R07trEUuHi4l
9G8e25Jb4uYU99BQIcqjAIzPW3OT7MEYeqgd8gzalNqyLv4ceSNp3NZLT85VuJTS
7yEAGo3nQdpL3aLZoCw9jfqUZnT0AQxZAGk0BrwA6cEzosySYUSnImN7O7vtr6Ib
dIusPyWXG6b9RDYD8tMCdcgG2B2DZSSz8Bnv9PXx1Pr1AdJ6Ey/oHVawCORSh1EX
ItBzYfXPNAPRoAI9L6p7UYTwpsnir0I/HpVTfunez2Mny0nsmRJuKCyaob3+0/le
8akDt2+UJ3iFj4Hh2QPctlUA8DCxsZunEQQKVPVLOwwsdGFs9alxUUCcLmn3sdAJ
J3Aek4qr5D/QvMXZxbh4iKzbuzPR86R9cb1aQjajiS2DoWFMKpO7p/IELDAmlVqx
BEWG+7tV2qIfebZFt3mjl29EO7kjyE7jv2bF6b+rFAQkUY8vKa1FL4jRqQ/71kPH
+sN5QnWDzkUA3kkkVVHAb15Nhc4/evdyAQ9bpe1dm0IRJU1fSXNh5CSipgCb5n8a
mVkIjp/ytfv92SUyxpe0ZuaVzOgqJ0ykKjkSRYx6J/Tkqv6jBNF8ygMJJjpktMDv
/sLFX+VaA+cRmb6RpqnaPzSyEztIzCUBkzT/3ytetrsn0VmcUS8x+4JyHi7o0Lyk
0RtvrVttFkeeb4hwznWWwXcqeuFHnOmXgffZi/BGhLmead2Q+LnRiVJYnXqktuRk
RGyXjYoLKVY8zKGvH0TUMlVfqbVBxjb1ceydyhCWQgezaNTE9KpqbFezKxMiZ1A0
tM16GUHZDhcOhDooXJ8Lsjo76ACbheprsIW1Yy3A8e4TcTrfAnZVKnYW7HHfqxSW
R8llXIDZTmhxGeSq2IlRkhlkGubTMXM+Ca14elXmVjQZVGHfA77zhT+CjF+VHzr1
JNgy3LeWYZ9MdMuqHQuESBzqN5AzhTBjV6/vkyOf95kEWneTrFomFBW57RdKXbpN
5ljUkDHhPsTtovzB5SgUDCTyZFWWhiBwpYfxEfYy0yFAmfWzz9MCZRQsR3lE3DYx
pN/nNAgg5qhlUYHawLiZMD2VURxgJnYqNp6IuMT33bSgKIYD/jGkKNDTHZBpNOfU
Z/v9FwMJilBL8pBUJtaP3CbwCZzWkATDzxV5KuCXvfVozp1JFw3l3U0P2i2N5rLT
UbN5S9D4fH+N9zs0j/Q1G1UGlcnaaDm+C67g+QiiFhYi1Kvfc9vrqioKjgnAkb27
UfOJBA86SlkqQlhAXxDiPGHJyBPdNG+Yhx/JT+44QL7saexC8BjzryEbylxwCy+R
naBf67zqDPrnyamgAj3i/V/XhJWFKcxrZtc31lyb8OPanIykoBQji3Jeuoumg6va
nCzVuWDKX4uONwuO9Cjg9+DPi3hnI+0bUS+hr1mBzXKoBesaFGNpOuoOSHI2kPWK
tMWTmSIw+8IAXLXcyH1V036mTKhJq2n/7LrJont391/TSAmgneQqgv+Qew9w1UFe
yjTRPfRKLfmdTJfIzKnNOAhGwjVw0phFCbMluEEp/ffTTFZxWkKRcmBYOznmYzn/
/yP1UnXTs94wKIVOb1om6hHTkgfMb/Wj9CWCCD/EjJrTFvj5laEaZHDRMyJbV0i2
eMI8SQRwzdfEzNiifAaEeZ8UZNeCFJloBbiGNlwZePmGEWVlRRvnJiSa916o6e6m
UEilULlr+jdmW7j7qNie8hPzQ25MvMxGnY6freNhdp9/dDBIg2CZchFjG691DIZd
l0pKdTNR0Iqyv2P7P97I2RdAf6lNpublbui50HqoIQjsZnT4/aNVBnelpg72Bamv
tn8qRfZ42ht6PK4nqtgrzqaRFzeuvhWA+Of+Hp3tzJAZrINXbMy9Cy1YuysrDoln
HUblHHURbs4efRqjRrkeIDtPB0S2NJa1IIaDYR3qKMZvaepnQkVXHoLtjd7G6iPQ
sM9VkLZuavVYZJ3NFlQPWLZIHT+Np+vZNjjYFfpMDcC0zaU4xSgaFJgHRSzE2RXi
baZIhgQzgklII675A3PQMbOp1ASrOfr3NLUBgfnC9nvE44QOXOUViImqc/WM6OsH
tCzOjMDgQAQ4GEZ2R23EO55BG34YLU2xQywt8p2mGxEKQxUhewieaCFlkTZWDF7v
etgJQ6BdOpebfSgFhqJBd1s/+USESuKj4MKWlz7p1b4C4P6dtmlK6/etrxENIYuY
wZLbjq/jW2C6GboG8HgibQAmt7PHDXkch6T43R4HIKwGJ6T9LqRMkl4Z7RCpVKfq
AF7A4C2ehwdCmvHONMaY1cyEqlK9PEmMTNJ+jNzK/2qo7Mv27R4CgpomMKiiIsbo
dh50DwP5/aDqEKVM3bTZrl1w8hXPX2zwg4W+75k0S1j+JrTMleInOtU1N7zjQMAf
2hPgjdHfcai4JGxz/Fchk7B5PxsulinuhQYpbiW3dg7a4nK8QakrqjlLXVqq58+e
kcjKNZIbr9eDjA64HpD3QWyBj8lljAvqWTQ7GDX3VeCtTBAQlY/yZu9pleiMGHoM
imgqobdMjeYelO0huKKpVMsNZ2Exsdy8TeBIElNwyY9sfaAWIBU0lpcdeclmLgP1
D4g3RN5OgLvwIvovCCRxN/IICAPfakYyfSiAVUGTmRjbZT2V0bBHeIqybjXU5+eX
tHZZIykmiFxrLAU0SqvMmWyYOpoYferA8wDgPdBN47A6uoY70xWpMkKAtoQZ2fCX
nGDimjSfVljC9CbNIEK9buG9stFxWuq+ogtNjSE7FZb4wVaix4qXNUoFGTBileRE
DiWE3OW7IZ8zoTWuqryhAgvXpEN/+01dk8DL9kyEN9+tuUzIgJb5nZX12g58bFFU
miZYUs3GdBemuQA03h0O7CddQRa5QL2jo/rqvHV1VjE08vpHBIhsVVAs+hvAoWCf
i+lc1VZIL4jWkAyScj23MAkv4e1mJnV9Qo+j3kdkjNgvFDQNEH+VlnuQt2TaBWRL
77C1ysdoXTvLsPmAcnzkIbQp+v8j0OXhPvqDpbnmRsPyzWVafijuSd7C2FQVghGe
H90pmc+Cmx4SBP+T3csDWhD0kxFz7l2B7ZzTQiK+sSW4/QTz8a3wAj0aEARNmjSo
fU0+wxbsbdO54LgzKn/iJpUZ/qGZE30P2TmkyEvaXxPGSltMkjkOuf+tshmS0bZ0
3Q9RF5/bOd3iS0ogERIKe1+OmwANaiV6z9lBsYUEj18Vq1yc4/W7xAlqhNisaWb3
LsRlMARHtmziYy4e2ALf/YNX0u+KcIqwuwMlacdeoKi9L0EyRhSlAOnHuvfuVHt6
vtfbSQ8Alm6Ht0gORUFFPt98bAQGboyYLHayBKU+9XMGddcmin54QwvRxv3V4Zsa
y1HKPG09AzbmsXeCyybTKJ0ziAvDOBZ3JKysZMvXvS2mos4xgFK/jnfFkiaN+hA1
LrlCVUUJjjVMLo9HBKuHqp6LfKTJZF39/TO8S10fCIF6cqpOW3HgzILCcpHIA8+I
xLZQJ2ov5xxzo0Iv2TU/PBJTieEvM4RwQ5H7iMdZivH0FhGul1Ytudi7XIz8OTsn
KitO/gXzHHwxESEeAuWRoe+TZreoBwyXP1KEDeiCyiEWPUbazEojrBToey9hOsOv
+T08tCuJrTmCsNdhGHjATGeEjRWQwusOht5MJ5k1cZYEALCZAcI9dVErX7nR/1ZD
CUETwmnNLo6/8kuEpFmveL4MuZCUXrEZZMapfIp0Kby8aYBid/RcuD2srZSqV8CU
tDfYqOe6tYGV+h09OOuOEiEohSkS2IetFI4TNZoCpVSDZPKhyaOd5x6TMgMc3pcz
2SruJj6e/2M/lKeBhHlt0q8JeT/5dSAv1dzU4pa4R/XZDNpoVpa36JwNEgY68w1u
kD4V3s+TnM3pO3btzbrmQjGgwGZUqMnDbCoNnuotKro3POUNFs0HrjugKZGx3Jse
i9Z4bxCVCBp3/Y4ItU8na/58zxZvHroQDFg3zx/2EWp2yapnX3cgXutE2seR8NXj
HHvyq3pJSHmmdkUP1JCVgr8aZDHwxScDCUSEcYjQd7NJv6OpnmbtCu8LBxm73Iqg
/7+LccT8tfaGa6ynWfjM8wKcQHucIGxUs1Ez80nfCrajQcJ2oURCyr5xPhZNkP3A
+rIYi/w63Y5+vFuOR83Gpv6vY4/fKzcARsNIw2YQzTc1unYyxqNzrDFwsAJV+uWC
EsIrlMwl7Sj/NcjoUVDEwuJu+ttE5/ln3+4eUEhJyRsAAXylTdkI1QLi2k/tc5eR
VADOxRRgquxqaSIPlMmTZDdQSuMOo0WS39BLF0+eSj+rxl4ZFzxx7Jxk8goy3LC2
sxK8gEWS6aDjvmhRRUbqY1YailSWVpH5ZiNmR9Q3TBeUK8KY57d0Rc/Mjw29jo4q
++SN4cVB7qNXlA9IOcleZuyS53pSsSltR7XOmpMjs0BOg+DaBBCFg+11LeFMPTw5
oRxom2GeGwTMVaBGg2/LiO05ZLqKCt8Axm7ZTeliBitZ/mCAJywcUcV3RQLE96Bv
R5QD4lOBv964LIelq27ggJxEtLqtCFcVM26jpUFPEbga7x6gbAmTBuLT8dBH40BJ
XvYGMip07PahTdf3xHx6ZWxFE0ETA7hkY/SIqxiFnykNWFp8I56Zn1LkAz96rrUb
86EVLo/HieNYiNgaXDMjiynzXRkpzcr77Xy5eKizzyavWUvcc4o/XYnz0ohnwJoE
t68tpyT2rM6OcEI5eMxgilkjgbmZxdfBR3he5G9+LGjqGklJuIfhfiDSy2YaBF8h
uTs5G0I6jRWe74donzeXpvyYRB/6hZitvh482vyOzweOKLJC9VAxDEYEVODnVBJO
qEFjsteLFDTYcv3uDQFo+jHmFl8I+CtYL0SN6/b8YGRPLYrFgvBjfmewpwELN1ah
wPs/M8zb23wfZ9+TK+LEKj3nvlYRy3sipteBTVfH3mZv8fl20rodeE29YnxgrHPk
WiOCG1G0xnGF/gOQwjVPEM0RIziUv4Y01EXk/dvEKgRDF2zaOYQhDU55MPLRdfzP
MY5/ACrldsq5AeT/natzMJojXgUmzlYiQYrBI5uLdHRyo3vf/7EnBCEtRr71ybsc
Ea0+9na0AHBcbGel3LWw9iQSGfwPVSSRZs+UOOYit3BJI1K5whbfq6uOqH1SqM2c
NRI92c7fzXMfCsUpl23Q6O+oTgcR9rnW9Px7oQQ++vGqPbtmT17AhiOMIothXzIb
7QPzuMZCVPyIlF8IvfME8K9NNTC0kNI8qDTXjybZ5Ux8bCUhpjlZEwR9KSkzbmYb
XAfwGB0MysubALzULHvNQf9wewqtWbPZoD+0TJAP616HZA8K1msVqeDxyOXC5dSz
lA/kABVtz8gPeEVuw1TMbdSg9+SBjlMaYYDtvu6ULNoq/3cEkVMxt9C9+m/8kI3i
gCpSe40CedRMbcv0x/4DmglY6LGp3IvGkoFHBniTQi+SiEofOlVVszWChrt9k4Qy
+20Ao5VGwbeLe7MNerse9nksa0RUh1m9xZlKrth+kuEwezj5IeNMc06jbX3LBlzx
4BD49xxHOaPzozNnZREbXwyRto5J2f5XFRiXGdV9/kz8Thzr6twQ27EJR8afs3zx
f1PVEHnxzDem07p9GUHjIdI7DoPZ5ck22VTjnz9CprWiKWg2PUA2kMof5DqbKqbi
/FQcZtX3KRYJXojGnfTd+OfafkBK/7lJU+RGTE9n7alwx/T2tvy8Unu7xJqt51K6
FbUWO4P0eBC9Sado/624cDtTNN5Z16DKWMAdaYFKPB5sHO734FLv3rnb6qDtUtTc
neJ5r7iwL91cGXa/GDgFecz0gZFpcpqWUmMSbrn68t6+ETL9rokqYbL347F8QL4X
pdmwU6BdBUvUqoQS606k0J6fnpQiL5IrGNyiRHNBLywqPMGbfJ9NOKRGMk2HC35d
e4ZNBsDQ5XuYB+x/lFLCQwWKUSNjs4Zysn6kXtAT/dxeN5o7Gh9LlB/hzPidGFRE
oDE9y+zIPAoN2BAyYUJZtaZPrwdcrtvxkNs/fqJ556aH2dWY51wHyMpw20yfgUZz
C3MblzDMWXmJZzyYv8oVSrXudpSB+XJE824Fl3FcYbS2gJquRO680tJAQGQRtogy
NVon5kid7mL116pnxDp+DFjx+T8S/DpQoxmQ+mRqUGSb5+2A7epZWTTQl0Hf5ZBO
L2cpHLnnx+5OoAKIWQu0zV51grGM4/4gWtKgKnjmTGxv6tQjG8c3GSWjg0IEaLbQ
UKKpHmoFJ0Wfg8il1G86XMPrGXUBOMrsXTfFezlSfIQttxNxYtunEI7CaE3XV3d6
eAHzCwm1jGNZBZhXz+Vr4EkrMtUNI1/JQmq8zlLVtD7UyCEIWHH9hA7vvon03NSp
1bQId4UXsQbzb0UYDULppWRGtqsbTlgLhBiuQvwPTGJnYd5t7DDBRONHjd4tC6X9
qDI1YHYKFYBz725UtkWqYG93QxmNgqBnK+EuXGBf5Yb5reaGyjkgmksf7O/si57J
QPwGN9pB1njXiVBMSZ7zJ4YFuZyjX4jnr7hVYbgGmWYrOTFjmAAN4ceIoX0EW1/A
gSsZc6bfxazj1JkKJ51yX9+0wxfxqmg5L0X0YtFOPGpkr205rRxPUjg5v/dOk3QV
Sd+yKxjFSJ+2JcPw5SeuHj10DF5MxEoRYjYjshFJf+ak58WO2kgnsk5yPxb6uebg
iK/xgImeYtKcBFeEVaF0rR97lv6QqfG/dic14Z1L51ppVDY83AuCCt/STc+HWKCX
Tjdyj580XOhmps2/Csdi9E1gZSVq9Qq26PZvzjNxCDA5M8QdH2+fbtnwvLJKy+Zc
hLYeBT/JDilX87IFQ+Bydh5UXtI9FDCLbROmBZkeWusOCGelqxw3faYWcrWj4FVW
yYaeejGfRQNQwl4pzQhLuS1jusiM+5GLhtbudBNfNwhAUbrvWu3hGhHSaDSyEHWk
HBbGBdPqYx4plaM4OujUnWrKxcfynvN/5SIpFD83UMMn5YK6auOHZRb4VOOjFyS0
NJRvfgB+IShLuenTODS67p8h0lZznddyrxOdRxJ5Htew6BpmEkaQGa4n7U6u0pFp
RwbdyN3DYTVXe1WT8k2Zl2LW+fktiJgvTyliUuYvMoGRgUTp2nmn0q4/Pogv6za9
IebjYiW9MIUuZvZhXVGjyD7I+AkdjbWycV6UVSpF7h3o4rpvsKbVOMIlbuiAPt2p
qfGjXnJvYIVb3Gt3oMvLbvumwpUBVQ96Px/kU2JcYkEzxRFFHXuNyME9h2WUqqap
rQgRsHrR8zzyvn5Am9N77W3T85GLcXZck1twV/uR0T5tK7gtsCHUapHZSmDfd6Ro
6IPo8foDUqD1oYJp8ZCNfhsaWqxiGbSEnbBR4nZQ0/QeCh7vpPQmXAdsI3SbyN+F
d2JoJW5kghkVPsNdRZ2F4dEJl8/WxDlhhAkOgSf+byLBIIUJ/yj/n6+WKiHQfez2
cW3HRDesN+lAJaJwIidHj2bT1zX7v1VE3Z1YVAiDdMJwi9+vbdbHImf3f9ZTgQO9
UwKT708h/wdVEuA7k7z6Mo/MUUsC4hIxdbp2s9ZQNBqSgSNswU7aOCccwW7nMCOg
pm27E3YoHYx8bQfEj6SCGrYVRpaFC9p2rYDxWm/kQExf6MKCDn+gljpzRX4eVxL3
XDF3tgCtFIlNZRcmLnjB2mN5W57JKN38FyKfF8KVO3EryiKBMptoRGmhoKTQwTjB
daDVLlc5L1oEqFnxF2+SpOa8M2AAzB4JZqkueZBtog/6NNzXu1ILfzdHDSf/AOr+
vV7nOEHv9gH0WR9IohNWgRgCuxa608Pbw1mDWxjNx8haB/eiF9jYTGa9Vmklvzfo
vc3DK4HQJQur1NegXZ4q/CD0jp+x6oLW7jZ1lD3VGs0v4HM4wMFCHuza3+nsUA6X
J3g6jWvityo80FN94VSJPEaVigOTRrJkGZdvx3ifsaxyZ4fZcL+OTXPVkGhi6hSK
z2NbSAl9ZAK5WfVfrE8SJtbpZIrOve5KmCWitIWlF1tpEWYbiUjbMPFqKSkd6Sbt
3/egD74I1oGX+WmY9WDdx3RFvwWLettUUAi9zdaXTHYX2yh9ITQuHZMtbMPfnqEf
xEyNR94QjDyCZ7aWB2/x81etXC6OA9FFrNRN0yGUD/kGXHjllf6B5CdSwGPkdh53
8im498nKIQPu9avweqqkExyEPD2p06zOJjzsEUZrZwylBOn1XBMHww2LBV4/2/sh
CpLgFTXtLtEu/1vP11mNG5pxBT/po/T3YJNkaYC1V2o+fjpWvJlXXkBnMgXQU+kw
cRxr0qRdcj6qbidhBf2gu3kKvZmpkKDso50/cKsfujvVqTfn9MpcBoHuA3qrYmBg
vFM0ccK8wCIEvk0J6kkiT+4XvmrubWV2nu1Vl0NTfstnHcWw+5HCAEKHXX6Mz9zK
hihfB5KO/cF0rBLhvJW0qTCuGkakpoEraqxzOb9G1Nx6G6Mj/WmFVKTGpE+TaGAO
91LZOLsXLOYxwgqt0LQwNJrB9nWdsmM2/QhxI4qaHXq6fULThOliX08qNfAJ+VOY
PyWLqoHOhsfvR1jeHQn/HRQR537lsZ/6679GgBx0Baq4NwzB1D1x9CMH7zbZn4CK
ap8XKTLL7qswT/mXqBYweFJrFPquHVl0bKeBkMdZagBHJTEQnGxqBA8PqPF942rU
Qb7+iGFq58IOXctQEIF+gU3QBFM+zzLSWYAXJ/QtXS6+2VNjiCFR6dU4P11clh33
ArscsGrf8NjlMVi6HpzwXCAmQew3A7mRH6mYiu72qQ18iFPVC56bWBrUUczDZRX4
fwQHSPanEzwZR1QaFNxohQx4qsRriYo3J1zUmeF5GgOIr6REPL/7rTEZBLPQUnAv
Ki2H4Mub7/34x9B6kNoNhFp2m4YeX3TiXga7qGozcEla+VUcbF4fPeqaeOepuJxY
lS5gzEg8VY1VY666fco7J6vUGY5FDSnSJUbuphMAhlAvB2ZWGJpTzs+QIL5KFH0l
SdS8WDFSJvLmjrI2bcrMHp5ZNxbd9odPTIgNronhaIg1hYiY2nSygqkT1ADIZeMu
Wuw20GYh0qBqt30NvAVjUoj8SFnCzONmlFEKa6MpSboD3RjSwefUksmnhF5e1J9V
jwCHjXCQbB/K9bmxESvAY8o57WtVAoUDOrx20s6gUNP/z3qgk4A9iPKAbTNxzuI6
hLNbJ33VsPDErnoO6FoXBZz2PbwZnAkOK4q1i3GGf7gvyfO2fKE2VslaD5Mhaoxv
pRlZ3tadVwfGJSyb5p7XbzpTtJ/qMUdErWMP0Y6xqeBsu6Kk9lg5kvUK0419Vqn/
h/q8CCnG527P8bslNzOnhZ4I+HVLIX0f+G0ma0GWwmbQNYgDj/Fazn4VBQ8MCyca
wK4N7rXhE7GhTe+Vgqdrrl1lyvRhgkjDy/NH1IOIRCN/2FldmHkwNlLKEY4fydCJ
36FRE5bGxkhSuNnSG76krE43a1Woi0PTTPA4tPY0URk8fiNuuRNpd1PmsK5/m8Am
TUtyCMUAEjyaz1R4AqwX47dRL83a+E5CitGoKB/RPTFS3coRevey64hz5RKdhO5K
qzYQbCAJt989IAo8QGBWlnR4sDcu/A0mXFX1Dthiog2ylPlYyc6cDvHFr75ZsLgf
7D7M46uh1FdSX0L81i13tbXr7Gri4LmSQNcn4Y1E+xLS16WhmBToRbBkpygJn2/+
yeEUuroy6eKta24v4NPeaUKdF/gq/j522oX/GDKuwDCEVHINZzEFPyNXvyK8We9F
cmJJFo+ZlboSLhdyLZgDpPMeP+0j5x3LuGoWuJ6fFUwGcn1mE7F5g8Wk6AySy+Ip
k8NuxACVspzPCouZIYEyTNNAl3kwx91lQ4h+LvnbUyegxzoIGBF4qTsXob7o7B05
5ichPUfhdQV/34o9C7e9SDvAo/QQUrlbE0MKNLeJEtzZgFnKgBi7lPNOax6EnyQf
+s9lwyNXPy4x6HaGwKkssXiUhWuwKYfW5pbQCN5xhC2Jb0jwgJnYd+ei0a75IiC5
uz/BJ02O3c8wZKb3YM9ct+OULv0+svMeovrJpXnntuc3UKvxpK0XsCcP5Ne7fxyC
q80q2ojICi7U4GpJLjK170qU78kA7s+a5gVl59Mh+CkwTTbEgjEKgK7WzGR8uvjI
dbDxqRMiLxjpQMhOcjxP5qOa4GgXYDD8faYficnILLukHvwZ7XfvHYTQCrbKlTBm
lmqm4/KRXXJge1xcHYFmMOCzgQE5kSs0X1R1GBD2wgqJyXDk9nh4TlzK0S7JHdhE
wFXUovOWWa596z3zXEZnE3xSO+kpI2uEAUrKlSZ2UMqUPicxgd9ei0CaAhPjHXm9
qEms3AN5/wXWt5DDQO/CPJ9uIRTo4K5yGhKE7TD3cIAu0LgiN3h7UHs7W4PbABN4
+BsX70ZW37Z9N6pi1VtWN1TyDm+VwXqrdKJ/Af6NiT0Et6CSRdCmZGdJfnbkG1B1
Hop9cuS3IaTveXjakVlBZ+CCwfppJjcpFbO6pWRB1WsnjLw1sAQy5Z0sXx/GtDSm
fgElyW55SMS0XYBEAvE4kS4BkMcxpoUNGJDDedY7Q30kUzAUFprV3UZbvBpKVBRp
0Y+UcX02Kl004WGWm2AS9ELMh00VNLwzZ5F0SUQ8NW9tGq3atJvOgfyjTw0GnCcL
R0vJc8xxA9VuEx1kqDPVHd5b7ELaWIWTiNLf6/hcbfoIUHCz/fqO36POhbZAZQvj
8CeN8KXqkiMTkBt8/e+j4cPBpLLUbWIp12Bqy+3G/XmPR3GD3cI3L0G7exDb1utA
GxNFxGJSb4/ogSiBSOx6hgWecw6s3XXTLNenVQWmCPqkfLvuQW+tLOgGAi1pnt0K
zfJPyQKm9gXuj1px8yMKkF+k22LNA47+VTHPFY7YmDiRjAyP+5g7Kq86c48yfU45
1A+l1G8k8LjcaVsG80J+VJ9WZN1skzLURlDfpmE4Rkl+5NjS/dhpL8jbspugTC2K
OslVj/Knjkx1MUjB/LIBplOhQ1qs3Dr7t3PxvNYVhM87nsvsKlHAJ/FqEv8faCnH
piWxmuG5RwuxZfsjVaicDVAXGHLPzMKXivQT6nuRU63U+vGjZ8J8DWa8qu0a5P3V
qPv9THscndsAYtvuDU9i+AJFgwBlt41Cxcye9TfK15VprNQ/OB1KySbm/Mu5sDza
o7QqHyaKzTNTEsaDrCc/EhaZ35YAQIom+MTssE2S39psla2ku/r4PiAe8tSyY4IH
8dKqlpIBGOeb+5vx3aqKRvuE2Cj7qJXeR6WiFGOo9dPVCP4tff6gsOGQwWWe80qQ
zbpSo2IevyBNVOhh3OeZJ8ufYoyB3J/v4xCvtINMCqvr0NRAFYjGotSRNgc9WiSU
zYnc6iCn+/Uacpg5Z0m2VmvOvi4gXd63+XkaccnypSoLlwlbe8AoMzmish8Msomr
n2PvAf0oMjiwRYzCk2t6ulsY3q60mY2GyMkNOG58DokRaW5IrBFyvju9jCeKhBpz
L8aeFZlqT6YFckK3U4aqwJph0A1fKr5WKbmgZAPO33T1HrESfCn1f5pX8Qsx6a9G
AKSN/7+97tXgUT3u+TEIGZWGi76rpC4Au3QA7aOUoi72BCieTn3b6QqMIUSAwp7l
17oT0+ETOQ81LQhGthCPsTtaWYtM256gbX34ituhd2kKqL31LCFr62sIeCT4EBRA
qxCFS/rVan0amgIEh/V8H3kTwaF2VVIeB3y//JRY0e8M6WQ410ueCeLLGLk9bAkv
U0uoAAFRZAV7bW8yaixQgZGmrmEkjB8M60UlOvsgX66p3Wz/t1gJtQj7MY2Lkjio
vAJyAymv2qKW5L93B6+ljM3rsUsnw2fHQrCVddoSZ5PnpSDSbRnwFfr9Yd7aZhSp
3Tywf0a8JffwlVC3mNJNS7XRU3oFuZsel3zk/GIxgimWfvwMAzEt6GhxI3ymTrSf
dL0ek6pqKg4YIeR04VpY2f+VrwKP3XCuOqnRRy752cV0BkhjhoIqKDBUEsh4m5XT
3K4t8eA8MsbAet22vC6//Zk+lPIzI+Xp23hJzsbWGReRLj2ldtaofokWJbGms4t2
66p29S+aXJQLIVGLJmRzQNWCunpZVLQU11ysQtSK7jcL+WimJR5/NCEaDK8He4Z6
/FJFJi8c4KoNdNiVIyRrREle1ccN8pazpo542HBjMMhnqMNFdKINJKYX4pfHFzv1
42Du59sRhisak2xuZPKb+/F7zkxqxn+hK3jtAdZ/+uRdOfRsRNPWwN1UQUZ8Mfis
Fz3daZR8N9gzijGrOgnq9emdIGQxvB/OWHEwtD6WubrsMFEtpP0BxK4y4vxLxNTF
pq1xWhMAuzVhW4THvuj5oJo4tZehttrUwvAXO1ptO2lEMxabMuNg2eslC4nU/2WN
F/ZMqGSXK40eIZGQ6qLfhKgJ9M1pBBUL/kuJirrLO2zAf0xEsFaeVkS2jMDoA3WG
ikBMCCVVKgiP4aBPpNbLkyKuFsgXGE3xktVxfzitdUsYaUUqqfU6TnKWXB73rje0
Nk8SkBzlMoSzlOoEoMJVL7zbnYaSNRVIv/0EN082dHIMv1qBajB3A0F+kTo/1ZAq
GN9UzxLk8arF/WXCLJbCoAUkcmfv+vSfViVvYcmYH/CrtY29qQEqx140R0jsENOW
aeZVrmCgHtsLd7uozt2UPZ1YOG7oES3N5rVIGnXEke95DvX2FGjdVmqVWK7kSe8D
C07HsolJblWLS1bu8jKJ7hzQ7GsbPRjWFTxvTziYh7ouyDz6lTXkP6Xwbsj+0Keq
y2d4+R8ePFtgcrCJ7G2kmKlOBYKz2rjXAgYYDNdApjq4VD5s++AInUH+mwN++dh5
bxyt6PYEcpIfma0ue3LXZXCFYR/HZnOaloCEcTmOMwTYE/d+reUTX4EucwHsMbeX
aHPsw08nqo0mYfjcOHdnQTQ7uNcTQ5i4VN3FXA5nvXqD8sZ8jF4JwfFVhSwc/+cd
0R0QNwCZpEPDF73DfD91nCYJyBsEV1wTb/hWuXV2R/tzrsHlY/oBjEJ6lEUzW+Hd
GtT4OAx0SIaGPlAeOCrmUQQFHNnhRepcVLQhUNWlJvuoiZ2vEfbMJmaKtE0nT8gp
zzmWWeGLVy04xLUAk013zrI7YOQ/qMe/ASdJ+lzunhi8LqUK1HcjCuLdKuqYvPr2
Dq5yi6sLc0QChbF7NvI/K8OAnl9LhnHziq3qhz9lkwiecjVt/8NiiVtu/eO3zm39
Thl8WsEiP/hMtOGUR6ULrdMdlV8++Lqdst5ZCKntnMqBGUeQ0+LYc8vU2VwAbr1a
df2aeYlGJTlMQzVnQONE5EfZnz3WT0ra8ZdDrVIww6wPTGgAfSsAMwo/tnGuW55B
3Qlrh3ifblNiAixUDj6dP+8Dl47uTKI1YGNO6eqmE1Zd7RvqbVa9x83fXI0k0slm
jdt7mw6GJxolpDlydBij7y4whBElTJutteok814inFOpGrMtvcri6R5YH8GDlntA
e8mzm5HAvlCEFVP4O/JMgcHqut2+Dnq5vOUwL5+dYmRIQH/8h64IM9YS4C7nvzWk
d7mY9YSu/PZOq7a3MXnQnpYVA3hxhuOWsSemwwn0mtqwusOKOVFaChlXHK8g9tps
aQ0xkd2W2HBBnCceDkpJSUWBPWSr7mj784WLoMcmBdOnxhYkcP6FcSiELOsJH77B
Neo3a7Hy+QoCA9jX9LuIzeLZmKheuifDL/0Zuxr85XK9FZnRQeHNDOs87njsERVl
Sm/A+ydD7GuC0YMQJPoUN6n/uWvLUHPUJ0R2ZBUxAaX12ngNVDNknXobv25hRhbj
9bTnBEfnu9AJ8iU6nFV5s2DeE3XFg9q7k39UTS8aAunt5VGrhwRWmk56SE8UtZ3v
N5J2ESO/eEBzqX3B/r81dMdnBjCZjkt2emwCtSSgmAfQkZPKR+WD1Kw5HJUCtX6q
vaJ1uxll22iWIvX/VvUSVzXKYdE/2oWAsDzMrAvszQQ9iH2mlNSVPBFBXjJh/23T
YQ/osru6IS9ze5icUfMjsxzQqWyBVbtMiH0eqJF/j4WYsuf7UTwW5sxD37OXmkZc
IgF7d2U2n+O6T9koFh7uP01W5uaeAhk9TVUe+3v1AtZfczSS0HMbi+eljzkKMUbT
ji8c0TQdl7HuIYlswJqhla0huqN7DBSKYGyZtJJ8GgsKzeRO5sF+cbx80k/A+8bK
eLgkFJdp6IITqTopP33eQ+/5xZAP5wAT219YBxf584b2zn3K3L5anMryG+iToTvj
79oMeeDiXGZa5Esf8MSmAvn26TWqU0jpVmjYuhb4wUzj12HQvEHlLTi/6Vx2LTyX
7YmgITOHoMY/xBIv9N763HO1MtnyADu02fPtxV9kUpFt/Xa7sIV4F+BytogWbDss
IHIIgwhCrrV/CJiVE3EcM3CWqtTovl2vrJlfJJ00wfLdAqec9Ko9M55CaUaVWRvY
DyCvE/sjQeDYDkTgRVra4457JslvI9IxKnNSCYB4lH5XY1CN9Lhv+OtsL836vlH0
NbFmNBR0wl0w2XzajwrKOGDw8QbkqJwbGKLFnlut+irMA/AzUuUoBpq2msKmN8o1
/TyrMv+J/jjwQr+4OGA4cGI7NLqqCm1MfNVeT86mczp7oLCYIR/UqGCviOruibOS
tVU8ek6vAUhEa7FjsD/o9mxRCTf+bWuuWdpNf0HnxrN8b0nFxK9YxG7spKVsb0x3
slzMMbbtbuSYHqRgHZwFYVLeW9TbD1hK06do1Otnt96N2vWBXsE1Q1jEXqkgsm1+
GVte48QkMhcDnM3IqiKxejbvy8WzyjLg7a2o3W1s1pQtIVJNH13QQ12f1SR3cH+V
v2WgdCxoHwP3bTPs5l5fTJdEjZwd9ydxBlER2PgMUe9wCWNSkl1qMDIvodTGSV++
wcAtlLwdGqUoaIL9mOPFVxOS/AihrzIOIuOd/JPU/Ripnwr3Tilch+vd4jV+xnLZ
bgA1zmoIOlLIVWMbdfUSjzjWbz+nS+rRmVV6iGjHKbS/T3JQ3pr8tKQYG6Mj2mDB
8buOP2F9OLBYGKYksjWEW1M8YgKFPXgiUQq5A9OyK3JFcTS5SDGv9VaqFzRzUlaB
Wd75SvciQf60IJtMgkoVgvcrH9nI4/gDzGnpg7w1YCeS+mGwKwkDPQu8TX9in5lY
jHeHIUzq/4bRg3AS0K3ULpw3ORWxAIcSfFOxdasFBbouiWLUpc4XWB3YDFSXwNVj
nhvk65kcsoEHtsc60sEuPYkAIyl51Ujmbs7xsJZ0pPlTYQZhp/CDeZ8BiU8ieY4z
XONyaIJMqgpiHNC7DVX8FhoD+1GLbHOBBDcZfdk7bxz0Y5nl9N6/AHwHRahiMVc3
rUug8iTvan5+5eTntEDPmGfKOnGW7jMPGRmlKTSQuAW1RoPXcXgOi21fSVYTPPvo
5wF/EOZaVGnHSTfGPBvPaiVryMdz4ALDg7eWchojyiw0GfTesRJstfvuxWzynhTb
GrgzlTXzXcxYmEsJbKpA+tU30sUvhr8MG+YJKz+zluyWgHdw2jeqE3n0upb9TdaB
EWcIu1I0HTFKmEUKTd8+P1OJq/qJLBwqTCY92Y6rSO1KXoONre6zcpQKp7VHOL1I
B1Kjnd0FIGzjsfkPNmq0TTPZrQBjr23Gxtg3B0a/7c99zjA44Z0t8vQ92HzoTpBJ
BNVJJ9VtZ8wT2shUYlDTuMyXrjpbw9gNSb09tEDJrTIgf6v7yxIbAl0w8X6mXV76
BsI2tjlACcwtHZHSi1tgLU8zeYM+rM1hikOXf1U1GR2aSekqnihdLjmt875mv9uQ
Sqhp74IESFwRKpRD9+dY00q+JyFlN+8mqc66SDorYp9oWbtYJqxBVXwXpjQHRcne
ipQEyB3redn4Hz5A7jbMCIAIQc6TDZl3/pGI/wVhafuK0jNupEgqAxtivFK+Xv8n
o90jmSOfBEuKVJ+cbWeoFm7zZ9tD8g5hHEw9rkcRBobfXoq6Vus/F5LXjH9pWZd5
Rdz8KI4bxKlLSt1Db9uNqckwHUvLnNiJ3vUMAq3v1XT2dRWltG/FVWkRlapY3a/m
3Lgaj/h4WRFOvgSXPygsTS0Walzo5ZUV9VgOQJ6PeXBjpJHNElYbp+0iBTL5nl9y
nBx8G/Y34IuN7DArRrtu4At0XGT7IO2YpLmrDLdBknedCmePvYzVXK+ES5RiuOnJ
Dn5gHUUKSW2UZyfuQXRs/Fg3dHKLMugt+4knbRI/3yBd82iI6evMzBAP3UAFXadv
Hww4Twcbc0+1+D5ijT1XViZbM18EEhHlcJdtIRabHUuvxkojfp1ioTHtFIx0uM1k
PwxMGBFhp4jk/jIl/E3EP4L7ccNubyTol3HxzQ3P/MVOQwgQyZoI7IUdRjY2tYnV
GhTypBnYFuhEZZdaLxSvq4GMN7tZnxmulFnl6AZMrMwG6gb02/WLEfg3XiIv/+XG
fCPaZwMji9SI7cg+4ZXyy+FP8RzgFtQrhxrPqGPzoL/JmhTbgdhauZxfIwRFwbek
g7m+VuFTxVrDo9ryimOWMUB70jw4WmSJySS0AH5z+u1iXF6tHKGOOb7tzLcB5NXS
kfYHxQeD1T7rDc57oVN7wbX6OnZ5LoCSpRP7MLmN5fkoq4BVdJU/nRRHbLUw6xQ4
skjlqXT0Ax7y6gTdHvOXJC92I3IgIsc8IE8LIh2MkC3qounUFxnQgqVJ0zlDySLE
ySxk+bjFKJyYe4IeSgbJBzUpG3/fRP6pvZLP9VE6o/MeHn+zuIzv+Sw48woW8nKf
0UZW8rs926VgJvZBNw+QxCAZ1+2N4ZphfyrV0Lj81xYs8Xh7i+y0+q2XQr4vuXbt
VBxMui3hXeUiC9hVi2vrveDqKal5/nizkeQKrbbDESRuK3PsTiv3ZQJYgayRhUiY
Aw3Xd1GjVdzPDrH11IdSvsh8VHwtiLolwEgCXazdweKVeTinXp8gxRlEy7wOWb99
6Z4J1na2jMFUdKAOmhZSs+I3Er2y+X1eYOHT3HoYI16lqcl4h7epmG4amnO75vSx
3zuWOI5zHgT3zLkUvck6FLrMC5K3oEqTvRh9nqNfUSMl8GmjbltV9NrVHiKW4paJ
z6s9sjipiGWiqBNJHoE1uYOYlCFlrOmQnyoE1eI1mONbuykQcDL+7B3Gxi0d0QcX
RAolsVDRwnIAIKZAt9ucVRv5iXlEEvZOTka+jE3UCQ52gWlTQlAmt5cziJQFIsuN
rUCLme6Boc4WlvOfVzV5Tj71NrKWgtGAN0GNO0yBTZu7Xu7c9/uClXmaSC5IVLG3
avpOyHmKRw8OkGwnsP7cIlt5bLkHu4Ppa9aNoWpO3wZi9vXwm+zwl+hp5hKULZfy
CEiu6ZgQ2HWrbkFox1MslO6e26/X38/cxe7PtRZZmiHcy+comLJ4vF9TNJzFEKoF
XEev46aQu3sI4mtuUYsG6WPmloPURxXq64nkCQgS0agK98Ae/AopnL4I1Aw/KthE
j2MEPnhPy9v5FYhom0Wz+pfrSsWIlVShku0M2H1bx0vss005GyuHr7pvDYXf/G5X
RpsMrf/EfMRhGnZJlONU5fb+rI8I4jeHZoZ4gBQKEYR4h40vUl2Enhe7ltvxGlDW
MEcEhi0caJsaHAqQQhKbRRUsUjgrt4lqm9ohXY/OT7vk/WYRy7JQYwbUMWmNaBLQ
7eloihf2ZOu1wObdOz5WZNs76E+bIS3HKJSs7dwa+8pgB6cFp1SktGgngqwBJV57
wLBQ2rguhjRKQRiA/InmXmoFOJWrMqUIFQOjOSESugPnUGUUC5syn79y1aDQxL5F
ZYarsDF1/GOhs6gn5N8SyNF/zPk7id45VpLdrLjPoznbPCVqdtjbAngbTInbbXL6
stPXYuTV4+XXzFjsYBrjDHZ9CbLTunaFXRmUo/CFI0k/K/6bhfqQEo3l54wf0vO9
5fjqEFMZ7rQU64it/Xh9NuJR8qVqFeUhn899EVCu4TdKlUNmDlCPc7qTQ2ET97+y
XdT8eUufF8daVJRhedp/tFr18rQLHugKlm8JIsVE2EuTrol3P4rS4IC/zUi8HnFJ
qWFWOcchWCaqZgycf/pKwA71nW4eKUeNRNwEsfolC2zWicZgZ4M2y/WLOEmuHxOW
6e5SO4q+5NeAWiwZD1XNt2QianuR2uH7ern7R7G1O7TCpGFBoTcT4jmrf+xvuYUn
zU14JWuLz7L7Ty2u9v5Z1n6c6SJwd4eJu+jn/kq2XxxuVeIFQEkPepmyzVBN+JLs
6p5Ty+YKVQAZT7wQH1GFwPDkXix/QvW4tE2klEPsRBjqEBRDdnHshp+HndRbcYg+
G+MQxbCheYH9JYnOqebcdQBCi2Xeq2LBdv5Y/rwt/BH0YH9+hVzJIbgA0gHYzhnh
duAsFA2Ea4GkY5dKKyS+SN8SmDRFKBLM2GPJtkaraa4mLZ9CsIsRPcJN0Lc6wHAd
wZpZiVuCnnn15lYaTagQnJ+ouOzbi2dJaC1vhGh4nAQCpTnLq3SMxLExfwkuXkYc
fbtDnPRARDSuyjoXzugFGGGK3a8lWg1piFLra2OxlxXGI3/14WjXvL6lVkB58ikp
08rviXw78WGxzgOnXuftjbx92Rbbf3E82m0bZXTQUczjb4COaW3ehJMGes5Ggp7b
388qRB/Ew5piyZSrrzhcBzL3N2j1CIS4NB1QLzZx5OjHSOQhZeavsC609bEH6sWw
Tyl55t4M9N9MOxQPKdb/+jLCvNEw/pzq4nyVmqI0opq6Tdhtkwyqpf54Sybsqp1X
mIEXCf/4rJPH96m8iYbJUoi0HEy5prLqM/BlLdiSCLobfDBfFiqP4yAg72eEzmR9
w9zBMATKY6+Wjr2of7TOXd9xa5EGl9I/LRkxfrF2dCOrhno2rzvgiJoGajcPVBl+
NKE+6VEJJfH2gBlOaUMv4sO6aTvLF6eSCA50c3fyFFfjjlqGRHxy07Epn58aWHSV
q965JJVA8aIAxxO2FgVal5m7461k5DvRwXbaSJx3QdGUeleetiicg9GFyIPOnK+N
YgPoTIJpZkqJVXY0E1K/sfMT0PEV7r0yHGhXokHonJrPofpQJ5zltIs3AA7dienj
WbCh29Dhd0gplz2RiNE/39F53k9OSQG7uEA1Z8KgI62nmc+BHY02+AqcK7Pa5C0+
JBfezJR4aU99GY1a/GpAtuezFS1Cv4/Tz+t4DG8Gx8lNwUG1NKKVOxKOU8gDQ6+m
xL68XgRc18Ky8rpCiXN7LNbMGsPQgV3qAh8kQwSAKOQNhAgGLe31o7FIj60ysDth
/TaJC89TE45bq7yCv2zXm/AZwVZ8h676IY0/Eqa2Zi7HbJpqGpPxJWBS7Ymn8GwS
cDzm8wkTCrFp7UsgZ2QKEuXjlwsUPEumBrVtV3pGMhkkV15e+NvQHrFEsy2blWy/
bfCNOwN4WrxuG/PD3QRAfG5GkZeEDzXnOVxxWuhen6F8FcDZ/YWMlHTqd+Luus0o
r/yyyo/WCgE+JzJ2KuqzIidmiHkbB0zI7WMoJcDu9cTIo+ImShUjrBYZuT/l4mz4
auswq7/0oxJFZ73RoxlqEIia47r84bYkQh+PQgO1HYbfOhkyvqCJfqYpagBLJYfD
RfseDHQbOGAevG61101PcbkUNCgN0qiRsQrKRFJ6HCs9d9BYJisxI36LM9UVI7wd
FGpV6sK9Yuwd0xQvqHPq5ftbKsHhB3cgHKz9XuHMt9GnYpDkwLAQgrrA2Fvy61Q8
4/p7L6RkRnCsKDn3rDEceNbY358cmf10vz+P9/1JOxpP7ej69YRSUnqzcAikJCgv
qNsFiDQ165zer7JvDTLj/NKYWAX1KVUsYEKFbrP4qHRsCuPI49hpdI7IToMQnTLE
/LflZ+77O/OQ1MKd3WhYomQNlJFE2tKr834v+bpVKHwQxX1ORkvc25JMQo58rA6k
FfFzEBu8IekkHAP4viz7M2uTGoLwmDthn5yonHfBGZwvfbisyXkw87BhNRZqQb05
K4YnG1f0FZSEvJmk7pgof0oAjjF9ghiDSZHM4dDaTLC6ihQ4KiCVmEbD3GtQud49
wSnmgPqAUPNVfV9NaSKXBlp4Qv25yPKxvTdgGXQFKbNzKekJm21S3p/XSxCRW1XY
RANIDsMD9xQQ7l6yLfz2YBN3W5AvzIv+oo/2cP4RPBxo0/YEsSJx6Aee/GjHCrYo
7X4NY73WBRHoULK90jO93hjhHsCB54Unn2F5MLF+n5VrZFSQnq6/FEjkVSbxtF32
keURrXCs36MM4GFT1YnWy+iW+qbQfN7/RTdWnNlrslkfoApdO2wqNqTeQj0ORSLz
muLVctVZXBP5G3GLHVwMoXao9/kOXe/Wor1mUoqlY2GyfxerV0WSVM52Pur8UTSd
flQSXF8BAsU8gcKBZOvw6bIGY99IxlZczcLSgYqo4YyfNllWdcmT33TqACjK8ssK
Lr8NDRAFE9JR0sYQNQniRL7al8WNvs+PWW84GA1TDxGqIcDMUiSystbF2L66f6Iz
VkrTuv9Pr63giXFzsLhDxet3O5ftGIZ1uuGxdr0DyP69fm57Rwwrc39RlQgcbkZn
GpzoJs0/83ou5KDlWo/gAvkFJ94223jc1pufIjV81XN3Jp8evrSiXkSl3+EdxPls
4vlRrTR9bu7zuWSQmXcJGBKX3km6I2wFsUjOn/7t3I0lra8my07kEPE7D2YwK2MO
1TmPbPjfoCHqFH12aVflKrZUPLw0PnYljFskdRfNJY8yoAmYNv6/fZWbj2jla6J+
H2mWZnXvdfaVwJQwOObbMKFuPGWgmsaAm/6+kX1fSOdiLmazzJl2XW9cx+j9YCVU
W3SF4fUDsWtVUoyqSvvoF9v+aeJaW7qzn6yrYLtPQdQYDJBIxz7+k+V3FcQDFV57
kJF83rmqeDK7vEUEFw7MVBdQZ8Q3hmAnKZTMrEfdx0ETIjVEDQ1+wgZVE+KOMG9t
klpqDA7Mr6ohwpJd2CoCJbc2XMaL2OgqE9gdi3SwZmDYI8wwbbaXGxd+DhMtYWWi
siP48UgLB+Soo/Xirfugu4FVzEceT+CsugB+NlxZAqMEP0eDdE8dumMplRJV1eUt
+hHYs3d325MlitzVSUbdw3F6T12dhMnoUrqyqgfzGQSWqXSM0EHs+0eKQf8r1NiM
JwJriHjENsEew/B1CifnI6stFhD/wc3kxWp9bdbTnIRkvW/Uk7cZQIInB9B5YdCT
fL8kLWQnTm1E1M3jrtiS11ymj6EhpQfNQSu1E0K4sGeEwUiA8JavV7/M7MPQ8TLB
QTfZjmfEUmyOgaZz9uJRmbZ6gwmjbsCLVxlR5kP4NVPcvNmPbATVOXp/6KITFJl1
toH0+mESx+vV/LekjLsYuJtGmHDC7ffAWkUV/AXCRJwjz9hvFwENhZjC+x1cgAyL
0TMGDq10OxFtvnE+3R/kUzm/Sbr+rVS8bAuF5/Qyzl0Kp3lCkadKviNPhnhnptHH
QwqDwfb6OQx1+y7F+/M43uFIpSX6BLvkaJofF3rQaMPGANXFjHI5Neli7kGNp51y
K1AvIUMYqedvOf9+1aFv8QBXe8XGece6fQBFi6bzm5+1BYl1l8vd/198FIliCvPE
3P0xDreJbOQM+6bSNUYe7Liju4DdcKmQhvashMh5bn6MLfexUn0T9sWCpaYUo+bZ
TtkeCziTPH0MwXU5hve7gZyXIAhzaER6fU4hByP68I4fHuqko/6MWA9YkkNQo5yt
Qvu6DWueia0AXRHqKjuqrTkyK5OMbw/A9acZ69ixqoWIUhN8+pGWtRd7gHxetG5A
fhxzUAIb4FETUdXGHVjPbSab8SDV0bMk6pFfH+Wbhm8PYr0Oqx1qNsUuxqxd47EW
glnrnfK5cj12vdU4hvcFZMb5+tfhKvp9SOmZNN+dYgLxcJ/QAWeKDOXjGylbA7By
vybX3HeZNnj5j1Rx9IZtpYN+8qPVI1YySsFhrAyA05YywvCy3aYnSjP2wDbMKouF
/BTRr9lxDrYOJkFT/GOgOMPhECSyHcs250GYIaPc8TEnv1JnETCwrgrD/dFJY7PI
fRHkAoAyasqiOUU+p6HyHEbGagnrmj6IPsmWxQJ1qlr5y3FpxZWdlarNdIyp4rH/
e45kLEbkdc1B0vzhN4tbuk52W0J0tfnEhFSQY30IbLE0gfNrbf/us9Ub4feE2hFJ
3dYURzDjwgbWhsAZYtki/rd6oy/gw7/takkAwrwuk+ybH/sHByJu1SqZIEr7hy9r
Gi7gneodDW34JLXNZnWuxxaALdYK714AIVhXvKSknGWs9UbopjRLDMtWnyy8b6C1
yYc+r/qP3rRiJUYDE3x4CUWg2513UiApv0RiKwJI3g0v0P+GBdaJAzDgzb0Zv+Cq
MSarYubMk5lzct8LIpeNPlZn3H5GRfOIG8PQmcuudEyXjP5Y3f0Q9YiwSvIQCq4U
U5F688aAS8tXBOaHMTiZ+VQXqYW9J+Xf29ZGa/JmPyVLl365ePz28Z/Sz/UJ/ULu
AeBVKpq9Xxj0utJbWwyOC4kko87H9ZNI+Prl7ERM2QTmly1SzHZ25wUYCJJjcbvR
3BVqW8ahbMQ2Ozlk9EP3Ohxf8bMQujpXy+adrj3OwGQiIQh836hbf56SwbhXeheM
C0uWfdfIdz8NTrR2GfioJ5RWt6aZjj97R9yMfAG+jilWnjpu27Pb7i8kCwkiPpeZ
Zae80FRBpcP4G58lLMKCdOpLnNu6zTvPZe2bdbYeft0PWiR8A5zvNJKD4IfofvxS
pNL2sV9EU0bEpB4dKbMeS/xyYGi+/tT1wUD1UjH3CE4E+9auxCLBOgvWo9MQ8KUb
J/RvDi+l4wmvotCMh9Q0+BA+zFgagxTvbYH/V8wxcEHv0BZa3Z7e2xDa44xzCSwx
LwnQd0kSjpw2rTPCE6TQjOV5HppQ/Y38BkFk8y+qnPJTJLX4uK2xy61/DgVrD0xD
QqHTu8qi7YNXXCKw19BkGHTpfDlqKcsQQ1BbY2+kqwjCpHsJeSOiiIZyywdV1ESF
8wh/wvpNq2TZxQD8YpWeenydUwVnM8olRv4cNj7yLqiMYWUlEl0s8v2RzIiw/s8o
HIpOOWI6FHhhspvyy2kz+NMSp3eRSfMemG/CCQ+8vZYUtR0e0XfYfd9do4rqY5Nh
x1luMgwPe11Mv5gYepnqXGT4zrltLnNK7LFCcEekZsvyFjupV07vX3qCQPRYcE2F
xMbRfPELqlnVsDFoYL31oNP2wL6mhhgll6Bem8OeScmVPzH1VpfINa65nw1a1ttN
GpsahfOVkR+Q992eeQC8PgJiLALt9yT0Gwl6qr8FeibngSKt3iuYflez/LyxyIzi
aGWWiY2vTJU4jQgNUXj0rfD9Jwerj8r5B5Wz7xsutPHk7JQH4ifqKIWxt6Cy+TGN
kcniEpomK3gtyAkC/IdIXhT9krZDMRP2m+TQJBKDSllH+U8AynxKBoXX0Jw3gssv
GYqDf0egSQ9kduCG0+OTKbRAz/oxOfGkuvNjXUU8EnuqdKvXd5+F/RU7ILMw5YN+
iEmdFdNk1hegR+iiukRaatfOm6OQE82SW4vEFNpCl2DTNILhc/dssESIMWqajDg4
WY2TnGPzLs/iVk72qqBW5+V17cLasxaPJjZ52mKaAs/+Be98a+RnjOLM+zHpKbtZ
RPK2xoXwKc7zl3A2pInjgR5ryFGvlR3vjt7S13VPNQgl6MDJv018F4kPc5iXPY6S
h+ezm1Ig89zsb/L1zh8rHXoO2f0qYOdA067EqIpr80UtLTyNi/7Iu7McdHt/y7jR
JdFBreLBLUqE9ibkQ3qEcc3iviTpPTkSfhCU6A/8bUod/Od9769OlUjL6IqDRb2v
klGvvLrQ+SSjrgfv9FWf6SOyL5NtXhFHZjJS/YNjNoTKhCzwfr7/pNrmxs55NT++
RnGAFrO5zcYq7nEtIT4i4tOPpAx9UW5bSEgDY0PG+aEZmlCFR2NuFP1OzutlvgxA
52RZ3r4WVtOGMqXJCpCfL2SH7y+sqPe4AYLjlIGnDb84nyb7vw3vA0XL1bZUMvnw
9W7YdDJiZIZzdv/+aGFhagYuBAUkrJTAK5Uj9H1PXt8Ec8WlRkNNeN8VBanHAPIO
0WsPGt/vSfoXMfc5gYsiBCPHk3ZRW66nQQ/2wgeWeg0a3XsgzL1F3dCY6R7e6iKi
TO4sH3DA/k4JW9YtYOCxEjaSjhVSsj3BPMaFD9ysgMA3gg4FUlkFtNmA2bqHY0Mn
9GWj7yTRXVKqIHPcpxnirwvYAb2qw20AFmTNC8PCQMuipPK3Xv2xEQNRkR2q5NYU
3nWXnZNyuu7taITCbdySQy5Mj86nCmDDyIOPGGM4bUWezVuffbV6ubXivunJZ/J4
8PwFvAaK+F1pzkCUVMSxh20tSCOeRf6f1NxwC6qq6RYJkt3umgW0WJqmu0E7mxn+
S1WT0w3ynZhoiVwwsTRJ9YPiMOWH4TGk6GZ4TjXhTMYacnhaTLheAlv7KQUBP/4j
K8jiQw7vis02o70tS/+xUauH/VWTlb75hJ77ugV6d/EMILCuzEEID4XJfXOVj54U
g/zEyxqUXbca+iCaaHDMbzI5aKohx0lFP7rX6eKdFoZnFWhT/fxVfLJ+L6wXoegp
TLEBo9Je2HINL3wUfP3iSKG2t2H7PogG8UffqEHFd4CwB5t3vtDI9dg9SOUY1+AE
nCik0ohcOFxaZgoL3i8Jbk0iljO57qH/FBBBGJVaR790zPsBUsQRuRkyBjzjePH4
GSxzhAsAhC1TCF5uWdBk0vmCPHGUYq9d5OEZIuQiNU2rO2a50usajzbG+DrgcAT+
YYaTmWk8pKEs9JHnwA2uCj1so0vmzc+HwUxdSzDr1Zsk0maIm/v6dLOkGWivmG82
xZhW6dxnEkRNRvHR4y9Je0Txr3KuiJTGViM5G5/Mpga+6bYhFiKcSnLVnJ3EMOcw
is/fcSWzBgCtrottDM+Q0JJBLxSKC19hNrjf7WUf5AdSLkt2p+IiIjy6FEkVkgYl
nirDgIobXrOTPFaDqrSeX3nhXOT0KvcYQkuHx81723gYwbz+GniW4i29OzZxTPw5
ndggTr8uqwf4CTXdTis9jVMQMWonYYLOaorUV4e4JpN3hnd37csSamcHXby3f+xN
zDy88crhOMrL0Uz3WfYNACUSGG/VyGA0zA5hrkoUHet+xuJCQAzcWzlK4SBxwmHl
ttCP4Qp2roiYXhCz7Zu4DzCNaT/+MQ/J00+T7MHfCuM+1NJDchiNYgTJTqBBJjSd
PDxI0ioFPNzJ0ZUkaptuJBtTGStTHUjswZWKPvtMOc7BI7xX8s6x2P+oV3RaIW80
ANZ0zsuyHU28ukFO+OaLpnnjWql4fOCf8IQGgXtdzVhRtZJyzZlUWl7qbjC7lXnY
k/rfzsoBD3H2V2kOg88B/XmRXD8eERECXJr0siV9u6EzaQDAwV7abtdkdrMe/4vI
wdlPbSELvsZoqAROu2ZBuo17lxHHQ272CkIJ/pHc2VlKl+uTl6wztPDq6FLRvCmW
pw6rdpnrPB3Q0e4JR79D5imRnJY6djBLJZ1CThFaeyxajCuQHgF7SBxXxxPNLqWb
bf1GrjNFIzAIY6nOLq6RiqbKifhydpId0TPpWkf8PWkJKs3nPxA6Oaa5xD0PW3X0
ccN1GOaS2y+TMO5gADYfnoVZOfQRFagTKuxinuFl8cEjt9xGczGYOQZ1vWthLiRM
nyDA/DBVrI4ZoK6V69xYEPouGh7EXIEhxaW2VmirWngelc//+5U1gA6gLkH/FhBk
UdwloHkmRX9z/0FlhzAzwaiDCRzzGY5eSf17L04XwEqLC7aM/KQVr+Tgw55hBa0l
SRMJQRGp/tNLSfYR1gOf3uGU8V/oVvHV74lyXdG/DdNMTJfIKPmufAkANkHRe/Ws
IxfryGYTfct2ABVKfzMqxnfOSWQ0LPFQXMfe38UL/WFFXDciVQTaRn++fIOBXIE5
Iv16/G0WdrUEh7wqdTQm3tlUCeX1v3HBoYu6WUmVXgeTRfwfA2jHK6glOK1JtQhH
k9yip1PsXNuQ7Eq3CvQsvNdYOaMB0ya7Te0w1rvv75vV6l/WLV/97sa1ZVEImEVV
1fmPP/Eu2vzmZV/vu+aEnQcC2bV1cjKBhg9vS4WL9LiR/wYK/VDwnCSwUwKLwb+N
+0OgwVkbt41QlXWG4Rlt0P0BZIoW1nZtSntBhe2VLM3Cb2hu1JXpLsRCRie0Biot
zP9Wkp3IYJS+H+2o4KSmfF/3M0aEYiftHEHwCcR1AQg6HA/z3ci0XYjvFFD/9z0S
qN+Pwq4K7lwFJo0z/R46JwIstY+7oTkJKC+U24icLx150Im8lW+CeKC7dWtx1tYr
B2TndFf6KfZjWXW2Ne97ZOVfEHH1tLegUPzanobw9Q7iYrkIi/dRjNdzpfe8YlgS
HwbppLPYRlcXvT1MBsx6fKkaWCOd5ab5t1LOW2A03YavWWSyC7O0E5qzJRassyP8
h51lGhiAC5MTLYetIZXwHjPHBGmMUF5g1m+Qb+sksE8vukJk8N8WYCqAcZYXvgoS
ndmfmplcw6jvRq/hXID8I/C4YMLX9LUnOYCQAOyRgrUL+hXYCFO9J/Jpt9LPNPoh
aCh1JFXILmnKlyZfhh+p3Xx0OjpGoR3A9IM8I6XTzZXSNcpeEl0PoUv9IoHW3YeG
T7T7Uosn6IvZU4m/ijHNEUt9N34pJjFv0pq6oFR6RmqaIdvE1P5f4HGn8R9aZ0KY
HFEGUhnVNtPvsGOc4igGMzFsXSoilAE0wiin6KyR2pKLkYdcVDNLhckQwdjbmJpX
MvtEdtjr1NS4BXdKQW8jSmcgoMJzJol2IBpti97L6X0NBQJMlxXrWDmZgOnJZsJS
TUprt8C+sAv2gAVt2gh0m+Pb0lx7T9ajJGcMs3vDioir4neFz0mRYHJQJmdWxA2K
8ivUNkGTHFHQlnS+J7kXlQQSKkpnifqEkAPIDlMIm65b0XcPFje2kDanAsaX27XY
xqATZw8jKWWbMejTIUSVahsUjiEsLlL7797obJUAbndP8P53iH7RdyNOm0rjhprH
Dc7QVZwHFH6ZWKWZxqKE3YGNyAoAe2DRa6pDFBz9keKikHylfHk9K7Ryw8Y7aZMr
g4Oc947CiRIBqc8ih22H34L5tj1jRLRBxMSpij11IYQxmATvg3dXm3K9XQtX0bVz
hFXyX0trt0Md2b10tI/Zj5tQTCPKJHQ3Ty7kzO146gg4s7mB5atV8MnCw6VQ+uce
i+TrUYnSoRwuYDMzx0mVbpn57jbR7KsjBI78tDwmCRWeUpK9vuJg85T+Rx6CiuFk
9ytRHNMPepveo5X0tfZ20jTOfcRqESn8vBbk5ryLR83B4FEFdC9aKtsFm5fDN5n0
6V4leZckQvsJPIzpRzO99v6owrcn/Vt6NzCp5fzmrd6fH/dhm4BQBPzcLla/xoin
EXJ0mLLuyJ/IKDfwm4jhcL8FekEJCDLls/h6Zbs44ptDG7Y0OEs106Zf4I41ILBh
gHz7buaC+PDZgdlG3FAy8PA8tR9EhDS9J7BwpB0VYgUoDREd2jSH93eWovPc9MIC
q2qHHW9JoxXfk0UUGrikpenppO5441pH8NAFPTvI+5Y2LcatW9SQGCUr+jZqgOKi
4Z8/ekrgch2DF80gc0EdLPfxHn8qkV7+gGWSNJyyC98bsGzsxDI46NgE9OyzIm6e
qG47VSwOHUuTEi2y6TN+oGeMdckC3+jxxatkSfg3GwpfBp/4aXQlCCjQ1n6iOBDW
4aJ6hl4Hmb9vQwKgcAtm4eu25AxwZxJcwJyIJ+mLPto8DE9wkJmeMwvbP2CyEjPK
7ADNFQV/HigGTOJwJ5FuzR8n2T8FxDJ5H3waPZkhKxcpSM4rT1XXYKTfxRqtflOV
WkfhvinGYevjr9s92Tg/MGWKZaQ7iejpZFVv1c2UgKUCwfMMpiqu6SPnLq4KGtRE
Hic9z/aFgq6RExucOyf4Twzjrs0PIgKfC/F6NZ6hatek8TNnSlxzv1Nnq+afq4X+
pXz4mQFhQ1Emk85zzeRbqAGUTMLtPigDiohPhWc3Ri9LfiTtLiV+sZX6uO+vVsH3
GNZ2/Riz5zc9mCVWnzBfDay1silVZoDV+cmpr2ujYc9QLycfSpnY6wTU7ZYmT19w
TDaIDryK4bz4F97y/oCAwjPevQMFka9fEavRqFZPJhi8f+QcV9d4hURWRSosKtdN
qrvwnyWhsYWO/PZ4kCEkt/iSNYpZIWjuYXE6pBtz50JayJDj7Dg+hCryaM6OsfpZ
F+X7RrrDE6vIAzteV51Go8wggOsxfp43cRpv6+uea55JUOuuNyJPjEPEAlEksEy2
jMmld9Oa6NQ1wPvlJCU+hRm3K1qePIe1GrHkDNzi9bcZ4shfdHf/QQRgOBDdbztv
HeIBspA9XieQcMms/GvLlI3TXYQokn7u8q3CFacSA5BfB5u4c12uTuZx1tsti9dR
5A4RDyy5Uuc9PFH1qjSChwGF5LFvuWXvpkSR0b1SNIM38ENyK/1I0qv5l2xrKrvp
G7K4L1IPBQVPhgVuWcq44aIyymmsYWPHH0ARBBmDaFfafSb+uf/Ii/PxA6ISXtUP
uFbA+qY4YdGZuzAhR0QOL7560iNeKhw9M85SVJ76zfOhelZD13ZQxpvt7Lm4X/eJ
iymPWDQmHbHfWFnvMktOUy60sLnKvHqVDv6XzCK78XnlOkX3hDzd7kYQVQoMqTFX
cKI1N/ADFpCd5xpkgVGd+omPVfn3N6bzZIJ/6hYKVUh1u0VCq6T4AxCpEBDvDdtK
28zSMR3/Cvug8ul5GmfbSQdL1MQxwJm4Xnc1r6hQSJvnw+TIneOYnlHx+BS6P1u7
ltXu4vnioGzhs4ykqRpVYayQh24JdjAHsRRA9GB5UmHflXg6UAWHFZ1FmKnq6S+N
QUQ0MQLEaskB6/yqPF6D9yhikE2ohgM1f81OF09voNTpb4uvvWAVNHLAgMCxLbOo
dz72snBH8qRlz3TtF0aQaUt7aWBt5wgeKvFCgBoD1cRbYDuyX4QK2Zil+59QAp5m
5HV6Ko5vO86BOZXdcoons59cL++LaqO9mWV/vx4yoZoCSlJHiuTNOQx7vs9SZf6p
1N6CnYVi0S45QAXTEt8jzSrZFJQuyp+PQnMfGA0kXp8bNMpOb4JvdzIUXl9i33Tk
tze7iSFvhfBKccZk4QIXnToRccScU9lnuoZIDTwrOqWsmYAVLGQjaJd9lolTqgBI
+rLL/kxwqyaVjxgmq7KTm1ETA5FyxbXDyEyRM7Zt1u5wYa/GfJHgJP+ChyDqAjqI
MFqnOA1qRt2Xaddwz0BsY7t3hvVUtrL+l2bTdSk8G/feADX9V+E/guyc0qTx+PrH
PW6EtwPbisVUdhhY7H80J1919owhD5Rwj35ZMwb1OWHPK6II4QZA9/qoX21b/lNT
IXy35o/RBz2QBcfcpKa1tAD2y+z35Ioi3XaE/apCflV7jjMLNHIDzciD6Y3R0Xxl
0icm8wwgaNkkusxoPtiqXhVlwNY1ikBQ0HyCwfwhZlRAU/uACNvXBkKWmhyZk04Y
Z373+U7LI6VxLSaUtQLdx1+9kM7JSdQHo4kib/D8LfRn49zghHc4zisIrhUoGEJB
xfp5uk8GYPe7KPJC4jINnUTKzCiyXnMQ3VY30bue8YtOzqWxIdxzlzozHjXxw8PB
8Smqlr+Fcc7RWeaTDGzr4JN4D3+tcUHvVY2+2s+RyiQ4e2S096i7O8jsp4y4yXQu
eYNG/o3d9gwfn/aCBu4s/khJGqSc2b2HdNjZ04mRyGUAOh6MC4z7E5XljoZ+ySRi
fyhxmYDGCYQmqtoVXgFdfp1kbbsE9KLvwoAo14JKChJ++V5U6sQOcPdh6bnD5ay+
FzkayoepWCB7AFzxkLEcNFT73+yumdp57T2dr71JAWeANTaIVFz80zJYyxSZdKFm
SCrwee3od+4h5o/ecUrqGznVtcsT6GocgIuZiYl3kK+OvzyM0fKAamty1dzvsvNd
sjUTOduF945f6URmPIlrtHRdjqnBnhsLwna6vX5zu6jPIrsATNbT2ADJUC1BK11V
hVHT0RZ7QPoqR9ty9hXVqvCl5XTaOdMmedrwE6ZWvMqWNA7qK4FwF4aLAZ66MWfN
FFyRZeKjmS52y5H6XDfBR3o59oxJhGVGnhdOn9Htejo9bIaG/r5T/Oe5z9QTFClT
N3KNwMMgNpM/YrqQ4MN5X5ePs7gIAjzBkJsrQ0MvZ/SIpMQ+rnG/0oq4H1M5n5/k
6HwAQa00+rwrpuY85+vcMNKVZl2JKbnNQBC0Sa153SK781HEPM0ZUF+MsxUy2pP7
1Txm5bdwvuWL1tplFPIDhCYKN8knz7b3t3ZxW74g+VEqKMbUK62GuUq2QR8O8oHD
mo4TlyLt02x9d0U5gqTZRfA/4jl/21h9NPQCLDnvsvDGVWuqTSfCaZ5YKSaUWihx
udptMZzMnZRZ0GXKOOB8Qd6Rl8B6s7+Hk0SCGIznFetKR9dNijveMynekoWa4n3F
BVZQ/ISPQ2JFs1Lgmlt+VjsHR6avkuSwu/8zW7vZUuWYzKIlSrXO5e9VF6yUrTPc
8ER/J0bEWFSQ3JSfMIWur97gnZ/hr4glZSHO4j+xJRcCeebd5R3usV7ezuBkvRXC
sl8aTS3V5/1+KfW0NwFNJq0QVDK0TikuE2hOaDjQuates8GVPhcG+z0oh7FzfQk7
q6vRHHC6ny7cMnAlSbpSxE9kk6pK5U1dBbYq5NKN38Nf6ym2ZLlqpzeDhsFq+sAr
lo0G7swMsPNqX2eMIjBDPdInabKhdFLmmH+JrlJsLf76US3i/1ZtEntwfQDrnzDO
ZKT87hGunw5IjSw5oG/Ik3d7H/0SiXevyyumRy48YAJhTzJ8BFRKbiD66NPjzEDs
oIAsLX/D9gr5XGa97Qaq9SYOK7w6daE0PfJ9t+waZ4x927+tiGa+B194aAbc4SZZ
8cbQOMEkf6l1hwb60XoIK322idfdAwzOh2nsK+PlDzPHRu8yQnJNRV2+cZ0p2Zrt
HaeZQBNaYOCr6nzVe+3ukKaEIb7DEnk82tWeYXux/SeezSrmCvhA1vlv4PCieTi1
Dn1WnYwFOq5gg1xitK/KPL0kYEF31eAmmCWHOjoCESGdIFRVjjJADoNe4mHUP/Wv
Nfnh+7jXgtqISNVHCIb90Dxqaw2jpb+kDWXulADxzUoRkV0gumy5wL6PEqNaTsFV
YJLj0mphBd0gmi+3O5+/qB6VHiFc6vpD0Au6Po1EPKchkSGc1EM+lkYQ5DFmRVUz
B3xu9mm0QuR6QjEEGaS/0ZW3A4diwLvh4HaUnPrDMJNkIPVwKUIvGbGIwYH5Prfa
g57Uig4Gx3fepdTLfzL5LQ1qu4PjpsZ9oC6vKG81/qos2aXWgr2dqU/Tl/natJsP
wM7ezCf1ndx+3kLTUWzmYEAUuweGlAcxHqrqUaEDClS46wU2dzajblA09YwXxt0V
cHCsVdRK0jcyXFhULdXFdd0dbW0TadiewMRIS9W4ZylkAAAL/G2AQEVJp+Puib6m
Ss0BZMbCg9RnGxkm/G9Dp09/Mk6lUaOxN66gU5oGAHAcP1bmEx9NRvsSBabJJDHA
eDm0YPcF0oUb5cTlULzO8xc8XE6XOp1+F+qQIU7P02TqEroIEERbg7AyGMROifAN
Bw3L8UWTcfBo28j0nBl66Bzlg7DJhzonBGRda7GfydqrYLVFg2RtPfkRkRUTn68w
Sa0SG0un39eHhSgsrSzYLVb/5BvgK8il+ixiN0vuKVJhOPXLzqsIZ7cmBolhnsXu
u6d3/KjFhK3Cw5kIC58os9Robn2D84qEV3l9Wc3qB5ejrhythWRajTaBFXKP9toB
K8oJMBMqQE90IrGykzVZeJyQrszlRtILA0fEiaSosncH80+0fxQ51yusWyNXTAab
cdx9ituV9iKSNutqZB9Zvp8MNTO1jTBH6yTTRCRNMc0X3tj71MPbgNCJtfSL9lWu
8Fu81RraUK+gZRS+bp6RJgqRNLzWFZxsvKf+3RRnL12wpXnUGsLi3JdvcKaWUXwq
WmE1dq0Fb53HuVb4v305VSpLeiXlyvdWnpREnFi/8qTbWLabpM5lKarw5RwD8NEG
FOWJw93HNWMJHnjKWrRh0NsN5bWR9ylvXCeEtuaqSqAqgh+e4BqOqxTFRr8n1UmR
gwKppKlSb+sHU7Xs7NK2vYt23nomgmtsKaJlJ4lAN+5PS3qBVOFeEJZYcirRPpym
3m4cPOjuE6fFZMtunbT9Q9NlOF2uXDQmN+urN53e4h31SoKDD/vr4uvZaEHbUy37
CUoLrYcTNQAvl3GSMH5xBKH0ErkpI/EqYfD+nyc2Dc14u/+jDS4DVN7GhgcuJAgA
/SXbjGqR2fWsR/AFfAOCQTQm3AqnMSC39G61AAMyXpQVGc6d98AxRp8zwA2Z280o
KQfkDzAKAUIdiheWmaE4i6mKPSJ+fsJb8qII89Up4ITQPhWshB7BHsds6aPGJy4/
6xz4YGSmnXOBwNyGd4MgcmHXLRkLLUbhxaAh6E2hVjgIKIAbe8oBUgut6bzVZWSo
P0cNoxunqOwnC6dmwAB62xR3uRnjBuOK46UvpAAy6JZF3wu4wMhA15ryMfSGYZpP
+1/1Ret4cTn6qQf8YFbPqdbGrle2MDiZ3LWfW4dHhJ9KIUWSx+DBIfRzzs5V2soN
mRZNnApO6bGhWdCavMgC0maLA5ZgioCUenwI90U1rX8YWVC+FqbeU1e47kEK8te3
yfnzN617110xOZcktLDMdVpNZVrCudo1d7obq5k5GGNTgA5IhZvSgGqvrHrJuTsz
0HJ6bRvjFAyYFIl4CmRi+TEncVMre9vPKZ6NwqToU4eFCZdpUfqUKL0Rk6fTh2Dq
X+1ZkEJuMv5ulIg27D2RPi0IsTFL8bcHrXuP58WreAmFDWhR96hEiT3ZyoCSxTxX
7PJanI+LZnDl52c7u+hccacB+ODdSQg74HmoyoiBcpnc27vjZF/5Wi5P/U1uV01w
sP2b/bnpL7vg1dOXbNkNdrMV0quqoA8xAqe270TmqEtpnvXANq0rE5ndpGVCBCFx
pMEyHTd2Mmy7O/psLdZxP05SK8RuikdiHZsn8+VU6SM6lBMS3x4/rYcFGnCDeYDp
orlvh7RGcp7c/j+Fg6RgVOfEhHeLug/6eM5M3OfD3S6PXgicjKFy7/vH/5onRUDI
tbBgeMfiQPJ3lC5JAd7OERhiSrtEL6tq3Af4ZoSncxqATueFe97S4MnNQhWwjm5W
VqWFf/u/h1cm9Et7ahY6uUIBrOWCRFLxSYvgyCxaJE1LDU+GZNREvLSuyKG3bEsl
o2As9BenfPSycq4Qz6KWuM+PSRaLkwQ/+duU4CXb088LozjhvYpJGY42rVm7SQzR
rk4atBIoT1ExtXyIcSKZCypvl3R83j1f94MN4SWVVMmHifjMHoV9awkxgTCw0myQ
J2JTDgsRyCZtQeRgrgsb0g+heYtLHw1xVWyymQ4QUBcU4ExaN7LMoCHVKvIjouJi
6MgxGIG4DRhVMOay8Ycrg0B0v/0gb8WwaoTDN5LMIKKe3WT1ALi/gAVBs9AOW9U6
jZw+ztwjJsnXFy+gxHLcWCVWKXH2UHjUHyVdPebrFPV36E4gNM4qTFkR2FS130qF
VUZPmW/SE/0w/24ir048PYTdOEeOLcCORR1rz9m1zH3Yoo7zyzsHIfFhvbmwldYB
DLvR7U/4qeM9fMCF0oeiUxEQ+d//0OPY0MWDCHj58mccNOzAUCWQLzxfelrhtJYl
NaPHUYb7ymGf1ogdcd/yZTAGu6Xtwdh08WSBF2eFLt1Js8oFHgzJ2AsFEipdrykR
gsEHzkhZPONz1pZdiCOwGV4PRWDM+Fpnhuy+kZJJrBcUf9owWjdyOeUyJtcKWP9l
4lJqWt5tGyIr978qIZ8so8be+0ttxdIeytSMWMsMFrzlVfr5AJXurT2Uqr7tkDfM
R+tWPFBR85y0FR58OTgtxHgq7lsbSEGDqhSyIHEDV9FQM6fLFNCY9ehOQ9UsL0p9
DenNnAp6ipebKrHB7YEdWvoMtk6KYdzOUrddG8Pb7oWwPO9peq2JGWVu9vYazXYD
1xzQcA+19zPtI4YdOw82VjqFqJg7rY7F9AGJADvsPosg4XnfoePe5ETwVQpSQOBB
yE5p/y7cHliNE3/Fz64g3mH/XCVc7PQojePFO1Hu4D6TFJmlOGFlAjdyig2Z4uIR
mqeJDAIiI1vv2MlBp8etWIw6x4y+S0pGB1vaRYiEQADhMlHSbdqgENfeJnvDUyl9
YfepPrPmYfAtp10mturL4Ue554pVS2+nZhjkHUgTaCthHG0TrWYxqkG90UNvWj6i
xNdMEIZiNrPoYV7laUB7bN/L/TJCHl1XnsepHBpZn2NfvxG3uk/1KUsNbJdk/N74
qLa11EJ8IZMD4yubATxA1/BTSB/35WF0gBAxCmpXmdnDRjqYqnR4HY2Lk5zNAlqB
qblnlzQyGd5WZIPgEoTLp/ZghhMQiN16H6fjiSO4biADEhS8BTZCikoVegCyaFrG
PJPHjL+cokUc1ScQzYUgIXfTkDc8fpA51G1z+dSSmXEcUqO1af6Z6DktaO0pW1qU
LdWPyhf7yUQFRFzFAklTRDGR4kKr8D1HBpCgj8ON55ZA3pNlgfsP5aQ2/pIfkdl5
rU35OjQZmzdn4Z3OTbMOkn4zZw+WyhO/8JzN1adzgW6lAectghklWXRrhVr+OUwC
yilSGQwn+5/YAmGU77YPSmTw/Fq3yGJvG3CYamaqxbJVa5WVkc7qUbVBOFFvz1KQ
k0v8J9jBjwH94VmGldt3WqRqFgb7JxK/1LkrhewDMXLAq4+Ve9LUKRqZZUvAL86/
C7SF3nODuf6LNOlkFuoi0vZuQIrM1qo32XqNmH2Xz1tYZMzxpIIY6CLE6tqzCoth
HcpiF9dDYIOCjM4rf8utPVUyikLRRmZ+q9gUI3rbJF/fNNc2AahEboSUUJoxjjKf
BURCMJZozWVXU35u9W0DDPzAOFM5njhJqqNi4KbJT3JsNhGEILeEzW5NcJXEf/bJ
2cFodzduZQidA8g1LEADllIvYZOKPCV1zilq4FCtaQ8wfj/kIjj8NZmELdbvDDdo
iIHL/jsSahriE/OfXF7/KWPPXCykGCsBMqvnh4gtH/xjL8VU2IPrDoHhRYgRf5qv
R9sbRGehPZBx4oBzRBONwe8BpozeIhiaRmtTPasvynceFVp27GS4DLYtGP6HTcKO
8T4zSKHnTk0NsN/91CYwvg2QO7+wTG2LwhDdXV9BhshaA2XvPFcGouk00roNnFxy
OA3xD9wfGAdNyxpvRiC7XJG1H9gWIJ7uQEI7/1NCpaL36TSu/nwIzaYc6Zvv4+ae
vf9bErWOmthVqWKOZuH9vN3Jc8QICCVplWVlOSPk45dZ5vhFN/+CCgxOLapXIYmo
GjTTj+9NpCwWBKS+8LMY+5HuMWBj4SKI7LEgyQMfU47u3VmxD5930RRfDjkkgpq7
kDLYrDvGj/UctRaIOthq0vqfOtSk0B1D+SbbEwKJopknIWouGB11lb2e++9AjdIR
O7JYvRF2HV/4MzSy2lGgzc1rQkkVTM4ufDZghq0AFKf2Cp71z9nUJbAa4jQw+BBD
ZUPWcYCzoxcSZ4qE8E4WjOtmyqmZD6NdiGUBPYKGUCXmJijvNnckdGLlwk3sqVKj
0KEIucSoktrm0CRQwDOZXYqk/DhMBkRPIF2FDXKU7KEejjat5CICprRSWVRp5CJY
7ie5OYOlr6MpvRS3hwGnl3ea+8vAJ1IkdeGQaw95cTgYLmSLFvwyP+hZy6O4QNF0
iLo9CJ5YqFee0SAg/oCBKLyoO/tQKjlHmocClSN8qxHnfRXZWQPeXjzCodazMLt3
0UXlbdN4SIMcDpn17RW+5GmpZ10uajT3dyf8NO8zYXdGQ6LsN4ln6tMvxlBA4hTC
5cjmFPxRoW65QlRTi9Q6y9bYQDM60zQeLe34fzxxGHDPjVDMrs9X/z297BLmDcOf
EqJ0V5VPpynVoyU6wmQaTgubiPxYO7mw9jz+lkc+U23Dm3YRaytp4jr6hI1Z9Aee
UpV15dWlJeJ60bNMR4A/7mjsu0WNaubGxklKOctzMHQxyMq5JXCb6J/tur4VzcL4
159tCCs+WbZnfRbA4IVBwzLubG6LRvFYAmw8p2kJ+k5ugiku6w6Ths8ldyCxe+m2
E+cu64j7eFhF9dKRnqytoeLN8lK9Lj1OGer6Wx3cWXxp3BIh3Q6FU+DF1qPLXP/p
k184cgA770K7vwPH5pOK57sO1Kb869CTC7MrXmePaWZkNGCYv7akoEV4vfHOCV46
hJQ+ogruaYb22uZ5UDkFA78wNrImAoOYOKnCQYlnMcgafWMAHA0eHzQZ3yWux9RF
QyeDv4xOiloROVDdnmuvPc+2lkeCShdHxITNj1J+ZnW0lvTaZc5Di7mDRoo+JCOS
VtKbIYktICHJW0kXms2kXqAb0085tXNkw2trm2rcREsSVC7lfS237YvWqyPU7QCq
5w8VAJXuPos9r0+S0aFHBb5Fbbo50+LL/7mIE6T48snwdHM9eh5zkP0E4FveKYGk
hGSImYPw/wASshEPi7vCWDxlk48vMUqajzf3oBs2vSRc6q8dvKEGn7qJa5SxWUzz
sVOIQ7MzJcnL/3W6JR2nehlkUCFa8vMcbr8By2/LeB8qdMbo2jOfC/YQDm1YuR0T
8by3FFmpW5gGZu5dqXsjwCRI+6PARyUWhtX8/IEzO8S8wrxJK7/ZAhTsSo6o9068
fG77FS1T1cGZvhGzh1OJVhFTgxhO9ciQQAJMF1w/MwwTyzkf0YGqQxUuNPmTHHsB
QC12Qk19lutPqu3m6yrIfIjVfTCQ1QdOkMOgpUyZPX43mp92p9iOxpg2JX3PCrPd
iV4b2PjU5Dd2cfrRf0fDBYPlEoeOPqmxJHlONijPGs906ls8sqCEXoSb6hnfsxwj
y9fmjh2XIx6kFXwV/ZtTF+1ZkgPWIh1WpvpOOp/xqHogC5zrE9b0H0AAaAtfvlFq
tCgB2J7mBMthSYSEX9ZxqKkPxcHI0nA+ormGNiT/Y6Pol5oORbSPQb0sIS0vaVTF
mkM5zKyQqlRTKWvg0v7GbHC+P1MqrmIDkVSUnwsZyLesxsHNggaYPfX0KJMhuPGD
UWRrFicXOEA3AX7Bm0Cg1rB+4OMiNoOrgI1C8/ab/0z47DEAU3ROS7odQaeWESJd
K7ZUfCCwvmbJRYZBiDFI1RDDdfrGcJ6psTWJA4x1yNNQ2GczAKRLJuzYrYTpyDJA
E19ugK65DiSp7lmrDzPis5u3+LO2bmSGlrYTUYH91jSi3TKN7ellmBx6dx25t6Z0
qnWAWDk9Rccqf5QBiv73TFwcmCQ0Y9M6HVYcbraMCDwSViQ8XsJ4rd5MmzTsZa6r
MW8C7nycVaRIN/77f91rTmhF5fxQKngloGnLKmG/rvOsswncl3FeazZjmoPvJGZt
NoCbb3ZWGzxLDY9ejSqN2lYhuOQVuYwCUuLYEZlFIgR6wxl6nRz5zxQaWTl4934k
u1qJ7kIui1dxk0Qs4juThgUW/mtsNbnCX+5EtH+rIF7hmovLdh28zWLVqHNa+r6q
AhoERvUv4SXlXOpXEvRIqT8fJgWFyljAnH8PmWVPXLQXL1BXEsTwQJkADT5HS6Wg
XKagUMUDrD1KgoxLD1utcZFrZbAyD2ymGXi7choeEOIi0ROG1Mik0QhFegHbHUMP
pPG1MfSu+iIiQWJqA6eq3c+y+q4qOi1MfIJHqqOJX1UYM88j+fHngMLo+pFYcFsz
MesPe4h/zI9tH8QNHHBbZR6ajD5Lxb3V3rPVLtoNkH3CT/3oxYueNlfji8Yz6xAT
rZXD1t7ank/Qwr+SmJ9UElCbOlaJL/yuknFXiMtBCOgFyLhFdhll9deFXTvglKwE
IHYemG3sg0cFT6OHyYpUzIECsfo2hyLWywOKAnsHKwJtPe9oFLjVKkSR8+HVCJu/
OAXx9s/Es6U+6Le2/ih2HSOKje5XG39RQ14APgnqYr9+W1EERWlVdActEOrai1VS
NfSWB+pbid6Bm/ZJFvrKtNlZkMHHD7ekLnVrAuZvpjqR1UjGGOUs/egp1xyCSxCz
i/15GUYxWiWZni+ouVXV8M5f0+5T3lHygb4w8ooV3Sx7PXszmUvhTBZkYuvy9Uop
MJTlpBaccMDJEU+6C0ZQenKNWpAMzsWp7pdaCyVlf3DZSuIeWbb+9GyBly0wxvNP
Xj8aStVsxtjU/n0TQcUvQfHUsVBuifrJVLDix7cxVV3XYMG/j56MPz9NFJYNvGj/
YAU81N1KYelTa0ew9QBcx0jN+h/3woqZUabbXuQbt3Pw7G3JNbi01J6rDDVnRNzI
fN1cTKUgo5Kwyz/o+GP9IRuA/A689sk7mOv6F0GEzMVgBjz3btfk3ZaRTdJzsn4l
TnH4voYXrv5MXdnv9TbWLdyFKCdT+S5fMsvCbW1N3rRolZYa4cG0rCyaVmQ1Ts/J
gP7bEzVhNR+A4FkIRXS00pGyyNVrxapyojqfT/1S7T/Kx8P49sMgZoqNUuZXl3Ah
y1KEk8iMrpH0maM3mx8nEO1l3C17HTGQiuCUo7rWoXIzIz+xKaRPtVF3vMzw5s3z
/I7q5WfiR6dtx9NawXccxJEJ2yowxb3TOLs1D2xNuyuocyf4b5n6nHL4ppqhoBrL
njACoMJmz9avNkk22QAj3AOeTR+KvWj6KIkf80Rh3EXagLIk8XopnEf4QijJ7su/
YjblxpdXVP0x472ppep5L0KujT3+rtMUMC1Q1yBMeSBAr0S1SmEdHW9jhZ+VQsQD
L+JGLhToPaztBvubzXEApohOzxo4m4S04gdqlGAkHC9R61syf+y1vk9jhHpCeRJx
m8GhblF7Mrr7+dh1x3mkwBxd332uhQirzUn2WKUFSTJwHnXUU8UCDEUYhQKc7wfI
StcbCZwWCN0tIk8aHvxo2nWQfJwigILt4/YcCYeGs8F9KWaLGheChpUph3ldeq14
kno1qT/9vWLyLNbkdx/GhYAMQVMK9TjN6lQR3GqSRuWSVIuMpenZpgcy4xkX5nsi
qpeUMuwpLVw3cJHGKosLPqaaHQwjoRUYh9//b6DF4krYlmSYhW8OoaNgCh30aZqS
tlaihXBeMojHcuqzP1sKh8My2AA+YuThBekpI/7AT5/gJei1CENcpdm4cD4VBzph
6nIvp2dO5DY2hAtgI7at4a39Z9+Q9DD5UvAPf5ZFzbn6ERh7MDbUN1nnPfMYPDF/
FTMUNTPyGmWYY9b6ySp2YpQ5n9KgKa8/S1vugs+BVC68C4LLv5hrAR2m8f4umMaW
I+cBIB+oiurBZDXUy2VSOWvjhOzQLgC8C+WLWgJ6HEUM+1yakStuQ3QSnqNisLVW
ksaaXsXQsyx1GcNQhlOo/B1t/aqMyKGXGVCPcP9DONQC7QeLKMUZNvYt1uLTm8T9
za1wiFcwRxGi+LALVGhLg74oU6Oxmql7+sXDrdSMxrI/9EiE90qKTrhMMdvyn3Zd
3SJUeih48J/UJxJPBUBOvqNomXbLniYypOJe0dCJXChXOjqNC5zJCC0iVsp5BLNG
RyYfHzBKnw8Tc4SIw7JUQyS6o+lFLpNA8eG3MfA5hPbfTpULHNmTRW+aZgN8qY4q
2z16Lhc6yuCpmsYqT8XC7jegil7bW36dSOM2sob6nJZIc4p2LsZZL7Gm4tyKafxD
oVkERtefnmXI0QPhYGdwPgHnx1Pp7JvAN2a4v43EOwdWQlb+nekOb/09Db5uA1iU
HhTdFGHplRZiCdZiqPvEvsDJBHmDBOK/dPTNMGLAJH+qicUBJPKQ1sdtVWuEC2LF
x3C+8HEYhorMrkKl89iiA4wFPzAElxkZiXhLnmq8pOoLoER0dt6HlJXmFbkqQOtG
rxC51SIXkkrs4dS+LN+X9bQbE5IPrq+qBfL+E2YSiTvD8ty2lL6QKgAfHAKEZBG6
/xnSbW8a4JiO+o+RjFAqfEk3atcyyZHUxiizUyvc5qfF0hN7GX/yrI3OzBZI+oVH
EiAMCqAw1Ic90J4+uWuP6Lg0DyZba6tpO5P8xxjzr1eAnGuBj3D4wMf9u0vD0JfM
Nd1sY6pjPHc+Hho7vVQ641M7l6HSt3kAD2xifmqXabDj9LfuKZDvPC0BrmUpv7WP
V9/+F9MysE73IHioCy1OIohyxAmblwjFeRbyp+C80d/kW/y9UzRO4nVi9i9gOiHH
q09WHpAljFJV0eghSXzTwLIuYa3wc1vrMskSId87wexPGNNEHCorM/RIQazP3FOe
8QfTynYs8C+bAlT/TNnNRBXWdSnmtxQeCurY6BgAIDWin13LsO9zrJvHjS7BQQ7G
ORYXeiU8DaR9dPSjy2b0/gHtZYUIsBmP79ETEa5aFGFdQpC0+/l6hHbETwbvh9ZZ
pzqYrFpyCB3oTvW8q5hZeYCfgWBKl5JglyA8c28tOgByG9cwdScScwtwSyKYbvn8
3K+1OVB4vPNv50ZPJL/ihfQPSP6zkUnR29VNJitJWCCXhMGOqerD6QyJjRuLAUjV
JN8l6vF+qirkgKYlHyEZnamRh2jKiN3G4XlfB7YHO+JUd1KirV1J9RsQUK9vUqqq
bbhEPnyVtA+unOalxS9CNdmUS+OOQjuPUqBpMePCJ2inddFCHJORIVtDDHV9MG2C
3zUNJz8/LthTn6POr0F8fk2984yDl9fr4K5Hx0ByYEY6vUDtTZ6eBRd3qpwmkbOI
Unq+9iBY+bK8dLNTGqftyFJDzS+JPe1cB5vFZTDNRauTQ038uPmXBI9mO6D9V4ue
PhkpML4fy86Axg0dCr495sGSmT59MxXvnNPwY76O7an+7ZDEM2sIyB9Ifqo9k/Hm
sMaZnQmUPNkHfsHo36LakOIrwKBSvjHk3tIUrIUd+uCkKonU9IuDHl7we5xQ4ySu
WfXDBqMyc1gxeuvdnz1IexUzQd/o8I6O80mfWOSOHaRR+w9RsuAoT1ErsSdETc2e
i+JqxUtWsXUSkMXTwfIVCWajNX5fiFL1J9Pf6AmEWe+8RrZJqO0zBtAZBJZvzsVu
3KYl+vDw+ogOcAnhlK4CDhVz0/JOb5WaA2ExqklSm8XUOru+BLjV6nDNaNaF9EA0
TOg09WKJsjrD6wOQyb5dJRbKwHqs55CLAtPYfrDmXiG9UZ2wbOlkah7WputEMRWk
j/H8lxqFiHTKRPl36B/RtJSxnV67qPURJ2A5tq31UeEzzyj9trZ2I29dm9Kr2O8W
MG/erruxmxEfCKVougbj/fyvJulTJIiN2ktwtIT5PTiZ93VAVm8AUxHr8OglYMA9
8wB+Oi7p1V7ZfSyedbe9zXaT1S19bmNdlCeCfVL9n2Bn6TPHp+tpJInwlzjqmUnx
gVcPhXPMLxesmDqPQ2geNVHdV9czBCCoiVOLNYTCc7lKbU5+CYCxlG/HYYrvbJdE
/usyZzfsTb4/bfCH67X9FKLL+PsBOf+W2eb1FC2jvzNM7mC6WtOYKQJrDI/Lapvh
s0HD3qe8+g+B6Vkxv3ZCdkySgT5kcSJLkhASqcaDACKdkKcnnmXp5QhxLj5b75qV
ZV1EMq5NSQ8rWL6+RFul8qZqZ2r9ShObsE5BGQr9vtpsAwVDucrsWpCBCS2KlHyw
e6yw230Xw/IqoQ2BBia1TZewSUbLay54a/wm+tgtYGvuL5id8rOh5d7hiXcmliQI
2JJ5o2gRSudO4g/4jByG6rNX+w5MUMm/Ut7jTsrIV+ACNpx/7S7/XGVyDgIuFdzC
zEWUWRmpJiUvQPgTPAGa9fsr4QlViqyRXAwlwpI9F5ZFLm9m9m8dAJmAaI3+Q4eR
1+84V2m6bZ3KuldGmQ082taPB6xPnQq2uUUVVZdX99KfUZ24CGiwCGAX7Ju+DxyD
oyFYMnrbdl6VJVl0ZN/0at1l4Vzr0yAAWckX7sQ/myZvWqcL85xn03N9QQ4vMg+J
mEK5xygsHZbPhGwg3Uh3lI+hJc7Ea+3I1ixDUFVMELCGGWgBD7oyeDTH1HlX/aWZ
bHJ9+IkHqcakXU6eJdcRGYKjCBIzlKZfX+3QfZS2HxQhQNaG+U4yv6Rqhnvdip1a
+6Hxgy0I5gJCpUIw0zYOobl6+jIKgjGTjTWZlvjVvSo7MrGG0XB2zFVX/jTxIJQT
lfByAJbHB/LvBfKya3UkupNz1J21n7KkDJeV/hGORSLJElk2HuIiCJLapcgdL9Ip
Ic4R0fA0CjuHbn5iwFi135xe/92zMultmOEWTVD82pVZHTxTehnOHRX1ewKKtspu
iZM+dhhgIgWIf62rFdg7y1swtcposgRZi5lHuD1y86kA6+03ANQgxRsNWvoAz1jg
UC2Plxx0dV7sEQMAnW37V76dLl3SSax+SsNEr1Wz+a0PzElCjFx86ufyYc5VN/gB
1LKlZK9YgTcHuvVcRPoVj9vR+ZG5g8Qp8u0SA+t9i+dsa8DpqqRnqBx6YqsPRQOo
enyNAqS92iAOxArIdXmlGV93TPnzCx//vDNfxQ8+c7dt8FWyY7iRDI504uM8OeyO
6kLnvdA3edNfdYRRjuTQ2Qz65Ljc0pQyR5MfPKgSocpDODUrxGddgg89pmta1lEZ
h/84EYm+6PaKDjTRn6e/csbW5MAXWluXuYbX4VSkTdDeE7F2uS95LmVhpp/tiPSP
y0WzYRl2rqWx73IayezNukxwMJWFBWe9CoTda++gekap415pQz+bRd4DPVOhk+al
YrNr6WCzN4McFIKaZm1s65BHWPDBjI+QIIC3b5QPLt1PEX0zz6yulV28+CEnj7az
0OXZm0+qDQtYR9XnSo8wvHt8blrv131R5PTwfsQqT0IqMsG6kZM26uGBN13YaySU
a7b2XX6PsqQRInGMr50r39eA7++tUx8VBCSSqj14HSCWwdEZBSNNJ0gHzdhBdrAV
SsfJYGrewB8ABlWqplkPOLaFzwZ+vNUHujTqTzc1zwyQja2/g00djk848CMWUU2B
/Cgw9Gqda2vGlmrKODx2HuMMtd8FK/fXv+5wM4oaAKgpRGuPaATjzQW+WxZxkCrj
QEo1utGEtSlEzHm+coRa1E6tHS0FFUJKhS1bDzkHu8E/x4x4Sc4cCHR8r9lDZ/ae
Z392H52+TNG6MXL/D/J9JcssfKeJ/Pg3rS1z56bsgIOOboRdox7WfKTUNm9CDM6E
Rgx7GLhpZ/LHkFkZRDWltI8zM7K/j3rUNdl48G9WmIXAYBG0dwJPI7jkaTqXFrV7
UsUbbDPF5RewrT1tCaqunMDZX/BZTqqhxJPhNEWtZTwS3BifPB8AZalP5S4dvA1A
TeGNKmRnLOCkD2FK8zJJjS03M6PFhLPCemgs0HPbfvs/RHWi3OIhI5962CwGBXA4
JIZTJNgzoFivDxazDCCWzvhYqj2BjksEjznFW4RdiQ9aHs2QgDyEC8bY7LGpOBVk
m8iqzP8L1AW27PNG85ToEizMUDCotYRzM0HXbwa39nKKerFeFcJPoLDjW5n05So0
GDnjzrgu8y6lW3LxUfbM5To1z/YFgyCB2pM0jK8OWVqc//S2OKq4NP2A6o+UxMrI
7RELLT2qesgT2/35O32QBRW3TZZ/qnWdxBn0um7Vxh83hPD9M9FQTC/OXoQPSM4/
hGwsVZYbc6/uIzBj95U7fnQ18vfliw46hpM7WktNaL59LRsuImk4khY1hNftR3iN
UraEPAj7ngmGdwvkGw6rJFJS6/yxWXtfp7KjQQ1EcU0B/sFbgNZLf8MIyJcQEM+c
K8F0xzBgdaSroQFSGU97DshTp5sl4P5sT3iJ7QvGPa81kOucc9TL1guZEH1/ZOM4
j1Z5p6pZM9pQytW7AGUvpnft/J/C8eOvtCaKivPqpIR0gG6kB2GnInMVpMk61feA
/nsNLmP9vxMSkUu1JYcFFFFoAuKNmJlpZ07W0SZwSukM7PnVT03SCo4PCTM3lMCC
DD3TBlIYLPP06O/AiqYLk+Tv7JFuRFRVVa/yD40z+zTo3UTOu5u5uB5HCHKv7Nhi
C9yBj6tGyeaYmTcbSsxJhtJigkCq7aLqf8c3mhdmtOr0iLtMW4X68H8qaZWIiZc7
QOVmbYra6D5v84m7RN+leBFznlegSJTTn3SdY4I4BfpCSvxhnj4Gjrq1XE56+edW
qCbPc1mSuLt5uhV3ArbIukV9bIT7GwtmH8jCJ9OdoS0xyxbpSOXHd0IjAWzVFyW+
bmKW72RuQZVMCELog2COB1Ot6N4p3PKpUW9JGjxmUzS0tCunAomllTBJQzPsbtgN
kXcr8P5bnzvCLPTpS/NSmsF64aEd9qhVyDfFdRtsC1ncGsmD5xhTD3IYY3166J3G
RvrY8+JX0b4n3jVO4KVGD1JEh4PNntu9SnxVZgE8VlLgwZkP7l6z3F4+xxxRc3Cm
EN2gUIaJEBLnUmsgj5wQUEV4XK87HCxlh5C601WR1fwzQ9iUkcAtUHgKQdwOi0ET
/b8PrhKDJ+qZTlQPc5BS+28GxoW/pLuJtXUa7wPgt/agTfjyCRZ0Jdwic4gX/1L1
L86V8tgYnCx4otVALU5sCVr8Hbpodb9UtS20tiZDm+q0DeHBlTQhnKi3Blq5J8ZZ
ueWXkGKxtEzfsL4V+2g9cftr2m09f8xPcVyCI6cjQeDwZw7AB0LjA3x2SWpcjObw
Q4I2OeBtgsdg77YlBCFisq4MhHJ/EQ5aPh8gXh0PPnQkGu9SYJ7GVRVCwGxZowGv
dbwlnbZwPoDRac4aKCmh71Csr5Mebw9HbmSp0rOPpJTFtdW1tX1M0e38MQU9+yaM
KubL93fKrWegQvLx4FXb7rqtbqtBKFoYc9/HXIrt5hc66RPLcv9YqRa9MvHBsMGs
Hthk36f6go+ougYY+DjRq3oDSI8p79Ki5//TfiVGhLQuQ3BDil2kL1MNwvwQg9hV
s5dTjXFhQpfYc8BHMh58Q8C7KI2yknRtyvkTM9/SLLrK6tlI2R/vC2obQGMWfm0m
xWOXK5jc2SA7rqinIQO3zKPbM5SyZ7d6Je/LaLWck05WgIujfHbNapPd8h22ABeI
Qtx0wlIsBx+MK+aKOK5R5Rgzt+U7n64JJGPOHljt0Kstl/lnAW0ybAgifZ5pm5E9
PRTnuGMpW04I27T2lfmxPEYzgAfmesWXr5eok//CCkiV7QqvRFDoZXfhaRRdUEAi
tMznsOPblSe34z9XXJqiMLbHj6gn7LeWayFLF+pd+DnJS+g3Wd61QpdKWyVVjvJd
pfE+ajXA1un+7yNzQuAkQLVuh1xCDQQyv9WGTs+zT7LpqT0u12zAeNm1tqrCL5lT
rZerCg0ikY4mcxsutrBwCR+V1UuZfHeIfUb8U9mLd/ixgZf9RY4s97fanFBg9E+K
/Rkj9R8H3LBanAkyYk7aNwazC+vn4nbqJMyBhWghbRvX3nvLOJXv4wzU1ZJ1bcCA
t74h8xXcBs5n0s1xAIlJkFmx5xrU9PT8RWCFfQ3283PlBUtLf+p2Up8zvAxC6tYt
K3JAFGcMeR4ZkJWsEZ6TCLiHvL2rrHSdBbCwQhN6NRYFbvP5VIxYrIrBN+57WFJN
Nuty24DcxlKDaZlOh/XpMjN4+vPeloTHNYKKTbZo7RKlWQzQcCUrxdnVlV957x4b
fRGXec6WuuVFeD/KpoMc6XRCUE7ZGawWGg0AUuJgUd5cwH5mKESBerSn51xTrUbu
qkrM2CTN7DLlXqXNszCGtPn2RmT/z4B4nIXO2UGVYU0E1kLhDKA2eN2aQp7RBIiE
r84aQ3X01m2bWaf5AHvJtm6CqOAXmyW08V8bPgc9cw6LKgGTGCK1fZDZrj2dLFo8
z3FpDjRTgO6kmAsQi3gIKYOkfuy3xW77WQY/4efIycNzk8wMJkmuB6tT8OohTShG
2uYAnl9aZYzEfD/JZh6r6Hqj0CCME8I8j3ZLJUyPrS0wcsrO+AvyHAEiazDcsS17
xXFmYGpuGm/ABjuMwsMYPtYunsHnrsKGEERP5RIipPljCtfat+0GexZ2Nszaj9Fq
gwzjPaNTXvn+rHNGr52EXvKWVW0NQ1tGJmf03HOGILD25BJS/pY3DoWiFnbaO7vy
5AFFZm4NDPTJXdms4UfaEF0LyeOGBpOkZxU5MpHjM9Ro79WjGlxw6vEcR0VRgHIG
XtFSFQtensVgjmfBJVOSzNao/68c1mSIwLUlV6bdXehRUiJtzpqbN1FUiJlDroH9
5JQUFNbUdxEi0lFjW4x3KGaGIA0QckmQfyPyyZhqq6MNwhhx9qncFRsNVq5qzEn+
H+j3ZLLLIIe+EM2DPPSzSksBxBq5dGtYKYoCfbPPvdeOy8pa1IYG2S9HxVS27Tjz
cSGZziJBq4MCeXdDWxBsWlF6+COZlSFvjaZOrWOz8qTsP3PsLdfwbU1myVW5UKDs
OaoLFzgqXKctxt0gkfYEqEq9fEnheS03PNVzjNrawVYc8U0ebCStMpTUn6KzP6yI
BKTYeRxUJY3gUyM3Y30dsAaef4mnweUqr/9vNMStJpzcJK+B5TNYgSejpFXDAL3c
W5tH0TU+Vx/Ups81iof5kjL52zb+pW1Uubs9W72OcIc44TxdlwUeZqnouO73R3Qe
+9FOmAXkW5CfGRc9YZzPHUyxODjiI7XN7il9YQm25F6HzTbQ9oa0if8Mdk3OINuM
gyrgAyQKgGykH6ztN7qqmUuMTjStZiTm/QskWrHRn/e4+pSrCiG7QdxDF/YkHdKp
rdY65toko5xt4L/YrMqOySSN1wt3kfHDaxzkcgaNAv2RxkrDr8EPdZwK2Zq1oRs1
ZkhhVRiS2D3L6w7EKnGPFknbZfl+BPpYPOfIDDwWM1grewaDb23JCBlid0Zu9u7q
ToDrqjhDPU8JBQ/jfZ/Dz4a3SCdfqLo29uFGx0yMbTyi2258x6CLShSbK2QQN/4/
CS3EgKQoz+gH6uN+RlasZLpIlssy4tYFpa+9w35/T7JSVLqw5lKj5DW76rxnJ27r
AUvsExd/r58QHjWeL+gVrDonbSBfm94dJABwUNZnqVDZZPucLDDWr6N1R0p49/F/
8H0ZFlRE1dY7X1Hj/KJw9+jIMa39vpUEcWy0BvYKBRQL+MaHPNFbWn+MrHECrix6
Igt9pA8NPmxJvuR9N4cC/qnyE3IQlxUqsBFjkHlQX7+/kbu7mgEal4odUoPkKOUA
qccQt8CauxkzOYCaLREutY3jHtSIeI5/qTx8prpYF/OWFf/QR+ZTrfMTSVRjptnH
2Bd5lQtSECxt5JLMPLHVR8tek6NKLfoH8uby5vUh3vD6j7ceDlJkVjTav5OybW31
sZqzCMGcupxkDdCiYBB785QWk3v0etwnPXOs+eVp6V5WEb9R5EghrqSpPv0dUYXB
R211+9TTXf/xi77y4cQNu3H6hUu7BmHeQZnWGxBJaJaFODC0AD2rKOS7ncfL0XMg
dzP6hPqnoH1QT+XkND80icn0+mO3vd9WccRIQE2fRkvACooZh0hms+kjNZ3Avo8v
wxuJJIkHuqs9S74atma4FTqIs4Pc4vKFw+qlCucmP40ul1AS564WNtrUBJSE0Z26
nA052+RiJUiWi0Xwby2CI4yNI4bQFiTo2MNRQ1ZcWjaRCV9U6tVEabXC4ll34FdL
2AIHxDUjqwcKXuIFPf9gE12/PGHUBqt0nAyl61E5h1OJP8RvgM8jvWgeF0MpKX20
Oyc14sz7BDQbAL1mn2zVLjZbVByFLY0vSGFqy4D76TcDXaTCKyOZd+AZvqUlh8cc
5YSWmdR5bF85Cg65dn6moNXY+CS9laTx2B79A6IzqdUlm86ugLTCFK+sSlhmR7WZ
HezP8nFDClioIREaBFcs+zQvlphJQCDqebOfEABrcNpv0fw2nKHizitWPXFoaWcp
7wrQpiRvx/eMb90e3g6R9wnbcXbb+DFKB6pi6aOEzCGcLgHm3djDYkX27/iaghnW
KyJirIfl9iqaL2nuivMn2zkP7yTyvei5jm01CnqdWys6Q3ICEcNLhQWpSzvff5VE
vpP8rPVNLchtY0Y6591l8RWotKJL53CZEKV44HyqCRdVHO1rIQ8/sI2b0gY8SIqn
QCYoRV2PfyTZp3MT7OB59L8mHZiS98RuI7Lbbve+xD6rLxwNBaLTDccd3v6fJ4Vs
HPs1YGU139s7Ftt15uiHedJfYLatBBXVwllCB1pZAqeXHcWTsbiN32nIHXQx+FSL
lx6b2/uj7Li6rOpGAVj/z9uDHaKXLqJjHwHAgsG0RnPGyeDIgM/6PPdIB8SQVbnw
mUsx3TFFGFadPOrfASaMaY+6NEW6Dxb+c/WolMqTUChefTK1yBX4XUadrlkZD0WB
ws2TJq5b9wLLhUW7GPLPIxdnTdqvIYbeeJgb/mJkslVX0SdV7eCpW+p+/BKX+lEN
wGYp2P+V8WF2xpTqDvdILS+PlOTMxlSAXZD7aHXYrdQR/b6KUiY0GElYStdX8CUm
Mr75+g2FVq6LJFbw5A4Agq9qYpKhgbcYfC6y35bcv0EHplWndwtkmC2eS1I4WuH9
5ZR2wgVgoxUOkqnlv0pVWZROmiJD7uh2TGGrqEV8j9FT6gqvZRaskhmw+mgXwnZ2
HrZGMjtyAIVaYsvNGLGfJkiJcuBKwDDQWeVg59Sty+f1WceuHLshZQum5MxalxQN
r0cDokF6V2vdN90rnlYqEYfVTwU/4qqX2gwyfosDG8abz4w03yefTmxy5iRZAOfb
Ek99r0+VsrMfHCFtwjLWe88zUEgjNd2u53Cbx1PVcg8BcB4LZlSQZPkZz0IgO4+R
NzIefywQ+mYMTVk9XQJBHTzpUe6LnCdGe+5pp9ImXFinkgCFvAM2bANymIi+Iqi+
qdVawoMtlPx/ZcLb4Cpomycf6cTQDiRBhMXyoMw0gv9pRGu7n71M2Au9ssdkwcLH
TkraGv3EGmzqSzdOPsv2jzMBe2Pp8e+9t5Eanwmh3bKgX6zIZMhOsQV3dxbwkZ69
NSeYUyi4i01cmef9jIWdnoTVq4wIk+ZCkpvocXGpn0Wsghqlq2IPAE2nI3A9Ipqh
OhCk6x0LV5xMl1iW6AkkhT/xOvntdOk9f6Z0wy4lvCRImMMhP8ctlyq/8zMVmc9B
G7jJHbKogO/J4Pnamxkj1DHNQmFrfLN+0AbsAwEAHRPFtyvP53gWV0iPX0mejJ4l
8NvFWihBleOyNer9ml1YeYUUi6XYS3aAxGeA3wAzLFsnVyyOhVbDbDZzk/j0y6oS
+qvUWLTy+5DGQ1QCjjFs7tysbL/mxfwBw9abdU6hMOBPmHX86YJpITb6iafYyKiL
beNax3Z/uicsspqS2SDjMuNnIYXP+TudIyFp7IBiMtQCM8qC8ZD9C3M5ChrtP7F5
9sLaq19e3aR+915BsTC96uBdq0N0l+gOLRPwOKib2cQABNNlCWzUNqjc7B3zFHr4
jKqtInTCA3fzQrldT1p1qokSq3mLUvMM7XMDwKr/qCNHSYMhsPhPBfET/IEgVe2L
ULuhKQCUp1uftu6FzRnLHtdvE0I7wDxbzvvUEvKT5vSkOKMFpxq6BTqx9C0/bUM+
tcOLFaM10kvFj72b3VEf/RNEVKzAr2qRekZMrsJAmt2V4Dm2BWxuRqaIOu/OC/vc
loCXSJDaOi3J2DOAAl3ZX8crLNJgPiM+GNOLtzbrltTKuD2r+ViHPYuc9Qj+wV+Y
DjK5PEdIvSbTnjKiaPg7k8y5Wbv814Qq96cuJjkxEiTBoLHuAUHIO8/qzawGT+Sb
J829aYHTaEroAsfwwdDqEICZZ+MEiIAESwSnN3HsL9ucH0xT5eHsdRCDxyhPr2WA
zPA9gbMQ0rPHpRMxaLlR7MfE9UubZizjn9pcb6I4f91yy7/1VmFw90Lglg7O+J63
p86wy0W9h60Yijn6m8TbAdn/RO689ZPmJY5X/A7oEj8zYGjwX3m/OXCNbZjuU0eI
ZRg4Xdz+7SXFdUhxCaRFE2rTiYpCdp6wm5V+Vmue5mr7p8g6cmOdPWpFmMqOQ4PR
EKaVPgPG7hNUfLEzH626iPtTI86jHLPCQ9gFE62ZznQMohs0s/p5xfVFh669vEZj
WoBrjMkZp23in11F+ugZegN5JUx98Ji5eMfuqqQmg/jO1JCJ/yONo4HT0blLP3lX
iScEbgnuy+/qN9hArs+UTvhzD38GcWk41cLS/nbz6LXyfmG+9hDWpfJpWrM9GAna
XWd6bDuUp1WAmk1+o0g99VZvI7T1Dg1s5amwmcPZIAsGYy/W29/V/hKQ/IQPDaoh
qvARZkAXipj4sEneiFeI0yGuC03Gm3+qy+teLgGp1lWtZW+u+NLZHzTmg6mdiwGu
ZuTY/1zM4UT3EqJNlc/TPV+3T2VDGFTckrGd75TjzMZed+t25Jwfd28hXqLR6OIU
Da7OqI6ybY6JgjI4cpjD4pJB8dSlZ15j6Bg6fw+ilQxSUCKH5BuMldCCrzkLXBFv
PfDXZLPWgy65vZunWx/RzwAPkonpEOfM9THUFQWGazXdUxvl/LHYT8MiNlXVX3Qj
9U/Ag6fYVwurCRhby7umsrtsttjJMLkFKfVhR5mJAmPSX1+52pnFNnATib+TPDKI
XvNFO39HNZZIQ5rUonMYko5KfdR82hM6de8ZEqVgtznzPH0945dHkrTrCgL0Rlhh
tmLl72BkoPTK1clh3arpW1bkdFCiV83rUKhs4B2TZY68lEZ3HfnDAq+9Tljig53i
HCT77eKRTiGu8j84Nx1fN+eaFNxG8NaiTKTunCf/lIo8X0SWw90joRMtTa83JRuG
1rkEdZt+UA0dDs+80dCj0wTvI+gC6uA42COdi4LaxLv1Xq0x231rEj+53/ic55ph
C0lLSTkdSD1OzDNDpbf//q+1cLTuyaGpg7DjQsdwvT/COL368wYUZN3yxSx3uY1y
64DTbxb53M/iLAUGjNzRv44G6WdewwmL/YW9qWu6fA1R+EcWChbYIJ/W6vyL9Opw
9S4MElrpv+ML66ZCgX9fRq7Ls14KlysL7ml2UzRRjJtGmwCC3Vw5EXkmkHXs210l
oLm9p+Rd7h+LT98s4j8XHcVqz3gzCicMDbKOUuGTUnXXL9p5wjzY/CobVSkStPPJ
Wd0c/Y3TcOjsQJu7cpNBM97ppamozuQAof7txbwJgyPPvFEWVE2mNWoxy2XTLdpj
u/0iFBuk4L0JBoRyVRmeDu8YjZq+STM/it5oHAppgo9PTtb33o7KhK7InjooglUW
IEeafqXBQs6Lh1vUQwXy0/4BxY+J+3ovYc/l77iKy9zQEMs30qOrfu97fk0tM9Az
V+j27ZZx3ontMPDO7vxu2bzZ0ZiwwygoBDFkcZCZyv1r9rCm8KMUwKGAg88byI07
WmDR5TE2SI/5/CPpVjYKYoy5SqhPhDBsNegIQ2cxZmztMTjgeDujrGnrLIt1UfTa
W9GVOCyFAgBvl9tySURyICZ079NbdEcjWphegLcUj6SYRxvQDAIdLvMPjbrtzaoK
+TUFCBX4/QCnXzEkpKJL+x4qwM2ERNAzl3Bbs+RBMlcF3aV4/3Qb0gbTg36ABrtw
OIjee1WYIGLuPXbQNROCYSp3l6vH2EzcnsbWSenQTVcbI/Fkqty9qf7HpqEh37uw
F+03QtOaLsaKW2ySuirt5nXYQBnVIKKr69DJZSi+QBWVvSXFqWCWsSiwkEJAurdg
Q4aFjzBg5Um5CW+naoeNSZmD+te/NSmQvFfA4sT7e7deMjKVbYkoUpP7IgXYfDsb
MGZNv9qgfzGurshkdzQih/fgRQ7SSaVFEXx8nHDcbzCwSagEodVx9RoynuAK5yTv
n1qgaKyWF+gqPJxFZVjl+4ndGAjyHxuc9PxawldSv274C3u2bSBF/uSpmnI01J7N
JJI6Gr2CVGznXodlYc2iRWO4DYKg5Cf99OP9xiKDsMPSPDHiBN+iDvcA+noCNNey
wHuU9Isbl+IUqo7F9pPDmqw9vAaGbY+e/A+YMcM69+ir0RrGghWe7FwjgdWoIBb3
aFSMCf59wjBd1aGHmTzYc3NAFhjfTq/Hdt2XnctlDr00p9Bl3XAp1VkUHdsE3wHX
Utkslm5IBG82fllOJrSfBDIy5XlYAB0M25Obj6nOngpJE310LaQNKufQTh64xZK7
8H+Oucx9vpbp+GAv5IWi2LeDgt7lpxZmn8aoNIBA1O6DueZeVvMGLNuWMr/1riry
hpWx4um7GVWo3tWNUohfjz1MsVSIqx1MKo97hrj0APaxQtGSKadjW6ZngJ+eVmO2
vKEzlm/mYNm0jR3dBXJRO/kWLdMiB0VuwH5HUTfDy1zdKACAbkgNMehOH9h8dg+V
ShsvPQD2kzZtqIaR58zUSDZUfoRLq4a5nUMIHvntYs/WeV6ptBPsJiRvqkr7fgpL
eoPCJktgQS8DjugARaaNS34j3YgaG4pQ2t8XPSASHtWTJEDj50PldhMbYFEXFedd
RkUo1GgISAvwmDHF+Sj02jqFs20D3Q2PJ67PLCiy30sTsQte1oj7CGVGzcEFe1rk
H7ePmQKjozM3kB8cckuNKMq58zUS0jzPDbV+uNkWTvXeXN9jAuI62L7t+K+F2KCj
CP0hD6+qNTg3eeAEKcV1gvNr+Fdf4K2e5Trnlh4sZDic6mpuwYXGkhEpcYPhKwFW
ZTw7bHFdkUKG/24YSWoqDWQg5qiECi6JYYOblWIRznU3RHfpi81HLRwx6KkRtD4H
ONbNCr7bK+GKeoJq/8Jol+oqhuRYiLopCbYXJ5PmHEbRP1y5ZxYQz4E6zP3KmY3o
dG3faoSfI4yzbYqL0KOSiTiMfvEBdzKpNjr2M4BrGjdOOZLi1vqTKlwK9TDti9Mt
vXBvqRZ2KQ42+TmaEYtL3P/Cp2jlAdyXDKplGeODR6hKG+1Dg67qM7naJMLiuQAV
6sesR3RWIw/zf8xrjpXNmjYQkJPBPV/bL2he7BcK9Vx7oi0M9XlYazmvv5z3cWK9
yU08e2Wz9Ap5iqanzT4BR8u4dlwtorSDpySiCkgj8MNZvW00vbIyeVl2lDPBR1qU
h/BajDLHY5qdwuMiT8c4bBf6f4UAICbvbelmgSlKlqVJ5fuu6Btim90IsRnk9rk9
wdfT5Knfya36+u8G8W/jmgzFR6nL3oLfveKQBAEZdzHQVwMwiqA4K/+WoB8a35tA
TuhE43hva6NQTVQSZntg0HBXp97wTDwCUrVCstnPhBMBnLT+1IphRfCeY1auoaQL
ed9U1QKwpUo2OHiuIHw9Uugkz8zrfeV6LJe1a9SiID/p9obrtGK+1dTbmvhLKiVM
JCdJpxUIejXH5s4bonSrYZLKWiwtdstXdv0drY65lp6V7LN1ZLQmkJxhkpGnRugN
S2s4ssQmzjAGqRMF6+wx3wImz4Za+FuYP3RTfcFEOJedXAz8fVyhc2aQfT416isY
AYS5V3tdag6oJdU5HMxr1R1wYOcL29zCjeWBi2AzEMlvKeyxiO961jV/lDsmWS3v
2/wO1n1iiN7SK7jnR+rirNwCiIhaWN7Kj7ZDm5jTw6NWc9uUkxYtsYJ/vR6uuFtz
yQAn3Q1wJihZNcc5gCHMqOdqwPZvOaDqzeNh2jpuZfv3941OdO3GbaMcxFVUvAIY
evLI0VXnz036teMhzZ4xoqFBr0SuvQq7PCSxhARGbVlw78P0WyjwoIG0RQaFEAvs
r/vwC/TzHPIKKQjCguLbY//b9j+lBxXaF0jl7RFKg80QvrmetiaiNwouUscn1V20
F+C6EeJkRMK+Hw6zIRfpxz3GvG1R7HehJkUTPskDJX5SwI4a+H8JxJG7+a2RlG8D
FPqHSkqyiQ8UJOyx1JZ5EUi0Tj/cMRYF2iH/ZEqWtUiH9mThpEEDrsh1EzjqrZQn
Yf8UjfvT1Dw3U9RuRiRJR/DIVsSX/9cHgcZ389p+pmwINzy4q5Bs9eGJdhxe4qcX
O6Ooy+a2Gv0cTWBno3+RoPXsDg1Us4pK0NLiRm6+2EsiAbYlImug7FSfFYrfGIYq
2zfuID91pIqdmHIfuI4uCAMMS5weAA8q8ADAGur3Zn3LemDsMWTS1odEq1O4Vq9o
A9GgHbzxlk7Ehd9m37YWIyG9vRDQXGdZ2xaQpVKXxc+hQ8PnmpajJslALo8I8dFz
41wgGDPXKfZIy36bBj9hQgSbYBgpzGHmh1kSEX0O4o0ij97I7Gv4j9Cm2wb3j3mQ
+D1caTzSyV/NT7pmF4ZWYyXthn7k1ucIej7nijRxzodQIa4D6NaLWwpZbsTXG6UL
2B2dkCvrLDRxk2HMIOskV3eKv+N55H1bjbNYGnipiW8OyfFAqfLCZWXlEuyn6uaI
9DVYzZs1WPYAOB21z2Pyb+sNGwuK68p9hZ5VuIUN6HLmXVhdR1fluxa5/G4tLbgz
5W2a1lHXi1Ae4ClRE+5LTA2ihAcb3+w4Ku1mf66vbMKbXdyVWFRWLkJltUBWHedm
s8XwsRY97qLDxE/QEtBclOGjYZ9zOxNJ5PqQcpCrMI4h2p5+TSDsb6zX3Vp4ZCSi
njfZhKv3dWG4lqbDBCCK+zLKFEzLuew18cgfJs10Z07t7MlAjN/2QmI2vSJ8BBbf
sfMiUIWPKosoQCekVE3risYrfHd0t4J4L/xHCQ0Lj9sQt0F72gZHGS7wmFS21di+
FaJDS20Jhq90aIZyl8os9uuV5FM3CBtO1+R9iFcF59iCkv9IGLVOeRU+3QmLHlfm
vC78Qg4uw1HOMrfuAau1+z+avPJykF+RWmzIJtjNsjGe6w4EZ+WM2dOdL7jiViQO
OEpw05XdDFWokHWpNMSRfXOD5Y1Nb4dcEXFEme+g/NxIvqMaJ9NaNONJog1uii4Y
P1XrVV4OmvjttK10enZdBMHm8xmf2UeYcZnvoUGj7LE+N7StNhVO+qUT0Zd/GUcL
THfYT1+Gx7stZvDkfXVAsMP4gdn3dWQ4pcDPNsVofqCGZm0U1e0kgEcX12doKH8F
MfEKTSQgyAoX4J6aTZPAY81QAJX6swyMmXk9olKAFuLLT75nrcDxubssPT5qA1AO
zIzvlm6dd+M6eAKASlcWmTxgereUveAMrjyGMBmhlqwr1NzgOZYWiFdR625fkUyl
grGJBRNH9BuJjUsZBPf8jjud48gylSzX8LHyLX0k3o6uRBvtbAKLV3E3y39HiKG3
qlqiazGH7xjXghUVl3wNxBVjoYcYEZN08e+ey53SIuBQpagVZoofMBYHa1zNuxip
O5JwWcc0vzFx0g8VBn1jJu/I7tjUN9lM0HbCtnfjz24eh2pEr+txxokBhEwzLoKk
GhgpUcnnx8jG6oQZxxRlliQuiHwweVDotFyAgrQAzHeuxX0QD5GripcgD7d8ULSQ
xhMalNKFl+Hr0JG4fT6sBwOIU8PrOxMHpIfPbRsFTrJsza7rY352tj81yReNOocN
w3i2dhY6L2N6Ma1VMopV7+tU+S3f5OQ3rizMeX6KXpUl7XqDEq79i22JM9KWjTQ9
h+1l1MIlQdRxn2ykPgpZAjNSHXUAznikTLAc9X66extyrDr3QsNLqTKwSUMO9gMt
3OySXvM5lYfgAbWRcPt9g6vdAZ7Nfr0LERF/UiQOT9uvndsSXVEyP5S0x6kntRpL
MkrZsqda1qVnok2LTtqACkCl7vBIKT+dViVYeQqX2jOCzliP+HdDF0+6qWEuQqfe
2HatpdiJVMzmx4gh2oarp6cICyuCDAsWJBDoZwSeWJiV/E4ItX28gSktXy9OKHwd
d8JVJv+baww/9X/k/roH5SCKYQrfIWbX1rbOfIn5jvPOqRcTWvVxB5nQQC/jN547
EvGkWoqBCNvbC2aH8gTaQF3qbZRsnUQ3OE5bebBBD1yYX62OkpUQgloWnoTOulsk
g0Y6/vsr6Pa2eIeECyj2ScHF3325HFiSj2NK65sL0kjz2bgNGSPWYR2m3FuJQHtu
1eaf+5/fxqcXPLNP2bWaS/jcgqDhltyijeMEanbeknE23ADP5gIC+TDFTAIQ8b2I
f69ap6IvjYnPdXKErv2kbn9hK3jkN0mGWqWt6BkMpLSLcQIY886xm3M0iGWSazaJ
/Uv9N6kunjf/JI6RH8kKOFOz73mmB88bg38PBd6K2MaSv1rc+/bqRS2UsFqiFqzh
08N63jVy+/U8+W+AIUy1LiTvg+3tSPn0SoLRNBZjS6ZrkkSkuleu/aqZERiZyu3V
yk65OdES8LmAjLOMafFcKN15XSXwButkJzj7AjB1XgAldeepdkwPRNd4TciuRywr
yGJ+q1geuevyu43ALPhgIjTv9Q3PyAYuL+Kk5Ny1fA+xTrZWTBy6Zl/pxAn/B68p
ymyv7ub2gzfgRAKF5+wpnecL382zhOeiXtMRqL9e6/ib3Uw9/aq/1pCTZdfRaks1
GpqmfLI1g1VVYuMzuX+rKC0ULB2pCd+oN9eOm6Hb3lUgYNtba3fL4MAZhEUPVDnw
yOslIg+zY+zesjq9wb1VxdgsKAD5Eg3eRb68vliEVQLEJj/e90bURD76Qxx3UsyA
Tx6Fs2K6UDimjFv8D8xXCmGXvudBUH4cMDX8Wacv7oSIXPdPgNlHGLUUoeW7Sh0a
GVvVArBnEb34HYlG5bEuA8TujSfCLEm4Ya+B91bcCld4HNDnCNZwU/BfCWDdbPHk
QJCPZAIhPjKwwDmtdNGw/Zfe9STjem4Gw5b74H2c08GY6y6Vy0oq7gx0mp4BLX36
PZrllPr2Gt8Pnjez8akXRMPcmcL4ClI/UC2hMiwd2Dn6NqU9vUGy9kj23Ke0PePl
33dRAjuMqIGTLFGSRnOHGzZCjo7pfK2/KOxB8G4Li9XLYqFP9jOe6gZVlRqbNkjp
9XlbwRq8nmD+Rei5cXEN31XyA6IVubS7WrGSICJQj5gHtFpOa+sXfb4ZQvvzXFkD
OGkmoAhBhHg0RbTLa9hu2Zz4FEFLHF2t823rnf974p2r8T7PQ+v/dJuUkK45MRaK
8eRKP6+zGPw7n1XgAwp4Uo3JU+2RkqEuObLS1qapDbV/ZdvYd4cHZVPMlmvCT/FI
JExt+IccPm4g6bQSn/tPjhkLPIhnl+3jyQpEc53fir1BoM2BdRpFUEnoPMQBA9/W
D5aDb3TNNz/S++SKUJiF4iI3xlH6usHfGd24UCxB6YfhChv1yVRanV98Y3NRhU0g
i4C/Jg7CNBilM7xCDA6l0sUsfElPjKQ79Z0qCWTvY3+LK0qQG+RxzYy1MwkyTtcc
QvZI61E4O7b3gRER7tIFAfpwdPIMbfnCND1bh4MsIyj52nnzz2sLcst+BOwU9r31
EMtN04x9s1K+s7exHPh7lgnnnCTzW/yUYcCJhc6+Nm/xsW4JRJ62mUfMbyt3JTmX
lGGMuUU+uuMzh1ujwPDEmLCYFsKk6IgDkGdPYLEl8hjlGDI2wOCpVL9oPB0GVDxC
69juIagqU+23q9eZdVKBBtLDcFwqK5QteV9Sj734BEMlRjgnW+xUuuK/Ip0/KgBl
M8x3qGTUxlsvwlP9wlKYR6RCECz7L4yGn7hbmKscUZNldfr/VCWKiGbSJcCL2ZOJ
FC3LHWnds5hVuPTxs8JsXf4+p8r1ZHRDENgXOnCgJCfArHOZjDw0BXROlAACxQoo
cc3nKtMBDrSadBUw8aUu8iMgAv/j8SMd/72eN2++f+naCgLwpthv4Gk8l/2eqTAd
skF0Mpchx9Iz72K2RNmkRykXJhQY92RNloQUcqD7X7RMZ17wEQDBpdgIJO4lxch9
c8PIo+Apk0wXkECRQVmxp1VvjqTM2ZEBhv9F+N9LBnT34wOuV9Wq7rAsj7MdJm7w
i+KX6pAwR3OOPhSGn3013Ka1sn9YcORE0MQNGmn5OmkgBzEVnlg7rSqiMX4mguO0
ev4iuJsDJnpA8fgOravSd6ms80Ih0rI5hFpYR/Ic/+v+0h4lHCk55zflvcarUaIQ
2cdx9Xml0W5bE2iRxk2r+aaCkOvk+WRbuRun30nQprhHNWLuQsOoIVZPhsAnI6Bk
Ogl4B0MuK1BD+dhB/rAb38CRCCjQnRkpKNjW1vH5r8f4qOY3Y6g5e+mxrFdP9l1L
yL1ANUQIjrikLCedrV7INgRkJjIBlHFCGqBeEeDzUTES/MiuSmSa8rGvZj3yqlMv
0BhVal7EfmyUnsrIfNMk7d/QLvvXATxDzXYewxa3Zj9oxSoCjrZzHQvy4e+NpUu1
IoEhqiG4BxsvboVN5+vAkJOR/b1+QT4+vqC4DA0UlPAyGAAp67pd+CwUNF4umb2Z
0HbwBjML0E114Pc1HO3lLVcGZC6xFY66BuiT5IbajcOOcNtCkAR0JO3C35KFTLx+
6886dwkHWdzdp4L//P59ceUI1DpG0xfYT+q7zM4QyZbv/4uWvLxBDblfXVaAahSA
rkA45UKRyiayUzvGkFNbb79xxo75fBfoh/N6rZgeSMGtWaAYyhbtraUL8bEU7LFQ
jJrgVy8bwRo5fBxzFZJqTbt2FuRnM1vcklDlbz2oXjRclDTpv9JIjLcjYFRN7xi6
hkaPLbrZBVQpOAHDABeD8mmdgmXoFEDJ/Ez20Q0ZHQWhS7difjnFRWjmX5czinBp
7rosPBvPyqgHHDmteua1mXZUARgRPGroP4QrNVGdUmYPlcEXCRE1+X7snPncxqvW
m1/siwp80E37OOCH/FkQOIynr5mwkw0FPRQg2dCSOAY++y9BJmL7vwkfVdUSy1NR
nsgwTN1/phvtiOIOKivYVRk8ch3knE9jdXMTr3lIweOTyW39DjQHdxsXR5WCOvSz
R8fx+sHPglAMnAKpS1DT8dalUps3kGNRzYhKlg0cLUzf0F2VWAFeG02I25vpbmfR
OhDxEdYB7F83z5g66GRQW6ktB9vRdL+YsOWaNNM6x9AWD2DYHhhxI73Y2jLA9qpm
ViFmUNDVB9CZGYVg52wb94JXO88epJ0Jr4H+ScQjUwlTyrxEMa05oXrvp9dOTTVh
dadPPy0GS+f1zgfEbDJlpQv4M6DsxQtuHYQN9aoUeYCptHE7qiNzONnHXpQ+5LUq
93xYASzjnpFJ7EXGIL5XW20SANQZVNa9iI2a0UDeejfseILwHE14kySBJYIB/iJh
qFBY6W9xDaVzokmUyJ1vxdDK21rpiqutA81xJy5s4hzKr3pjFqvAUVbrSc+3WdKV
LQCQjLTsGUGBlCRH64bYGpz/XLRzt1lGiZrOSQ9/Iw17BDLQMUeklNu5m4Onu5kj
SCNAwBcAmh1ZCJRYEzke7WA0vsyDWea4fUBCAMbLVckH5vVm4iMYM0HjWUuvKsef
mfJBxTAaPBYE/l17yk0MPyfI08Wbqvn4sj8tg9RwbfIpnjBWL/s4XNTrnkvJ+VZV
x1qtNol8GLw6CLOqEFRxOY/yfSbkmCC+mSngC0y9GQUzfw1I4yQWQjvPD9VUlOwn
KA2bB1a4ZvBIw+rOaI0p4OXfASjMVmMjATidC72rAB/Gf2bXJNquF5AgITlbOTGH
xfeAO5B5lSpwzfhd4Xjou57w9PSl8ssa/OUfSBBtGejVabS++MWWYiM+ucpxhykS
E3A0J7qNmQUiDy+DVaxI6M8AzOny0YZtmUbgc/NiVz91Qe4cde8RvuE+HpsGfMLB
oIxzeTdCAy8VEs0OyVb8/V56xwbWgjjfBtqfay6zJjj0kQ0Gf5P7yaZZwYXM1H8L
JdQ50jFAgznw9l+Ika2KpDW0fKXYn+EMvJSnWhWsiNtZrDFZFaNM6xmHEoI1mZcH
AFQmQ9VA6TGGZ+hMESimfPZcTPyzgDjx+FGAZWI8W6V93HLPFukCaI6LpR56GqIl
h6ZI1YTtd2ODZ6/Mj1qHAqay36Hu8BoWtQeHA0ZBbLfWedaWIrvkHdkPzPofMtPg
X1jHRxyiyAQ1w/0BJ/Z8t94PPpfvJR86CCtAIbkvItHRgC+HLTrDMVCMnjxgjDcD
vD1y7aLyBHuGOz1jjbXpmatiFVLGdu8rj6OgfZTaYArifAdQEN25C7EE3TlKr4t5
XqWgjMbZnILQse6Ee45X6pOij3gRopwRhG0RO+6IPpbMTW11Zx5gwgKkt5b3Ee6w
NiYg0YHenGoFPvhYUv9U850KujG41m5a3KhICZrIQ9SnTygBYyI089ZamvelfV+B
3PiJgooNk8OAOzsm6b0xjLH1g8nr92R1zaHVjRWgNpy6ZyBj36hDhW4WwDaUW/3H
B2DlNF86mQrSUElCymOauU1O3nw5u7BpeBep/G75Dpr5bfDMrOVPb/XjAK5DiKhY
VVBVsKFSCcLQ1cIXt0nHNhz50is1v7t40/3DtpQvTCMKPiKcSgOUuirU920zO5rQ
xgKJhZ2oarpo02oaFsMHKJtu3inhSw3MHz3gW++VLDVd+UZIm1Yluz4bC301CwhP
O0nyRyEYZf1MDigEjnkoCtSh4nPHw5/EBxDUTZZ00f0ojX7Ff+AJW34SDJ35LIDG
E4Sso5CfYGKS/RyVXN3C1Qjty12i82381G3zSTSBHi5knnM5phD6A5hqfgrv7T7z
LorLxG5Xp3njMVUfezR0hSSWMZI1wMtLUPoWCGbtivDlQlfRT//Oz78QLJ4Ms46K
ssQb88hGV9YDHwOtWwirTkx8T1VPBtgWRlXaxc1OxuR7p8GhP3WklAlN5qsPB9e/
SMDG5quzOAsFVfCdim8vFZtw/x2tjnm7z5/kwc8V5eFg9Lu6LEwFlZapNvl7XX/V
ieYuRI+f+y3HNw5YtWpPjwg+yp+Dhw6h48/514+oDxDvWynvSOkT8rXuP8SZI74X
PztH1uU9mMVFTLBPcO4uRL+a9nuEscrOynrJWgUsjlKTpFNckoMvMPdNqlEbvDRH
JaETfsr2wq9RKPsrgU2x1RaB99KaXO8w1sQWgakOBTL7o6zoya+Gy/QYwXJTZF5J
qjI+mEXR8xV0Wh+FOWQbP3WPbRCLORtzwjYgOooCS/kK1BHnOb/HsVSF6beZuGGP
Hz117fczagimAatgPolfd/zv1+IVfm+VmKWANH51lyM7LsFz9VLzyQz4cIpk5+ss
eRX/bgXxaTnyW/Y2HAwJMRXtkSZiDMo0A2XgQkFKSjoW6Q+YqIGqybO1Y6bM3PTY
Vq1CAj5mHj7VTcBhOnmOiZYdudDeM7MArnY02YmxEb2pC4WJExGpRPM2vDeZuHom
Q+4+mGizuEcZkHGM0cQZpfyf5WEY8FGPz2cjMTuwWLLrXRQTQpHceLBKfUqG8/jH
H3GdUAVSDaExjKol3a8oUeReK5TsolCjmjp9msJNLHO26VHTxIGvwlLaOr8D+I8N
9YJTCn3QoKI7l43+zYIMFVFb7KlTzUc+OdAxCAXq83ph3HD++BotOR0fTcku9Cze
BCUmezZ8KvGz1TXTEQf1GN/UyPYLWFnauvV/dQUPl47qoHZrH8fmyxTtDhH7xQXu
RFSR9UpKDR8kJyUmjPzEHd8Fr+YXAakqwQaSodtafxE13xEbAiEEmxiR6rIHjpr5
lJMytY7FM8xqtHcVdhOwIkWQ4N4LyyjzGlUvo0Uqimb2l2T+tlO7URk+ZUoYyFWu
QoKXqeA+XAU01cQDnAVy1F4WeIFAhQYI6pGcR3BVvQdsD8IT3UfcNRoB1aueHBaG
6MgdycDgbPbFQXatKDy09fj5z/YdN3AW6am/J4okELbnANR5lQ34GzS8LZUKLMlI
U67ifUGc0Vlfh66Csmg9gxUzykOIRULBED6iEHkTF5pNODO1Q9DBi7XUHNVTR19+
rKutyxpqRkrpcu77KOPvOOv7pixdGdYUNQs6TkZ447ZQlXl2KfvUIHsnOIp/jfOu
9cVgJhtIpHVjpqNz/n/fz2V4TJPNAGCTEyFzbR/Qgwas4XW7HnKVOVUy1OWYOChJ
758mk52GHd1SVxrk2S3b0Xo906/m+JvmakPLUfS1RWTNHBtdCYvLcpXyttEB1BLK
QMUyIGbNZbb+L+oDAa7SzszzqJ86sN7qQB/BRqrclvE299U3l3thuQz+2ig3MtGj
MRTDF4o7I1nBCVvas2J6nIiauKgKl+YS4NzMmU2m4EgHC+SYUubQcYZh3Khl7x+2
CoTmuwGiWfqHYQtcviv1IEaqK1NWsei1KzGNvB7j8W5tBKwgu8xrE5iawXzygH7J
RKl7O7K7bQV76UoRaSHBx+beSPpkQkt33SlhlaJ9eRQnCbfhfUsYMH78MqrizAdT
9MF/mrUs/8y+fGj9UWRR9GLLbcap8adTd8ePgRy6LmXPNglfLVNBuQXYG1KN1Suo
BKJIA1zN88RAWFruN9IsI4J3MbS4fR4aqHejKZJFUA2ioaqWNLZbBy8ra/ozJv3C
oPq6PX4uNxvzXwqSvQqiXsjxjWZpZH7jF4RPBKheIjaiEu5KabiJu+ZeWSu5OXiM
BeImXIpmE7GGhPH9r6QpjrKXgPcOdL5ZWpWOczJFmMvmrGaiH4d+XLXVgm3aknQO
8mm8c+GSjr1Ot1xLmdcZdnrfhMxp7HOtluFptjMLm7tUaQqLJmZAPHnHttC7+x1Y
WFugzjEhUro/rXCEcHQ6qS3F24Jq/ht90SbhJ6k1803HALGCO9Aw/XYTOXVVjyW/
lq5w4/hyrxD0lh4NpaDgVj0ezslo6/Vadfp4iUE/ItD230W29JEs4cNqx85F4Xcl
jOYyf0sjcO6b+0PniT+pG/TBNmOU4Y13ygA5usgb/8GgoE2pEGHpuOkplIDnJHES
H2819rf1hICGUaHk36WSP6BBKdg65YOM4QaSAkSbGV3LSw8gx5CDoDcZvrIVukZq
G7cWdUxF/CaaOwabwM9SyOZG0qFBLX0uW5kRKIjAfTKMXFi/1dpzqGkTdglUJYTI
I09mNYfT2QYDdcd1yySFyh3LSPBiKSBUnu7Fd9ilBi8HuchoBtXwAlqvmV0OJ90Q
OXTkG7lRmurULBs0/RKUD/Z1Li+Zv+2vml7H+eNuO8084yhugUflCtXB8Za5qw01
TbB23OZBdZCUaZDc45X4jUS3qTGYyZ+x8pTkutpeymOQly6/jTi2PgoMwaNsPVkE
l2H/GIPqr8ruzPL4jdd3mcK5LzKrLeKsWypTIeLo+I/0tK3DiReOnVgyAhB7sZRU
uY9WMvde1xc6YujPfBQCe02bpIY2ub6H7YeI49Qt0ODVEqJuuN7afKUNquHic+Lo
zwLidjUZX6t13FVOXA6QMYaxWRyBs5Y/na1DGXoU5ccp4BO/x3VuN/afCXEc7elo
Otqh6Ub/ucZp21Cs1342PPmKPB+icdAoL+4YJ3FUfH4Jbx4AX7urJnZW9zVW+zeN
FbdxOYZzz3F4XLTfBts/WDF5i7mkOIfQkk/MQ8o8HMYlYAI8SH9tsjkcB01uRGfh
waH8kPOswdWfKuxvEEEMTk01z7wdfy4f3iFzN/B4jrrwaXnjqg2RSf5oiMfyzCo6
2e7pMYfjmGQTkkV/lMf6YnKH6zO3FoH6LF8aDW94HY0BT57Yypt8wQrKJlJDyYND
rP2sI4pDiR81fOf9qsYk9EDYdIzszHcBqtdUAPiifH/xIpdmy7/n1OI/bZLPR53N
PWZmiiZAVG5xSknfjyEZGBIdvP4kgQwTla0DKryR141UM8slQdUGrImVgzmiTvv8
Su0W0ICUL6cNIyYO9WJ1yQeoP17xZDTG1+8eBpUB9yvdrgOvcZ3PCpFueVF2ABX1
uJGSwc1jMLcORxsSh23LFK8d3leZURC5QsehvWJgDaoRpLu+t/YBIYzO7xMb1oFg
rsA+IahY8gFkJ9yDrjj2VkAt8ijv5tTS4ozOcSD9H/xS54LcWdj4d/aXiroZNAnq
ZQXw9kubyOIXBkzvS+GuiGK+xrpDnOR6rGRVYEGM2FM7vj8Qe8xE2kwrtb529PUF
xupAROPWHct1xxgB9WtsmFCv8ucYQuLBEW6jde8DECEn68ZRYq0w/dScMpA+I6aG
Hp0LLrG7AJfld22U4VQpZlZwiXJpqlCHV/qTZNwJzZXGZf+16rWDDgU+3x6vGNUQ
EqrmKjbQVeEmJqbJsBq2bwTk/eSSBU2IYR9889Xls4xOw2aI90Zqd50zsgMPS7fy
H0k3h/9dFtRNaLdsev3519XWqAflJnBzdS9b48dQwopH1O2vP8kFjKEKVhfmE/DP
Sca2Z4xF5GoJlffca4Yxg/frssCGqxPR3/Czics9kpQK/QMVDPax/uR1zXPYa2R3
2i4smfmBpErSMsBNPxm9V9QKJD5y5pKnJ8VD2iRTgbqU+VKJyhG6LKmuFUBYNqrJ
6J7wGJvpCOtd/C0O89w7yKoF6AdyQExVNvBwAg3GI1Ysesw150VYSoG26C5z29HZ
2nBLscMpT7s/jWGajbxPJVEXLxtUF/q4slLY+HYr4XNp+JdzPFyh54rGqBEZKbr4
8B67uC4JCIbG/Mw3knnojq8tb8E9ugiJJNnD+SNhLK86xBzt7GpRa+R0PG/qa4jJ
UXl7JpnqCNGtE0Amwuj7elVS/u6gkO/lqOeOBf6eXbvzu0rAPDBZVpOSv5fvPh4p
oJo4zb1iQFU1daX3P6Uj6bX/nN+D1vLa9Dsx1dUXFMWZ8fSkAvUWttVqUPj334/9
yKuAm9LC/pdmST9/7bT7/Os0pH5wMSyWv1fMYstbqgHDeSw9xQqIiUKoWAwg4usv
+4th28EIK382+KdyV+gRQlLTUvnPdfmOV/rNh/Ry+XyALSrBD26ovMUq0U9UP+2T
Qzk+EoUvoooS1ZmDNwweUUGfgLYshXRoSllXgfVF6vLxWzm9Q3OB2QJCOnmB6+fQ
iIZ+PedKzr5ra2mu8PrX4uUctecCmQICCYrvGJYAY65QIuTRVc0gSAzWOtrj0PSr
39cjU/MZ2AOyG2Pg1qUa6lfdn8tFgGBp5G0fhkBedfAFV2awqMtxlH9FR9ERQIgX
//l31+uPkPE+5WheWY5DCUTILv5TQfwkDDreTpxFeNxaWvMqg2RiIyWoKLtP/LZs
dbZctDWVImxriXpO5J2EK9EXj3Ibs1V2MCaQl8t5hIxroHhU4n5cshERGdvjLHW8
XsBHJyJSfp+oDIFwQpjfLzrZKz9qpDz6ZJEyXyhDrrQwmsL/r67z42FeGhnp4wmK
Ovy5x8HMGB4Lo4T6Z/gPllDdBAJ+lS9ge1BCnW/9GSm9KGmHeLx1kIbgpCGAEJ6n
vxrheoI+n9yTnq/Fcy49rgJk7TfOit5eKC6LNEa9JRCmmVDuilWPa2/ILI7e67fQ
KHSAAI/2BdZxKVQsCZitDBZFSwbddRnnC0acEyOks+4CnPlbkh4Gnw8cZ7Tq15rG
OjWxOSf1YDjVmDaMuij21jy/zzImzv+mSzHZEK0kS1vpI6ltr3slmaMtDIW2d6cs
gMi6qvY5eH0zTOG/Rqwa+QGcm4GTjvnBNi7+C007eToCBFXiRtd6uI7uKAfcQuiJ
BtRTJv4fZoSageHEE7c7/pLNT5qfqI2oPOpvoASM4Ic1c5SLNRhAQ5QS2xy7Fm8F
hKwiJRuOD6yifsSxed5IepIIdy3G69Mbcx5F7GHkW2Tim4Awxs4VcdBLfDX9/luR
YvZRrCpz4yyD1WxgdT05WHNI2DfuF6EA0JsFLItk139ASIyok/4kdx+7SSW9AF3B
c0IcftVLpOl91Ra3t92A9oCjiBTwv4qejXefp9YXAbgloXU3WLl3yX143j0k4urt
nx3JCetXfmvXfyMHoKDjePIQeT1pOATaS9gKxmv6Xs8M2btF4K09Wuj1TK5zpewb
hPGjNxKkJHNQdcfw16EZ71/VRCLEkmwJ+Nf0W7ACz/Js6o4r5bZLZJTqDvKu0QbA
KvEsW2rcQas0Ao43Vg13u6lc7gYNMGFVPaCONrvCinKFluum/JeLhIuA+WvpoQjd
49YVvNe+mHlgybgTnAnuyNF22xAuVXzNzPM0oamDTbEGjMEfHyXtB+XlIzvzvvk3
PLUbErNpimSZ7mNqK/evvymJvPvdKYyAekpCrK8QxY7T6cX26ZTeCk6BgPX3Nppb
g4itmuVeqv0tjBodAFi0nJF88VzCidmKo3tf2lwfsRRGWej5Jqhe/maORjbcJqHu
xHyhLG6arQ/VVRCEBunnQ2HFuJcm4Av/vwxcwq41lfXUdFfj9Lv30d7mll1U5p2a
X4Mc+J32kLzD7tO7qlwA5JF5YEk+c9L2NgXbBkcHEX2/05qm+js2IdjSLEreUWiu
cQaBU77HnzGxO1Cmrm2LcjuLDtzSmlaIByBVmYcpQUXv8dPLeOPuIOTZWonW2794
s+EwVu/jaQVrjpYOA0BNO5SmNWP2jQT/+jU1MzfGCsnGz+B7E08BqjCHhkGCzTKv
+s8Cm+Y8pWn3v46ZP44iejo2ylj/Y1rLHNDx3u09g23H/8CHa947tpTZgv9ZE7Kh
EqVeDawEo55A34Ckg4Agd6h9+QNe084/QhKc1jRj4x6IH/AoP33V94Mi+OEX+mh4
OSXTD2DhqMYW8UL5gFhSFMyxHpdB3IMRJ9m8az00ulaWosF/IVWdacuqV9aEDlPO
9OCVFZpC54pztc+ZM3+GGWtWKsMcTGW5T2+lcloKPM5nO3WTqDnyvUcq1b4IXJTi
dQ1RyV+pf+h4fc9/j7BFAqlz3qI18v26X2kwEWazPgitmBrAwXfsp28aa40xNof4
Go6HNks6UPa0eeL7NpB1ZE9/ljp/DVX68YNVXMJukL74+d4QO4+DWtvhvuxAmOb6
2m8XnJj6xkJuNHvx+zUfTXKSrIyHgEoTpy5TUM2nlFPE5jGKEr5H/QJCQPgY2NKm
KMIAeQJADZtpwbDJFMQC22cKnyRgdp4ud7IvhtBdu0m+joQIbcXCnLmM3ku6GXiB
eii8CI8pJvlg3XpI6LlcXLM6J4WfEYcgQTMcmNnuciYhPQlqmM4eQADW18nzIwzW
G+nynRSCmBZw9eQuWRbnczaaenGBToeQdY4uZBAZQB0yd8luxiHoXNQEHo53h9hS
0N32P6+xqFsHYQ8n3HcTyr5cwLROuW+pW24Q3rhw66tK1VrnZN1wyrG29kciOJ1e
+kX69v3NMiQICVrlNvvJfzoxwuOQoFzvWxU3Q/QYooBa+zoHWH96dHoDcSfPQfgf
Hp2IDrbG4i6oSzZXHjYrwjb/OmigytGdPaVWMscl9Bl5Cxtvy3nyba/kBI7VJX8C
Tr4OaH5a+I5P4k8iz0jrsYfbjLWN2Dohaom8zaomCs41BmoC8UgTgHMK4fja2u2h
x9NQfT2URCC36LOQ6/g3mejrsUNyFqr8n6M31mKLzmpQwzESw8Vp3nVyUu9cNV7S
dZDP7b2LzjQovlB/HnB6fJXHQw3XZQ5DV2XtfEvUOH6VW1bwxgJgaxVP3kEa0yq5
yw71eaClCdyu1yLxPh8mtebruOMa2Nrb83CpJplbpnMjtYiDJTjSmSUAlbBVpKDN
PZ0ACO+vLLwsmFFqvaC1OPWYiyH6Epl/42ABCbGacy1tQGZ0HFWDlB4VJ5O23q6Q
dkBzHDRwZzGEBtIaHwNSQ7Wlj0z6bvmRA6G2FBOndrM48HWqQNA7nQY+6+hCZOU3
pLWEJGvu+SNBeZN28goDxdlCpcrQkgGTuBdgedNBF86d2BoF8Xr3R1JJV/5zoQ+m
L1NH84QMQoVtV5gWyVOBYpKI4A+CakjnxWupFAGHvFQ33MrXpanHSyqeZKmylELu
ooDMmsyR03/nBde3filK83fCplLk0EAP0nFabGWE9BNF5ZtCCDabzv6sw323DNue
CcZvPk1K7EEnHqtj7fiU8PK0Yt1oT+DJHuYI9QIvgauHlSNuVQAByfdXJpv5tHnA
rjOFXphCzOH4NiojUqeXf41ulAozPJwhm19vKpraFPKdAkBfQTMgS8tgd3pRR5Am
Xa8UjSj5vVL2oLUdcsAcGh8brvEHJ8eMWRaL74iPEwLwndhR8q/2swmDIFVH9LVU
ryfSvOar2ifswg0dZCg1eqLe57tffa8TtKULg2ROSSVK9rM4iYX3JznDxUy8XoTW
1mmbhs7J11GorUs510GlmiLBCG5t+H2A4R85u0Bk3EV1XPkd5dinI3/YEfj1ul7B
vBtYPjYegG524fgOrEO/qtiEu7UV5nCqjgG8rnrhiUo2lmn8bCj6DhcV96TWBs1m
ZBQZo9skOrLUKSg5QmmJwEoOQEgSwEbSIYE8s/ibxsL4vbFz4/fJnBrM0/KEvb9A
oQN+kGjgVNOSjc+kUC+88p3+nlYGKppv/QwVN7g1fErGcm3JhSMH093rM46d60lb
6rUgZryTJPHh7xlurjh3pWdsc9zcHQXx8jBxZDluDwuZMprFS+QFGwaYGTAD5CqB
PbBL+k8VJeuZ9WQ5RoVz6vWC6qubNCwPHVt4G+98mvWFwR4Vfiko+X5kxTEzriU3
8gosjB7q7zvimWojARFfEv+ge9IhqPkj5YtSAu+eazMMu6gJvI93unz+00L9j9RN
8Gei+NI+Ln/0Lx3RhmYHV0Wi3AbjGGm7qlNPwRDQKaXH9z6W0qJO9IP0tJNFFyT3
VbtP4sL2C7btS71jDIu9piUF8V5yD7ib1fdfZK1LCuVHs30W2uFyjmgWbE5U5Ypl
2AccIl9zEx+46XHuI1Vy4nd7cX0ctU2nNihgkhkk7CqUTZQ5icBEfdejrDQZnqbX
fWjeWvVayfCQl5RM8/ST59Jb5YNqj2mAvMTfOiIpUH+/Bw4951burAljB/O09ljA
gvdfR2oBOPahVH+B20iHJHslhfGW1BvptVYB07gLAbmd3P7FL1QtnqRraJBu6SwF
HwMSv2nRpHWtd90MrJQOu243ygAWvvbazFlDolT6SsCKespaUG+CzahFQ5dL9THv
4K+5TRVbnbuOswxjayFj0mxKvIJ0A5la3YEwB/aRRS/VaGSYMwgMPntbxjV/Kadc
lcqd3C/iCTbZRtC36yudNRNziS1PkJ2Qo62V0lz+0nHiD9Y7pbDl9OhwcjVRyqLA
rlLfRySN/GDsPlGharO138CxhCkKq3IAPKCI4akVY/X/Qx1Wklx37ipHBJ/VKyip
dO+khrvDtnITbADvwAaodkNwwtdHPfvy+KbzaUoinVWnpkjMfdh6vB/7AZuJAh4z
j0E1XHAAWu2gGoqCJK1qsuXef9l9sin6DAiC7EiSrCBOxyJVyrmiqQMlWMU9Zw1/
sbucNQBJ6I0+6KDWaHpLhEqbpLJprunvMBW/DxmwsY/Eta+t55TPKcgaYzA1J/JK
5ykZwNstawg4/hw0nqsuOv8a9Isos5ZQYYnsQn0Y9la78Pp4XJFZCf+2nDJCpo8U
V9Rf6NLrB8nGbE8Q0cGZNP7pNoy/wpoGhODJdSzi/B/4iWcC3tyK7udoOL1M6x7v
ACSjSkKCFhGiSgGmabmq9TxzzOnOOgm5v2eH7PyJ3CZRYb1evld9oNZ92DsiFeHX
qR7kZawCcWACXuVe1k65KHlRL1DIoqR6O6cKpl3Df3tmq+yE89CS2bPNl5KTomQD
X5jRqkMz7kXKT/L9XaLljvPrxeCx7v7Mom2zTlyTcPn1SS5GKpkyo7ofh4PbFUt3
GMFG9AvRYbPzy+CteyyloLmpNXGbgLhWZ6OMuwLopBrJfgTWXNrcA0q5xsMK8lgp
JN5erKVYsl+dC2seN5kS+q6FZENXXfdFlJY+cC+UQEhljINg5xt+u6G05aAlHwOs
mDwrrjri03FbI/jYpuushET/KoX9d11r4shfJCP2vHS4tENWxXSa1w+9LWPjULgr
dzykQkgTUTbx9VZtPigQNf7HTxrHxGZMZ5sfMVTKfO1uxCKo8Vn7knVlpkUeWSza
cy934ASwWZvLuEAwAVOrfbigxNo54NVoDqqfB4pXxL383U/rX1fUQKMooKWZ+ZK7
FLS7/w2oi9R9k80nhuv/vtpQSJsOA2JqTPsdI5o3fHLY9mcn4PZY+slt70fsr5SK
u5qYQTtJuTBfY3/JJ8AsKizg03SsmIL/fxO4pKNoc6gFFg+NMPceCf2b1sBH/EW+
Lw4ATm9LqqqKGbsNmF6Ac+pRqTE5wUrgbLsvautT+HSwqqB60G3k30K1IvqFFlI9
Hp4dH7lkkISvZ+qZv49gAm7gto8mqUqvto6Z45s561VPcpb3w1ot5apgo5bupPmn
c/X/85HIp3mWKJcdRmbyTmCtAJl7ZQblDt/LSw1qDv5Vac6eu5ZbOAXUSq7W4pw0
UEjeQ2HXh7SvxsI6BtqemjBQFK/WOAZR+qmg7UOYaWAI2lU/JYLux0YQi4Iw93ov
WDS/fizYblFt8nX4yM6NUYOkCBnPyR6bA0Lu3vV7JpoOYr720/BAyhVPaDOQFOu1
Qo9RyPpLYFQM4VkLL0NStLtufsthAj0n+hE9bjMzie47SpQvD8kNfSo6ZhqjDLm5
8aUrU02vqsWHbex3uApHClk8UTY+2Zmt6lgz5S06ab5T1UWmEACymH/HDpFoPPP7
viH4FKynl0nnNsATkpGFAhLiUisZvqYe5Zj2Ch+/apDXzSPwJAWwBj9OUFkd6HcT
Oab3als6UEmGzx7abVQPeoUG8mcUogwAiqgytQIV5p0CZCOHjOC2B8Ah1552gf6E
35akOnHCRsZDaI7w+lguDGkx6848jlfMbzYjfcz4C/ZiBTA/pa9truXUDcOPLY8a
8zBNj07ACyXP/p8NuFspcZj7W6qWDmxoKp47I1fcKlorz6K1YlsSaRpNMenkppDs
umY9ypcZ+8YVvVO6v9Uam+Qd9vbsnOFXwwVUrfacMixnC3NkZPOTrjL0WjOWdqT9
CMCpfvJ2ueuf/kcSvvy8yX0vMGXJ2BZKZAXtG3/LolflxKyIx+1ztEZxOUrTrBI8
D0ljjrzlzZrPVrgnOJFC/I/+zo64aYP9vmKqjakjo9bg9br4i2LwD2+TeYsHHcCg
PTN0Gm6rqvIoGKsXtyTGYHUTr2ExsPXQpF44Xw6Out9+MJSrTkBpFDC6JqQgR7GQ
1qNdzF8SCXpvC57AvfbZhlheLADb/zRYCs6D3hMIRW2yEJajijIpxJ/5XRvLzwC6
3Kl8K5U/mfg2oe7kGTZA0f4HCJOguI5MP7np46nUtWjELOt+Ass5ma4j9RjZpHgR
SHZOhdDDZ3wyWNJSuK+zBgNb6XQPwsTZ/ITtK1kT5lxl6xZt1LLsW3IzWlJBPDi9
bm/9WYylg3xcbIz1M6OjLDdbigko56Mfk+/cPt97aBkMZYuU4uVqmE31+INEcuix
IUg06ymfxjcb5spCIIF4l4jedDZ0s6gw24wGtL9vCYOKjN1A5m7jdcdoB2mdVaL3
T5kgB4/oQnoRDO7WutT4aFlNM+NkXmcv4Otor9+xeL7feI1OHauF+ZGf9655fB6F
Liy0M3gFipCXhUfFQA9LJt/2rfD0tz3HXLymKCkK8bv6wj8sgovPdYIYdLCAHbwI
xwdvaoXivoGOr01RVzHuTlfBXjDW5a6PqAC+rMp/2NVXJ6d0Hg+rm0wbcQkUbIaA
7S5izgUUnkcih6DSmV7BUnlR6pFUeX7X1KuFKPep8lS2QcG+GHpKsxSNMfWTBX9d
J/Pbf9iMc07PIPvS+DmcqJB4UfyUc09gZwsnuQFOpRIICYBYSpOTulLKIJ0qhZG9
SAZ60hHG7j0b14OfzUmMGP9L1AvXVzRM+vH17h4nTxLbNBaMTMSSSgwGZ33dHGmk
9Be5ftG5i4WOqaLC9UifdiJEiykTAcq9Y8VP0/TSiOdnkIfvPWGCraGWAfGKNBJE
tJZJ70AcgpDhU3AzQeaMwSpqTvsH0Kc8DIOxW+TxPFFvE58KiWuk0VX2Yp+8f7yF
RS8foq4jqDjMsCx13DC2yTLQam0BtPRmoKliuKUCvDb7y9n2Rywrm1taPM/4Vo1/
vuSfQ5JVsb5vPrO4XjffX3+UVSBIVwmgC/7ttSobTLYodr+j28rOAttiFFKxvQ08
FzQdW0xYyhKll/ZRVUx+Cv8+h7lFSXxcN6AXJPSlegPeyUVn7NVuy56sqOU2d+k2
TDll/KWvmO3AYTyTPfL6beGHUQwru60FU2VWoQYHwkQjUKp+BUbCQSMFBC9OHXQ2
JRtQg9QOJcX3gQ1lv6z7g4alSWMJhl8VX2q4Bg0wOYNNkdJbPiFcjbgE87PBuLlj
yJJn/K+rZXjXuPdpfQRVJelbZQAe2B1knjCEhcWWTHVklHH6sRwdGBsyGln5u6ji
kZ5kh7t1CPuj6ak/o3cY+Qn5e4lLOMbESyPlN97AwaAAyEKModJ7EGVll3i1acQb
Ja1lQquyUd23nxPdfGyhqmQ/SwV3t28CTEPiGJ3nO9x+f/cvpLAAxgvnCmO0zzEU
ZBBeSsvCyq+wnZki/0dKYKCb1QDv46uab4MENPoXahzGWQkkOyQFG+Dmd5I4GIat
xmEILWlyQAWl7RZL1r2t65uexgHsGOQUNUTkcDPyVoP1T9CQuMwjp1t+bsKGQqzA
Vnk2xxghUnXtKpFb/quqLYlBX2CPebvfkU28ASgyLQTa+39ERSAcXxn5o9oIpRU8
lvUbSKsJ5vJua1BoTXRkWaclCfWRe/AFHkYp+DIz3b/olBJZMQyhKjW/XmofROC5
ntmWrfgmraxucWe1ZsvEJBnbIYSLwZRksM7fVqkDyjjuKoL1dFd2GM3iXxntLPn7
+BylXm1Sbbky5VvhkR2fmNdFp+nVJy6FmjTsybuD8HjYO/LrMXvYyYu7d9z1DXSz
nm4RtakOZsSQm992Oueml2Ct6j0/5tEp7BIYwm4oJkM1IOf8TITpO3yRb/NHznwk
KgxjsNGvMoJ0jfKVFq2Zun8sZjFYGL9MzZSO4nixKhggufEB5bkRZrNhpOUHrY08
wZa53scqKhDIY0kUTVh6rH3y0bGdH4OAUQHMjDU8sYW/xSg7BrOG0LKsLb8lVNUb
qWaihZR4OVc7czQ+XJacJqnU0zsEQM2Td2CDCTPT2v+CcdN25PwRB1hUrGzpwybZ
loUYzTzySabrGO+vLE6gnYy+kIYj2Uhc+ZfIY/n8NlZgVDx1ljoGwlUYY+/N/4J1
77lZJl0n80bz4c+pg45yszanBIvEFCmi9g6I4uHB7sXQ3MHQ1RHq0vPPcbqr/x6b
5k87dxALL7e//+becOxjokx3i96lPBz+wrUGffRcj8B7AZF6kSU0yDr8kzzI1GVO
wOd6X05WGtcwGlcKjiV2M//wzG4OlkgOxOqW2arvaI8sVZ2iMV3f1PiuNfaMBfFZ
6bFQH+A2bH5xmVAsLw1hgNZroIra929DZo4KV763ja4shZLeLTAfuRGbl2oIS1BA
U4uUvdzyn08d70n8mlI3XnzSBIYu9u7vtA5eqbQy2T0nkespoF7qV+DZLjZzx0iv
50yZeAz3PpuMFgAGkwU+9T3Yqzx++NoMTHbRZW7+6to7Gst3fOx7aWQduGnBMzui
Gc/OoYz/AY7c+Z29W1Kq8zqeXGSGE5TkKq8etX8Olmjc3cSzPFBTVYJnI8mg7rFo
J5FB2namBYfXZDEdWHoxaGtSkbNi6CbzhzwyMz4cAvbKvGK9EMqNUvLSoQh8kXI8
wMrid8fHexDOBHyzGCSykDIT59mW1SKS5/XK1uVJ1zCVBTp/bE5QaHfcjlfk21VK
Xqn+IZ7Bzm8clc3xVsxlRcaHDLFbTNU4FFJAPnsojSTJKoMLnSLVKyBSuQQzxCwU
Zz2JGwcjokOiiOmudJpuL8XaQ4n4r4EDrvXjm654e7MP0ldgGZdge/uu7JN5Krd1
ZkP7rG4YPcmdN15g06cBOu4EsdZYD8Ynxdw9t0O8krmxcHdPVrfN6P0iIWfsy+zJ
0N8DK0jtNKkMDEjHv7184tsB5QrVYnkILbbdmTkAFGj9giNxcO8OBy8crIMjy0F0
PiROvEM9n7Q/bpO45WVkn8Zjl3fcJjA375+RFr5qk6D+FL0XcBvUdOT+CniREKUo
km45I7dCKFYX+fOYOKcJ0llXWN/16fN1ZLdd8SHGNPkbRhDvjyS+GjvIt5n3i302
8yuMURkLXWY5UouVCuY73jvOeOP0qqCQTItd6MrEoGm/AwE696LL+5YrhwRBi/NY
Qkbn+629bGbHci7IBXziTaYjB4Wc+jbyAxrrh9A7ut40BB5dGrriwn/AYTWyvYFa
OevaUjmpKnvHdm8d2EGLSgvUaj6V0gbgkouNVivutQ6PUMpMmJbqr5BtpWFnjTeG
UWHKG9jnHwuea5nc66UFcGJqQcZfm0PnP/TtIZl1gc66tGgAby/MiSZ2Hky2mBQy
qTSZl++5dxq/j7a8nr+ViiVDW0Ce24P2Adqcbh9Y1yWVAq6y4BZ1rQZfLX+qEAzQ
MRkkWNdVyK84ioGnKc3GK1+wVuYwclHwu9Dney59pHy/F2BPuWfxLwxXxFF/NiHN
ROhWW1Hxp8028YDdkc+yTaXyHR92FqiMToBHTtEd5W7OgDl5WrrfM/FmAtA6Nc1r
FSTMYd6Wm0+8mwTkm8F+K7GaNZ3K/mdab/J6ggmnvVt0BZfM0BxHXRQyD7O3AOMb
SYfvhvUoAqVM1Cwm6awPKf4qL6ZC2l2fIgnxWFCsaYYLWvwG9PSy9ZFdge3j7CRS
oYQSMw4fdpQ61BWZBxA5yBNpqvEaFFR7S4T3Z5exIXhnPftOwA+nwCmEXCZncENp
kdKL4vF0KQeKN9Ubz7M88AV9BghVRYY48pWCNZ+KE6ijVKNHVRu7Src+R4qlsIWW
mg9Zkml9WogVwwlArwoV9zVUjBrFn0c+M/s3Eor5/TxqJ4Q8rNkrsEhWo3QCOOpT
5JJF6AcWE3bR+NuUH5WK1FCaxFYTyZRFG4N1nux1kdk6K1EHQJKZLK1f/ffViu+n
a8MFsHlLQIU2Sj7jdOTY10vTFe4iNuwBQGGdTRV0wdUbH14dKcKBAfgoK3MLzbKA
qPGEmBeoqOS3k8zhYC8vNrkP2T30IG/zdzCsblX4SepxshJ8N+b1RHoE4yMuoXw/
e+LCb5j65l036Eg9o7O4Vbbcan554c+eVHU4p7K/RFWWpKbC+lYAg1PsiEpbLC9r
I0AO9GwFcqaqLbGzTuPAJv3eNNYqDqUXiVqUf+q4uuaGXifzVs+FIsUSWhJZK8HL
bBGnlpf4+8EGI5LD0b7gpv1Ti1wQiVQTBTSLlgm/Bp7cBqKquskYbZCEBBN0afwt
4Ohnl70jV8JhfUHEs5PbzSmlhzBrMd5HUioFI8Uj+aa25S6hTWvT1Z+6h5CNcBlN
AqWmkZ9rnxREpunCWCx6jiyHo5od7Zptg+h7krg1x5ZwQkn1LSp+WtaluKSpqqcl
s+4Xxp3JXLoGhPr31X+3QRYhEd7zuWCXVckWhaxwCziZKA9U30wZfIMmQ7VPGfLI
iLRDE1lRwqM4FSvoA/xQYyHvMNdqSZW7nDoW+luOfktLyWmkJUNlCFin/TUB2MTJ
dlN7M+hPH5sKEcWOjQ7yYsS2YdN4xjgtPhgPQu8miKWP4A3/SHgrImNTymgs9wkk
I8rYGJY3QddxIA7xMuWG69i8be8WLnZPPIDgingaBxBLVMMeuC/kd9ZnkHZtqWl9
XwLXo66zMw98CSetk3fSMNir7COIdHL5Xa9UxJVc3It9coeCcf8+nGiBgVMs5HZG
W8YLMT9WnD6bs28EykQeloO7jP4ODVKWMgpeEnnlha2buODGq2i3UYmNifTnF3K1
SE0Yjpl9/jQUXZhukyPZwMlLK5Ik6tPjcJnXrGBmOSfERvaqOQxzq8YS1c6VPbA/
A+d8Pnji+hnLxH+Zt0E3YXLN6vazPoMXhlGWKLZcWTshJuisiGwnU82gYH9+Un7+
N7fQb9iHcNFX9eqK/g5r8MB3HgjTYRlZZbbRXUgxUguQCs8K5Z/pAxa02hcTFMBA
4FI9ayFACI6FO1GTRleouwuX59X86m+0NKkUfTTIN/ssS4MjYtjQ6m5pWNa+kwYi
FhwMNg0lukR9nUmW0AOYxAGemdNI2K9Yc+MRqDxZ9jRqxvUFqJW2bMBMZvF4LnY0
Qah5xDWQV3MWrnuCFDvkxbvIYbMIKONXN24Jp1kb3wLPAHpajM1jM5/PaGzFpnlk
eykikkViB5fRDgo+JVv3x46TLDml+OirJreFOxkYV5ozoRecy8SZEz2dzemY/bsd
6N8GOS4/z/FWL+W5abUxASHXi1mki18lIOOpjocuPNEMF+R8ozkNFr2j8HN+e1AT
Xegtcg53v704yfTkVCjRdHaESQqLymUQks/HwXz1aJIyCJ3BH1MYMG3tfShTMzs0
MPsY96BYclreMMR8pJSouZHDuuWShwTC4CVR/1WXCDunoMZjCy1WUVf9vJ44g4yC
+/KLLguX0825hFplGNdp+7XQM+/vkwEeBnYa1OAlIy1qhJkRUuukvXMI2u9hNtRn
k9Tl/q62bTmH/8Oq1igSNJ+F2vcm7pcmoouOfywJDE512qJz3jOP1d59AxkbOHrP
aIFDcTPQKS/MPV6qnY9CJbEHrcR8EGhh0YrbebtHIDfUL/e/BGwegbbokVvKhs2f
K6ZX0c5MedZPD8YRVxGfeR7XELBMjbswIqXyyDRhOnK66M2RYPW4DTSmv4U0XzRA
h4vp4UH6wKndXluxXNEctgfSDjKPQGXdIVrd4PQpR2oawXRTEi143VALOZbo6HFs
c4TxbT+mVfTVvO2kwFRerc8VLiv6Wwb2Ff4Qkzdokd+H/7ZyP/+uv3cVbCVfq8ZN
5rOwQZbeNEbDiZDm8KcTigl4HV+k4lVKqFoIgbqJHT9EgEfVTTfnamAfx4I20oc/
NZ+fFdLaPdxHk+fC5XhO2hMyNSFm8SN3k+JVGJAhA8Gmjs5ltANQ4ndXc1ylj3s6
Ymx84tLLeMQUa4duuFaqYamA9n7DHQBHyXRgiup9H3AruDKP5b8yogY5+e93LE8M
hZlYvATPS6XDNX74SmdrLCs7MY9dYd7sDiwQ+vL+sIWAq2/TySg0d7PDks5vDY1o
hVFVNIREbg+Fxh7/saZ6V/87Hyrjh7bJ2aR8FU46LApHGGceBlA+UaYuxFzP9lf5
evuha0n8uN7dn5Mpcp4WvPvxPVDa1OBVtivHwuboIbj5NYaBhAwJFQrGrvgARfKW
66InfzPB+eBSkm6X50Tuhi4rAaVEmX1uFMiH1EQS3/UwMxMrASzFTt9y6lVgAShF
o3lkfwPSd7lNkeELjF5JVniRfr3qbcn73wIds1prjZQNGrpurp8o+STwwwJA4oHq
Kh8JBg+h3s7byjUYNSWdm2HaRDbnKLl1tGzfJSyz5Gbx0yfLi68V2OE4MyHN88cA
0KDgmQkTBN3rPNV7Boq17ttitbemKTW5X9qQiQTZKhICkm7EujQFp/J1MRnVcl9b
CdvMvhHK7UljKcK/3g/TaC5G9qc7RtU3esZDYs/ceHjB6zo4MN5W2PoGMpPdelML
2taQSZj3388gyhTIdGzqFnCLioooIeYGYXMYkBeITwLvwyZlpnBhH6RWHyXNrjpT
wLEJyqbxFdjoj0WIq3Y3FXbdmmrp7g156RidHThw96Ejt2Js19K/JH7odg3J1Q7j
bgGq+Tnxdr0STZ+qZfiW8RAK3UBA6fXBCfHNYyV1z+lFeRW1ViATTJ++ULEKedNe
8zGGRomrNdrGI80blv+slYZEnQjOh6nxn5fZIuHzDl09LEe5AxWJD7US6eoz606O
NXlBqhYGTU53KqwV9Gu2Lup4a472HR3jWeffB7aMGrIZCLKn4keSp4e40qmE13VP
2pteJb/rNfsNoaGzptz3ucIuOt/Q7/uoYBGqw9OniC364jm6gjRsmY4VGrvbCZ9F
R4IPPiW0PPKholdYc0QRo60unof9ow/sGPq8KKjTKtB7NEztVBokY0lYOfc/Nwxj
dgTRxXA0d+hdPbNJBu73B8YDJC5C41dvbJwgm3zwbJBgcbqliWpVxVzc6h84dgDS
tW6iespzeEhX3rRTC6UMaYSYBjU7Opksca/2YPDm98XOO/4bEo/OUCMjNevIe0Nc
TINC1kmzLrrcq/AA1LAWG8pqTNGUBOdSkR/cghDDUaC47PY9dsewwoC7P3NbDCqH
/VWPASzeNy9hQWVFoteXYQMXjDzuXjP2KPzReIw3ZtUueTJCU6ftrd5C/6pnvRZX
xf+lfR5vV1yEMYqtRDyZq09biFLxr2lWRIYsVxaCYkZa8ymRKQaCflRMp/Uc7o8P
Y6an1xfa7/YXzRA22rQ2zVsSQisWgphftDR/IpoZkaNHi+jxuPZwc1l5bAqrYNZ1
85omf602roqfcKPB1XI01zMF0kxUXmEnN5S5w0QHqBh7JhPSzo//+k7nKzkBhGI+
S0O6sKiF7rHeLjc1DpfgLYxMJDFgQXWwSU5ZvvQyFzvOVyKGdT180DJzCswGVIS/
/SNXYMza9qoCOf4yJZpnfCs071TkI47jH02zrbXSVTfh5Rn8Nk0eHflEwheeo5XB
WXWIxIlRGLKLB+xtDG35VTVdWA6ceuvTcxIvAR3RUXCMyPSLcyiFYEQacdKzQX6s
KbnLCtaLHZR7GTUE7zcRDv5Yhqcqhv8rUBr0uqvB4mmWjNEDQoR3HkMfZXeNKtnO
5oU4L27Q1pf6P1ZKtUK0CFK5Ssar77KhzNDl2x91Mx09QDR5JI080tgsSKhUQAY7
yzJcAqVtN/Dr3H+DoG45UvnAyAhf1Jeb1e3CjViC42duVop2fZPcwerVg8bTnS7f
SC5P9k3rDhEXpjC92EQj1kv1jcmASGWBb46MFjYHf2ne9abVGDG1DM3KppyiCzxj
Xm6XQs+pKJVt/VPktmTL8IZcorawQEhNSSTvs9SbuNmpNOLWwAACNhJhYijE0Q/r
SxnF4IIcrqKmfBQ958l/CIF3YANi/KrpR6gJGWFzXL+8S+JyUX/8LdsxVRbQTG2s
VzTC4gAKKBIXJzFQMlhKD2Oepzc63jdXjxXkYmykU4mRrg66OFpvRULjdSZb3tdi
1S9Gon03lYnV/pkcKoqXWm8rSkY+3grVC9aZZHc9HNa89JYHT+YSHtu6bquNq6Nd
zjiuklaHr9uEwWb2EbC2rGXGa28t2OFsCZmLEDgsfVutieTNvohL7JqYQ6rVVAiV
WOrgVfEAytzgfIV08rx0vT5JzTM2KAz8a63RiYBmASr67d4Rdaa59MT08mhIn+YG
L1DIzOI1IJ2q/EMETWWhDC/EGGaOKWT+k09CpgZtgEl1vaMMxMDfCTzHDRUS/eKq
k/CyJBi8dQuAmk0IRYLn2jIvqZooxfnFrkQO0abjEH/XGDTXply0IsRJkEXZUISj
3EwGTjP3dnSJ1zmu/HCd9dOjxXyT82SYqCXNVCUNSmX88Ib4zoFjFELQtD6Nf5rK
37CesCPEcbiUSTMWPyOcUlF4gUvF9PBCs3tSoIrz84WfmbpUNa5Cw4/hJlVY8V6j
GUqUx747gtmnYquFfyRoiqAUmuQSMdFPP+LUwlZir1X2R0jqNAtcfVR4Mn7hEHxO
jjPGrxf4aljRQ/d92+SjKjPJbf1wkrDfhBRg/lyecebnXlMyF7j81+r7gTQ6l74T
RDSFiQD3j+8Tz2OTYbjAGmQwT/9wRNANNWIXE9afnAei1IVcT1YavWwL3F7mNtTL
eyB6Gv+uTXOFmU3SybeO3Qbeu8ywF8OGny1+PTiwLjwzXF5stnruPpmTHKZALaTy
IveWS2lvcInI2UBAnaxU1y8k/UchgvUv9MU4fDNiPTeUKdvwQdD9kJ8pQ/EKDZEZ
08q9/sKqOX261FQQLvFEMHBXfI4LnE1MWi0EtpEW4aQc1xpWOt8VwyxxTeupe/NY
Y0Qri6RyBhw/GxwfRzyRDPji+/aayrSRv5NjLnB7gCHs5H5vrIhlGdM3NjoT9PuR
/QMUEgid3cjzXQLjKSQizvvU0EOfItwfLVW+kXDLHSJFCRZjZIiaWVoVNaybGxt8
Ce5CUrCFsFWMswmFtDEzyBhri/WeWZj8imbll/oa+miD/FENH10O2a5ZuCOpYVF2
xk9NLIOV85iVaJf7v7Dd8UTgm8cykBJoQh5gxvEjSMmXFIlT+QNnSBCSIR1UkZyl
bGeFC6OYDMOanyY7sKJlurThyBfBdYifA9iZXD6jA8PQE2R8GjFkRf3F7nTMrK5z
ZULtNph8mrRqwoU6iWTPCe41O2KBd93l6zKG9mwkwcII49XQQn85BFW3aOtfTnNi
QfIu0vGGhCBS9hyfxXq2W4dlelUD82GQE0aTcadkIY/zjO5vcFABQg7r52LdnFXg
80WeJSKQ1Qkyz670Cz0tHFrzA7zMq4AUtLs4HmJMeqk9u/7gotWVwLFEtMJRzqCs
ooFRB6/3KFICjST4w02f/OT/jbJBA08BP8YSq6YcTzfLVHbEjzGF/yg77ZOAUbjE
SZrZYlfiTPIncMlM3kP/ywTGW2DqTmLKyKM7Ub84V0AVdQK9uDjuuQL+0dh2oxNH
ln19wv/iEQmeDXE2rnes9NGsqt+jlolxOfEdfChuTcSAHb2tPuomKS3xjzNb26vC
8ZHh9pwr07vFGdnU0lWrw6BNso48/6gOXsZS+OeJiDSNzTjpwSIv7ZeqoxOXCF1O
01o1WtmG4yKJubYrMfrf8fzDK1vhz7YG1o9en8XLaHatnzVJg+bgkefSEwVF6rvs
ZBWh8N5uddQ6ZQiqtJezIyyW9ALDk8qTZ/KXk8UJ/KxAnRW4vtHtB7SEAMTOdSXn
ewk3o+YqB9TAczV7XseEQ+JMHrz9YqL1LXyQxJBi8gcUrir865YfE0glgjWM/tgB
Ph9MQutXAoPsBcU9TwPVKQTgEquAF6jfSxLNEO/CmSAzZ0+7nsA4F9pThHfsYx0z
9eepCSb133R6wvDDBQjf+lUyttuswfOCRsJMR5UtQ/zl7edjjLTdZsA31UvOpHOt
1Ggc8z9tswio10RtY6K27hndTHPddZtWjbJ+h5QwZAMErmkJHL8UcxymVuQJxdpt
1F/sdaDWGeGBN0kelUffMVusnG7bnTsR/ePJERcr9ehyWmmrZA97wa4b2yKYNDzy
KbRGnz4glX18XFxDJW5tYmobglrIhXfrheN4+/T74j2LYqoSRxO4n6um9TiKBsQO
gjZbmJIihgrNvRp04/J6LI0CBwtEli5D0TFYn0Ow/1Wqgabo1i/RfcqmCl5eGyAm
PwvPIL1pc+p/dpt7fzZr/uieMNgesIdS7VHLbWgzJI7TVVMw1M4Iuqox/Nh8DCRl
ao1XD/T8dH4P4LhqhKCaVImDFZqrspJngaSPbopRYoKmW5ENqBpD/DD4V/W4GqCR
2qvtiy/pXL6nRfAigMK1M9H86yIvRIbbnEjqVeNA0gdhFAPlvEZ/uGO2xvYwJoHR
oZD7Rju/FoGkJBL1rggJQg0jLlgN01JQcz2Sm6SfrxEL/yZSZaG6DuL/SwAA6LmF
WKYfPBGd+tqqFGKjcf9DEc37WswIxAuyVDxD8bOcC7Jt0boRnnx/Efu4aHuitTLk
HUUtJYecDBHOOr2hNo4ifAnBsuVJbziH9XDb5a1oUI0iPxonx4v4gOI3/PWHufhy
/U86WCl6AKghcn+CRMIu+0uM+6B2DxPBWAL1ikQHpWAZWgM8nzt79OUAP+R4tZfZ
tdNhq5lzzyfFyMR6+F2c/LXG4V5AwKhqGpIkF+6SAwumVm4Jp8fB9DGQi3mBHYhP
i0asT66Oy/o4v64DGgOaK7kOhisbq1t24fS9Umj96rywwVZLkcKlCGFkx+tzQgnh
3/HsI+BFDdy+mDzUgCxiR5M1vhyGirG8O9mNeoPL7y/QVblBzLIrd8/SL5/mQS1I
RyczujyCUI1qMWn+M6LYGAaHpwpZiGke3TmeZi8kDQ8ozzPGZFgNvmh47LHZyfaA
H05d6Djdz2JFk98hUMNCU3dKQ7z1ZdMXpsedZGdJvfVMzRiDarB53lqVb3fSHs3c
RvQUAyDo/Le2ewJXMTngqAihHz7I9sAQSxUtfLt5LF1D6vvJ7b6Km7Zr6b8qyO72
T6P25Ym2x05elEXp1PDwygT5S4EVUWeg78ydDxnfGHom5x21810svOtKnqcMsehq
OPgyO+ZB87iV++noH7kUkfvAqmW3Iuj47jiP9ZXq0J2hOK1nkYNnIhXglo51gw2E
9uacgP9l9lJj8EVDV24bPETMfiAcSwQczJ1t9B8U6oa4jZk6scAMInQM6x2SkBxx
+KCarzjHPVmG8y4E15XqLjrA51gC+U0eWIjUTdKePkYCW+UMEqj6NWND/9vEBua1
qQJm2jgDrDrhmooDOBRlgMySu9T4zQ/o/sUyyylxuM29SdSTQbB467jtO76okOWl
tqdC5/EjdkyOtkd0WusU3D284mkVZsqSmUXMwRH5c/UuylDnch/6QQUQAj+mLTuC
vE67IW4t8WCSzXcgdF+YrLVYE0Vi0vc5mMvLUxkzBg1WPJ5GXGxLXUG/YZX13Tzs
bQe6V+Zmwo2ScQ9r4okEenkFXfTbzMutLN5tQD1raOHQQLqO8qUc8uo1t3BrfGZ0
7EFWjz7dZUnY8wALKC1xX3gtSO8rXj4DfqVFg3rewx+pWzKJzyYP/vRYcG0J1DF+
dpvTiPZcAm+RMQOnkKVIypAShj4K1v0BTRANJAyz5VhD++atSShzPvICMwJGzCjm
kIxTgpggQ///6TpedyLtqKSkR7JIV+SvJ23lu6D3CUNAn4jH3ZeHOMrm8a3bIkYp
4Kqi+cKg3VURU3NquAeQCMlzbYsMUvxpv1U5WNsa0ojHllPC4QRDA0hSWwWGrWfY
YuwWhNS2T1ajPM8fhf8EloQvrmwhTUD2TXu8Tt/dQfWalX4oplyhHHTr+jo/WHSW
OI/XIdmlWJDyKYYRbEPxS1w4n0o3qmY+mBzH1yhMgMFYgGlk7nkiBXoYaDK0/8mP
reCUcE2R91qCjbvcPLiASuLDBJ2d2CoDvcfhRGiSTPnqTO27eNLsugu/UibEmQFD
VmlbJXF31wi0JNWpaDthEjlqTkkwFCx/eT4DcR0YmVqoyZe8M+c0p7tAD7TYhuZq
ZD3R5Te5miIeFU4aPOYnKupXrdjdM584z+TnY2D7EH4DSpo4xLghITox0obvrHa0
mkzOAobPKjJtJltKis1o/wSY+txJck2TDa0UDHR6num8I4UUPj8sOiojzT+fIVAA
tXwU7sW61jLoxczdPRaf378QFkRTQJoiGEjochWqCHsltyQlPqHuxy2rUNgmbe8Q
JmNNBqQES/8Tzd4UVInwtYnW0Hz4jYfiO2QFz8ZgEDLbV3WDbLgQJgdnsql2vEVe
PTTqrBllM4D17vtAKxtCb4ao/Uv3dGihD4/IQ9QWQ3yEJj2p7AGv5B7gd0BDls77
kgyzb09wN2/utWCWZLUmFZgNtoLU10uaUQ5fKB1K2TCF2aQNrpjqDGOjRrl8YQ+M
G5+dw/NcgDfr95EnPyvjXM34+HfwAmQuwNu+lA2QeQX2OjjyF235xdpQyxjoJ47G
oWTGlYwM6kTIM7esbwDoqhamAkRQ12SyA/4BNjI3P6gQmvCxS0A7N2dMR/3S0XnW
PtstOwemUQLAUPQn3N/6fSXdxs5HaWuQ7zlsGcI93VTPZX7hzffQBrI0K4WVh1cY
Ke3fs4aBsk74u8uzck9Gfo64M8w1ZO/1vgkyTPOnTx8e+VYCaSw14B2w08OoxxPI
RAXHGUC7ClCfIa7NazsZRgsIUuHC+ZA85cutdq7e0uT5/EDDMBb+iNOREtZCcZRD
JFNJW16zH5zvyqjEeQXdnB7vNi9gl+nxy7jQ5TiJPB9POaC3jPafIL/9/L95dJuR
HKzW2EAmiHE+en480s99SafcN0aaHqgI4mV7pfhRfHvJVAyN7RzweSyLKFSeb3a8
s5mMMddQWSGwpxtoMIrDI+rBgZ/PJ2vw3V+FMZHaBrzvm6ZCwPHKiBwABBk/M1fL
7VzO48d3fm/u7eqOpLPAmyGZW4SLj2ttnZGY/Ysd4agAfi0/MS99a7OiAiVyNZJR
WxAecJ2qTgLuvZYMuwTl2SlZabIvYJYpdaLkhx7VesqP0tubS3Ss0wb+AgRMbN9t
JdORx8zjNwHI9sVmZl1T+Y1u2MUq731q4wCKNyBUl+VSSaREGvjAs6gjO4IACnHu
AWs3k+lljGn14xIBIj97pRzH/tpMbuvmvtpjesH9FGdGZj2nW08ELvuzAJfbYcdq
9KgQw6lRNN/P5LeZIl7APdYE+zcnIpL48Wtw6WKpuviXQ1khEF+OSjKfiGl/OT9r
GR6zRRR5xkT+I0o1J+p+CH8/pj5vR9irjzcrQauQYu4ANUWGghaB9biTxEsc2b2V
OKIlq55lCwyppbzizN2/j0rXLAbrtECWJW1RTa5yZzwC3M9SNSnQyF6eFeKNOtd9
VxDMhiaImAi9C+OjFrGLEWF+wKsKLEwVmNNfRUqHZPFT5IEKvLTCMNj8P9zmMIML
Uo9pmfrDf1B4NaMGDg1OgRf0I6ps51yrm52KB6JOHnmPe2M/u1AYn9JXbglZXbrM
my73EDjpkMU4ItlezpVfO694SD2hzIaTulKFVIjTVL50w0ywAF0eNhi0f5dIbqz/
xLfGcn8qRsTmbk1wap8UBQcrL7Tyg+bsHVzu8a3ZiKNDIJsgWV/1t0w/WjQz3yb6
gMnuunDSRTquIBbz92F/ZVhxFnrEb7A9dRHu6dqkfRM14OsZfgMbnqRrbpDobzYa
7S/CkihdUV+PI+rWxsYyk7yS7sNgHz+w+tTawHJZRZY8H/owxDB5e6GWiBv2CH2t
eccv8EuN4H9zLn96+KAGtZ524mG7O+3sf5Hi/SCF3KAUCpx0rjIJ1ABcl3UX9obn
XyP1e70y89z4dS2s2mrOeKli7F/h/VzwTRdFAS7ozlsiHmc/sxkAPnl3zAfIknXl
N7q+3qgizjZn4T4NNt76WvCD73jXJ3KpM2DSKA2vFCCkIyoTouhmCAZInRWkvfOh
QoX3j7MltnypCilEt0WKIW9HcLQDb5jHYbUqy7Kisnt233bbHqj0nH8r7CUn0cxx
nPYbLDKf4vhgeGmmV6pTbLrOTqfxLhSdPFm1+u9KSwngh/VPk1rRLg1ugOmKg5vo
fmUpZciQjUmrC5celSSqE7/8tFXjOdPFlpKzkYNdMuQ/U+SqZOO2UlNrEiwydiyz
2tGvU3kUryCo7w4c1/d0Kr49hC/PpfacIFpOMzQYfsHBEkqvQ3QS5GOtEWdmb//0
lE4OdOvXeulYWPrgRYLMjKkaVgm8VFv8viZBn/RzddovBS8zCQQkC7QzdwmBzhT9
zqdWIyZS+GWPFdMcWuXiNT3eznyE4wXnqStC2U9NgFBHdOpQUDHtnrPqHVErIrys
1cfHu44a1x0WwxSQTy+QQaqfHg8P1O6dr5RYTlpihXAiDegMv0JcZTbWmXZw4Y8j
lGGE8xGdPV4Cee7SSBOoOmHwRHp+OdUUI1xybBEoB90TXq9nOxuU7PRaArJ87WVI
N8r6zTywt4FBCwSPYNGXSZvy31CemXWqgGg90awdiO8+rl+tK7uiDmJkV9mw3lZU
CVmcoqFq+avjLhGnG0lmznl7fIb2dGR2HGpRX6NYYMwvPx/8oLC88UkOTnjfXF7R
pfirx9+lNd9cblqxnJLP6j+2bYIFvCAOo7CLDlBPQWfpIxad4cgopo/eCkiQUPu7
UM5Q9aV5S8t+rCwDlnOcYQK0CfM2cL+/DB002CdLpFXlgy7nmpMXoCA3ahITjNsL
7hLnTE4EdSLU4CTkxBgyhHtlIhEmoJMbQItc0rS2j3m131U7jx7s4GJYYGzbj0gV
E1wVcO8ywV1Ev5FbKsY+xw+Sfbt4tWkr9XJWMsen04rqwNE67stIkE0yHKlQ0QcU
AyxflM90BqPQ3eO+ssJR8K0BIwQJAaYhGILEGfqYIVIZugOL0eCq9FnhmzmYoPcv
n4lHgH40mSdfJWF4MCGbxBsgPH9e9IM6rjQSP2McjNhS20HnwSHvdG6jQeoIsu6C
Amq9y1E81QDIS1N4P0KeeBiTXIO4uxZUasQulBCRYRan+gtnWpUnSjqGHqBs98ea
ffRqGEL9g9fY93zosMHl3bgbOcKVeTO3OUUuQ9qAmX5j2BVYuH/b2lCM6jauMP1M
XSRB3+l7Zh6j5LZiI5kV09Iqnkmts5OBbyLHdmXcTOzhuX1psK/jgqIhSfw7Lok9
xLwyX8eR6J2KCJEIKcG0AlFQqGGZFXHlQaGHtbS44iMLjsQxyysG26U1Jx223tWn
2/FHsG8qKK4IIojjJYdeQuOHfmAyS/r4dOJdgpDLXgcT3748HQUmYZ5PBlQThDH7
PS2oprmBocBPlidpYALOfr0ZaF1EgsL6msumcMNY5ueurur6+7b+Lp8ikHcFmClm
iZ6LrQALuw+tYCIYUdMNxCd1V0VEckmFqxP8IEMTs818GyM638sxX/SKsi2g/20G
GZPIJEtJG6Q5WDDu0NyvvGhbrLCxBIhzZxfSGfpYP9Lua5bLj/1vyyditp/1WzbQ
ssjCBFOMhFqfD4Ku/01gExeULmaGdNOBxyVbVLJyeFn3A90BXn6EHV7F6Fq+NWVM
KhvLP1HSTKFia6WTosQTOrmuV4s2/6FHt7xK2V/mx4zFYGiSCACmLXP9I1XOaODD
XVpii10HrIfiFmP5jcXhp+d6qSAxMsFa/zCdiqcihj1TgqkKXCrlCXYw0XqxRf2X
PsJzMk2id0iflGVpsLloABdVWh5/Ey5Pl90xytdJUavwjrZGuIZtfxGrtm7Q/5rU
Z7UUD/hPMZ92bK4MPqLG4vaWAQEPIuOSMKn5Vd5HGIp5v6jPCNxzr1BJETb2euf4
nY9PJQshJxKbygfBedPyDUfolsyRrL041LzehHoDJzCIoaqJ6o57rCjGrFXzFM2g
NqhzxUhsODZGPpmO3u36+DoKmVfaosGFo9bLoaFpiRJ4eQo8EYkk1in+tZRWKLt1
Imp6X2cLr/MSv6QxAg5enm9Z14GJ29qL7ch/Oqci3XbiLc9UrLiEwMN6plLqCM/I
EqZrNCBQThs/HU8EK/uBgrH3q8kTxwoEW50GZwdDyDirVEJbQUyo4f1DYt10vL7T
htZ1eWjcL5227Jo16Dc2qplj8TNrf2Jm0MeACtRMMz0YSq57f6FVxXWzlFVYRHS5
1ETFQXAvG+Slbl6nNggyl61/WVoAuKawE6yiSZ0HHw51ZcR13kJaLi55k57xo18u
4RPsMekBcFf/xsRGvX1palFewwB4llMGFtjJi/s72Fg8ydJy1QxcHulLnOEaVR/X
l7UNqp5P/VE92C33I/vyrpIxsWn5j6gdv82Gwl7gxe+vVAUDUL8lQkwdRbv0qMKw
nxDUAUycDjCB1snpMxrpvlsUbt63/izqCaMA6YfLXnQ8kkm8z1pXoHGB3rZMSOOw
e8GjZg8xjKWhQGi9aq5Jn+eak7qQNCNq1/uTVXUgt1iIXjMoR8JyOB6yQboivOPr
yB+y2tkp0mEovb6xDr3DBHp4UrbKwkAAXWguDwSkook6OClhaBD3Vz179wtmWUHq
xDd4Zouyn5McOg0F13TT0YNC1EDJDQgCjRWsvkPxo3He8ZHS0Zry+tB69TBF7V55
/sb2/5+doTCRV7GA+rAAMnKlw+arXhKQ7wHUNJ8JXSSuWbluYzjd+86pqkXKznEw
MjIBEVNkFI8M7aJ8IzlvQxY2b7VNozvcRoYlQqoWzs+g/BcqJ8LBxIhSiO8narQM
6IdSB8tC02GPHh/oVSAdqomu3mioV7FeqDkAu1UeGNzWUpBzL0xfIxoGCOELlmQU
Jja4uBgPfj10D9svoc018ZPVgCZKpT2Q3sHnlic6HGcoCtDqmGxPNFUXIxpH/1nH
CCGdzpqFIUPdnblnPGaYdmGwHQJpGEdulpKpjh1CrEXxl878t4ESwBYcvmRtshBB
Gmt1eyXXT3nZ8p8KqV6jfiZip+YtqB0LzdpvvGpKzyKh9WQCWZdJibXEKBQtZLPx
4HyQ+A6gKC9cjlWd2UJiK5ok5BhQrD6nzKcbB4bdtftAMdQQsq8MhAjl8nsxmzbd
zmehVN2kDG1K7WPwBQ2xxawJWhdNeBI1Gge8Xiyy52tChW7to18llB/S0IrfHxRc
Pt0ySm/XrGcL3k+rE8D/g3aLfkQ5ZdU5XovTZq34T9pN5sSHZHZEr/GTFyI3tp3+
G4Lng+3IaGSwfByz8QZ3Qlu3hWoFzUZSLqGwpHXCQTFvz6rPTvo9rdMcdFxNeB4y
xBBe7HIRlBhwCdwRWcgXJ3E4ssdOjspQ6i9agibg3ra/b6VYenreiifRU6jvrJmS
yFcRwzY7kMikrwtOKUKIWY8UpdNQ6u4+0cNQBahAljXYbZZTjxhA+frtHub7i/hK
RR+7V2NC0aQ86oaU3NQLo03/1oPXpqbwsagLnHPAGeRXnkV/teuyOVwvoeh8JWLp
WYYzitJHV1CauorNYh98FgnZ3QnjVKNsQcmKrxXRvC0DKHJjwlpH1OxZ6KcS7ycI
1cWbYMR5+6ZWw7dLgiRarzCfCleuzpZ5UKjB1uzB6XkAWoocl4rfnq5cUfqyzDcV
VYFq7/E5jkF/GoR99DKcJaIMWXdNkoLgtwtkzAs2RMVM4MMwozcXhT1s/c65vVRA
x+atlWOotNTwG1BXC0YmOWRyYmxzKYDooVZkqlskup5FAUhpznsd8Zk2FMXvxSw2
BWdI+h9cu52jE76qcOab30sa9Hs5K58Q+9AeN83gnpzbVOPokhM4gc1HdOn/cZH7
VVrj1aN5BGPWpIe+VU2hE1gb30U9d03PSsK/rSvrf0fvNYWJNvnJAS2GaNW1wjdU
jo66LA6SWWGCMne/vY0ye/4dJQ0sVHk2jFKIoLEGM5EGZFsS6RjKmpzJSJ5+/h8n
KWfKp6Hog2/yIC5yUEJ8wFeL1CWDMNbOSHtrpPRPuPgUiH20XdBciG9Lm2V1G2Kk
Y4wf5Vc5iTmKnrOrwK69sSLlS+U8OR5D3bhmr9mN02sGE5k82FvtIE4e/8dGog1/
lVhJ3QTCqOKtIWhSzEtWjoXOvr1cHly30xBn91Omhk4LZCmaJmByFA2txC2qNT8h
EFq92i75z+N9ujv4aYppNodVxsM9c9Ga6FIcSUqj6UA11PbAmWw5MkYkCNjxXSyN
+2Kq4P5dzJCWvmPH63h6SyxECA1BwflVmad+VZYtLTMnEC8WGpRz8mnowCo0K46Q
L0BKhXR7vpWeYZC1oPfNeaJsgq92XKTYjMXog7cdvXTq80N0x8uH+K4dX18SdICG
N20IHHFvUHK8vwUTvIJPBlo+eQ3rd/bBb40idxGvs0aSvo53zAJ/tF3rG0R3Bl8b
p7wCieWWhW+9OSH4TH8qzDqhlhBY0H+ZbNdT1CMCvsKpgeN0o2wGv4hqrCzPO4qD
8YDHT5ul1SpNwhUYOqB10Qswb3Y4oHwE0v3if1BmZX5d3mApFCZVa0uFy/bPRgXF
RGO6Mlu3OBjYssvrigQ6h1+ARIJK5NJjtKb5x8fLyY7CnWCo1QfNK45lCrHHOj70
DOcdBaM7mAGyVzt9i55H/pJ5k7VNC5qYT59KguzFubObT49tCBAIteHDeWps5kd9
W31KNxLI60m1qSY6vDWkkKmkPUeDWYhrK0GlIyJCqzC+KGF7yO1JPMf9R5g4NzHk
n+5k2n49zZL/OxWe6WZBPYmDbQ3+uC27QAoglDWGFnGYJRERweqsjU2Oywj7Q4TD
2t+GJ1vHP9uNlpayDbubtwjmmvPkXxWOB8yI8u2igPgQvA1zALu/l++yF5tYP2hy
lahc31n2f4d5iLcTfdxIo+QvEqqj+2ngsGOuW7uf/Pgx81Kstp+WfHD21M2dhxbH
rmydI8bDeWRJrlB3DqmDcvdUlGmACpFh6orC8NQVPm4JO/VSWDal7iPF+T/26UaQ
NTT0YLyuY9r8RkpBwprdJ57PumrmppsoxqAJBiGeNKlf22xAWBwT0GXAicPs6vRy
uUkZzOHUxcYN+z5I3hwoOT8YkElp4ZxzkFKDBcH9szFWgQkrTvgDDX+gBrSqz83R
4eM1SWlivPjwY/cxL7jyy7BYJHo9fDvM6mTS7QnWcl0gGcAyDgSrahwgqXTAl8Zs
brKMiRXiz6yOVP6Yb/YnV/daZZMCWSOVviwGYsWv7tMTTfhZFOBT6+cG8nR9AzEz
HqBzQHEbeUj00ibwhq5sa9oFzTGXK2T9wL0gLNS/eyg+4B4iJso/3+S/bksAX5wz
CMtZ+ZVHFVu004Y+43Ss4hzAJAE9mUtKmPryUWUo1L067bBEomvxxoPt+NuOiwt3
33lPXT8ni9xsfOcS06ik9c5DpzhlrtmhfTZmMpPtpDx7Eg74OZkpb5UIubYxrnlK
erZ6/a/azh2YSOq4ZfYiko/w9rhG+OeTA8l4FU/8CX/MtD6pRrSfJblrmMnIi5nz
D4UJfMo2UN/MYrRdGTkSHI3lifFwoGbifcrZR3aD4ypXrKjLhMO/He3iU158S0y6
zvanAPOp2nwhY5yl9a9QR93N24XW1nC+7RrPPfNpQzuOAdEZ0RspjAHjQzA/ztLM
5+mCtw5IOYmSojJRCgQOjzMEETFnVg8xCbyyXJw8NdEpLPXS7iax4W26O/mdWtQo
fuLLZifnVdL8fqv3+APnLVN8JMi/nSeSxeRr7xT+U3akfSBPo0NMq4d+hLDc7GVn
mtnY569PW5H+RsUFZlALwrjKqgg+m1HI5BnZCg/JrgAqB/Ech9fS2ZsgHGiIBGxO
O0CrPuvGHtOHoaPTZ31ofrPlE4QzmIsKQzdmVQNhKa+E3U6AOqeyQiKiIMw4Do9e
69DIsNhwXveZlJt1E7fmTn5XI7X1H4TqRKL8yKni1PeyqQq2/RcjaVH9+WaAx65b
xEh2X2z+zWaOlzEbUsUEoIyKdyywJwA/BoskPY+AtQfQ8wBnM5SflADfUvNHCw+Q
5ynEX361erFeAWtkCpb6COjmYu4T5u8XnpxMUFzovHUemfxZ3A6XpOZtvWBPcTc7
i9cQlfzmG/3v/+jvK1IG1HUDt/B+zUzXZSnFSj8F24k4J5vSJ1fl+BDq4latLhny
2u5xcSKmmED4Jl6dLmMSNg6MhQCzWkYcG9BR082F4WJIYX7DWCKU4dfW5zt42FnX
L68zB7Zt4xMjkj7trsHsjepr02+I29bwe419rGzsIuETbmZeb5w0arDlFcCWNcfA
kLERr7iMvtTazdYdWGF46Ww0nzQwr/U1wdWMgUYZYAzs65iISBmP8eOT7w8jjglD
GgagsC5KOrKOtsaYakacd892ys6S8qYOmhND0HYI54GjQ2EonoIQ1zs/jvhx9+bv
05KB2iRJCXEgE4xuE3q6v8GnFf4PxVi0CEKn9LfQMI58qm9RjaPV/F2hdOssNQLX
GkJLuWMCxJvnenKKbr1+m7R5UC8qruRvgGoDqQHg42L81sXkGUNFgln6npkfZgXD
F+L+Hz9UmMFHuiSTp9f4oGsgBQ2Ce3G9QoEtjK04bvFa+C1Mtsl5DNNrms7fw+nj
GdS3wFg6RuRWYfr4Jqgvuc6AT9aCi1T0G79TN1tG+KCWX0pIlOArINtqC4aHbAth
w9MywkAPAmhHYTqsDjLynxVBvc+Vv7Mztm5ZTthI0e25NGAcVGS2v4GgHj1XIQw9
SEhHcOU/opztWzd18mQJGh6RG36kzm9B6wPSdqIdYAo9ZxFlPPAXG4/zJNy5LHer
AbWGduQMt9Mx/9N7GDBdTzoiXtqRGjSoKGpVYhprIj400fB9mJH1Xe0akIltrxft
jTPFMMrTtabhjpXT3auk0+N+Jp6Uy9NbQ9kpiVRJ/fiCyj0/y3RyUTn9i2QDBZR3
B8w0p0QGQ7JzRMuNf2VlZ4+ZBvo2MxK8rZrI6TE4EbwwGMoXiS/AlOQw29f0V8Kf
jprko1SdWD6k14awbdtzvMydsYS+yVFF03K6VNoGyPy10t7QANTXNN7G5H1o+FTi
OfHdPZAzctGPHXY7N7+Q5zBexjIFn698d1pKkptYLFSCxyIaZOqEaNQLrPJR2o6o
bt3M8CrJpdU99ykkxai0stFqc9elRTh6mcRv9MOumCA7YkhTRGiVMV95ty6PqGKw
XHRvsE2OhC38cbmH/Z6Ud+sXZzLp1CZ/qKWQr6SlPSGwuJ60xroZVRTAcNga0tId
Ko3hNPTpe4bbcSoSVfSqMYIFbWawofW5DUS3PndfzbEx76Y7AbXRJSMJxiVaxC2L
cPV1b9JVnZplqbOSkixBnwGAArRzv4T0HB0b0oFaqn/dRs2ghB6IwCPe9JtpRIDf
F4wJWDvdfm6obpUqxn50TuTP7q91cobEriLtSrInRyoNqkInUAMuQVFvtZ4gCJW9
D7hKpE8kF+bBCjiMp3fVSzRnPHbjtITcAddO/WzuERTbn1HSzl2jMZ2o1uTUefto
/dp+7vj5ktb1h1NjOXJs7PUiaFndOlfVwf9pEL6Xsc35kawSmrXycRmvu5QDAjqV
K8OTO8rchObEP4lb4Aqh99+a/40wXwOmBBfDGK0eQaBHLEJleLsp1SlTk4VeaXlE
L1chxecBk7KEmGN4T5VUyg3vYfRae+S4Lx2GZ6xn9KNDQtM2dtmMAjPnb1s5rkT1
ZURl9PeqLif3T71Si5RhgaHd6cbkPcXOCkvl/B/8dJyQwARu3+blsJ8GQw/erxbs
M2oJJIcEl13TFAuG1m8ToqSC0oN0FjOltA/zxUrAXWEz7MxzrsaWQYv40HisOHiP
LhfOUcrbQCg8qO9mUdXyGZdOIwld1Ux0LXD+lWE1eSn9sdAd3ehK+5GZymWAR+1k
1Y3Ntuw4YgI9rHcALnW20z+WAyNrReCOce5wkC+oO3YG6Zo9XbyAnCgjijrjaWu8
uMZbH0E+rhMXc6R7xkrc5LFYKdBcpBNTbkvRFsmGntxmvQHnHp4MgaKe7amzffSB
4/Q70woosNKTd3XZ0w+/z8gAVeQIzJ4L/7ZGzVZfdwIdYZQNDbHMyPTHZo9VS5fq
jJ/9vBO7QpK3/yHPPk4SL4zuVn9erHKk4Jj3EQE6tPwUGJlF2isYUKsqF4y06yUx
ZWEPOgk5758JNgbr3T1VzePKXUXgWDUclSyu75GEPr/U1HWSDdvcstX3xPwzUQmp
UCXVwhqyHIB1VcQ3LOr0RFiYfwG3zcSBURehlP30ojMofRefdWAFSfwkfSPf+ZFd
QnmrvOn6vOimGkdMKvfRxHfr0cqjtbTHQe6nEz9LyUGOS3OcHzRry0AZSLHKr2XW
n/OJiNv8zmHNu81yQQPreqUOzHvXBXTaYkbGoSskCIfNtf35taMtrca0gq0YjpuV
rwJ19y6+IGCmb4XuaKBPLrp3Ygslg1AK4v9FJVIOfnUa/kCsQVmKwDHYQ5RbjRWU
KIfvS6Faw+uiD3TAk9s3vfDPaKfM6K2SZHeLTayA+M8cIq23Nx8YS533vvX8/Y4b
XtDYUlK/Y818i2UdqtJ9DeqaSSZFaD8ZOuq3uYbT+OhI9yPYa2iTK08taxPZVpMb
vpkIGYoHCdtEqd1ZlxVNW2OnK/1qLXDhgN90W6hrHO/g08JvYWye66lWbNdUO+Y/
s0SDVMCepNooQmJ/Ol7G4n3XtwfAotKxo1ROluBTtNQDVHtVwFhqCtzfMUL5ZQPk
WquTEekfj2fYoYM8eppmWsGJdvAih4PnWngWsOG5M+7w5l6/FZt4vktvy64UDYhK
VEfGWZ2Ov+1gPqssjgRtHihTrv3Tdu6i/iJ1qZeaHlX5OWuLgCnusw/NDTPA71g5
DcUv4lVet8cGV0/SKywQpPbqkaq3uAaBX4ImDQhfwDC1tXXFyzs0KLCoDxbNSm2Z
F9wvo0WKaeEX02ZzbSJjbFNs/QHB+ahZ2s/Jxq9NPJn7Tl/nouSaEsMf6R0d5LJz
63H8rS8KrvMPCOfX1Y73FnJL9kUCyF9kQ7lfs8Aii7xV0W59ffP8tKs2auRTROWu
2ze81IjBe9JudCHxwIpX90lBeGcdf1cHOphgnlseIEzTXo08OkJ8x4mXtqbDb5gq
nn0cQhbfzZJW4RLu+vKIldc2ekBCq5P5usHeaSskyBdlnHXvVxV4CWR6w+iTaw7P
P/MwJHNqzqTNLrFDWUcpEgjPg5OlO64Lya6bvXAKUSJc7b7xs80QqdQBwcg+36jI
+GD6fakCvh7ujrGSlJ9iEo+DN9d7AzGAEVzPsxscBSkniRSeD+WNrytteh46Usxw
nFJ+u1T3bnDvbwclaL/VySXzWNs8xMv5IlJn46E6rX+tkjZvZBoSUepLjjvLju3r
BRtdAr2ORtVhjfVxAafs7uzTwMVv/Xjuys2909ZYz01JiKp7L9gzfdO/NbAN7sUy
Jyf1sL2VpQoHrY593w+HMYvBOtaIjASbBI8/wWnti8UVlmIqX5M7zbqD40hZdczr
3g7RFcoyb32qV92xto3f0Mbud1XPegrfUebkRDJma0ybSKlHpyMACHX9waoSpNyn
r/EQPDUmJ4C/cfZ/W2OuGxcVTValHI8LHpyRfmJkkTNaJM5mkqSg78iJjSG2mUQh
BtO1uXSXJhuCyw1hognSlLQJugJLKU0ODwcT1QZAd0XhQef8Un+N97YiR0A3r5Sa
EXoH+oUO0iGr3GCmGI4KZoybkS5V3CKISodv2TAz4GRPs5QKElQ5phyyBqHyAEuV
0GFhKgX8uImtEhfadqrSKjlSBrPOdTYcwbBrcoNFJDDG5GSmV3fuy2Stdj9lGcou
YabZ63yp20QqYvsBP2cpjjr8tpG6vIUUCHjJpdu6+NZihYff89V1tCcs6Z3JboLR
zoXAP1o+yi7hdZ+1UvsYnI16nUW0XNzlilfeRUh7jlBxyAhbWuprzCegkpBC484j
TQCr1c/freV+7uT0z2KDC3AhfRVz1tnBEnbEUOL3cNeeYjdEmn181pYqOvRxdpzV
HXBkU3acre9hVMusPpk/dRfybUpDVxCFoYsTqH/pWeTOMp4m4GSxyNTykG58qayt
0m4fAP0l5B8bltPWIXuQE85EKdb/PrviyUV6YXNjUm4aD7inSNOM8blg0ftIhAGt
XMqyscjGcA0Ly5DDuNu9JDjpoigOLQ4f5DupwMlXZ4RlLMy0jZO3zKSTza12nmjn
4p8Ai0nWmcj3dmJgfy6VM4LkGHQM02DWAH8Bhd/z3BLH6C0+Oy6g2JHuJYwUBjc0
Vf/f/V0ogbWuAvHZ25dHR9rRK+GynlI3hVBYInJvvoB9V2z+dRyUL2Mf0R34XNsO
1cDyzN9tGHZMNq3GAFYYobFc1XkBxgYXdQc4Df8/e5K9c2xo8y4ewVJHiao9eQEy
X1cVerlAUv8bUkVGpImloZHhp/t/6FGL+NAVpGpde3cavGAcci2eAh94+3rRfgxt
Vvr7ZmdkGMFU6Zw/1TGxUoFDLSNdUpzzJ+5X94f/tSa6L5vMEesW7JFSyjXegFFX
2xED/SgTT3r7ftUK3tDNDSw0F73SSl2/3Cy4DsuAuiy/7jmqODOI6fWkI2/0keCc
dbAbCB3JllXsN6hwvQLRJndZrTzLhEvnIN7hZa4afgLM2JdrTLZThqJ4wZaSh7rB
9PzSbZYx8yebh27fN9wza+UVgmTE1UObj0i5YnXPnsR4rzTcVnJT5JmQkoTki6u/
G+hrS5v1563evxse6BZybrMm8UgG4C08n+RKx5nKPnQD25T6it7p27EGaGehXYqM
94Ct7mrfq8y3wAgxdAGlRb5eY1OzIbzkk01CYy+x3xyghO9rHqExdP8PnLjgTiO1
akBEM+oZZ4ynOJxWMs/7ZNGtL3QPN3RB2a+uYGDIZtt02oiSsOaZplMyPYOkg/il
XKMQtXnkYrytZ+iDlv1hbZ5o8EmVN48DT0mCeVe63+H5kcy9K9/N5DxqAJbKRCGn
C9Id7Y57/Wue+vDn8NaKLr1qEsgSzyxy7LA6I+qdAIc0Aa8Rpt2B8gKssnFK+oLq
o/LUgZZmF/+3ll2GpNGqY06xjKgF9Eu0GIMyEF0Xg/7wSupXiffVhR6x6zy/DQS8
xhVspk7kreTVE8Py5uhreGU2VIJzsGZ415clvaM9SbAayIrPdB0jfmBhq+8QzLGK
X+4yIgqpnpNl+nL/I3MeoDILlDqMQ5aJAA5bYpeh8FwGpEFgd2Sa49M7XwDS9epX
8v6WZRsCXjAee3IGZS96+nWRDdEeCBP2PESdjSwWeixioYYkQ2o+HgC4AOmjaP8D
CMnUCog8WPojwzDEiFHmcb5zZZ57DIunZ9eWcV84Ode8YOufVMcPs2kojyGGSZQP
5PisLhKZMGZSc/FnN39/mgHMiD+QVpAY/uvbS+abisj3afbnMGK7RmlYzIqEafNr
fE0Nzmm2Tpwm6OCd91y5CjUsrptTHsE3fAnfQrC2nHhkEi/wNB9YxCXr2h/SjuyO
KBE3SLGmhnnZaw4B6JDbwTR3mgRY8xt04ePOGdBS9A5HQkxaCduAzLBcYsrmkV9n
rSQu3kFChTgCPtn8YpEtkjl14xdRl3blbXccO5BuepqB4b0dkaUHsfOlGE8UV42o
nA+H2Ap2ZWQynD4f41Rg5VsYvm+HNULrGWxkjhCw4yiSRXfaoxGX+tdAsD5YKCB4
CWFnrHc13fXg2D+S9NtTvViB8Iu/8Ecj/T5A/+GlxVzXCciVsge9t5bjyQLLh7kC
foSQG5y2qxHwOwh51b4IiBoawRrmZcUrW6zOE3IBcZsX5lakcaXRYmJnl1M53Nb8
HV0tPOj8YWMd5JPWjLdSO5nGivp4NjXqaYj7MnkxsZUgSKOYbWMA163AEiFwsez6
aqWCoBsHV1QVTz8l4H5s+JhPlN/6c9lJNeQwHbnfC19rAfIlL3Icj7n6w0cv44gx
Z4Jb+XAXlBrNrmgXSUDyD3Dcbg2f+mIRjQSvqvhDYuV5JMVvbSom3uosu8zd/POc
+iAToqTPSUW555Il6b8/eA/oi0BjCSyehNL5guX60ZsKfMaisl8pWo73wJYWs1oi
JesUZqx64nGkdeJG6phC35lOG9jI0QUI6UrykICs2k0A7saxmFh9Nf8nm4DCMaT1
QvXExV16Njxp2p10RdrtqSjA2C/xIa7y3kUAwF5zS1AzQ4ELra54JQ1B9b6LDzYY
YDnj+mG8YlPizt1q+6lmkGKe2J63z5aEIVeW5nZh2/hRZFa5gi3d1kdgBX7VKrf2
HKsnFRno2eTQG4FU07vyPQkDnEzTiHUDUsBuvQpTwQmrtv1N2GjdSqGa3SJab5o7
UwqyuXYc7LdzaYO77iGn8+6DN+J36+v4eD4jwZpLKG8Vt4pnNJEpPV4DRhEOsMp9
1VIxmtBSwGd0Z2p0x++Gxn8mLD9XjsldRIxPdDkIdQRt5jAjxQY71I894ajKvMZi
17CxEMuQhkDmbVW9c0yCeGaqjpImukImvmXAlSW0wkNZv2i09BvXG90D4RQuGsPg
7SewoJOh6SYrZgol+9jSsZb4zgrPA5YmIWXNWJ+HviRK9b6VSCxvCDOovQKuuI4L
aaj5mmARmzsuY7x//LTlkfdOzJKAqGUey7r9ejc7Pu+X3edqoCYQdk7qzArGJN46
mI/G/01l1yTAdqg/xTIR8v+jvSBDtGodakfQ+1XfkOmjlbtVMJfFCVqj57Gtp2uU
9t8THu5vgtUi1cQ96fjseCRDn4LJrjpNnCK/mXfMwv7IjFIRN+RJoabetT4oukaF
TTwYv5qnX3SgwJyUj7dCkPYJQxLGU2rELIv4yDjp0qtO3ydiieQB4QOgn6Ojvps2
YY7j0VQVTgb38BTOYK2hgPJxxxgdmiiQHylDxglIZ0z2/isrFq7hnmAoNNktZJeU
opZvi2nNOksg3eLG9juuF1k4GoSu1pljj3WXC3ZUSUDodcdfWU6IjTgadEaJw4qk
QYy9mRR1E0w3L5QcM5mBnUlow1NaVWsOWDkHnNrCzKTNai3/zfpoqnuD0hFzYBp/
i8NoLbOvNnpd9qyCiyHHEl1FFIWMtBUInFByE0Pt6K2/OsYlpTDymAVQbONfoumO
20f4xgLB9XWluwPsSIho/d8XGghc4cFDk9Kn9B9SneqSYnFFyUVQYVpQJcpMLwqY
6SviaaitKePdFEI1u1R1t+V3vnzhE63CyeThCIu8Ni39vF4LaDeddiyTlewKjtj0
UdA05//5X/+BVRFhotqVmY2Myt0Mi849mZ0KqbvSKS27nHJaGvWz9u6TS468nOru
Jh91eQCmV70jltdgwpHWqB+gwSNNqL9gow/7/JWAblDQ1S1y4lyLAWJJt4GmdPAF
K1LsgyMpkJoHWozGvMtFnHdBysjbF7+mJ+FulB1EVrC7ObtkIQNfSTjTaS3kPN0f
7BoWDoaysU/M3u4vjJgeO4FxyMaEfn/T3jqvaDEErWNt952AHrtyHELsIyqsEBGv
ppHXf3BwkRAMhjocybEzrIfEsNUQ983NqfZC/dV+ZYCQdxQ8MmCoJCOqMoLXm/xA
0flvAZ+nPsnm+OBZBGkUDmmrk619AsUOzngUeqkBhDmXUBt9PJ7R5uFzFsF6WDLv
KvspyU9v6qylF0zFPweaNMYfJo/4cD0d2lC3Cxqh8vukcAiPcNc/uWng53qBfFvp
EBcSFDMTG0l2OdBWjEoX0ULFUaKIZRQORonfNK/nMWiVXBGeq/g9hAcfjTcDPR/p
qTXkfY7bhWjqGNC1JJLuxlvXhSWyy9UaBxXJ8bVg6Vi0elvTr/b9De7jVE6ZcA8t
ZnKXQIFxjkyVYVp97oVXwjypXiSIG2aYBBm3wJqmA1QcB1380sMXUzGQMQ0ZsAB7
OBFzlxRiQaaXfRUE3Rt+hi6qUD2JeD1VGify1IUlOGiX9bElOVf7vsaDe6GKzXHs
/bQdNP7soBqNouZ2ud5oqQ7vCSZ/gR9qjTuQZbYJiwHIxBpmZz7XgFVHkPUvdoSC
OE/uodLmLfkjfWbli23czJvx1b1Y5S+8Pk5sMdefkrYwkJyMbO4Hl7ukurovYQfk
RWuHlnLu4zn7JbBai9iTMIH9JeGoHoXMwfiMx8uLIPlUKJKmw3ScOPwWBeJHysN2
K0xXexo4zdC2MQ1xpjv9lyGsYkY+GUWQUiTPo5uhMcL5RTIr55+QBFRsgbkr25oT
6kDyBF78Q0nYBpBF1eaLWMwoanG+FcMhbToCvbKnZ/KsRiMIgCUmiGwZWGorWqcx
DD4G7IRMktYsDhjSs2+5AHoYNeK5jFNvCHnD10Yq1ee7kYiZ9wWgtpFp+dI0jfR9
o5yJztkSQ0xrsXkjbWEhv32cxIQcZd2faXiMzcxxFl4cITXHxiG7S7j7fcSgvuTT
l9cEjoGTcp5Y0bp4DctMagtBAgww/9YqgqyVztsEoneGis5jqI6ukKnqe4gPd9Tx
hpfTgkzEuFpwdJviKvrCRy+GvkzEux+k858lq1rZBud5DwDEKQuX+ZQIYlxEU2OG
j69+gpHRLSYFGhYWLxZXNmA1cLcTleebWGKul0BatUS/Abzui0zDt6SmsuL+2Cbq
YGwXzExWTJJ7V4MhC6DhxYcyJW+LohXBvzY17nao3OdVz6frYdevNIM5rRzpcPbX
ZmvhV5Ky4t3gHqP8B/BtupdFIOC2GyaqUxN8F0HDAsLDj0fjWSrLW2xHeQ7iB95h
P7gXUaL/+uIGjPCOifZ77/76vvdSeOlRA8I4bhn8P0gcp+E5ouWfmQTINJXyxWc0
k6R45q23Or1r1gJFzupPBcNx2Ono1HUYdAbuqKsFbc9C3R4pEdUJPF8ldrf1SjAe
ZUws0YXidmupb6QsA6l9NxlJp2dhcXsytrcB9EvuOFDQmXVSSX4OtQR+l+Hx+4eQ
Qz5rWh0yjEwNM4r5qOaEpvlggXrrd2ABxpbmykFSoxnTIy9qt0ZdFaFuQazJeVOP
xdM22eDhsKzWjqCm6utosB/PsWZFilS2B51Kl/y15UveDdJzCyMsOaf5jvPyukIg
islR2eiLI5yVA/W7le7TM6ipioj5//YQrgs80CMMKctLNmH5G2uZSt+yhPN5CEOH
Xj7KRnUXhSNh6afw96Nc7nqnPE861HJgco16TxNW5QKO4o/U+YZsy8S7O7B1GPBl
fFJJUi0d67wIR0l9uCE9bhwsYGR/IknWwVvTQ1C6OyrbU0LTtbYCbp2xPRwY738h
APtrRD0YP0dJFN1m04S0lgt//TLqf05kMU4dWyPiiNQPS6tEyOkAitcjDjAEbTQA
1aqbEGC/oAE670EYcIg0Nb7TjxZEK3iwc0jIUP+OURj6mRohwhbe6/PvqBTux8Dk
8sDXbkdL6VaQrh/ftqTAL96ziCjMDgafyk3gPNtZM3TRybDfw8zq3jvwlMHPfFHQ
J353izUj2qhrpEA/lMh9ZQDqwN8HEqb1ps4AMpJRZ8ndDmJQyf5L1Fy2bk8jz/u/
HySaR2Yvq2TudsrJDkrwH8QvKMsvH1Y2Um8O8t1Hr4l9Jt0IMLftnckfMoiynbyG
OWHoJtHSXU1pH3XDrjgJmojaKCyMQLK0Kkx/kEwxk6CRiRrtxzroQ+8vWbivOQXs
kkDxNJy9RY/uTK6p6Lp+EaM9gBBZ3hLzeEzAAasg1dqCP8dJIxtILMgDhWhpNWiR
nBvrCtPSXy3PR6Stv06WJN0ZmG7n7Y4btBGg//lA67bRrLgy1JmNMSmKyqTRqGOw
trNYYZ/PLNzg59fYMRvLQwcDvuXUhEVcrVEdsDdTSr81Nm4XRflKWhjvppXGVpVO
QgLV67xa6kBzNbqXnuq0GYGi6ImqmuKTtX2v7HKekrNbeB9K8rfVSM9IN0nJhRt6
ipwvtUqcI/Un7DbWzCtluN2sj42sEBTihnGfgWlEwdKH51opa6QqWGX24b8AmaNf
ka7QzZNRIyoZJL1njUrsXJJK/SkX/jC1fKsoXTydyYMmzYGB5IOecndL7clQpoa1
sK1tXOYnmBb/dqXrodv4EdJm/kL6IYbnjxGwjJr8CNXrnLhyfPGsNHAo4V2UdQzZ
WmfIuS+xnP9n0fm4dZxqonw/v9qyqbRT6EtCve5Nx6S5Us/VIQnjSJ+il3/QDmkW
SE5AuynZQhz5eZ8cqR2/7iRg0j+zqt261kH38PyPdIJdADfyu9WZRxjHBCmvC1bk
3fi+/nBfolZnRqNG8JTtYEAJ0aOt27aTuBXSa4q3HMik4qoRjisyeb38TXcWz2cs
URFFXeNqA60mXJwult/BLztDBYnALZTDIMNHXJcVfGTxao3OwnrH0VSwYaCfCIdG
IMGxrgzXpiR5rKGU0Y+vlEjUiFbOuTtlVtaav7QPzogIwXd3c+P0r0Cw+LvOjdAT
LYSsUP5ihi3J5IFRUvmHTJLAd4m1vRwKJboAV0FhYB21XmHnCbXg88Yce6w4FJuG
w6T3ffBweVHWCKOkHmcSXZuGpzsuRJLppAk9KkInf6PFn31u0znxBqOKE4wBD55k
z9fJ/gocHH4ZOQCaS8y+7O281ouaHLDNdQf9WFCFCWv7V3GakaJktvNTusJjBukq
rLV2BwhcqV2EAjGMhcbGfBy+wNCWrmJlK/ycfjpCzGrnvV3ZvHIbam1hnV99bQOh
qWm/Hqut3AMdLR0RyHpXT3bwv5VLUaB2gTXxeq7CcBxTr6/aa/BxCVxTy6kUoK0J
6qnf8WOAMh89gzmNoetp74u6ee9osnwRkIbL8EOO3F81pKB4M6uQ8G8CmHN5+ONM
PLbA9ZI+o7rR8xT7lPxxFbmjzYvW7jrOdHuYSLruZ+t71IT6sKO1E6r7NUdbFK80
BNLqKnfS1Zz9ZFoYP22zqginDxb82BTrsVb0ZdCf0E7cHBJIWxHkDOhrcOXxjUDG
xuq6xL81XID+2rfJOExx6qDibFqg44DnKKKVFjEPEirhu89EbQpInjHAt+cezN9R
Myo6MiuvMaOT1gfSq0r8n6sqA1k7y0Y2sG69B70DoTPjseJqAA8mX8hHZ/saC4BY
+lNkCsy60ExziDPmoJvdndzTWiY1B3SVPsFxXHeSnn15efHBzERRERjZ6909oc7O
QDgnzshg6pC+0HNCxpg7tHOTyUnT8hs/XJOP38xp5hdpwoJG873HQcCAzK7IKcib
ervaowhUWN1iDJcYq6wQaVHjkjG+SKWW20LHKk1QKNkUH8poX17fNJmtc8tRIGow
iFC6mSsI2PzFUSJQI2rFLVgmALC5SYmMzbi4ih0OATcxKEcuA5T1y1Pohqub5c9c
kbhyNtX79fKFnKdB0AD6uremKpRKLuKNrIuGL77nFpneq6aipRdg3NLhje+1UC3p
8tSH0Q6KgjAj5SZ8qH1pVEipF5f//aTDJ/3TfmkS4Rsgohom0SUn5HPcUdUs8d/9
IBjjKHmQzUkF4HL74TLMUQYQ3LLjdDMjJIa8K05OEI08kk3fFVd2dLSO07Vk8k9V
OsIgLpeqZ1DJGOI3Nlt2aqmwCBGOr9HkrxOSlGz8ySnB5FsuL9j9VpjnrjNjmfJ0
ZlD4URCack9+mhi61DAPW1U1pCGh9mxj1GS9L1s66HH6wLS1facLxMfWlFW4vxpq
EPxzznm7+kN8FaUyuvMGxAShVWbFY27yklCXhnl0cqoOXsc8DnyfVxpt8dcdM8zr
3ox8vzkry3c5xV6N4R2OUdQ8bxnpV23BoAAh/IU8BS6tFxoTYDOF136g2DNBnNHN
+wIZVwzca6yLcmJy6l6wdvT4kACpuo8YVHhHMvSy2VzeNcFTHI7MpQymPvuyPMOo
vo167QUs6OW5Xdx5Jti26/IlpWBk5Fntx4WIMEjSRljdTZRbyyDumfAa2HYh5ljN
nSsA3ugOGbnssIo8Zm+K0mIKW85HfYkP/zKvgK4EBvdkNdt6tFr9AdfNKasy7IUg
1eOvMAeZCHGbG7wyZrLiELmBRTkRefVfcFfMO5iFfnGru8I83sfhFgIwH2xAIIL7
aYsnusYJ6zAs1BWavKNDnV0L64fbtFWFGucfABbzArYA5dU43Faxb5QGmZaGMj4i
cZGeYrumMKJg58RI6c2FCclqcsv4wjJx7MiuOTvW0uJNbwzhU4L0ZwrXpf+YRCUb
A3iiUslidXaiq7ORjAUn3NDufFGFRzSs40X4S2S6cSVMsmwIhwiapfnr7xVjkQ/N
ayM1qQVjkU8kWrM8avMVcZ/KtcIlfK6AImIl/JxeojxzEfgazz1YNjuWUy8sWWgZ
3T+eltdVBEo8dgQWtI5ZWfEvek7eUbcwPBfy/e8M5OO3kFY1GgxezugBfompHnKl
YZgyzF3Qgg5g7MBCp3YWjJ3dPHythbNsI22nPqrGw5UHxa/mCx2dIIVhy0EfrVAQ
Pdz8A0x4ONKqP1cFrKP9aCh6UNrvDhnb3jqEMZWU37n0s3hWLDzA+F/qu6f1SIvH
01zY/V8aqnu0WBUfxFD658pRSFdKHM2dxfL4v7CrcXPvnc7U9n0xbZwif4B343jX
M28dJrJmUGNJRUDPyYbc91dIuwbz5U0UpLtXs0tAcYLbyJQIvxtWodCAI2ZV3+SP
LtHndIAmUTsSDJ99/cY513VegZehw1PFFUCAh/3XA2WzC7Nyl1f1m3xyVkBIgmFt
yGweTCctHeQAm5vtvfiuEhcSv52QrJEAW92K/3JOeGAhgq1mAFyhUtKrFgtLhCRB
OHcBYmXcMlPo9lHz7jteDA2LRwWIBO3SsomkUXciRTOfN2ud5B7uQ0AuwZD+ATNp
GFua9eXaEUyHFkjeY5cfcQPlS3UIDbfEkvlA6Bms2JYP+GCh6AV08uZNvfB69UKW
20KFv3kGmglLF1paW/cGCqqWTYhrzw064VvXYoalI5BevOx6o70gvHVseiOWO4co
Bu1a3YEekNDMMbFNSDF3vq2DfV32c6aNtPS8VqX5O/SrwPJUf/bbSD9SSDr00gZ0
yj4euwjRt7IZGFDrJxzeVHIuC+Drs/G8wQnMqloDrFtiDUiANZ33rRatAVJ0M/ff
9EHp+zYfBPHrDutk7xeNNj7WTe+B1Xc5BdZOR6VA9gd5/rMYZ6k0S04tQps92gcS
B97+JTVj45uVIsmwDuTXHMDbXlw2r8KOXmALoMd4rOQnkKFvhlNuX2W72nEBtt8R
SKpIjBIrMAfWEPkK6LEBagghSTtDEA0/k8p79u3RFKxqF7k+U73DTmKxB7ZBO1OE
OvVggbyzOAEvUEXVHsW82fAv4spHwSIHYKOhf852Cx/1erWzC36gqZzDFAjtrDYN
sa7CmUZzqe5WhqOIJaPE+cd/nwJRSqxKGxggX0wqRGfrRTqbFGqfbpOnFlzahT/R
J+u5s7V+1iuhC9K6RCh/4RTqW9X9M3lYaLigwln0UD6uDsMB3/M1CRCnglrK3PH0
lhQBoc8qwHT7jdLRoEbwRN6ko5ffQmkrHUmnTKW61SPNuJAQpVGyyEiBHp7MBcn9
DT/hLPrn9TUb7jz79LH4S8hsd31BY5OPYGBPQKqhb3h1Dlp5itbF3ndkhrZzXYxN
OUi6EB9+ZD5Pdv3/cntR1DgPgjO0FAsWB4NyiHp/M2MXO2KTuB5XVvMIMuqVDgrx
MRvQFkqMowgQHoG6TQdlMGvNkwIjFMt/iY+7B/Yz8cQEHzHD/xYlPXs5VQYhbOwZ
T4oaVf+mQJhrzXgRehXc7E9VpGDlS7QF446MGkOrGkpamYcXbyG7VcYZE5eNtKjC
1Q3EOx0fBNXET4kGskA5UzonKLO+FhqWH/Rpf6MBC7SwF94DDV5sFl/Md1GnHBE5
75v/XixoDi1xZiEQYclwKCZQFBEX7K697PzYmoSyth4dVCd8E9BdKTMnd73rDxGd
0m4xpA09NNi0yajhRYNfUa/y2WvdhgNpDCGXcJswvnbm7T4cy+0oqzGLAP/ykTcw
AhpqAU7I/FaFRRTHEyiZqHCHvCSKQ/Nrpi9Af2LsAbZ0wef0FSNECWq4zggYg797
LwyvYXX/scVbWQqh33fdYmooFg0CzZdOMZ5r40TT+B5oyrc/cKSI7Y8Qhe6IoGR5
jxxZRXwGNBcT8MFLRwPQb82WLGxzhWqb4j/1PKqrShDTK8ObCmKAF3ouw0Ixqged
ZcEOSDegFrx5qQCLWvFX1n0Ycbld0X73//FSLKRKwFmMRnm458/ryXJ7R0ejtfCA
JTZAcuL8usf4n48hJeglS/wto9rlAG4eX65BLl/K2REupJGAxS1hxbcg5Ghlm/+l
AvtvuquSjEb3mBtc57ecYrrXCxZsP0rN4oXK4yqSUfqKjNk88pIVC0FiTRtIkQCa
Zmz6QVbtko8fAqaRCex/qoN/cC+oUHKYjF5Mf+V8tk++uaTmXXr9b+shg1ZrM6IQ
2L66wgAtOL4JXqrIG3oN0FrxQD3DMoJV3yQLdPPmuyq+CoUIfmcVy2C8Fn3QGamz
e1OsE7tWagMakZyFMwNu19Kpo4WRA8ZSLJMNOramHlzTAaFmnqfIfhksKZtbwMwE
YJ2We5tr49Zb+2opI+gFS87HAn/qPDitNpTuCs8wpZDQhObwiXsqGx/CDknaT9Fv
shtZ15EQ3Datuy/CoUsOlBZJqbsh85+BeWUEY9kTuSlYREVyaDsH32D7yCgiH2Mb
HcVQZcOwa0n7cS/7LtvZRhks2ATW/zOENmUhFLxrxoMtURSV4e63DrUtxL15cqui
kUS3goZAluFBK1FGARjyHQmAg1aeKF8ZV1entB9cOO2Tm4bjmYUjg5Cd/NkeZ64P
MJLbkROCQOQHtEk1O9r1ZZezNaNDT68FUBmm/HTqHNhtRZoAZwXeVfiyHBW3CAzR
WTlJr9apphYqmzJp3PuanpiOMs09FJsuzg5347LzA3LMIbJaTmk7FW3w/hLhbIbc
4gEUoPP623qwPIm/wzt7bzlHtsOZxzjaUxh8IJs1rHNUa4NBThDS039tV+WDiU1k
ZYoSQoycgFrIlCN46mryjOR5gyUi+ISfjbSvvxJBEQdLMwvM9tRdmgVijnR6t3/W
qG6Vct4Tew9ypV+0lVj2c1mKzjCSAl8IhKdSzs17oxUggl2TSJfpKJRbiz3kYdIf
SqA+sLPLTnkcApbYBq+a6YndRcrpOKPI4bEGUL8hsvgPr7i5Ef0H3Jxz8EVXtFyQ
IUbrcmcNyVpHsU+KH5BDyJevtrUQshABYjPb0/oCZlGujQBPZbArwyGhjhB5iD3u
bccvbMRXGoKNCsG1BgeroNlpmsWVBtsk2KLrM8AVuHdc3zxp1UL85u55tRb7lq7U
BqArD1/k9KPa5RB3gftEE1wkD7GiJMAQgYxCCwM+FSBHSz3Rn0eG6/VYvkLtt4/e
EC5RuhipLhnuau5tShzE/yEU2US+MaCFAt8BQKCim8ns5W8STNMJXxPVugJOm51K
u8RD7ZAZXbFe+qAc5YUfEGFiDtte2g+ufUfHDUnO0XXn0Gh6/R6w0BJJAyPbA8sV
fncVlFRyV14dF3OMDWRwUNDok8PbrEfI9yVQnuetHYwNrKE0RvzRBxokrvmbUdvo
EDQJ3AevV1/tWMdZPbPI7xSh777kesEUJL9ssBQW8LkzWiwXCjo157k5lwCcElZY
bbB9m4x3Y2q66WclpOEpZGpHlhr69R5AnaX9gBtM7DCOR8stE6Ar4riasZgjQoUa
BlczFha1pf3/5hHn1057Y1LWXk/e8jLvOXzRlLvDvCRpm4doi7+YB9TbtxAYcOON
CCmaMrIWPDrjwRWfWqpX3DC8yaNZVpXZTXycFOjR9ibzXph6dVzo18h+3jv1BBs7
B2xR002+STnJqfkxmBdUqJN9wiDd/KTvWuQC6+wvegBdHS+q1c6DzrfEc/CQD9Nk
HymUC8+8zXl++buYXFDgUcWFAMZEPwXI3BXyV79XGjww69Hnsm1ECgZv/wm0pKnH
JGbDBT7X2t8k7bYA7RVQb+nyNsuFCRjhFiGWIs3yKhvecB/4HllBBw3TXl9xRg16
80CVJUgW1Vr6iDqoHCzmBtARS5aEukGnJqDwTZWLZ2Ck1NzhQ1NpP8l9iBVUeyyJ
4bp23k2FtYeOIoQU0ZrlxeFD6nTCsyQXOBxm9avq4oz+LoUDUrP2X+0uIHNaje44
GR44bN9Dd1S395RkkAwXf+2pv7fTJxT38Xwxv2H3cduoSxRO9hjr0SGHhIR2abeK
DSiHPzhKxJvtu6ZbheIXt0FvmndwoV/pJjI9oEJUiU2O0dbs7FxN2Qu0IJY7+NfG
cUF1capsJPapHTlro6lTfvPBJ3m2tzzbYBk9+VfH1sYqmFShwESmTc5/9lMAa52x
UquG/hBQXcRdKphd5z6qVvUGOcbdsEXJdyTm8QoyAS9Nl5QlOCFAcQjEFdBntngf
bbWw193XUMCbGw+YWuHvLYWJ0KZPAeEgxvhJ9w7l8TpfjoadHo0ss1M6GLCxuCHM
DE1gjgY0BWsakuKI03lRSy6YJkZkNIPGAdr880EJviQ5teQPCjf53DRKj3vTr7XZ
XUSlmvv5Gl2VWlsP5KMZ2RndXeCnWqMopqyT95nmBnV0e6M95XCQvjSqUjZoRJN4
btnPenZQjXhpmkGYzr5N/gJPgEws9Y4tO1w/o+KOVF9XqM9KSKpzfs+Bi5Xkh41g
y589VYRbunugtxnU1UyV2Th3TgBv/POOPpbCiv2Nt9gzJmJzN5M8v3YHzom1M9dF
UzDn9MxN2LLpiI+sWE5FApVh2vUgIJELuqC2MTeLtHOyVIn8w71mSw1kWdv5zfCc
hWPKB7QNv83obSRNMRhwFR0/aKk3+OnBNdMq0Q29Rwqf+cPOIFHuINEAGWtDdvAB
4AKR/SqockxOlJIWauyJwCfi7M57l82RtQJPqwhK37OiAgz16YW4GyLZO8ZieYWL
bxLVJpIYM4JF/3o+ZbKs9Sag8k4IL6ieroMNA4ExekhZ0AqRiu6bG+/SPovVWbEK
ZqxaHrZYX8qlP81P/VJgbP3tuSXfsuoa2SuNJrkPSpWtcCKm0q3e6f2YG3Q4kT4C
hY74I9XfEWT3RmL9xYhT2elT79+6BcM/Lini0Q0MZCMZ6e7uHhx3sSpjAv1iAtvC
cRT4SpPQRn3+Q2BwSAE5n0P73iTyCG4AEjQHuOlPPe5ZcF7bu/gAjJZVdRImUZKb
Zru+dsat7RXQLjgqfr8BBfipG7R6+cMCCmszhMbQndXjuK529hFJJ9D4OguJLgvD
ldM6ZpXq3BeeZ6Zpf9QZsj1tP/UfF/MwSXYSCRXA2L37nST84ql4cHmtVX+O0TE9
Q94xesYjGPXwEB2BY/eln24J8GTIVnxe6I22CYb3+PSXCYHwfhK3V0SkkT26VlnL
DHelv3TYxyoc8TVa1O8BB2UwtQ9nBXdxoXWd++weyhoDFGPSfSmskh1GJKNy7DOv
IwGr+Gtd9t0i5aUQm+eSBK8mJNW0Wu32EHsrz4GagpiloyIRoPzjr+R1lnVYLao1
jMuz1eWKjjQ+74ptBATiw86U+dDF5SGQPNSFFHiHxnWdV4hd61yntJLxUeZJEOEK
1EQWjjp7FWKf+3csEQr4/4DcHKucRgxwXrQPQDHZ2pWbBAVQsdMhUIFPuIT+cZju
uqVjXT7yUAQPxHFrfL0c3B2pkUg7XIDpSAcrC+MZB4niN91t3z7IWeErDCOYZYl2
rK2rziQkIX8PpZvjyHc1zeAC3LVwjAZHP3pAyAjb2z0Pv74+eAOr9jgvteM3hw3t
80R8u0ihfylM/OXbm9Qp/YRwh4tptymAa/nh80IQRTjX1hcsvDHZDsmxvxE4KabV
oe30yRilAbxhP0cV5oqQ1Hnlp56sJv8rFWLH6rpqgSeUNkjcZJSW5ADn0R+fRPFH
h4Xi0usw4Lc0Io4v678brcCrHUap7qHAs42MsHMyeeLTRgZjPI2OSx4/EojQzeMa
SnE6txpz3VWCEZeDerRcy/LCtykXs3hYsTvcneGS3PzusHGWZHDYO1IV7Ks+BH3K
m7FmyBjmukXNi7o9XC9WBpdxQCCavuj+zzKLk1LUkcz1lFvEYtWe06N0xnOL0jpk
HnugAEQd2kXRLwmbHmKo1e/+eTfrP3nWXf7B1ZStXaoXFbOWwVxXKVZjE6zZjBkj
WQY3dWVXDrqH186eQIZboLn4XuYMYgBUcRNz32E51myBAbXJ8X7WHatXNVScc/hi
hcCMcdRZsE2cKqC+HJfjrMKuOr0KNr8PpzZGTqpLzfUP6z9ndaVLHmslCkAAXJga
lE6oNmYhcczEN1w9f9oJkLMpTuz6WiEu/7jY/lQQ257/RNobs3qrQMYtKCwvc5Et
YTEWGiwNRyCrutGk/Wur4fWDOZywFk8s9e6m9uKJy7k0LUqo4NqWzMK27lQTFL8r
6M/SNtvwX20/D/73lPy7BIptNXW4CKngsv88WGmnlda+ZIfQ98RiJnJ1CTSVv/Id
+zo1dXWdUdrodaOwOm9NE5i5Ng6RXljIaan5BLuHewdK8hIUabtyiUUL3uRN6+Kl
4K/YI91uDOil1FWFP5U+5zz9L6ZthOaDYfQYLThv4WSWP32OH4DLae7UbKzbNVB/
DZ4S1oZdZojYw4I6FqA0u/Ifz0SZzYYGOABR+nxyDrrTEdUAtiQ4oXd11oFkcpG+
eVgW3s4PUhX1bDRh2aW1Gscp9F66ti74MSr5eGJq73W3MsG3LsW6JhHFfRtUQZhe
q3GiMONdWduh6lY3jjj9xMIZaWQUtBJQxxm9CyhAH/AaausP5A7rFhXKONAq0rkK
6Ua2w9kCd30Z68xfYqNnTJIDAyrDdnOfmxv2m/Q0BA+7JNpuFJvkxz93FlNE/WLr
JWmIjpEt8SDgSpxBlW6CNWOwcWbqO9OFcnXFTGVbyqkWTOdaBdbzfybzbZ6fDpA/
K5bDpbHqcyR0ba4vypAwHV1Sr1AWMA0vm6BIqwbHROz7i71XMdxVaKGNKt0PnttG
ieXRjcXuz5kxDS/7RTRSd5dXLZnMoKqggvFIxca3LsWJwWP+v5RhI1ppGcya0MnZ
hxqxdwKGaVpU2H1pmae57TVQ28pV1lRZm/pJRPz4gvLlAC7oMd0GLYiCK9twuSXo
LzHfDBwAtkMEumKO2YL1ZOCtMMa6mr3HbkjoZ7yOQ7bWv9iamAn9q5x7W0FirASX
Bkg0vGfVFfLTjkJStHm2F7WMW6pYzatFQ5VXbh0IRIEzpz7XlJSueIwOFwNUjkYV
h/QsD9egcRmcZaoNohl9vV05j90/p0r4pDu2umSle1XP6fr+SKCvGoVOlAdk7+r8
7LrQC9Jii7ZaHAENndRTs6TB2r1jGGFoUIa69H4f/8+UoAxhe5SMAPX51Znn1NKb
jsvqdxE3niNVYwDvoPxPZdhSSeqgTHi120kj4dvm75fjvJuykMl1ll79uB5+F/vF
QtRK6iC8vjTJyWPTFZL4z+gKSkJV+NEzJFYgsBQjORJf7mpHmEOl3Lz6UVhuEmpj
boE06SXSQfHytksrLyc5Dkq8QjHg0B7DM2jMLjEwK+8ObIGG2+MEem2qYtw1GCNX
gZrsuCm41goJZNiQn6RgQN+7creGqBRCZvFG+hiCupoCiL+rkwZ99oCXPouPm0R7
CGCb/iwh8e4LcMmkRH+MrThAM1clVjSdrk6f5daAaZdZopipK8L6gHBALF7t+lsV
MsBbxCkIOwfZdaS8IT6YpsaBFpFA3G9aOctG/85LreW+xec2lrzOLhSrRPHki3xn
Q3l7WzhQ3IYcw3ONoBan37rKIeIItM5QMLNPqYnBhtRTdE1xky693Wu94JTndUkH
62QwjI5ILQZUv9Ji44XxSETR/+B+f0f+T57+rjNILrsh57A46u8foEhUtTeLtfjU
AvcBv7Btfn07fKxOzGvpBiRnhDy5wnQNz08ZcJrC1WAsQs1855+854c7Y98uTfhl
/RiTsDfc6YVCAQs+ugkmuuXwzohdyD84zc8YSQC7sRWLQ3zfkQXbXdQ+hsmGAvqH
xqLdysPr2T8YPtZg2EanItz+irGXiEqxvp0uC9uJDGMAzRfTO632Ovrqb23nNyct
0itlqz7bxjHuOf0nLGrrV9/hBplllL2ErFiJxlKj7DdOBf6x0QI9zyIRuGfCMVHW
t5Kx/lzQt/n0eeMtW/GH+vGlNVB5RUSmsVfx6UfL3ZBYzlgX0DhyB5RqLKQ0zWul
zIHy3Hgi/XCBnN6EJWIM5/3YFXqEabl0Xfyiikzh6yKXOKFMPkI2ySPPW4FdPsuj
1QESlgzQvDw2e/C127+Ew9/PBZhdYJOMU/2z8bPGTlec+hqDW+5sgxqCpdcA4FQe
NsWHnTsNthH4SIJ2HaN2PdpLsiu4l8eubRIDWXAbP4fhJfVENAAjPz80jt/Be637
n1c/PHKUvImdzWLlrZYuczApOW+RQxwa8l/GtAdQxuBygUBeWN31BYpS20JO+hib
ezj/B2dLczmJotEFKJU3+LIYwPW74SoqijwhA8gI5xKXXg//0BEpgp8LbwmT8VT7
h/t2CPbo+tdwCavM9LzCs6rxGELWXpd/rGeLfhoir7na2udNR7xumnFWZI/ef1jH
Hz9AjJnyILPB1Aq4+ZlZt02XOHrq6UzZeH5vtUol8RskD1G1lQbTyNo/A+dtKaKc
BvLV0oBqFwPTg6CyVcWOkDGqOv0YZeeuoPbD7GCF3JMep5KwAUTAPLPMmz6WLeD4
A8+YUVd+viHMG8vhv/1L622vLeYv5G0oNlYQNh6UX6W/11RtyDofp5ilVHYyRe/B
bK8ajsrH/NA1qhvek+9tMO/92HCm/hvmzOcJIaUcoWkVvNnHE090T5OZViwGfz8s
gl8/V6dGnxu/onrImi9+y8oUAtyiHvaeZrw9S90bfY8+ch7q6Wx1utuNlGCxHn7J
0vwgVYg/HMj6dzmDm1JNfh94i2DNIQxP4Ijs7qVRMvqZKvojh4RxSwoA/AOn5JzC
khbw5BuAgaWrm+OK3sD45pes1gOsWUVwJP5K7ub5BEteB7ALd7nhjoANUej21eOH
vxbBV5Yk/EmHdcF7qTgP5diz1Yr1VnZFVNccjZYWHpsF/hBKefsTKG4i4oXMo4ek
NCEa4XT1HvjeVrW6rf8vYv1Mq3HhcF6ahT+Brwfax4KohiaPh0qpuFsucTGQifQs
DQEywtpECzQ0Xr81i+ZqHpngCEw+3k1wO9CavbWDeW7czssO4FjrJZ4vbdOY1o6a
tedPGafnAnQdLiz2ge9kG0Xlt0Z6qY5ub5dUT+ulXsg2jPOhJdYmKpRIN5lgDwq0
Gerbq8XzUT7wNv7+shM/IvnO1DAdfjI7LMZh2n7XQaeKfXbecxIF3iMRbZ7kmW/z
DR5LG2KKNfg3kkqEikz0B2hB950SHxsXcwfCFuXaMX6J6FlwleXQlUmjMbF6wBUh
dcwlKeeqw+Nx6no8NQ4hbtOOrJ/R3K84po4qhATKbaEbu8OHafrI9NlMTY8tRIM5
LWroo9HaJylG5bivy8Pfe63aU6Ai3SzCOtzeODeA3wDYmHBFfh9mTwE3V5+k0dim
SQGYaojPZGRdnOpgCD9pAy921Z4o6IubuM1XYVxADrVIHHp3Kq4YcI6Z/Lkho9R/
Sv9o0DVgplEHbP6LiEUFe7I0trk7HyYCoZOfpbgEfjWCV7/D+Lg44hehPYs5QEk0
eXPw+mriYd/YISZEuLtp+4+2uiXv8wOVR0Gi7tahqtjDQcp3GaRiMpCkBbqewOi8
zyfMdJ4mN5Yjst6/uwDz+ASSEs7C0loBcFB4N6xtp8tSNnTti1TKzwwOGvqs9aCt
yELNxONGEs1fiwvlrpw8LuEbQ9DAocn8f1jICsh6ZRlEO/xVaEnQDQGBzYQEZX5i
D+LmMH53liPPu8KSLT7a5kgYtnQiV3wyw5gChdaIeQrzN6Pq3qW2s03TwLAYyErI
qwHQ9PLgFlAyivuDYrt/88NzgvkPcI6M8HNIlisuzVP8JP7FbIFYcpdsoRMMngMq
fXOSUg2lMXd/ddU2emLmxuQWePVEslF2Ub5vIZwwpPDFkMdgQ824VM04RABk19s5
piwAfRFFF55LgkTtIghB1YrWRJ+G21lCI++e+pCNaXRBgltR3ryYj0PgWn3J40+n
9KTzQxnRcyw/1pw8WYbsFP6wzkBR8wRHupSIGbc/Uxw8aY9jDXjRvPGk1bA2w8Ix
lJzmAqI87FcAVI1d7fSiN56idtFYk2BTjYOV+TC7NrJFPvz8P1DhkuIqTVkX84wR
4DxqItan6I+C5h50b6NTMS9huA5pf06bF4bDbrlzCNfi4151zrNhmIjWzDgohH+5
0M97D1Ln6SzjCGgsIllwpkk+QP2j6Uz457XDu8paRA0IsGKE6xZHTMA0yyJMg9hd
CpJZI6/Y9JXjgNT2mJspIjjIW7VgzkyMI3VXxZSikvbv4oN8L1yGA4DZFLyocY2g
YYw/fIGjdEn3i85z728wZlOQwSwriPootQ+nBLPMXunp4E+eHXl/XIB0v1jLeKdD
MhMPCf37urpsZOBIpvk3gNnvN5QdWM3ZoxZdOFMCV9ND+dSCfoLMNO/KxoEsoJ4W
D60muhGijW5QmDuIpA9d0ZLUvNm8QMyhrtwSEgUBMT2s2N391yusq3adgHN/V90G
/cyymtLAK4pLj9Q54g/uflkmsypgbzpPfysna1foBZgvJTjgPBiOQRC5dxOo4Rbi
ILr8LtMxuMHjE58tqYtXoOqcMUsGEcERCbg2NiSj/utwigO3npG679GrOSd+OEY5
2n3qz15DO+w1sc0QcbHpeq7kHtokJ68+fX7cTNKji1ENn8XT9douwFKZLkGUiKO+
bHc/K/KPeBxCKbjHajUBdZiTZ6Zsx8nTf9f8xI9pZ9k7fpRfr8eVczsOWZdFyf6L
KeRN/w52FSx7Z4WgmryzaN+fgLghlev4VeP9lq84ZGFR4aws9ycc0/tLbwbkD6Fh
sIDuee41WKasN+bJPmsPH7tpVEpt1ldoLPrZHyuF2zKG0VdS8yaS7Y46fw5TAEeB
+dHf46szDxdFUmmlp9tzXgcYonlsKxsSFLVNEzmAkvExt3IhW9SFw/BIhZp+kkpH
AbTTjk4/4fqJZKAZ7eDTxpP5tZra/saSYGnSzUOuQH0iu5t+Ro3Gv1+3/W1qWcWp
mUlTO0vri14s63owm32wtu7tFD5dN0TELeHVLB7DX7j7cd29RuAx8ayO56ikXVQa
5Apox7UawL6ujjY0WU7PSyr/WHXdJZ2BSPpFTTBdKaguobLS+QynqsxjYbe+pygH
PCksHBAXJ2H6Oa8szOTOpOhJlv+CRzyXJixLbdTcJ3W22QO4s+LWu/4HVfMY/JGZ
Q/901KvhufkEk86oTv8nHqwMR9keSs6yXUx8IO3coRTsNyd28GbMVo5kznW6DfV3
jmCenDhQTDAMy3D0DVulVtcwgJzGyTfQENWN5flRFV9pB9sbeA2TQZU+slKiaaCK
W6jaJe2ahpv6s/6qd5y0tmlVx71blu9w0+NG2fg4u3yKw0PmmQh7IDOV/d+Pm1st
0fWiPLGNIvjMkGvqj3YOb1gDFeyG1oOGgUd8qQqgmSShKRjpR+JMJMKdlLIL2XQA
igJvY8tnI6qxO9s7QOY4o5lk6k6FXR9wPy1ohZ9PojYykI+GkFFUGSUtO7VrNzFU
Rl9u2FVVod0mU005IrZcxyLEhg35Rnfe4uGmtNjnPs1I3DsT5wbpOfINgBhwkhYY
y2vncf6RngKrm69wvFGIrHbksT6W2i+EHk5rJmfBGXzZzi75a5HmzkBIt35PPBG3
gMMHbXcDbReChry2MSBc4embskEPPrDz2X+yVbRDyT4cj/fNnMiGZg3nzi+eSrPQ
oE8VUzaThYSiy4ybyngWc/T2Ufm0jlYY7O2ZTzGIkHjPtLmdJ0TX9sv+gnS0ZhL3
H7w9y679ZTi0Nd6mflf5xauynCW/+kw3wUvW733f1/9hRnryZOoAiMpNOmfRfnp7
pMgBCmDr4rJmetg0EZXHU/ESMN3cSF8KwlYY41yDsl3xC/HBzlUClyb1aYv7LYLB
wSdrNyR3ZHSh3pTD/10U9amTnSZnk/EVcd2C8H9jxSk7HDYJwqlkuIxZuJ4fCrjw
VP5zsw1bmxrXrYDpP6R5qAYbcry959+a+mYU56kufpQsbf8t81+cqAZmvTHbXuDj
MHPGVTGY2bSiO3tnQmUai9YRF4kDf9gU0Z7EJ+TYwmxYW4uhxqsWOOCP+u8uTaCd
zF/GXZhKjDh88rCj6v/dG1pP2+rcIuLOTSiscGc59ePdiLD5MiAEiIAOCGRd/FC3
ySMSyQKQvx/oo3PMspbohrihfT1V2v2Ae/816bEfp9xTQTSBcy+ePJiI+IAIqKGl
dpDhg0MAgBKWA/oCkTGOs0EWcUMpVdU95ywDQ/ZIopr57aSG66wF3P0GWktTSNOW
Gt1iPJY23dhBJfV54jN2m3Uto6w7orSPbfL1Uz3czNNrNVYe+LsLdn2gj8BMUsx1
ISOAvNEnheI+ngZXZXb/wrVh4VPZLBTLstDsEo75U/yD7l/KF8mD65I+5l0R/iKy
4p1J23lrauTXz57VwTcbV3Puyam6cQBIQSk79+NUKDYGL0Ckf87z9pzMYNfImuWF
4NjYQBeCqIYFMa25X1Dk4a6S50xG26Wdd4c04mUXttJx890zg2XOwBvu0dVVjY8U
Dzm96SNlLXjx0SPbkW2QI9JeFeU+liPVtniAKzsR+mWTdRfkcdA3a2h98JuuZ3Eo
qf+yv2NERoa1dAm9Juk0BgJBNXX8IJ1i5V8KNIuNIBq4q+S5h2o/jANkll7SKsr/
xwojIiuaZGiL/YFVU09xpi5EYawt4l8MAcZ/+0pdJsCqZaff6nrBfrXLppjxj17N
68i6xoMQzHP4ccQZNxzapRTX78bPEOYf8AwYXMoina1oIhuOXHYMl+Eol9E1iOm8
rse+YPk144iqUI9QidLkGvzjISBovnpvIGahrvcKSXetwyDLXPLDoU6tasX+65c+
mxF+jxnF6FwRcfRAoiDaL3Q0pvcudkcRS4HzEOwZDa43FbqsffgzQ1wTVnc/kPnz
76Ox4M8EtneVM/RiPOG71gjiLU2ujPuzhoYRAExwQevOT/uvbLOg6+VMyMFOf7fM
6jueBLhxCfFmVJWpElfAsbL/Lky9+vDyRZVyph+4/Agndo40nXu40a8cZTxPlcXm
RxezO/8yMtyBWSvsefU0suYYLu8w5hq2eHHcMlPHsJcuezlkM3OeUSbziO36EXdS
HnvygGPBNUWDdy9d9b7KcFsfJ/rdllw0YlyPQ3Ga0++JWIqot30CHR2nGcGs7g4t
KkJ/BjnWRddD0bDwc1jvJkf2FcPJjdw1fqrzAv//9ljZ4NhTBOoDHUavXt9GR7zD
6G8M3Ok2c+N0edt7eHYwc/S0nPxJZOBk7eTteUF1m5nC3x+9F2HRkvGA3Z/MYo81
BbC2ll/ktFxzx7R4rPPzHNw3IGdu6gwo4dtt4p+aQT1SaGLnPAYjr/iZ56hMWETV
4iPvTMw91YxVAiS38m7OkUMuEDd/6b0AIACUgixfDhsx2obTCjYhD9ceJ4T/CJ6l
emXYhA9YomJLl5v06luzXerxSkIBP9P6uNrXxfLyDM+sm1XD/vVMYL4Bf86mHo5L
y3b6FkyFpBHNDBrjpFSzYFAISiRRnUWCZODOywSaiLLrlrGcJAXN9u5p5FynqKpN
yey1hZp+uPEiWB0ByiHdyqC3NCDapIGDoTkuGQ+FCBLNFY7wf2Fjc1hDhCHzMKNY
eCBtCPoe1pLNz5GWTz33R1JqkXeF86sICrtiqxdZZUnx+RqvoyTwIpuzfZ4sDcRH
YsDby8yS+ec1Xtuhg2Pd6tlrO3yFvlqWmZ6WU112m16tdbTyCigKlLiuc+PQm05U
uqBOsGny0wvJjBvxu/JSK6TmsqsNNHH0eLAnEckghuC5MXr1K0mP8E0TBfHqG6Za
ySOJxlUQY0ujwbQTtOggyy/I3quzAjmtdz3Ckid9gr8NridUXrIUNqEtuJG/3HSR
dFxMTnehEuSjXhcE3UXrSKRtFHzinaRedQ1k57TPPfLecaIGT81SxFC47MdOF1iE
yahaWDSujb5C7nb6V1E2hwv3hAAHUOVJbhCHdWe/+wLACRRr5r1yhNmvFLPSoFfH
MD3KIm+hXKw95D2TWlpRMRAmoKopiqtYnnlfCJmXBLw5erGEyCzr3UidPI6OkaBE
r9T0Upw2qqvmRCfgq2in/0Kb+Ztf2aBKrvvElfEpp4jW/h8xDDueR4JEUNVsumnd
NaiWSBFy7EgSuUChx2LrisoqeMRhBVtVKebS5NnTdzJ09j8ZA8b9ZFoxD88+bBWw
wHWR3R1R6HC1tA0XPmMWbkM3a6S+9tRKBxAxJFPW8/cNR9H55LYw/+P+rrm9391n
rM2lQ5r7gsgqP1ho7xEB3Z5gLb8zxOZ3UrAPCL6y8mqX2bzPTyCOM23wVkAhck8K
Nb2645+dA8AVpuAqYEBvZAPMpkiKNoeG9XyqP8u+DvkwHn/T+9UA00QDfLcKPcbW
nVk4wfcHKyPS/lNqKdmhni7tYxJ1OmGOxhGxD+medqAGmh9Z0fYQ9pYYspTJVjfo
FtP5JKurnvUpw9Q7ZgKefrItHMGCa9K1/aZv7vuSah50TQ4uJpn21rqGNqIoNx2/
X2LS90daf/LjvJTLZG3GyYk2Bp1UdqQlFcBgJFILpYTRWpVOhFLEkzTMY/BfkXKU
r8W41VElkptQN29jahPtjAxrcbXfMvab0Dhz8+bPT3h9pr8EFlbgtgOssT840mrH
aKcnO0yy9wa2MOGhnRaWGKBhbH2Iv7E7gfPkaZeajXutSowIvtCY7xEOpRlVHE6f
0fsd4eKxu5etFfzZT3PY14nQDasUT1jA2W7aFSn1oz50FcSavedupkvD0ArHJwyn
GudV2bGm8oHK87TYk0TwF4XwfR5rn3IXVPdLiswKdtlDtcOE6dpWg1kMybGG49D0
DlFT7STPK5W6kzaD1GkhvoGjkaIzd/DfHIbtfZo2S2bjGGbEQ4kTh3KunX+JL2Mp
z/D8Bm10E9iOccXLAy7dnAPQEDLgfyPVu5RAZ3iPkNa3tB5kvzAzFFUO925ZtmeP
YmMg3ylpw3zBbmPrqmdg2iGecU9MR3P+xnY4SdPjVjen0MHNc0bHS0eOIsrFLZ5c
wR3j88aFxHUD9nCnPtF1EJOgUhoPkFOd1jHhOWG5Tp9IGjakgSGgJwEJRdTDzbYZ
+ku920BSRPUjeQQrLXm/GWITQTo8zK3jKGOqll5lN9mNqGwkjVUWrzAMhLM/Ost8
p5obijhv1pjM9ZbvKrkxY0zFPXhu4cpccTuD5W4WtkC2c6ayZKQlqOpCj6rvBFjU
6ofdTzVP+gZtjSXyEsO4JoSHTfzISrtet5Jjel5b1rb2ePZ0faLXZ4faZ3RBbHFs
Qjk5DT4xRRdQ00rZhLMZg3Tsx8mZkh0rA43aMrnllSFoBfJYmVAulh0xcZOwkau7
8boS6f9IMoIlZnIKRK7isqAMpOnSyiR8bT007KSYzBLE+mp5fGQPC5mdzlitC6w+
aKhV9vACyEBDP0Ncb95A9+ndffevyMZXqqrdWrN3B1rdwaggmdCgQOgEbQursnTA
n6lNEB1Y27HcPCJ14v4yOLWBT3Iypvxjs/3PdbCb1p0ceRTHtbSOCOT48Tro767y
zV1r1YMBSS5ekmgM9ufwQXQvJxGzljcBzoQ8SjUYunXdYhEBESFYUT+Lzyn/8LjR
zJvagKvg2cu6jxZBA62JF5ETLZE+EjA99xNGco34erhyIO4UugUfdNsYg69fo16/
2nIP/dn2GRMAWV/Fa5lXH6Q8CtgKbc/DbQ8Ob3iKdZD0Qr8TzqTgL61qS6221Pep
kL2PSaRanNtOb0gIoM73cfUwoCmZ+vSHII7mYVuCw29DWYTQddDC/P8iS9Kdfwz9
+J2kkhOWNIUVyIJhUOqiRJ4o+wRcKW3CrjCcTVkQGChv8QtGfQxr3mf39PYRYvFW
roJGuU7j9Vhx/rZ3qvmBiCLb9TRqH2zYFqJEvLP/RMZ1/2rXRN/na5VKmZ5CnGz7
J/KIHPJCgACdLnN8fQHICZXuOgtEROMwfDJ+wBo0X8B17lv9Mc5LgVZU0sbl9yLy
C+tIxYORA3fLEtDdiuy+BwGTW19pFjSNP/WfoyZnQ9RtVFjCcNUaN0ONTvvgMyFY
7mKgG8rP9P9twxWy3g0lJsQeHVtS+hduGrHxaocX/nJG4ExG3aj3EsqYURq61thD
LJHOOvcPjs3WerQ9WhhT8kpkh1Q0F5aopnvNIhzg6Gorq56U0U5S4eycyfhulC83
15W3Iuq2/csOZoFEAPegy5ryVVsCbBfhG+Lm6AwcZPVSYpYM3XxANhZxBgJg2264
Zw95S9HZIPUFOEcB/hso++2/dKcaE0LpW8hSZp5RC26f64sxLSk1X/xD/8Xc75fY
rfvXllieJnIaZZUttqHtC9SLaQTm48fxreJo7obYcueU3o9FO3AUQAHOd9H3Mk64
VZ/p19LlQQjb78uCNr/dLiNu5FzGTGfK6SEq1HSI2TgOtkmJrIbCANoGRDKPV93h
a0Tq8UFnS8tQ4BbdVe9QVxIPteLVPRe4lg6dwBVcqLyO44MPw5sYHaKOU0LeX1Du
otGL5gYEAIcgCKpL9aYhWeULPZbuucyyH1RdW726iwFlhvtq6Y/ieJy2D0kwF01S
und3UTBnrs9pZpGBePM0XmQ2euEzwx7YKmqh2PfzSCmv7a5zykRooIbLdztvX1lx
P7VLlp2bCt33SvDp921XjCueI9Ni1uo6HN6en9RB+SK/52ta8U9wszE8KJanpe87
jl5ivINXswaZz58cBpgAZEIouNS+VihvQzQavV5DYtCg4blSU10SczeV+UuOeTqS
88DMT7ItZZqeMKE40kCFHeZJFbrWrsibRd83bf8fXWBzeIBAjQQww9pmZQQHX5Tk
s9/q5ZMe6e7DyrDv1WecLIfQFyeqbAMK3uvVrtFqX8h0Je4VvaLrMKnS1tcMzjJj
m2qyQeCytab08KkaW+HLlKGP6wKU9tp191QXZPSOo0tUWYDZfHws+5kBZ0qY3FEz
rR492FuMstU9LK5IDCLxftZXTQ7VlLTtW/DO1PCVB6f3TdbEG9i7LGRraaNifbdz
AqeNaJZ0I15O0E6XI1x9cAjaKMYTzeih0fZMHw6YlGi0VDuyiNvgrt44V1Fpgqpz
VWgdDfeKbeBhN2YnzEf8JykKtm5pNdcj3T9ycE5GeqbwY+OKZgUjIZ1CvOjo3y0p
NMr2n3v/CQUgOjJ7P4LKHZGlWwPDATHmSMPUOfWdnrk4AJ96ZNnBZrrNJWcJ6NrD
/6ty5MVjxDkixWMWb314RMiE8vc1yY+YQ/m17NOHM/MibrRTjvegoxCP7qqjLcnN
5or96Udsg6QPTglUKpl0ETWyPq+V6mXS7oM1JWAr4qinFDgj1umGVhq6CPe2AS5E
uxwBYixYyN0o83YM+xPpLFeLY0ealn1LspYvyhrvHaIFN8fHh0XQnHSGzkYW7u4D
6h2j2It+HK/G/6RduBHv7QNfs+Wbauy3cn3CUDIgZAKoMHrH8UJHOH/V7ja8CpnK
oarz2f2PjnVS/tjJ6+lhw9j3NzYEnW1ynZzo8tQf5Sr11m5IL+lxqZGVjGwAl91T
y7FU9jjV0fWY7dBdRf6yyj5yWAEHiil2s9A+JrVJ64ow+vWrlWYN9EzcUot6cCSL
db3utKy3zt/8SV6cqBbBKvhRaXOA66pWoota53TCav22aW2bhcxTWtm7dNtMisU7
ACez32Bgz+Ncy1AJ47cM+7uTYI9+ixpH8cEtYqM9zZTUhlInkH9uGfI2Wt4ag3Iy
NLPW73UpY1S9YP8uJO6wwPvjG8M+28HoM9I0OuwVzlarszIfB/5V4irA5vnNuYTh
j5YFnZpJ8UYrd02jNqCKlWT4Iv2JyvYXmH3y3pOWPgj421jqHrXYdhQ/6I1m5r81
sKqRo/M8gvPayUxPz6NXWIFXOcybGLntgL8FgC8lxXgWKT8+RkUkOO2qhGf6Zwte
8aw2yzrtq9brpwof31AOYMdkgjgIXEuWUuNC2Scz9dco7WgVVsstjjpMCvpEeSh4
EE9OfUTy2t85ZiXX6dOKNiidvdrs6rx6Ay2H1EI9wzy1+acOHLfozzCx/yzlcgVm
d5xUEp1qSSfXI2th4azjM/WlL7K49BUvJgP8IqEKyunjaj2sSe5mNQQD514H7mXP
IriXMo1BSAIzWT1aA7u2dqOnM+SwRvbuLIb1LjWlZEx9J6Ofw5QO9UtPa/19Q9IQ
1O7Hb63nAe0rzEZIPf1b3e1sqy44Ce0D+9OhVRuHLOZ+BjkO+GAvhzQLrRoFivSL
nokqwZZMPA+T4JigDOlYEzgNwsuMGGISKFWmGSyYMmn7bR9FPUb92lLVNQailOH2
6pokEUHeMCyT1BsW2s7bmrH0zBzxVepHSReRJJb2SP7pMQG2Oriqzfkt5BJWhadc
U4Tn7glUBgSRX1zOdjM1IYMk0NYQXqv8qHYklTAgJHHhge79L5BB1/Vq2HzR+6Gj
gfkHieg0jm9xMhrk0Crpm5C3dsoy847rbXFtjR2uz9f3N/qMAHByAWRWQ4+RAxAR
4j9yzYf1SNx4Xch053GZz5XjiffLvhNCJghKmNn4R7LrVbXplDWUQM+l9HrgnNtg
+4OQXc/YL68rC3fP8rolU+23V76vJe06BeBk4uVjU2SSmC+rMcSF8mUoBTVGTYsv
zDHPoS5PatuZ3FU8E1Y+ihXA4/zAjs3fxnAkC8QdUJQgPCSzIu5XBo72/WJqOtl8
YaYfJK9zolf8kFFZAbg5ztxrHVoyR5IPxvbE/5t53Csti9bF3K6klbvKy8f+LLu9
fTfcBMFoO3ltM7dhf5hvlM0gSgRYYFwtdrQHW1+mzokrzr8r9Wge4IHJ6/wuY4l1
USvWfILRKY6lwqJ0vbKLKvy9/I+npao2VPtRa+jThxF0MQweY5SpAdbzEBF5cEWT
u6etUJbYL2MEZXsu1OVObxDY8bXihsLqlE30Zuif8XzODBf8EfjUjF7lTxe/VmaN
sfNdrclFMn+bEH3AcLyjCzGg7l9Y3W3hpjCiIOBy6hqPCZ5bZggn9Xd9ipFXN24a
pxyhQ5uIh1p5+EgOYvJ2HCazWt8faPUx1OI7umLPrbepuLkFKek5Tda1WmeC9QoT
eAQLf3VjLv//wMlC2+dnpoVcRfplJfpwgR4Jgx6wpvB56Hp1LyeNHOk0yFUrmwYC
I6ZjW3E3IX1AeuXwzqdV3APS0X7fB7qKDEcR+fDc5AH/OotbYgE1Zt9ktLgfmPd2
VlnY086kAixW61l+OEcA03vMfxyaieF6mFjWqGVwEA2DBQECRplDTk+eWExolhOF
YXnodBcNxVnnzS1/Ju3ZUJ2MyJJyzQCCs39Whfw3LYfu6a7bZiRy/dfc3jV9unhM
ldrJzCp4xEbT+HrdE+z+zfcvrtA3H7u7+thMARuD132O7fzqpwU7fpLnbq55QC9v
aHzRKhsJoSb82lfhdw8JVGU06aDaHU1KkRd2aFORM2J3zyET5YbnPcWSMPtDc/lz
1mcaR3CHf5DjCNimfQHbQRWFtpiggrb+aMUb+jSTpSKMq8MfFKjLEfBY5VJqo0Y4
sjpYclPcXPZKRdUgwJlymVcs8QEWpwIf2IAjn6Xy2n/9y2CcSs/x3FsK8hTuxdGA
b+84YM26yjt+NkzN19CdH6OAkAZhPdHAe5Z13NNzbBs6Tr+NcPRePOIMCrz3Fxgv
UaZ3Dm60Pqt4hXfpEBScP0vtw9fqmAF6PW7WvMPvwSIw7IphELK7OP5lPEwsZy02
Mik5PHCIWqkXuWlHstc4/sufBlW4/RIDspMBzpzmtQR6dDfO52rJSM6SlH+3WmdB
xdMIH3jIi9m1k1pQPXgidczxuRH51xyuUfbJka2tqpY/+viHtee9T14YfS44earH
Y2wYQGo5InaZFP3SXFZxUQrDswrTzUWM/LzYlAMNosP9oqkC08AybE2/pIj9z7t7
Juiv4SNaAP0RDvutOA1KwVsxhxVseBdoM26buEjHZtXclBJveHl2P7PMhcYdfjUN
7n5o6CTMTdBzfmJaG+OduHa/XZyJuAXO506Uas0KtxhYfmxkhXAPpAOsf8rBbES7
bpLmXf7ThKPASJg0ruA19clkVuV9u2dpCuzglmmO0IX4vAWQV7pyMK60YKXnpeiG
wljLjsDTbOGxg3bthgZGmUPcuAScHgdQaFTqa4eqXj7f7VsW/rZMQOQXobJ48VGn
Kz7pSAbWM5xP+ZP0oAhRibM6Fit8CoZzMloP5RImhF/7Fo7CGsU4k64T4tjJ9Wdz
l5qQyxNwisTqg33lv6tZfgdZZe0wVS8HY5hJyiJgegdfgguSEyZtY1gS69U4FuX6
LgvXWC2ILTHc1vtLNHKa2LvMuHPzv27gRN8zTFFK015ubNnmf/FSSHXTBk8A3jR/
VjjEyegta19nr5D/SQMqN9hwclvxd3kbbguG58Fch7yVhRrFIwVBKQKFTczolFr5
vb65JdVF61WIw7K5zIMq72V6OB90qq9X1zQwKWIKONFkccLEOCOxu0ZLXhg17THy
z40T9FrmJ9pBFpH+lUFKsLBdu5ZyE8ZwOOCxBk1/RKJw7t0/aEyV2eeGf6gN2wds
hdCFDpgtMFiGyHG8mIiiMnLKzvbrRVbpAd0TcBe47KJol54MH6eQYPxZ6O2cMt5K
AfSHUpyE8+4fphK+DTyCzQI6eRtd1JfD6G6ntVJXO1QR0cKRj6LkbTk6IGFQvKrp
MTlJBU3pS0pWxvYcmmojivJhfCAB4qvebLmXUPyH+f2FQsB69qXq+FtB2uLcVjwy
vRr82TMO6wsqM+NutKaRxREYOgGii/SOXu7V9n33SuzTeMjdF1Q840w3VikSFwZX
32EeZlodXvJl37tCL9niTSFmZx/I9IxaGmKLfvlr/vKQo/9bmw0OLYgfg7haV8/g
dCBJILkBZFrIOn7dTsVuOVxqg+urV8lkD+a//9vSt2EJFFsj65yRfcZIGIqThkwG
PjIUJ1vlUXqUvYeIwx19baENXrlQqfjA1WDCip7LVSAtR8bv3tClsI+aXH7jNuAo
qIq+nuoKvzXjpIj4Ou7m8dGt773vJJDv5buWeBBjboy0pEvi80d8ryF6HmXitHpH
ayuBVaJUQhCYq0yl29nR8MolPcXsKxKSyvKD6LxjMsY1+zkkBZgbCTcD718eEUik
Y8BcpPssJK0ugawYq6JgJGUW5gvi/i6q0qSeFYhP/nxxhCreblPR1nEbOGbcOgLE
owWTlMLqWUsfPuBSNeztXedgcLS6pfH7aIXl8KkPmJNlbjg0LUzeK49OcZk5p4pt
hIQQlgifESXBY69ZTCg4/AeAHSewu1p3+yEmUEjOrhgzIIkj4NnedymooqDm+kbQ
wjO7cIpclLU9KZ+jp7XlC79Rbn4oFZjMRn9YKgMBC46hY4YrY4Z0eHrC8zWbG55M
G18KrkzZ1Xdywh9/xOVlFdjulQCknktD23+WwYEJF5HDTF0zeJ2TOQOdk4NTM583
M9W0VmX/hRlwIBdIcTI86l0eMP2cQjHIi+6wogf653TlgHosKZwjSxKw1x0woepB
r8I8/T2BOx/DisS1RVrrthIfHDIiJUGaBo/2rzEy6jrqGaYrv5CD5rYL16HHX7oM
6xbmvGOFRhQ9DmBNH/O+IoQ85ar0Wc0SlF9pKkrqwUdhKUla39ABF+tc65A1Dbdr
UHWIn18TABk3OA+Zz5ISYQKSiuadRQ7lY0sjFjKDZ1hcQK47/B/4/9eJ+zbnU9Vk
vNB9VrlhbMpAV22vkuXLTt0OHRAYxk7ojV0TfUjc75VmioJQ2ttXUyY7Wf+i8kYN
Os9cyOsBe9cfRx8GoX8h0X3nSi3EdesAzG1uJ0Z2ozMWBfPQ1/mZ/iQ7v1lTBXYc
30tJX7OJIfLmEF+Es4Xe4vkd3wnJ2j+L5m3hddy60oMRFmaOMascaGYaOC3aU8fs
RXI0CiqXtKPV69kywL65rBvfM5sIyLyvbvlHEQ58kVRaKCVwYnxS6tt9hrCyN0wl
LeiF4jHeI9AYW8Frv0XjAv1dQOYmUzuFOlLwDYBmu7EkvmOdeOeFwx7Wn5JCS0Ml
5b2owmCsJY5guncxYgsY+oAeC9lYCFS0JbKiJGWjZ8NraL2R8jboZDziTnR5OMEs
CLw37wID5KP8LY8h6YpS/KbR8DVGPBnBhmVr8/ppylMYUspbPbASzR5AdBxF2s6Z
4D0JGiiaJqVUHFSDUreX0xx1Yn4uLQN9VdzzFMjOzKo2be8s91pelgge1MrV9XaH
4MmxWVVdobjEZe/M8iazPAWdLuJkld80W312BS3KbNjuHoPVPhowz4GlbNoRu+jy
LjGIN8945ZWPrMFJIq9e3f/mwQerH/MZ/39tofnS7+Yq4ZjNjfDyW0UTWT4eawRN
HHSruNutQUZr5uIFoFWzJJni6Yn0RPX1Ro703/K7ddMHxYdcp4Hr3qBLsIzQ59IX
XLSJDMQ1ceejmR6Z0b9nIrObtq98jHVdoMjIGbzkjgfg1UFnvK9L57+/7hKi/3H3
e5tWCDRV6aD7tqs+YxPEjmwHon5KShNaFiCffUkp7tMrQXDTC9RACsG3UE6NOZa3
UeNH+sfN1SUqJmUmkktVE5mZ4Jc/kEu77kCxwMYDcZVl7gRq7h0RpBQMhUXYsnt5
AnZZ9Z88BdSk8GiRCe4kVfIgbaV9Sg750qG/9l7IMR9EAJlifscNXko6CvOvtbKB
Gh6a9Ml5MF1uOz+yvw9IMIWoKbc+2TUic7AJBXJIRmGxAZYA53jxoiIzOtZ1+Son
aYf6IiYQJjzOyTZL2QNdDLQKbnyhee6PpC6LyH2QHCLa9mrBwZ7q1HRfraFPhuHJ
61O2I1bJ95dmU62ao3LZiyowRXB8cnPkk9u+yawR86GxrgIwHE0CNvROTzhqFd3N
b+l+6tq+4BBs9p5Q9chbNsRMaYY050tpSuuan7eT3E6R3tjBV79EXp3R9uICPteY
TWonNI+mrjpZKRyUW+AmIAWYGDLEuX9V9fCKtxWpdrCHoLKL/zx9TbmrYFVcp5CC
egddphWz2l7hfmtJvuWg4sOB+zWfox1FGGcmnBOKTg6/JtVqTzOF5PtuUpKD0109
vh8s2nPBWaIqXZOOnSKzqA1avX8EmV9BIA0siD8SjVBuBhMJBSrF89OJkbs38lko
yGPAZHK0eOU1nZ8cGKBzEwmdoA74yO/ifuyrnTPPrFLplPqFHKIRnGo0wyofOgrm
eswj4w+kBwS29jb4MTTWzeC3S3ulXoZivW8qTNVOBZT/Ah7IGitR5mENWvkQf1Zn
Xbv0VkATOr2qHRgtrWNh320LdxJamhINzpHGIgkAawqp4BwPITz5u1vmGMETtrNt
s9UqRKN1Jxf/dF5q9vGhZ9oXsdVoFGcE9ZHTulbaqxaTs2WeYqO1S4BJSkefLXRt
MhAJAZMwKu9eYppTy5EmaWjKDegJfVnaUHklfub1I2YTGCOwaMlwLYeLLBwlJRNx
eqj4yOMRI3Jb6LtsQs7Axx/A1Z3j4HHyzveYygkAJlhp7WI6X0tDIFwA/idrUwvZ
8Ieze3Ctts5vNQaeIDWQ3PjJqSyHXSPYMqTaP6B2SL0qo0zxFB/NkYoZMNF09fKg
Z+B32ajKj4YydhLbIDpTmkMniOXtt0GkRwaG5ergIrxDrXLeHfi7C1h4McpOjv9L
YD9y95aoxjVADh0qNq7Kdjs4rQujTkhR3cBtZGlzRoTZg78P4j+AdJW2pd2Oy2kl
NTKfG/ESGTH3vYzV1H7Ly4YF05dGm8tJEcHh/oxM9Yv5F+pgI69sjs0zbAwSl2D0
NeREZBLEbB3vFH7uRZnHYGbOYCbrIFoMGixjMo2fBDkV5QdfnH2WOcRGEHiAiDjT
1VAZE3B3NHTT8PMQ3Qpty+5QINnllmsJbW9hT1LojZigiHGeP0/PfsctmheSpZYG
cQZHSVMKd6VyVg/SUOeKTWRc310ZzjHER95mIrp8IjrW4TfnZrkhJy+ZQM5yLM0I
jx/nNDpgiqoZA9N5saHvO/1TNsVmBnjXKXr9O2JIvla1I8HbqXIVWvioXNVTF6+u
vubbZN46EJINWSqJ6fHv3L1b1Wa8EkAjTZGERyZlc1UoqiYYAc5LQwnG3i4673He
koUqTB88ewrV7qKf4sa/dplmc2fVA4kSUuBeU3AHATEXtcBKP5PDHOwNuHxS45pr
TPjNy9al7qaOsp7UF+QA0D9GVlfeNMjcUxOB21Z1GsP8dsDh1UEo9WsZJSZYGrGZ
2GVuMPdUCrFfaiMZMEnAMpY6LZcatNTEa5TtbWsdn6vLJ6LXcBs6jyi+NDDPsR/k
i/gsmvG+D3BKoE/fnM+s6GioOz2eeqzLXLhm1XWi/RP8b/IHbOxmiXwFO0+RmsqV
mI1fsxnBWANWrdjoNlNs8kt5JQdtoeKSh1XKnL0N+zcDZp9cRDkFsYCTZU1lcZTU
O7V0Ga9UKfvmoETtEzxyMmYRfKbIdG26jp7dQDdK81hbYrZADrNqtcicRnPMiVig
V/qYv9Ke+wM+iCco5qoahXxqRigZ5iUeVLyZ60AjKe3PwYA4/mrmKrggAIeWvpd+
IlDHrsht5tjKRdv/bcqlJfiWejUcmHs4d7IAJLPgXQJWLSsOQDeZ4MLDJQd3D+0N
1ZCU9CIdX49gUFQQIg9JWjhGRP8pAlAh8eY4itdDD+4969b/zhT09+eyjX2Ma6GO
jV7SdxOGqPSLom8CVDFv9LNx1bgZvU9lUCXHCIerFNc4a9rlpNHjoGVvGAcggYzm
vfwTbUWf4r0fCalURH4Z4ugEQKzYXkI9dS/uHzzcO1pcZ94DwQZz5zIxug40VUdZ
KW5hHHuTLMF+5tZDwvQMnG/+HQ70RSW1376YP+i33urVoVJALFiecjSwRvUhZvbD
X2+kg7q5mIy+sA/Scxbv1Xu0xeTHQBlzhM5kMCr+8EO1xQ0op8Kbnlithzy/gB4M
//aWhBGOK92iz+D5bt2QGYF+vSFxMF1qbKwCM4vqXntZ5ZotJxBYH82XvxXC9T0V
77J5bZ/GrS8qlH8KuHqQeyUcHqbHvPFbtQpEkXHiBOlGD72kIlzJIn3HWI6tzY/D
2IudLc6JetIYq64Hr7pB7dX/SB/I04gn7LIgTEIcki56/Do7t7zEHA+C+szj/mJM
e6llmGRW6wV6G2/iWnVohBf7VsUH3iRSZvtSByY5s51L4pz3xGLkjPf0HA8yByYB
fTpJQNUTANF3OEgc5CKfCrijiXKg6rknmzPX+wp5dIix5eA1FJU+c8jSl9OFe/4d
QJA5EDbDK0DDYBLTHwWaX4smDBwOrnH9OMGrYrg3EXpqCBC2mTobPpPv5SOggrrw
pz/TEl4naWt1RaPbZxQ9JNIej4Pvg0ZoLdTtf0yl3ymLpWUDSdv6jAftf9Bu/nAL
oXYWsUi7U6MWIJVCgGDy8/mngOQ2z8dIDY0MSaVCF2X6j7ZqyBMXAGwBXOF4I7db
doy3W7L8goJ1ODACz1F2WzmYyJz7FS8Ou/sNy5N80Y9joYT48HCq2nQE+1yWVy+K
e/jlGLn+E2DsS5YaDh6OKL7SNMeGb97jK5G1FxGlhB3RQqDovgNLim9xN9R48qyu
1Vdil7AB6yMQvez8YFhz4RMJi0fhzKeCNK/ffTbMwhCMq448Idvgu4ixm2f6gKOO
gmcJZ6xuDpMXasUFs0hk5NVDyPwGxQ8M+Moq890I0bNJqhQXcMrhOcVR50tu39bM
uLVqYF/PLlLFa7kI4WVbHgLSll+jxKz9ak+Yt/lhBtxjjQlajyKnPeF9ahi1uOsW
k7Xbo3udvNbpYNm4UAv1H0O8KN2+DCoWlKimkBIbn37yXZ1qFhQi3NvNHB9NaUK8
XKt7FjUKmuYW6LeymCtlrmEsGM+REW0nBhuA/RguoZ/N1mvBlGyDZNOXQ7Hc4nMD
Uh62VUeKUCkfJWiCazBIqZsmShLhjGHGds8QYla4wQrfoqipJqYjy8WcXQyW9di3
YEOoll+iNhdCzSItndRdPfkJ1r6YEEFEdaDgIhYwyndMMx5WeQ2tSdKHEymVOzlP
DQsfog2WRHYPgJ9mNok55QfNWXaPPhZgvYoP+WsMBW1ZpvSe0zoF50KRCGsm0jCZ
gfCcOMhYagoptXnPN1W3NcjYUR7S7vJZac7/QMcnFOvLBSSO4DUxX5YDBHigSNoT
Xku91XcXWWXXl2TvYDakwLlU3KYOQS+ZpjOxPZuGK3dYIXnwBTSsy0a64viJ6/8t
VEK4tVqmUyDYsUho8wXzHb7c7tdIR2w5wXOGFwOXI5xYOnc+BHwDmrrk0EU2YhHL
B7t/39uEBOHISZ8zrCRuHHBPWmBzZKMVF1KVsid4fFm/Tx+XSg/fOT6CcdaeG1xQ
hu0fl4ya2opA5jui5PPuYmfw6C2tT2I+Nyf7X07CbWE8FihxqFaJv4KU7Jvtxc8e
nVBuiqyTNAAvam56zwiYh4Luk6CCLeN0PSYJaSBb+19T7rPgB0SqKB0YWwShSlRZ
mbu3Hi2ch2E4YMI+IvGzcJDcU90fE0pKRLhO/I4JRK0aiEoR1i2Izf/Vnek7tyA1
CENgXSLOrYFptcDe4mzBp/fnzUWEjZ7/h13w+H10H0byZkB5mNhG9G1FUSpT1XxV
JSRE6lwNT2d+Ljzos26z5O8ZI17M3cWD2NL1NR0eGvkw8CJGpuLX1MzprKtVYdLr
1Enx9w6cnLmOY5hF6k2caoq9COEEILr5aEQ8H2vF8CO7wwZqzVHOW8w7uvNVMwgh
4WYoMTesKo/WCB3NGWNEbcMJIv+CtuMWULxJ1z7IO10d5WCDIQA7LxuzMO3lPFgP
RO/eKSuVzZDTos6tE9PKXnD9J2jN0rKe8cFThcAiP0kP9OLy+Midlz2Lg2sRKH3j
P1/AQznp5vzghMtU5pD3nVodQ44GEDFjjj5A/fAGwKPihMzx/eiMucB9mFAZJlyH
y7noLqV69+NsIBfsfBXkLqqOv+71T8uR1e65xA5vvXhr0khNO3IeuIs4MhL2bd6R
aThabFVFVFFoB7WhaB92bkx8Fu6nbEJi1kINk0wnd56wAZ4L4/emBcHEP4fFPjD+
Cc9sW3jmntSHXUXpxcLWESsNa5MJUbZWpj/XYAnTnJMV4T58wPmtPEV9Yz6NsbfQ
o4PwVXD8pDAUd/DrJ0n/sSNqFroKbilZFHyl4YSiETBdSD16nNDSaFeWdTeccZeo
9WPP6QXlS4x97Bj7A//auJ+v1dlXVfs/V6alc9WJftksYDWa60KeBrvCwxKhAE70
X4YBek9AuBzeWVmpJJsCVivRJYoBuYuKd1hUQsnZa4nzpvYvgYqGhnjXsOa6vXwD
s2YSgYLuIHwOoH3P1DItktY1MNg4rSflvx5s21Caw6rp0v1Crq/YZx2bt9s0dbOL
J5usHsJSGk4j/YgoJ9GP5HhziXN0RtMLSNMjjC2RWlRnIXy1bJEP7ihSZs0/AHyB
U00+6wSy5g9gabv+ERCLB5s0qvMppB+99EIL/1A4e/D4Z85BQl5y1Ch4zD5+F0bg
DLWeBpgWruPQyZeYh84+X7iooS/s4s8b7NCO60VK2od7mvu0Jw74mhGV0iuK1qXv
cQs4xQBnz0gY6UDdL6mmcEj8z6wh7saY7YkFGJ5qgCqlF3nJBLVa/cPuS1fL9JAU
dO64884liGgR00fclgirFdpS93J0aBNZD+gvonaQ7jbeH5txtIcQMLg8zGSZlTuy
VWo4KTGMgzl8QVsMy89a7S+urYKPLmMQ+1M9sP/8lbxNsHOfwjZ3AAdreky1solj
asfXz38t0qFhOnl+UsyfcDcp7d5rH/OfHbHhqIgNPb1n6dfALF3QoS3t7wyTzP3E
jZJ5f0cEYZw23VYkV1vPVGwBVw0ca/OFm2aZu2ucSoAe+j1BDTTU0lt9nMlaeuIr
q0+9hBpQZJdtYf8RGcVodQuoznWqT1Yt4Jo1o97SpLLe0SM/ywi1SXQEFpfh2zk/
nafhhqTEkHz33EpTc6YLipXEssT4BXQhSMbqn9L0TzeqdFoFgPeuAZgeIbJ6LnhJ
He9oKV2ErpY487xxkh7mhvibaGpCPSgspu5didqEZi+9EsQLuKtEKVW03Cr24y7m
ZKcK9bQDxCxiEqC+W3Akv/0YCQbMR/OyVFrcBXIx5FTuVY+bwpuILnsN9WwKEml5
cJBjwkg8YdlO0COxbPKJkZF/UqnSsOBBdYkd2+sv1OybzvRUeUgvPXmQE6TJ+2k/
Z0XRV7WnmjCxajiF3ui4pPVw1KdGcpNH1fZeW3S62sO0zFyItP8HZVlPMxdKh1jT
a9ItwOahOyOouDFyk1NIdOXVlzM0P6cgQ6M8kPqkJlmrkobiTuKGX8WsIKlRD5e1
uLp1GIB8/ZwVxc4657zaHxfBN+tVLrdvvUO20FeOHPcGCupJBtYI84mzhDeTB1Dl
Q/48NYSzEnvxFybWbyMfnQC8MCLPdCho+Yb2EKTHAtCM6x0jpvapnQ49lvNuVOBN
2qJW9BpIoFKHsEn2CbwQpFvteWtK0V3D2mJ9kjhQagGW0hQxmKAccaQHu4myAFj8
LkyWBQS6BnVby0r6UPxy9j/PLjIV7mGk+Z4WOH6vXXJFOIKIcf4RCvYmgcGX5BAH
YIy6OezF1fzeuUuCfkTfcXu/J54Kj8k6bFF7PW6t66/91OC1e6O5CQ4YQ3OxnTUF
HZIMFcPuBtWwESRXgZsoQkPr4HGQ0u/3EU/6HwvJKK9uLLOl4ttvFZTwlPRXxUMd
sFiqb8Wo64Y9WwavxA5dJBqR7mYy6xkTh2FYjzlLrhunlba8JraUdUqeAsTyH9qF
hiBSCwCwhoYHEPwPpUhu+98PsLZb25fkK3HpRo5gShw8pDCAfL5Beiu9LsC7SYmZ
3+PehvFAynYQNOwaXZx+q5dsCjNGxEPIGp7IfefaWo/6qhA/IZDzRzkKnjCgDEzP
9AZb4d4r8wpbF0fl5UhmEoy9b8/cHMyDdtbRIhSE7adaKvVfizruJDs6DFOJ+WVP
Oq7eXLeWpBnhx5QO+G8fbm3EiinDEZqr22k2eEBPiXzni09e5jME61QIdEr5Hd2/
pNEUHbVaN6kSou60GKEa0/2K5CbVwAqIfMJmOH9G9QHa3x02yYk+q7QSrLLZohlU
+oTbDulqVpr42pw5BZBjLhwlclXY2+l0A7d2QWpxEYO4LCGvXGGSq5dTvNVUvuyB
yKxukiHRWNxaoxIdDepevIqTEGX05oFfNK0Z4ZRW3/1ZTeIt7iMWxjAHtBiG2Odb
H6yrz6YFkjWcBARglTg1eX21fpS5fWhY4S+bUSX6SSCHQspQW2YSz+zagVSVwJxm
SDTjrXlsmJI1a6Hy6zC4Eue1wOQ0qDo0B2Lbn35P4l7UwK8JgL3IMOod7basbNEb
72FI7X0AQiWzX76+AH0T9hKaymGei3FXeWsxncX+YKhd+762FGaie68d5teUyklW
F2WnBXmrnaRWpMUrK7i8nhfrwyuDGBqwJC5821IDpZq8gViX4spnwi4ZaEaAe21S
nR4Ob2gH5frPQ9IC9OticWlEVMvoA2ebC6ADXQp9s59j8SLU1VdqTjdFyq13pjws
1yNB/IITIN/LT7IjZ7Gb+02zAUuTkGST1JxzOjEujox8E3vyy1Vislw9pU7KcIYR
fB1vh9bQYLk9ca/d1oh9ur4KvXvKyo0mTTE03NqjMJsBtdZqQA/lLud6HfI12vsK
d/HC6lM6IrEx75LDTEOVuYxD8kGtxLhLHJ/dRrWwnuYekcxjUAgnJkFoiSRIFTv2
U9kXjUMgx5WvHmfV3QEhraoRRg9qcVFTa4R9MXrsBqHYzkvAb5FdzD4BDtCyx4/2
8g69qzsYBgugp8j0X9ESa1/f0YCt/Efa/F+983bPXM1waoY4TiZ4vAaWp+5Ve6dC
JSwK3sMrHhzx9wymKfsIsd7maMz6qqeXRJZLkf2+ddrareSF+EGlDBtLj57m1tky
2ELMLCk927idZbyb65fpABXZVA0HiBdofKzhD6uw2Ks6Ad4KP4LXfToQ1DwI09oK
fiNGF6R9rCXqLKlZZf686uKJNCuP3YVOHaJj2aj4F0IU1wwET7fXz4lBHLUjTBC3
GSP5Xj9tvIVaAsOvSAaKUHNBENyEf8/cUaM4rKifIfkCIpmNhqGCvtKF9Mh/o9vk
DiS5SAD+zOFx+MByFiDcIcVdIWqL2wlN9UkxmbNJavzuFN8gzMLYFpVO2O0Ue99k
YrQYTqKAxGs6M3gRzpjZnT+PIz5DT8UW1UV8LyFD/nP5sGspTXUcWOVTRsqth+Ft
jsN+iLAL5LnTDA1rjTMCMkhbPXMoa3zpOpTM8fp63BmSTxYKkh+RWmbgf2kTp++r
/KbfAlTe8TtkbTofq3TNmRvBOEjyVm0EhGWSag7NuqF/tuoXBwtKk/k6UWb8Qxag
1drGdOPghtLFrrmIYSPtZt7I2PqSw/mbTXC3DZa3UfdJgLN79Brv1mBO86xKpLdC
BxPNRMhhj9/h5anzaHPyLYCDN6RevSojY5ys9IX0qYSPzuaMqOtW24M8iZ1XKUpv
hJ3PEadF9eF3tKfZIsCFvM5lE4GoxcXDojpn96QKIBsaNgRmIo91sbQxDvovplAM
iBnlPTovb4QUyfT3vCtypJksz/OqcOvfqOzSyX16iP0IZLdY4KpzVjKiH8CxwuqI
YKM8gU6MmdgilTYXOmRX5v5AoybU/Kv9WGCwQYUmJwXFDTshp2ai7zcVV1X41yeH
tH9i1LAK/PpqxbD8hiyCcOkFsGgDGF8gIS5/EfzXmvNkzWK0tL9+7NlYd652WZJX
pbV1qWDZ+AA3askOLZs4P4yASk7yY+2HnC81hD/v7C8i3goTuwSWk4myvB7O4CyY
lATrtH1WFkqUKdxyxWNHxac0HUr9KLxyB19RdPuvITWRCS11r4AAf1pLv7lvuv1i
4ZbeAxOeoEmhtmYFuEB7fQIg71PyBjLZc2nRSIGmLeJW1AOnjZQ9znJf5jgE80ea
tnkzK8oZEd4mgwsNE+mYL+2R2sr2LBDWSpWGkss1nqBSYgt0cICEGtqS/fqOlAT1
5m/0fofHEqW4KTCv0MaOS6gg2ziSJ0bmgW2abuqtPRkFY/VA6EXjmLOHU9Pb2LJu
uILf3Tvidf6Qr0QQuoZ6Pp4dYEtQH/TiBjQN8hfzk53rDJRjGynthijs+7gMYlmi
1MPbtkmikDM/oqs/cnHBiEvy7yr+Ct1qBA/lbV5R06DyvC6v8vGb9w0RE6ZaPCkQ
parXRVgIliJcL3M4tp8NAO2Jx8Cd8rF8DXc/rcypsfsn86wPy6PkXBrP8oPpdoam
p8/MUxLRlbfANt8n6xMVJEtRiwvMG59RypFyerF8dMyoD2Z4FEGUkHTlSbn6ewAS
9nEIcPOimYAq+pGwaQgy0hsg3c4rNYejWfFpYQ07uWg50x+Afg72JaOdBCEAauJe
iCfg7AW2oeuu7ayAbOta4PFiUoSHyNOuADDo/nOPIClwu+MXqbSK8ig6xl/28ibJ
O6kKjjMgZT6vy0R4AMh6JQD5a6S9PLNTedQx+rn5aaVxiLqAgL9iZcE81QRiJihh
bgHUqP0anUeTnaGes8mQPAlyYk6FRRK8yhGWJbY1eMCvePcqbidHFseghPUZR9zQ
Y6zebThOqxDKujyTJm0rnSjik4kq1HS/I6dll2is0DsBT2lhbdMF/YgmxBU8CR6A
xiQSCITxUwotTykzqPtKVVU1O5brKXy/HAcWaR2CJZC+grYAB1J4v53M+m0HlVoF
ZJ5kuxCNmawL00Nt6Gm/h4OkSL0ofDctLiP9CSlJwQVgsolWsiiUEt2EkiwfehFx
CTNmOXFOXKuJ26d4O0q09Ea82k7HmmifDifAdwm24tObrlZSQs+cUj05Yps2p+HS
9g3rA4LwalUXbiYf+yRNfHx2DPlUk9v01+AmhcyI8VQxcBOTM0lfmS0VgJE9bHDN
UV/QY8obkiJ1JNvOLrbxMCMNdLsyMauqo4bp7seeIsFqRILyAnw/Qyh2LEEBN+X1
CwHLQ9ezUovqP0I9SF/GN7oHhMDq0IxjNToAAApCBUyF0lFSvgxB0U5710NOC96z
uDMPffncYxK1wCnSi54Ev+GDyDmIDLoaM3/X/mEyru/dhspvhnxsHW48m8udignF
C3GWdDxLIrTTI/lHK2kT4YsCJvwubjNCvXX4BRfw8PxE/765t0ZFVd14gfxEWrCb
22a/50nUi8dFzMslLssjXXW2uIefZHt/aFi6I85ujWvX2yYs5Hpud6tlzOuZ8uCB
qhEsYbJ5JCDpw6AJeOmBWqVN4fuXWOkVnnQFPdJY/pTwk/YVTlRsDigN6dsMG5sN
nur02gs6qdOt2xQ0ByYzGAaM0WuyBVcsx9JD//BKvBIkDGV+N8ejMzwHnQVm7Tvp
6pWgZPnGM4MDzCvO5DKKgMeKaW4BalDNXXm/r+/AHsgGk20HGNf9q7xnFdYLUU4h
HczNs4JgLHYGt/cUch5SrWmFqfI/CpymrzMeC+F6okCFBmE3/uwXypvORBUgexQJ
0QcIIfvuDCly/uNhD3sbAryKAyQDzeg6MLngNwHGGSI2qNa9vHCpSwFjNomsXZ4R
OrLNh5nkQ5LbbwX+YU9LZzZC15tfUpCG/3Xnq7R20idZwkHTu6CHAgyTEmnipV0l
xNg0LQWYLve3lIP/fBqlJzDZUMq95sog+mFjA8rJbiRCC3uFsmFdFrNSdrfosPqa
21ygrCJTLioTw0hlKbC2eIja/QGkR8ZJ8xojcia8LB5IgAXj8wBXAEX9XVV8l57t
6rJeRJ15VOGRCvPjlvko92qGIheKwZjxDVBLmmKNXTFs7Bjqan5iRnGMWPv/JTHi
/hSLH2Wd1qZYKIe6q//8xFlZuIp3DXFpTuT1eNvFm3FR++PR3eXUw2UBG0PCEPyY
Tio/xEbeyDCm+ZHcGR7i6UZO0nwx6ZeJKaE/hkmUjrKoqS/N0et6Raw1f9V5CImf
40GxwpXY6BdlT4Grv0fNHmEJIFvHhmrMHD26RURno+Zf5Au6/XGvsnJxXCWRFvq4
FNBYTWyGdpB/omsugbDMHNBNPLbOUnGZMcx7ldzlJVRRhehSDO8wRi5gmjqIlSFj
kiGhW+WZqEJbQdl0oGZaZKVPmel6A9od1B4TyKzegicBjt2NxUgL3x+9Je1mAJ3z
6v+II3O3ihJ0BqhrkXGFQsun1CndSYpYjEU+xZss0kVypO3sm4wuFzWyHjZZ+Fqy
HeX2+mzXFS8nuQuMfmvvYz8aN1Fmt3N2TLS0VoLiKfAeBMRf/L7enTquz2xQZRyG
4ucEdBliM7P3YN7b1MuNXGkeLsmMVaGe3LUO6IPNDRnLlX2z5lcjes8YqDqMychK
6eJw2DkCO6Rl45RA1ETiCbJ7b7+CHatVChLV2vNMIOkFsLWm4N+OPYPHsgD6Y7UR
bcY9qlayFiguFV+HnZH35OYBt54Pe/F31Aaeupg3wfo5cCSCmYGVxGRhWeDSw0HV
9kQyCKriSOJjN9KnDUgZLbRJx7YE7+S3MvlZTv5pvVp9SxzVU0gPwi2j7uZg2bjN
eVyBbMRzsvq8ZbPeyWYi2irvcu4nyccvAfzBefFWr6IrGkkuqIVx+ue4UEBpd2Ep
zHUR4gEOAZwnukrMt5IIBLtUmBUQVyy8izC10v9mbhidExN/05kCsWfswBrI7ibF
sb8fbeGJIJz3Jf0+S45gcowASaK6aOro4V1fAhn26N17jaQolL53q8Ch6va2e12I
KUX4tdYEDDATHzIq53IfWvx1H/5XxbC3qz+L8knh/mV6L3/1Hvow8MmbCbQYOlzj
Ozzb3InTKApPvCrNwb9VKFNaJr/2gOE+5/WPHjV3bnuIhsf2IFI53mCi1lXOG99X
bIjSB/ayU4m5EPS5kxh2PNVkburQSR70vu33p8tWEd0UKzggaKGF3yEqt1FhL4et
QQEp+zkexGmOHv8JQF0tDMQ0i74jel2EyPNkSb7TOHYiZv6iok2DSleVN9B9Ay0f
bQ3fez9O0RnKC8rV6Rlu/MV48yZ14O56kJxrH+TrYKcHNJLWBliYlVnEuhfejW5t
piIb2MzZ0hV+a3Cah7+SVb/JYhHVgLoGd+O3gSHlkyrIuZJF9fwIDWZnkb9Ozzmt
WHnZn34oZhpvoxc1NVHxjQqwPpU/i9A/neCIjIzCcw1mer4UBcMS4eSWTIAzWHKA
PEmzTpiqwBP84VdTzTLFYCTU7EeBZgdUV8KH/7SHLU+ZAtsbI3kOfCatokjw9TWv
+xERw2xeuFQNa6M4vTDghS0PR52+dGjSS/LNy6F1yrGwfq+vT0E9R2ZUEPuqGvhL
Yiw9YICbinlYdKddEgbpk8US0xkWst6Qgu/l4LfxXkHSprVo7EmZtyveuZTDeQN5
3K/JdAMXaabWB3qwnYFghRpSHfOCvx2ZQuI7h+CPuk+STiZRDqUbZehPliWCv1QS
lFj3jUHdeDt7p3E1mF5aZG0bDfuf7DFDmb9SiOyrPl+h8Xo0U2hn6U8+BqEWr/I1
g93LSRlZC1N4p4polCuDAuZ9VzVPyEdaG2Yni2Dqok5rS9Nhf2h3EauKaG5/rjnA
xn3aYUkpXNCMmdLHwxJ33Grwfogr1za+P41RDuMxK4c927ToeXZ8X8OTdh1LURJc
Z1XzILo9kChGmruvFGe3ixZDvgkDwoZBDB9b4GpA5dAmOV6ytAzSXABO5xQA/cub
HEfbESmiHtaORjnB0HkLt6bTec9yUsksi9O0ziuAJI10Cng5+JRRfyfGXtq0mHH3
6pHxE+B+gge4MuS+QETOwsGDElQNV+wwhLh0h57zy11oHifq7SQ4jAocbNXa8Nn3
AsMZxp9LIZspQqBhTWsaj8kGd2M3skskjf4qgFf29fQTlSBwo6jH4hFhHz58ue9H
GLn4B+XNJrLWFLhA8sOs3al0gJdIMvk55cwK7aS1z6rZMor0gB2psv+0nmSN+/s4
bqz5noPVxwXHgKJbPiBw753du8PTFBRxj5peweBBHafpsmdtHhbW6CxnFCvwPWlW
02F/nIsTkNuJHjJ+dg1GIyknhLYedkP62jrsAc0OejXaBePokSmiHqTmWzL9i4Hn
DyO6XIKtiUZEku3OeLCIPuzI4PU0uvnuPW1MAL80PBx0HyTO/mGodPOS5jX62lBc
+s/RNuVJmG6D0OfKrHpKdFKmYCIBJVte9/IVTLqTMUgrfBGoCrtdpNq38gB85C/2
NlmFqDrAibBZwkx6Z+3ckd0Ag1lI05XlJSW3ssBgx4/IRZ2nqdJqYa9ywESQQ607
tAKTHBuFFbBF+gYH1ltrSgZ6bveLO1uO6hG6ittkJdDN0VwsBVMBNSkybY144+N0
zoNBFSJA6RExj0Hrw45dcXssWGcPA1dJxNoclBH4L8wSro2/Z0RGSc1iyW62EL6y
1qXHvVdwBAdCuQDUerphmUBN3EZmypfdAslAckeEQVwukcPzOWuocQUjUaoVwW9i
1I2vVN+WkT0X1JBwkXdWFJcwe+vjyXZg9E5soeIoLcOVeidu9hAcoyB3lbef4LVv
A+1hI4iJqSe1W+Alvw6WrUoBuKtvEzLWbDWTmbppKry9HRVHdELwJrFCFfyY4yD6
PQqsaN6MRlp9SA2SAiBjij+HFdwqyH1obvEgZQ6iTY4tdqTvkdfbZ6IRSUTRmuT9
QXqhTntAAYqbWXfp7OUKvYdrdMZ1LR5O7tFKDp65xAh0Y25aWUBA0uSDF/esHxm1
xYp33W7HllPSdLvpw/dD/sro00UG8ds/GsBqhoDTjtSzzMIpVO4jRYcLrCEU7Qp9
pMIOVA8CaqZHHCz0x/ie90XIT0c0agJxlWGOk+8RemK8jaTMTP9Gb+PojV50Wvdm
hjsvimBh3Qt8ImQl92RTNu/TEeLLGSUrvkXHPoM9Uw2TzHlevX+N05UJ0VBV4Jj6
jSHRxRMOisf52RnKJsD3WhoFBZrkeV9uQEeqC8p9J/BZ0Ix/wlTje3o+DuGcH2Y9
vbADNwRVEXJuVjXktn9Y3DjE4yaU/ObGa269d/5t7WGMvxpLGfaLnEhlWS3rm5+t
dNyTs/aj2e6zlIr8SYWb/z6Lj1UdEbWjzD3PJAL1bX4sn6ix2qW+xpJKuae/VqWV
4CdjD9NX48an8Uid7RlCwd0fP9RokbxZeXUiOra7Tvb7YjpORko8o6ebN5s72Do/
CGbjutpjbNwg/vyPqZ6hqcrxQLzCdyXO2k5us8zRaFKO61KV5JFLsg0Eyp9bCGWN
cpoI0sHGqCrnqduK7BJZVCiv+eIFIoP6f/WLxknjwjrnthiuMxjJ1HZB+b3zh6dq
OD75KH0kNajOjKnYg1enjQy/yFIBhZVGRlSvPWEbNnIc8z59LJBaoDVsemqtY0MY
3wgnJdCfrPUBvGAGXOFy1FcSeSeieV3sj65XD5d3CSv13jdEBlcfbFkIv+JR128e
VygTVj7w47zVKhsASJmKWkW9tvzYCrpE+wF1y5HdSqYkAp3270eqxVMgIEpRSZuf
3X4RHImEZdmhrX8AtNDJHP/xC14IwhYEaYcPeV8U/ldamlH8qaMQaisMGRHY2qTc
6auzKuEV9qsckftvoLRtM+CBolW2Z+dvLOVwBfGw1SQk+OTOVgacAmTXM6ZgkdGq
/ogMbrICvu9rd/w0jbQAUcLYvPK8/9KH1K+mAfrFXP8RVwU/M7U87r69sIfgeNLh
+URCYVVO8i8s91Gjm4WhKpgkrY7VwPXglH8SR9LhU5hqIBNKkyTsfQ3P804oFO40
6TZtLvNXxIze+VUdMQljQeYnWU74visyhjIVwgI9HmrPedwdBDY0vYDqJ8bOSdwJ
zRjl4PWCe08xKx+nFgxqLGQXTZ9DoDxdv7gGfjGdoSZ7Bai+wEEHPuZ3PxJNVy5D
HHYARU9Yc+Yy0WNn2spAZcYk6dfFKY+pAJxO9Y5cLnAmWykG785NVJdt6OgOWFtj
uJHIgJcCOCdNFvO+/EM/aL0vW2yM6yv0hN5sX5eW54VjruC35ij6t5jHWKIW7FiN
xv7clH0SBluN9fr/xHhc25L/ttQ4yRcPtm5cM7p7vZZ5+1o8HNoQoxHu0EJhz53R
DS2wbQzPOP8ZLVDv39RwYFNmz8GeKhq1aOomw1D2ZACS8DJ8c2NS5Js2GLUOUb8C
QOxxHqEFztw6pH7tVJnyTn8dJozXLczLC7hviys8gd6bkWjBU4b+tNpIl4Bf8C35
q04IdABZEEOBryoE06SEJ1OF+2BNMOlTdCMRiJnKJKjYq9OOBChnELUscfihiaA5
CexRWhxC0uXluc/P6AOzvT1i6m0yYkXGpZY6nBjmaQ0+uQxx0YQEnmBbIK9iYr1C
FLjgjAsFXe1wJLoFdgtJUcEte3RmTpaM93o+eV1Tis8ApslQ1EVGNHqsy6wzNwza
y2+M2XlcqxukzclqnUqbp4HpfJi08CcxGDbxIqwEDOVyki86oitVYPrtb1wkyVKe
ZIOJlgBQFrkcPBMSiEtMg/gtXA8zXTktkXIyQ+tuqz2o4Z4hzEBrOUs711W/cLwg
L5EGMzWxHRc7Fn9LzH5VlPLlZPYkQ3rgLVmCyAAahrfwM9mg/CbsBazO6RkmNmnu
fGVLwvUqyt0TRRkqXDO4v0CIMsiXf6qDmF33QcLmIpDLQmkv9e/Q/5bI4qkOQo/N
w4b81z0unU9bKTm8i0FqhfsMpAi8HfR4gC1Gz4i4oY0H1jLpPyJgIkEO+vGvgVM9
kitG1BPAuL4esxJo+j5NFE2/K5eCqtivU+jY4Sb2B351JWyvDB+JcDkAHTCwCWkO
OIn//FJljGpoEACNAwaTjZgBvDyqg21C+fH99LXSuCBfBd2iyPiylS+CgGJGyEPL
57JDyx05HpKRKRsL2UZmqRIWXrp3o1NQgzAVbzvoqDGwB2CCpDV3/FSR+lmrqa61
JlDlUT1pXcI9YcRPC4FmzYZjsvYjmNDK7h3Uzbx+s9mGeYnqwQLJX34ywNuF4BxF
3ddzRWmODRRptXGWSuiIKtBtYmSqlzEYqItsz9mlOUXisO5sloSWs2Y6d1kJ/PuZ
N6ufbfevGAQ7RIax7gI46N6Ci6Ohrj9BPx5Jps3RJa3IvBQlMO++8Z6E5q5ZuOxH
8G9LDfYviLOnJK9EzanpV2yXWL//34j8+bS0X8rFcCKLAM521eGlTOAHsAS7Lw/e
sZi2EAwqpCTR0wQOC3bOlU/6FrI/7Gh93VYT5Av61r3gqb0mWToBSrCFij46IRM8
mE5DJ3MnlOGHyZIUOGb98oHwXMGf0LL2CtvCajR6ART9DBYSri7EM4fsZ4Lf161l
Q2KjhDWwPUTJdAnMP+OMkrU9WWvfPSat2ffDoIk06FOIxrQMUvJ98i3JBB+Tkiw+
ZyTfkvq2O2G37BhV93PXlIk2YGT1D4HJNHsF2AFLy9ZW4qnT0NiKBGRkejACwTYn
zdZwEONQGYivFO+oHGTy8B1eln9Rsran7OCVBBlObWFlTtFlgSBX9rtzGlNbsAMx
miiStHsD1B0usLfQjRsDeNkSn/Kz0yj/CyHvfbTYcHijZawKwUTnNDmroNQZXijM
8zweD1if6w9gQbXlr9Szcawaytur5I5Frmg9mUhSzgeKYnwUSEVNi5k0lL/GtbEG
/msOah9Vchz5s/xppAhZpkwbhYDNl1Q3B0i9eChiIfi94q+wj8X4Bp1z5++cj6vB
V4Lq7WGq6w8+Jj4k+hoiT7BOCSC0IDZA1ZEMq/khXym5+NpxX+Gyde0k1/xMa/qZ
/o74CbAVMBCO7rXZeiK8InfWlth5YYnEU7LXhxRwb9cre20eIomrJg343Xd0WcfO
tyY5b9QYBEXgiC01Ms9OymUqnhdK/NllNBftbmEuicK/k3xXnMDqk0oD9jurE/gG
AhLZAHBX+veFUo78OHUMQgxOtGnp10HW9Ma3R8ULhBeRdL79/7kOFtQ7q87XoBsP
43qhXlBFdGyE569sMmI0xs5qMmJGHhnXLFq/sDFQimObZ7U8r+kaXhm70O4ngJL2
ypQpJ22LZkrwzuYc3hAdMDgZt7r6QeP14yiu4QuJ5J9/S7UG32xuw7fEEt12n33z
/0UolvcJKMeF/ZhfuZQXjOwxOlRKyadTUeRsQbCelwjrEQydECG1WOHlGH9OJVy2
RTAsZoeCWUVb2REANf6JqG+MlZNouTq1r/ljbUr0cBZYST73OKXoce9hs8Xl5vKK
qxhILmRJflQuygdgfypiaZQJkpK2ctGmZJeG34NSptXqZAkWlPVNt4iRCNuLhwXV
BdhvycodAJBCcz6g0cQwObfbKNttlSwJ47mGxilNjrdiDdoCsmvwso4hq7L+zNUt
E947WWqgxilU1DR61yGUjbupSc+80VqSciALhX0a3SxIMSyGTy33zWREdrPByhci
rHv3u1eqI8aoEKUjcidEI8GvQvG9aRyQhwGm2m5NdCwCFoT2f2XTlORUZslC0+FV
R3Sa+HNGbyVbW82eIAiEqUy+N/0qLDX1zPJuoHCTvqp/W+ESdmzEFZKBqxHDhkXq
RMznwfnqVrXTpppvXwgNvlFyz/U5+kGKAuJ6otAcA/VfsiKgTS73YPbfOc7WLxJM
3xMzqTCSd+sTzJYu79YvLx9D2DHw/P+AWcLL7oPaObPEKLzr8Xcj1KBE7pbXMuFk
XUcDO4jqwG1hJJvYNvaMJTa3a/+OShYhFgsKtvEF3yK1M1REB4pGVw9ea8dUkDE8
nHGlQA/IDx/dECflRAAcXU5bxdv66urniU5oH846U2QCZ6/WQC1gamYV6xm0yIPu
zjfJLJ1uWzvxXULS/i/ZMtVF++9OiECS4lH5N0TnSeOGiigE7VwFojyN7PjBTLcE
UHTkkxVRSLuwrlHdclxjL7hzWsYlusc6+h09FA9YwePD2bTjDQKE8UC3Ccpl6EtW
jCrPrIi8LW6D8g2NwAZm5IC575LXL3kBimTfY7+lqoeT82AYxM1wf0gYo3AdZ/Uh
z20tSHP7emi2Csy2eWcAO1CEG+DLUboDOdjXmmMEOkUUEryEW1my76yR8vFb3i2U
iOpUvqhQsF+89y1xxB2mQ+HQLzLqTATbe8avZ0jDLEtgR80pS3jFPOqi3X9yV1iB
UHM+qzXWIr0JgKAVLzj0IypmJe6I2l2OTNiz1prGw6IYHF1DY5SUM8osn/Y0vn1L
W0vaog2hpnALEMNJGqyJsV94bVHHDOV78DRdg1VaNlC+CmnwVwUzAODEYP87XWSq
nHYPq8l0NgeHb3VMHoGPugOGx5mOgrBcI6TvXGHEVGzxPsjyN5tIoePlvA4MUGpu
1b5i2xReBQvE84mHHlMNzsm6yapyt2XR/OXwAu9M4Nk/uofLngkbEkMJ8wBt8bdU
V6mMQn7SsO/KId3i1MSAcqbIhDXZAbBwqmO+/8yVoZ9Y1KVMeoEEgWEW0FT3X0Sf
iPMKccXpWsM8bzR/Gv+n4Bt9IpQuokYtdJLnLScRhPeAjZZBOs3fz68+2DdL/DDz
x2PNrSyKRAc02oUt1GUgKcsijzrpRCWmNZ3Ln4qAc2sNK2aZkum/+QeaUA3Faa/m
7vKs6PoXdajr7/4YQ59LABuYM1ylKxBsk+j49ghzeVDazfpU2jbPq0m/LsOCnVFv
IxwEumd+MveL2Z2KybB5aT7pKzxyR5Uo4tBsGr1mxnY6carrk/AytQ2ILIE0fM8c
LP5MHjHtvjUtvWkwg56Yu8vMFoD1WbUgaRk/ZCLYXFAL7nXdNwq0aBvPDbjjhJmX
vDo8sSATRnbQri1qXLCBpXtJpi1pV8OCZgETPJosuhksmWFXW830kcMkP1jcDhh3
863EB/rjJ2EwPuq5eapRwbJyVdL2oGauC3ng36paLTR6rXkff6gGM9GQafFysc2I
1r5DhJmIvZEJDcbeHkLLEbSKndw3q0tCQN/kvXqHdilskmiVfG1Tz14Iu80PYDFn
HHvhCnU0mahrALocOlvzSNm/7Xo2Yc0Lj6ljLdDPXisV6mbCjT3Esdxq4YtjY1FF
qhWq9xrl7W3xmfk22G2AGHdF3wi7lB3EyL9f3vhiU308HOBAbvEa4tjaqtY7wYQS
ZVVlQFWQcERMtgpBII/yWhVZAnwLBah8oS/S5dUKxNKUDqLabN3fbXA+X+PwNTGK
0VSI7iROfpMvAt7PPC7uSeU9Qyi4CcQwKW1kOEYoLC2Xg3q1vuiBOfPBelEwwcZ0
cO6hXsfxe+FGaqCKIVTTNCJOO4xpB88nOp9x7DIcGGFwMdS4Uii96G8nFAptO3Zt
nqcS+GhwyAIr/2YLRwH5GlCExCwhZmZEI4IsNalEz/OFZ9QAPJ5IrsxMIuvOLoJZ
OFR096u7/cpcovj54bTE+LI8jv7mZegHuqRexeFiShzEaFKeAhRj/VzwmfgTS9ZV
GZe+w43llXp9BUHcJGOO8Zgo5VqAiG908hux/mj8+GdEIABJkS8Dlw/CSR2BJW0l
1XpeII4varjRee1IDEPVbSNMrV6NHIdUzG0lh/ZLzqFoY6XAcgNYpmvQYMnGKRZE
VM5BRM0dn2VxtNbiDI/v2BSLHzfHhEPuqNW9juoKTbMzxTOizuOArkXmQR+J5eG8
lm1Yq2EzaZiqHF7JBpeF2QJ0SOXeaVPDhY4RGALMcBKsj3bmQio505BrvOq60+dg
Bb9+6s4FTGgq6p0yIaN9cAuzdrtBGbBLRq8VD4I0Szs/qePd8tkMOELLAK1nJY5R
GXyFhARma1cpg036gBztMho6FqTnBz9ovyZ0dh06YgnfwYfnytrNKXYlyDhEIVWS
qZTJ2Mzm8RDBAxJntE+Lh8EJ5HqkWOLm/37trvsUmHzvoF30dyE8JEohT4EOsyr+
bOiymclsfqUI+0HCdin56IF9J9x6APqz18DBrZUqZBF5lwIVQdw3VZFoJvWcsSLr
xfwxAMQoMOmPxOklp0aOf5MiRsuUM4YqECd9QKcZIl3jTNqstbl+FVI1Z5eI/crC
AdZ87iwOBUYrm7G4jLeWvq20oGL0Rh2jhIpJvbswR5hAaKodzNY8PuWayIRIgwZP
F7vdK23/f7lRdXkeeCzs9QXIqxD+H0UwXaSgWfwqDITyyqbt498OXmhqbNKJEOvn
z2A+Z/q5rArKYzt+0QiaHI3Iml85V+3oQtJKQoIgOgZQhLWIOgoLN0acw3yMqPby
pU5e0J7DqOjHVlUhoOkTrUcV6uM3Qv+CZyU82esUOzP1UlbnILVphAenTl3zNwOV
0dEemqlUxcd3ySWaaRU2SgyDch5YNZSTjUPLGjB/vpOYTzLAnP50OIWdgnSye2pa
aZIik3F9Go2TK0MBDSpdu7j9uwksOp6onIDo1N5nl3fZHUSNbGMw/9JmNb+r0YXn
ld7EjzNGmjDHVQHzL0fxns9liK9/q8ZfiXrUJiuV1e9K3xb+/wPsbChZSOA4WL28
1SoRk5C4ZZpUk4b4X+Y8vjTWFp5F5hlw0ggusatXRAO8xz1EU/DvB71LXKT/jswk
6XlQCcFLNwFtrV9MOerfVr4m+JzL6jVD9Ki9PCZ4ANynTWeHhLlvtuZcDr6zwEln
5onXa5nnOtJgG6pK7m0fX7nlVXwkgeseIkKUW7uGlhx0kOSr86mzvqgOZeTQQH6+
QwCxNgdmdhbF3Nmc/V9bJeJhRIvCv06YfI5ilvJ13BitFTN6PkIItkOiA9U2Papj
dvMfs3KjP6JHF3v6+OWtU+iLCo9OZQEx6I81qF3Qi5CIUkQnVlz0xOraDh6tOqA0
3sq8wX150RNyvSmNS/CJudDv0eohtWZlDhMl5xzWBfcUn1lO9SwzOaVxjqDEzMyJ
Yja2Pm6zP2mkYRM15ODTxW80EF8doQJhSSJzNqj6Jfu1dZfcecPOn3YQ2W6tUpYT
/K3dzRvBM/TPCtmJf1fKPq5pfz1878QPIcvigTiy0vCsYrVOnyzOgIOWAQu5xpeX
HOcfkjqFmqT1CjOlHez8Q/klieOIhqzu/Ndz0hp9/soaAQZtxRKVJfynkCk+M3vU
iE6CIqtjfAnSxuoJcQ5Oh+Hhvju55GYRHGKuz5LCr8yMZ5CoxRonUMiVhddHG7Z7
fWyPFlHEcRVNdAqzj3To1h/iChyQkhZPeXzUNz8q/Q2K7vNNMyDlfF4ROGViKKI6
dc6/7pEEl/fcsZAzEGi8kLzfrnxuua0qYeQmM2my13unY+yIvNF0lfIRMnHHeJsD
qdUEg3uPbCkN6mDtsfvhuNjiJ0o5L/N3VmLFiXO3algrsFyft+vzS0tSpEGOzAXa
y/SjD72L9OHxIYQfO0X9t0sBOjzM7shumIluOUpL+Texht/oN+nxuvVQC8un1nnx
jagGOVtZoVSGC88KPxcdlySdd+wvISZmmQpgv7eayvl2SkQLSQj9dKuGzNBSdCbp
1Wei5kMC0j7mKYIdh6TZNPQfnJVQyiA6ck6aA2l6QQcFY02KYiVkjA/MFayudQSb
ix5eysrluZH6O10RFHYtJmXhdALoFTxkx8x07JDpcw7fMaqPqxsAgQqGfaazT7GP
ewFpAPqiQbhe2lJa4q/EHXc4MfKOdHNTm7lpb7QhrBWYogArxDMvIuvNltreSvqf
tuQhe0jZtSqfkgVlw4xgsEHKCHW9T1fye8PouDjN+tgwnmvwhFGXWevbMc7yNnKQ
80+7jyBk0BhGM7no593fhL0/tkRva31O9DOVW7Ml6ylnQu8NwvB2zUpN3j3PBAXf
KvUI3vM6NQ7AsMJEPfsdw7PzzLlLe/ZQoi7bmrXGanGlXtcccesXxW/SN00e3BME
ll33cm7MHMUl9ywBUEoLXd9DRMDCmNw2v7vNDCYkM+IlhSbNeZbuQpA/lCEdjvls
MQ3edrLkS6KUotnKhp1LCAfHW4W7ypzgMDQjWmXyCOwpUXH+baVpOWjVwvI/EJ4j
GL1/lIU19DS27jgdNwPUq8w/nRjC0VGgOJRBnwHUrwkJc80GUR0QErjxz9s6zHcO
p3NkmULsXt+Efe4A1B0vC3HpDlhV1uDVH13h1My2ohs86YG4UPEZMI78LBmte9YQ
i//7e5Z2isn3Es7f4bIlacefQvdTdK1eLr304KT+AwDNzRI1zXg2II+pYC+D6B9g
8S91ZAWu8D6wfJJ632jIJPLuTZkm/mH1oprWGGkgCDnVF6cEKykCDNyugnEobITf
N5DIGr9rSulaPIPvDL+pzOoK/yefDiz1qs+12VQ8R4qR3/od1D9bhKcqRqoAIFlq
dVyu0Bh+eNtlx3HC3H9NKxHPH7XP0/YhAG7JcUJMHJUH9xiCWdS6wUIiGSyTZumP
zCIWGuQKySq4DPP/mbnq/pGcPB1QursizU1cPmY3x3J3dVJbz74aeLJrsf/WMit2
LESUbRqX+Fu/kurhX8EGKXXswezQQkNN3hsnvMq/PC1EV6pDrM45r+pDdNZ8Bmhw
qAyf7jMQQrBOX9b5LT47/a3GeRdBGRqmfLKQzxhBVNFPm/fizgteV8kkzC1Bk8ob
m/pPtiQSOkoX9XKAKtT8WgC9AQ5VRuaLWY0SWVqIlseZgfcXs0xtfzhWtZtm/i4g
stI9Ep+/7Z+Pu67hj0bgqQT1w3jdS8pb027A3QIPYY0UVr3GV1YiP2TNmxd0dG0w
gKurQh9IfSs6NjRJLF0G7ZC/dsIRMBB0jxThtY+o19xrgH9jqaKe3RnpNVYEliwR
N2vGYNb0Bb415w3BcRj/xXTgcNf7nuaXWttJxlMRSmLhh16mA3plwEX1CDfY8Li0
FDU8rgAZoLpUZociScjRTFAnsvHGgxDP55tAib7qLNqaVPbYGzfQkUEuN2M/ZDFo
vXmOEvLSf67Z6GH2Z//PKz9BA1uYaNEaydPF9MEapGJKe4JSkEkqGzK1WftPNub0
EytMiKU6NudI7AWypOWX30NkH+anNnTvQsnjCMSjg1EjkYQ/u9eVkr+pqxfgFoCO
9ZJmrxFuMacIZdK5TKYZZWYCwdK138CtAm9qELqD5kCX/zX2xPQXyKr/Bu8yOFat
R4v3DyXUWGg1dUUA3ZAy1sxlUwt2HEIA4w389MZQdSOPQm10gf2H9ZIDnCrnOy+z
tRi+Zi2OsrlA1blT9l1pAbiGjwp13Nvd1NepiOoNOKgWHcz+/+WwuvZtnA0XPIad
SnKhyfBse+/cO8h+tJcvoNWjBevjsAmEREkctRXVfF1hyJdR+ZG3zdoaqx+Uu7XG
haiBA7yg8ixQ1kGrMYc9ehxD8kqScrwKFq8945p+q/sgcAJfhMiIxtLtpcqsHNNz
ZyxeylOekgqlwttMHUasuzsZYJnoUGV2MIlDUjFHyoczBiZd8+pqyCbZ8/kRVswc
q+OvTHb1Bb0epoHjXxlLKGzT4JRQtvb5XDhfhAwDDeMyKB/Oc4zx8qtc7o11d5BS
9HA/HHzzH3fJyxDls4bEANmJ+VBrcQ2kOqwfxUq6NsE8M0btswyVV0i3t5zJNSfd
i2ZFFVoFHD1NS/8k0Omb+NBrHx8g8OMcb8VNG8R575QA/e9MstOQB8CiewFa5xI1
pnJZbBCVhA2ZfJUs88Wm0D6AN9qpW856UM9/bmCAfKZUtZ2QzS4yBNU77o8JvYpx
dTpHj4PMTu5BV9etqArfKXevKt4TgCJc63UB8WpPUCEel2YfIaCgQczHRXgwNLNT
5OJGW6uWGCSbWCwdkbDDDGPPNiMGIAINHbzfPnXw2MliEbezPnZPXZeq1THQS130
0W7/UbrB3XUQqK7PB0rnHIHMtzzbhrnABdSmE6Hcuohkj3sLUuoXlaX889tVUPlb
ZdU29Cl05Xl/Vt2wQtIQpKLR7R6+KmLj4hI2Ke0HZ8TEKTWJVahFoylXtmTxgnL4
CRHC/daEqXtI9lBXsVVtJEgIs13TyyYN4EDFdY7MwttmIexJ80TyAR7FWOz7tAqM
wjvTNZalaF/QAo2E9MAGMhDnJktTWd0iQmiHKVgh4aL6UUqxzhi+rCMRf+FA+6zD
IUYs09sQE+NSVxDxaNuT4859wmRbypXm0a13e6TH8cUX4daV7ZTS7X1YE1PIDHTK
CgWhq7guOc86SRTPixPvVOVD0Nwbxsxho3W0aWbdihlWzRapji5Ozth2AzBZfuvS
UTok8uvUTcbVnxN1IRucWiBB8giBuvLmFJaCg6/dc/JRENjSphAR9Pwz2sSys3iy
W+Qp2miiorBV9Yxvt7bYQeLHm0Zur4r7qHeDDXneiQCBB2MyiuCgJiZaNTxC8oGS
bVNK1qt3Xp9lZVdLJtkTHt79qwivMWPCUtFqlGhGdqlSBDZ/V9VKBYXiNnAKEWD+
4kzb9RXZub99YeBjfJF7UT3LNBhq//DnIxBeU+OFsA6GtD1J+WHmKiRijcEBr+Co
MfWLWS8Nrp0m3vQ9tmukgONDBT4scR7azGD7No1JGMHmXrGxhytU84i20JhOsNbi
oeOSk0NT3dO884MY/6lv2abDQx30/PrJ4cMYKlx9tl9k/wPiK1d7PJQ/anjY2o8P
LGfObtv68OyYTBWYZCwuprxXlka4UkYj5mlHji0EyPlUvZOdUSrM6iNySiQcl+pZ
/fiOhMicvhE5O7cKF1D7DkN+gABwY0swniSBhkq4i73fmqlgf7T2gzM3xsOJi8zk
PUteeTtZbg5ZgAI/3X+rTUPu+J2dlQwgYx+xVZ1VXAJ14ByJ3PcPU9Po10481L4T
8+mF4Zpuzhp61pNg4Evic1iD+UbgIosptjzSYoWqg3LsFTwdMnZs56bKZpHVHpAI
v+cRyFbd87iP7fGVMP/VHRiEhojn0zBlBMFQR2PxWYTd0Am7uWYQRLYCmgJA0dA3
Swz5FDZZwmDsY+2Co75kdYaUGrpKKRdOME+W7RIeakyNj1PxNzs5XcV1cSN7sJXs
u/hAsrolusobOu6D1XFSaWHO+Enbg0PAXHkmJLHRTHk8zZ2lbmeO/nU9aF0kIFxv
pwApXJHDTvrvIFCrr/OMcKLkf1EWBi9xeGODN8u6g7UOWsa2C3N+uPEAzzr7E3BB
uBIKXqG/PWD3msEb5/gM6UJHpnCYTuovBXDDxa/CtHDFD3+QJMxvV9H7Ce3z+PHs
5qAx9fQfpR2UjLaKgE4cEebLJfXC5WWVq8qMa380z6ZinS33uXJ80p1ZgUUC2sFa
SjotlQQJuIvKpVwBlmURqV+XNTuIcdJskZJhU3HsnFfW4CHGEnDq06qjQQUMzx7Q
4Qt/bCxq423KcqP1BlUO4B+wU9LiogqL0AjY2FhN4TXOgxGSly/2awPgJkxjOdOW
4rZ5P5U5yjNU5RsM58hf9to5NdLtWdFEwEhKAEz6WnwNIb2oPHgsbFrQ5qXDkNzS
kkpJ9OGqpWGRZwevqs1TcqPwYWBdkgrBKsJcQeL9IjG2WmKB5vbIlM5Wz2R1V6jZ
f4ZRQjkkdnK4Vx6x7WL7u3pC9t/y097UQhfXI5EO3mP+T1YHxhOfxeC+tYg3uYz/
YpJnraZsa6muDHS1gxVhOg0MpEHKMHm4WkBwSrMHOHKH1DQWf9r79Pxe8y2tjgos
yfpA6gdiDd/mcB+80orj65kd00t75iMj/BnwMd/t0lEbEHM5UcY32Ozbfk6PFrug
cpj7837M5CY5GIGvBoNSU/UuxUoXaWOp6V4wew8YftFVJkqdauKHLEHN/y+zdsLI
8hH/HiNZELS7mSniuRs+CrJ4BWE0VMSF4SGwW8SNoN+zOwr6Thskh2DxeeMEFNXB
mkMmwEUNRjmZtOo32IF1/+0ugJme271MFv6yoA5W47vxl4Xyaod+zZe9Bv7ARhRI
BqzaqgSu2SnZwkrD/C7nbxfJV5csBCwmzMb6To3UvjItVwHtK3L7FNPuCf1E8sgA
K1JKFkqzsfIbkvYI8EZzJo40kehUS3EBn1t/a/TnddBV+3HwpNBAJU+r7p1CROWl
CZv7SeuwS8n8/ThricJh/rLfqzBxUVcuixkdv4v0cTSkHw33lfjPKGY+96PZ+W/V
NDgZ6SVaMZe33uealeTm8ZdIuZHiudYok6aR+qyCzcjQ2dAJMtGx2+Ge2NTQs/QT
1TGZzjiWY8mKYxoEkmAbA092eqjstUmLSt4b+06pnk0vhwkJu4luagRywvwuJ4gf
wOyDtUUCcSWbP9xLpKVGeXoL7zH6ToZmwOIbx6UF2Qf6LuzZ+FRqgOijd8vIc6KN
8e/DECbdfW2bLVKZhwL16G15DqBTADEzvuVqXqOGirvkp+lxCxhLbzeHxZjpcRMO
P6mzoTPI/hTwFmsWd9xZCy0MNRzW5+aRuiySojvJH7rTvBUzzjdFQUNRZgOlZkKy
yw72sW3GTg52chjLtcQsbijn6gkugt4YBapr0NlR4hQwSdNsQqp4zb1uRpw0ax63
noBvslTD4dB146jSFrscO9C5EfbFc14y0ApG2vaWBlGomOiDvD9jW0dJ33mcQnV5
ZeysTLnd1Aquv243zPjdPgScE1yVhCak4piB9MYs8XhnRjt9E+pUxJXr15wXSGic
SFxDh6+xIzrQZeyZtMvQFaH2JCEmIMZT3rlhMXdwk+zePB1qFVINpeLmJVCD3OjM
2Sr3XLy9uyyX9sx2Uwg9XC64If9DCJGmYriHqqrMGtoh11xBEqtD4PjOd6dKIYDl
sQX8UEVa4K0gC5I2pyBw0N0jnij2Uey9xaDUDWbR/LCx6ol3t/glt3TvPks8HJLR
H9sALpRNDHHKmMYcdLoTfEVzQwuqUAp0YSwieLgx0yYp92ZOc1HzL2oi5ciyvQru
vxNZqhqY4TwghhGDx59akjo2bEqZsA2oGgEzLwWe/GluiFGEt/SnTDIvda7I+H39
p/nusuP254mqtLyaue/2E0tqY4BwSOqjdVqu44dAzo9CI0UM4qo4Io1cpqlv6/g1
GEpbVfLbNqjYw+w3Br2otHQEV6q5spbsjB85l8xLs5ISND/dC6G5B+0Q1rNEWuT5
UutoDGXd7NBzEL/+S/qD2eUqc21xltK1hyrtTsrGKXTSalRsZwPnYXDn4ERXQwT8
7BYIpNdgF1jBJQQOHWLxQSiyJqjQz2op3BUddoBBOWZwJuvQ9LsrpfVJc2s0+YsQ
7LEPum06qJWZHvASO2lm9pY6IYFewDkCHfTDHUrKoAn323zeAu98cxo+5SEyY//Z
pFBPPDPLaTjoeBMB/LPgkbJg+aQZgUV7BRG6Ou1WK4hCSJBF7EoZjzCLbaEgp8tO
HNhzjAmOaY6j+w8n1CNCqcZ1No45/BQHXJYIwBCpYtHO5efJ4pETg8xIPNOclg82
axCzZgRdiY3ntNVNiNFEslmtnsuZpCpMePhfSj6muR1o8SPlrpOPBXRYs+Z+abEU
uBs+/dmmsVt1YtMYcWiYOBPAqIJZScfIp/wvxJdNyaZELoqAU9rG1L5Ds39l6UeF
LS8V5LFh0J1iS/j6yKTjYT28k3zV9PxtlZl4vWSGCHJtWJtQV4rTUJxIx6LHG0st
1oEoKMldIahwsMpjNtUllYgn8Q6d42Don4wifNaM1qzNlyYZBdZu0rJW2KFvTvQZ
1nAyfyGmSuQPsndD58fjFrX7SS4jZV4N7+A6cMHvyF9O+ivij+9H+O+eBAO2n3R1
skehYqdx938y7zibq8MfI14fozKonZtfMLWhWmgPUrcj9wQuTGUsq5wpVLs0tPky
jBGgGioRebBvvZBl7K3I8Rp0F0rOrgZclzf62KCeyycIfXin9jJfvjxoepig1nkG
7e5Cm3ScOp6jCE5bT9WdzUX3C7MVzAkFB922sArEFS0aozskvLRwv0pXQvti9C7y
DjW1nhxoyKjqhe4W+rcM0q/160ME10Y0gMKDboqG8sOoXBkWxjA2rWhT30/ybiWG
bw6G8s5BfnPacw9qKzQUmOxoO1zEpkCS4y6sErDNkcpC8JvAckEpOW15i6JSzXfK
Klem0D9roaQhxiU89+PEjJ+ZwDWQMa17vFIa9xUevtxaR4KlbCR36Joywo633DYf
ozypvLTkSjo75Tiait9Xq+l3k9rk8gbOQ5K4o14vM8LzivBtjO9YOV9GbKnH5naK
SaeQEtpdMpLO1QQ5Ct/8NM9hq8O7cwzumJRs5/4QC7Y/qJY0beOfsGl4JSBiZOnu
QvOWvRfELSxfd5LXeEvmtdLpTRGlwt7b8TZ9TD2ezfX5Gmmw6Hu6+j+a+Vwz9/r4
5m4GezfRDV3mztDYY5zNv0awrp6GgRhh47z1+jXw0NyHabXQpeNhSo9R00oTqlyx
vsF79Un2+jgS/bLPx2j6cHcB7QO8YaXQDzMvjI3/jTaaJ8h2qLTS8+6WghyRLqUt
w6akFZX+8Iqq48EW1mCpipxButw/3VXV/t2tTKFAnW1nt9m0ZV2w4euZHQHb7Po5
2WRc0gDCwfI797CvckFRgsoCifdNZZpQFmAJzV4o4AbeYnoS1e0XjlxEg3kiOiP4
uYo2L8fPeLmJ71qH0ubKzp1OBKsK9MS8x8OSFPgAd8W+yMwrRWLktIl7tKD8nn4h
5xlSIISnk3SpaPptK97+mOcHIgzims+AmITbC69FBDtVgehMD1+wUVw8k8D4teGW
tJ9q6XxkQ0Cp4q9bP4wGIWBbReq12Nl1b/6BL2gS/gkJg4koIjN3tb75BrQjbIzU
SsFo6Rer8iub0sH7j+FwdVeMFtW+INzktyTvyw47Ght6sjfIwsUwwcLO/aBxzUzS
pxn+yt92QoKjxsnp4s7Rl52bBQI+4GCPGzE+xM1MoRzrOklHEiKfj4NCKRahzCaY
XhfflNBEyeotcN6EhJROmOpWFONKeIQQbXMwxlwdyS4/+S/POnAyynO5vW7ezQe8
BxQ1f0coYpvOa7K9HYw74K2fy+Jvlmtqs4xV1B9dcsqDGN+is+7lNlfUTw6I3nVq
8Q5jzYb1K8uEMxD8BJ9GsiDEo7iJbAD7kIQ/cIv9nQDdEQQfbVuTODRIJuHnohp0
WslRSewXHj3CCIBOjRgQ1ph8doMxGmvDIdSqqpVP+gBtP4zd9V2IXU0Pg9aaIDpc
6sTer0uYph5X0luVwgu/WhzAFXXqatKwtOxSH8bRjDdqRxW5Zq8+4JOgPZSPw1Wt
SRzV3wVghOPKnHCObQGl64uppYRoHx5mEdMYS9di8iHVzvneET5KidII24a0qeem
EhstuEUhPp6mHzbJiB38KpmzeiwtzfXt1DZc4IT7WwPQ3J2TdlXW+AdDzg008Eqi
6K7uvyPq+3pbPeCG6jSDyjnoL29JB5seN7a9+fWqPR6WA+XDQliRLDkwGwqGHp+5
lKVd2kfoqhwckz6b/wfFWMYOHt1zFjW9VsGT4L5ez2zjEPpm+KcXi3yxm2tbbw2U
jn1upy1fXVAZ+9oD0wbfoJpX7oaSrnRglxQqEYq9UtQ4N3vVZPis22qWArnXOjvc
KVS4KyBVPNvVSG7et5rlx1aEqlIeozgJoIUWN8raU/+EAO3KmnSx01csZkccvWwv
GNUcvXDaunGiZHC0P5S30I3xoZHqkA/yJjcawiMG8VzdUB8BMkZ+dy3g43qtjy9q
TY5P5PR/PqIczY7JOQCIbOBtPhA+9p6FJP0EWqdASc3V3TQrLKT1x6OA1+hb+jON
KbFfaCtPkRVsN/5IVem1rdSV85c46Ko7ASyfRzQ1rp9GsdOpv5QNUF2QNk5cbKND
v6080vupQO7MOnBLSVuubijluKLJ4w0gfHI9KSI2FIGuGDMexvCcQxU0ebW9Euer
YW6OhiTQOAZ//ipjPNKqtvUqP6i3cU4W1QnotomZcFKUeuiA2Dm7bosB/42Gb/KB
EhnyTaF/nOMrm+HH2mQL7yD1RApc/MmJx5yuKO7TBvbsVcXpcmMEbcatoBTGVc+K
zeRg7kxqJIv2TkNDUYt5AFSRzPnepeeSIu/a1ye9LvLzpjmlRXqJgnDVZzK3JWmv
EwzJrKLSptlBxlpeKwlalWrm6GmtHH4lHhqPuJXasNi6SKOj7S3G/fOPtINTd5al
Y2fS7cWL0IbJhqLGhGIJ0LXRKuGTYn6+Gc+VsnGUEPo8GvX9m33ZhoE1e0t6ZDaY
9kvj7i0cbv+oh1GGfD4BM88RtINc129rqamQreHc0knrGRFvZ1bmo3DMFjwIisWv
gHNxzGX7QY4Ke/l7R7wpEXChX8x3g/uYozVOWjACImREbNVW3BXi0zsEK9vfugGn
y2Q8OgtZwz2S1SiQFaBv2eEMG3lEFKYoEWPGNCyyK6iv0iBqlWxZ9Pc1SNuWYFA+
R3oZYgjpgwX/an1WG/1ZUNQJIZknTP6NSOyyEeEYgof3Sy3uC4ijdY0QLhiD3rhr
myVKQdzoufY7KEfw0obBL6YUlYTFcExOSZKt80+hrcADCufBc27hFwvxINdPBGhC
SwibW5iEYjZVaEVqtyENa6NiarM9vr8qwX/4ccGok7WP4YUCSnWLvvvDU8P7yJs5
TWu7VWiAlnxKR+m3O64qHvkzWO3z+bGQQIYg3kJ4gl1fIAQFazK7fwUg1rFokOBD
XFb9uSg1ee+Libld9b50bpYjnvTBX9M36VaRS2bxK2JtFE2BeVXvNFtJjc8x5+Is
r6fOyWZ07PI0d6SQP4uzm/kFED+BNhx3Oj4p4ZKx6zmuaC1wmxFsI0jOWT4mNM1r
dj1GOMN6W6FXjoZkJWoK/zvVpg8P025AdLvi5mqC7MZL2A65+g9J5korquskD/qp
DNcuFCLSM8fNTIjpXMSG3/MW9QHyTYFQ9qpq1BEn873EAk5FiK4Ygp/7cmVYQujJ
Tw4mOZkT8WfqJ/CSMRtkUvtAZhQ2caMYgkkezJ7kW8cayJY2DlghiKZvm00mqaGE
Aj+FRlWp+mWg6/nIIJf6X9OTG/193q7wYVj6dFqOGvjBekgKy3S4SSJo9l0scFCq
fdu5iOMmN5dP3MyIfDE3mrc1VGSEg3zDhZxDgFv9X8R+RwW9LMoTeAVB3eZd4gbt
rAVmZg7TN+1TAxEb3Tltv2ilMFNmAiX6/c+Tz2YbaH/eTIgkS5OaWBv9L3aOIqR5
dChYXQEk+P/1R5vfkHpUyJX7+5akHyWS68tPQ9pW/rIHYiaA5NcLl46KheDeZ6Y2
3ghxZyakrZcZNkkP5gikhlhkg1k+n1gJZlolEHz9Dueyf7b12vubgd7dZ7P5zaiV
ANx1JUmay7jm9hqxiT6oQ0aIl+Wp6PLYVtGeqa3uycTLfRF9XCLAROXj+F+4Y1VL
eZgMCFfy5vZBY9YoVcHsTm8NfknYtR0UAlGRi4AMf0mKhxx/MbNszmubf6+Z5Ddc
qMWtyYBrH2ja3U8CQWOztBADNqToESySD5TBVYsrehUbDpLpiV4P+a0z6s6E8cgN
pBhhhF1drpeUx8oyiF1MIq+yQhyugX0P/VMLjYB2AzilqB2ZMKg1Zm9MdLFuwTiB
UmbmO2RZ2OFtV8qgZ/5bijCsmjqDqI70rZvoPPHCKVotNinYLS01HJJGNYMyqH7N
RvCWjzp67CzwNoEIXfqSvuOvLhvs9W0A3Q/khBcBEnJ8X4pfcoPTDmcXq2hoJcri
DFU844UQHNW10nZvbCBxAQoU4CelzoEpk2F3dHotGv0bdLrsj8bMN4lq6mORZgtP
sH/1CCgvsSf1dM/WNYxocdSGVfjRjHVAfTV7j3n0nQePYfUyrVGyjqbfv7w1/FY+
4gwsJxGlJK3dvOhbgwaJMQ2l1laIEjj5zvQ4kzkOpbhM3c7j10nwQ0xlsousLehK
Rf329qs5cYX4NmGgoJN1+ht0icCCsIn4uIDn37uuvCQGlT03sKpxJoHMHK4Ya1iP
Fw9IyLKqZHm3YdgecCa8f+e+kxFHoqkJsy7N94o9G8qldk7D4JH6IfieLdr6uPP4
MyNguNlgX92JuQbDjuOAb7WU0LKIGRTMRYlo2J2Os+LObWE8f2aaRY64KazOTTtx
8V6qQUaev01TMHRfYJurk6xxZ5v4BPh60/5qpP8SpjYsXo7vLI2lQW73nXCIwUDd
/XzSuIOkrExbOOhn7QpfR87BNREXTEI78iR7Zwbxe9WUXVg0ZbQu+K7/Ya1udZS1
qAQMcq2uRMRnAdYX6vNtCzUv8UT7CcPX6fq5CCaVaifNcR4x4XVhQk0jvyaU3ZQ7
RUB5JXir9JcqRrcxTeJhPv2Stvo2HLqXcgm1MYMKNpHPmKS/xs2VSYYZA3MMCgaD
oe/Wuv80OpwmwX29zHmeYT4Y6Opr9qqvJuuq2XB+4XcQ8dg0qQYZp9Ztkc5jCeZX
YvkkHpxkMWk5qOa/TtQWPGzFb1hjjJLeEB/kQoXtvr1E/BtvM6zjcr8h76T2P1go
LIlyMf8g669FaHRo4kr7cmjIJwul4vwcTvFN78ZTKnOx/419MRIIAyOWmgqxbQtq
1NM/z074bNA1NRnWx0QO2iCP5f202exabE8pDml+/aIxaghjQxt+UDnFLfz035W4
pvfPJ6tb4eSUK4w/tvjnl8Eb1zBNCuszh5DGtA/0DEmWBxEsu6lVEYTCooRm1sX5
5AiZigWqFaEgyfTLXYUFvWIcJCs1M8YOVgblICqocB8VgRJSHbWmrwtaRyzOdm54
g1F7X4hz5AI1OY38bp2siFRrLid8t4UAyFagI398CwbCZJa9KRUSFY0XgicNAkFj
A54ee5ayE1pRgz8a7CDN5vZm4SOZ67eeUSkivdLJKrEBqEqLs3UsVzm0P8ODrqQo
l9Xive4qfxae1/And++XuyihgiND4oxL5eeMfykF33PsaWBzFG7BiMta+nmiGBUL
WH6ZoXu4hiRIxWBP7DfDnp2MBacMebNqzhPeBl1RhxXoWE+CHxLEdevK+WItu6VD
ZnCIXuwqYKOuXCdwaHj2N1hWsoj01fOrAVb3BO8LyWJxoW/RfgtZS16DyYlyidMu
oiE+/Vv+V0ularkqkI3QEY6i9JpyVN+GjKzTBP2N117rWic32uEsllZvMOBlAw2B
mieFkCUg+N6LvipXrau317MI1d1G0ynoWOncHYVfmemCgG5YkrBqU47JqP+IYkww
JidZUybKJvoTwJMwEOWJbFY5mqvWQtjOd8OhV1gDnczSyd1F877yNJjwfGBxCbZw
2pc318U7kww2nmAgCd8nHrmTXIG04De9MKCxtJ4XgRfTrmHDFR0TfNaVcbjaEamM
DKLVCbVn3jg7ZMKRKHSzuLqFToUgvqlH4t++njfCMb7hdlOBK2gWCT0yZolskal6
YjM2CBWcc8IOfnVmTqcbtuqV5N0mTZZR/NU5W3NiYCMJzObFt5wnlBQhVZKPdLgJ
Po2YTKNsnTm3L9r/CobNPxskf82+kKY8fF1+IXmnx3XbHoEhy0MgIT/TzkTD1JUr
3Qy4LJoGfcoe/3csoaOMPGJcJy0dQ1+0xqiSkuAKGvSgPX4kP0Hv7ooAv5emkAjd
/Lt+lSOLV7wKOExBFDkZKIEvpC2K9JRnNI+VtuYfhprdjmMP12h1LhQnJluMjUwz
7IpuNLAn6+mLP8skb+9Oo+UTVemR03VZ3eU1GWIjfs88YPoCN++QpJbs1qpbBKwd
P2DIRCrdNebW3ZosVSTBmNhMNRQdS9Dihmzb/4igNWrywlTmZs0klseIK632oEhk
OSRS8t8szVAZBiOentDkruRzm1zwEcNZFDD/7hoqgMzGI5bAvIRL4bNQ6YXsW3qZ
fqnlfcwTdba0DqZCGpZleFWukMj83orXlFBi+yZVbG2r2r9tXQWv3qPK/+BZ/sBR
gmJ2VdnEugiSKP9caAPtR29Ak4/Wq098llV6aL9AGpiOegzN7j8bpxKZwaI0zR3O
wY4aEsZmwqVbpE7SJWHbS8RLNFZqrI0ijnP4lb+YclAamL44Kn+JFU8IdZpCLXiG
vSG/L07uiEvCV+ncrjVqWysQNuw8RQs6Y7zl9ezXHrx3wI1vNWvlU1dA/uQIapin
o++DUeMdXQ+TIpWb/YH8eLzDcNzYTnKorSKJDRLC0B30PWqoz8dP+P+UoFjUE7zb
/jYQkav0fMUoRFpvZdTW+PxWasz9Tazg/KnaECsmIYna6FATodMWvARJgG8TUoXP
cARltksNriZ4v7WBRC+MN5pmc7+P17s8dufNAg93wBMfllkhgp+L+NSgDPVCltNh
cIqwvNnngVUOSr6ydknboC/nVaRPp6c9PFRmZkZtF10aNgHluum3gXlH+JCtWGQd
zmjKoQvaib0km237+mCm7ur7t584LrWzD6/YIdZaMYzgzwAhaSex6WRtYWR2QKVo
gba7qPfH+0iBHU8oAnSR+oy+2RQQWdYebNEyiB7GmB0biRBTEiq6rbn7YXqUUg2P
YHhl2mWELIxjb3hkX4BbBp8zwccUh4ysfXyeFRQZO95Ofq4164g/Y54xzs126BEt
B05WqboH2DthNHgZ/uFimCnFZY8dvw3Khvjwwh5KOty7Wr0xy9Oplwm9KvkUghnA
spqmqfJ41qR/7jP/2QSg7FtfOBBrPwzP3RGndM3TD1lvexwcF7TEmhZ64CgFosVU
AEW2bXxEXi6Qbnr0AB6ft0VflCyvJeTEAIclTixCOimQm3vGZnZQdTrScMlcKKUI
G4HzLy/1fDDubEAmp3TVYnis3LAzJvDwftDnSjYWuR/vr2jZIBhG/xSf4PwblyZ6
Y5SRjd1Z9DUiMruelPSYfoaIlbjdeUbAnq9CV97jKqoKOEKrNRqiol+Ib1fXjba4
PEgkoe9nEJQ5jR2fTkUoL5c2w1kXxvLNARkSyY3Bwjfj8LDb5GKeM5jlqTZTVB+5
edL2KdLAHOcQi0R6beZdE6kZLLY3KkbYll4RjfkaxFrZgwitdM1kh1is827GhKQ9
gsXx/sDEmuePZrzeC7rPcCJxCaI5TkKWQrKmrEQcMlCrEIVhgx4+mJMRapvy8q2M
ozIQ1h8JSzIw9lKJ2QBX68pdgNeIN6WkG4ULcIZY8WJWBvxBe+zGRgVbLsMUolqa
d5osNkk8moV8D0xmY3pZYpELgOZQuZ8JarezhiwvEocOqmVttNTn+wN9Az3+FKUD
c7YdhCamFjsY3iF/YXg78k4ekHNdCH0E0HavGkBimneJaG96hdKkcyap2pAR3QoI
qch/HGyh4KPcB79Csy5nDYPF0szT3TT20jqLuHZQutLUMB73QsJ0tqNatvmVyCEK
6KwnIXfVsFGkXLaoirx+3UJQn3uddaIWmFs61+yzle2jkrxDCVu5ppz8WqsX2KXJ
GaAT2zMnHHdMx8GwlZkNSrh/MDAVxCHsm4A61CTwRK7kaq7iGdTTt+sFENbq13wG
tHX0oqcYwPeB2ewUpSiP8HK190mfeVgbO+jtX5vxDbyW9IGfjncb4ODbXL5IwQlG
Q6DKDfeBXbE8s3bqQUqWD51yELV23mbkDgnSvjXQd5gaMSUHxqV7p+BD3r9rz3pW
6yzjKXTb+Lb+ITW8WmAeYrQiJlrvRJr1vU9wQ+vRH0T8I4gRIw1bbp9wnfVVdiem
nYGf1o8HwKjprT9Vl2E6qkoRwUAaTG6l5N1rxtaSA4qX3JECiaJe5m5SAa4qunpb
edl+DkgDpPo1gg1m3gFLiObTIGMhpExbUfEvDqF+V+DC4WQneyGMVyMmk3u72ohz
W9qujiciX+PklDEHV15xAqW6grOyUXdR80YTJcWEoGhPnX5zuT3lQhQ+60w/ZlFR
ZGxkrwSkUZVsJeC0PJXSIpmKjJnvSvyctCRgPyHtsw5mcjKTuzHs7nPHf3zlfFrC
9DtJwl+PiupminHZTdxeCLimVS/20eIOK+m9GveMyZQTnUcxbCmknPVO3fHjJgtV
K5cV3c76tDKKptgAhU8Xxj76swCJt5UUH+eyes5dNKvgUrMQdp6iUZ/jO293wRU0
bSSlPqHyKq0ToIl+FzHGZW2F+BXoS1p9tk9UJ/OIpjMjzLBFGlE0TuTJrDgo4nH5
jbXI3Ix8Df5dSGf7FMnKk5Nx58ebI2TFqsfGDsUzIilOaKiaD6K8fEgITHnnC8/6
K8XSlLjaPncf9gL/ZWv/n22CLu4r4aHwkAYffMGeTyiCnWCfCF8BkjKV4wxGmYPr
Fp6O8IHSIIXPVujV4MUWfujK1zLdFLYQb+JR4ubbZoXy+wiaJyX23YsxWvFkDKym
qPRF+SuuzntU2tMbDoKco3JLkemfZdb0cfoOL+YSFcdjR6u/sKj069Hgik8OOjUz
ge+6ukLMuFxr6NlEKCCusswknKBh1djcXa6A6AXItiflTnjSRQN+XXAe12GKffue
c7AQ2fiJGLkQt2esUccWPDxX0zbVKdGAMY8xlQ0+IKbID2otzfnjtbWGYih1JmK6
1wX7KR9TwgttOa9I5NoAJxwdtXH8OyIBbJZ74yHI+wwyEgJtWA5HxxPb1cvfXxX+
liyTRgg0LH5p3tX9YdCVkd4DiIhH9COo9qXDc2MbmZql6OWDMpGjzwth5x38HoeE
rOo4blFPkwid8+xrjOAeJ71hKNxC7QUFAo/scgBYIzfp/UrE5JpfYpATVD+59ZPF
bu/rEVQ8JuUJqf7UUBAVzpvtPDP1bHm3XEpFfdRa1i07nwpXUJJo5gtzhCrOTzZL
RdjZBp98CMDs1qf5euoyh4PQN9eNafwgdYSE1ADX8ZJ34XTt2Fcqc9JlJ8FNnHc0
p8/g12DvUtcg6zAy7K3WUEqOFpRbRay47CrnkekWzf1RHFTuOHxDAj8eHnnVVNGZ
Podsx4W3fjown+4PoLKyrNa42SQ9G04lXXYPhA3UlJfyAPKxD3PJMHU9jTlaaI7H
j7MfSJGdifj9xdLjNQBKl5JjLPxGYSi+tUtAlIgvkk/jM0/z0bQtzqtu81iNig4R
HRgSOM6SznZMn5W0ZnG+7+L4kqVWkCbAUvHHkOBK+wQFQ7gzY+9wHRF88zxfVIdk
GklQG4IP6oHsk5E1VkyQ+S9jQ4ZWntQqid+ywrkGOCY4Deo/40RSI6l20Zxg7K+X
3yigqjDoNlgbixw1VUVmFI/q9+1hOKzGiyD0KMZyWSU++6/RfH6xx4iIhJltf7cQ
dsEp6rEgA1KMUwLeNaPii6jAw/qdEuXGdjvbq8uhbPH+4VlCToJEoI24IFVWRlch
bp+TxCii8DSliCAL9lCrmiW57tcS3qPKQ285Dw/cJYDZLz586RouP7COVA07DMEL
yvHRe7miGJZcKmfA6xfoGMUblFST2vYrkg0qmmqdaB1w+DO632bD5DNMHX9TXY0H
BYODWr2zL3Bt1HelNkcZ0m8ZHHdMEqMN9QGjSmNt/LPYlxCoYUPUSnphxXmhWrFX
QRm8nOyIyem/H3DKc64jRJNQF8QyIvmL7kHMJ6CBp9Ceeb63SxRvaq6sT6D0X1qb
VIuiRa+bBR9pFvXjOTZSWZXEJ5sJJcmTEYL6tR+2K5EoSIgEo4uToEjz4TzTAq7E
/SyDe5pLVf/YNyLCrY3VirJ2qC4ZGhHjIW+FxnU0Yc7LrV6AY/Q6wv+omXDKFeCs
yEPcQ7YbL8nHhxM+g731Fz0h5YogI0IpMwHeZozH0BPUmTuweInVGmSG/kc0ohhE
UlCj0ITEgVNsyH8BfHNWjCt0MnlHoYvA1+xUmM3TR1+OkFoEtGYirv4ekyGQDV1z
SQAG8t4LmvMCZ8LdDmkFk5CUvvQIn5pOXHlZRu2Qtud3XpgPwwLW0BJgMZyv/QSb
r62ozrKvIPxhAVZi0Z4lLNXgujY+mTNr0nsS1kyFuuHkJP1bC9Rn3qL1qLE8oC8G
Bo7b3aIfpYxKyDK/Cd59tCrSH/smCRtjWu0SBKv/lT8xHoBZVdtixGIReJEOp8la
iB7FDycai6diiyoY6EfUorGop14SDi6kIK5/6D8rS5NUk2+Cy6va88ek1OVA4JCu
hKB9qr43GLMdNtPeDUnX00VPymzwFCnTDYCQy5lv2T3GrNab11qsRWVTLcDUBuCk
qCBZvQYLYDddG2xyoLgq3sxPTMC16w5ZxP3BOavmfO87nr5vvUZTbW18RIN/u5XG
lt3NGDG0xw/O1CF+I/M86R6YTM9EWRnAlOMbrekQOPPwzFOUmKGiR83gwC5HZgLU
M4jDcKw/g1umJmcy3Y3ORsHfWOqoKaNjUh01nT4lFtvkf5pAukigYDFJOrG4Fd8M
vjKrhFHVKyO9E/kghNNUB3qaa+JPV8mhzORGdfOF29dOWy7iJqtWYi78q2mXrVzA
+67z0oE8GNqrHilmLwOYXk5QwXtUzLLfCb8yVEmwXvUlce18hyVWmSpw6i2MEtyO
fbiD0vTLAjJ3s0BCO5j89h16yj6pMKEAF++y332WVKDGqPPm7Py5KXknMgTcNaLI
KfMMFU+wBQiCIv/JnJ8VNPLacKclyzWwxlE2rWelTI+gAQmgXyRAw/o2yWqlWEwB
KLc0kS3a+mNGO4VOPDe1OIqgXaJP/jTeIXZpBqSwvwsUx1x4RoEn1MgdqgxxNkN0
Qlt7aZQaGm03hAA9u8nr8Saw4f9uO4qSZslNX9G/F7mMYIvAC5u9KCkjGQ23/11T
aX+a8v2InPIMICP+ga5rirZx14GTejGF8P+SDnIZE7zlmRJ4KrdTo2zQlrLexvPH
A7BzVIfzAf/ITB5HUUAUlehfeR7HWFNfayb/j2MdV3Bj8aitCpfCFayDSfpedw2d
RlAW32BIWbVF4AV8mDMHmn49jVOYY9zF/nL9Bxe05HeunDf+MZEAZTaOp7q1anw3
QbUEv4KGatmPZyTccm3GxK7cHYnujPuS4FIV9yh0d2GJYxRYWbIsZ1RIoBNcyXvJ
LdiTXg0QEV+Dce8bt5s95DQ2vly+djh28GKKNS53K+pAOmq2TMglmXGWV5vlYSWM
HAdC1xIfyLlcNjp+BPCBXenBflviAFHMa3Wi99ggU/vEDvHLZA2obZFby0b6jKt1
8ouSowpIuy4/2L3tr33SEWzC/KhxsRJD8i3R9SGAj6wRoFfiqy2uAKtXqalyM+Pq
sHMLiKEfMZT2ngJFwA9Q0Wb/c2Yo7ajSS6gSi5d1vb7qU6bmiUepTuW8/K02I/LK
tik4hNwSBE0Ws0rK1hQjUfE7XpggN7axOlCN1uh8lB9In9bEL01C6++tBpjJiEFC
6aWN75rp++6mapYbYeJWofAmbDNekJrH0picpliaJ5AyG9n8IA7gJwOW099N91p9
x6kg8GsJuW7IYhPVa5NW8bqcT2FG+skXghKl0gnMsBJCZxnZeKCIAAXgPWmP0Im3
N3i7GIzOIZLBuMLa+FZaTgeWi7crazh6dAp5knbDAyplUb8MFklgX5jTL5XK7msS
ohgopRn7e3ql33N6EFZJ3YpLiLh0tA7HKSJBI0wvZkA/8/uYSq7qcmczArISDBjc
+v1VS8HJJlmNMEN0+pndgycQKAws4I8QNPeaNw9VMz1qD5Q4qmPoEagQMuYHdeUX
+A9AcxFViIn2t72hzn8gtiIjKvV6MvvGDMv2D0duMhmwDScq+UFOBe/rmy9CYWud
F27X0rDURB1+sW8IbYf8u3yD3ZaNUO/U95WxQSnQJJZHOFRJubsI9iyqVFI1X1dA
A2S/rJ3BvRW9D2lhOcEM3J6KDsonBzvhmapKmyZZHLYD94wh57jlxjR3Um4aUeI5
EWIe+G4/2wImxZn5pbSfnBarMxpeUzV+jEDKoSLcPBBvk4vt+Yc22DqYqkp/Sztf
aXenK95EseSMgmpyIgE4yhlq0lL7wLKJEECtlciprELJoTRpfqFXs2cnkCaPe+O3
D78xKPoTFwhePq/fEZ8gI5wDAyA4WRkFY7Wzdw5FbnTRWaDGgNeSKIt4jhP4UG4I
zyPf07L1XJsoVauiCPxlCzXAUmmLnSovmfzuiUmb7yCuRLTmWnHu37iEhlzmrQzc
j/YAQh0n0syPbssRUpU7uoPZM8qdmdDLMVQWV4wf9GgO2YE1RjuAUjd/mPu3xcnL
9qTThC1695jo7STD/0SVPUVTHn9X6xdJ3ljZcBZDl+Tj/h3h0/y2MkKNJ7+sLBDK
uFXSU1wwlVWc30md22R9Xza5Gh1TX400uRXk+s9jgpV0dZds+ykT+GXuRTHvaW9t
WsXGKim1ei5mAXjLSqFi0r9SkgCQ+1WV1elBXL837yJovyd+kBvHbOsOiG99d/f6
fcC2irPeBQqL7rk+MPafA24fEg8PTP+k+2ZPJnCwErp0Ha0cZVbiTkW27z6eLhyS
4MAXxKbX6FyEuD2VpQRazvJWvohYAVhV2Q1vbrVK/7UAyBf/BM0m+S57dg0GfYpJ
rSMFI2PkfFJH1qSYynTvY5tKfwQUhJITtc96XiUGFCU8u2RfNsPYh+2sagQA/B6G
E421qAmvoATMhZCdJ7J1jfUWb39s525KtsQHEExuAB2koLq/PFO+VB4Aj5GRR/xP
dBj8DUWr+ctysN4U85lun8eI6GLvUct8zmY/2QoxIA699Jgl14L+o3ZcV9XD6lsF
ZTmi0nkLmCqUTHNi3blnCydjR39/oBvNZkJcYDuLORQWqyyvDKlexG1DkBtuRdf/
bUxmirKoGe5PkgPAc3wdqzTUBh8sLjxPMiFSTwvSqkYQo8MJU1Vj6BebvJ+kQnDk
vrhJFXxj+xK4nbkm0oZFe5p8jKOwxIJYgLRYHE87wQOJRsDU/D1ok6ib8znZBm6h
3C5hpdaG4h0hjR0WtGWKvaJ01oovW5zsmmWN1PY+IXi5UNe9feme/iRDvJcL03If
3UEFxd0JWZa60C+diMJ597aABVdz50hfPUXkpJlpeYr/9gPC5cgU5gMFT4D8BQmp
s/OqoLowUVHlduBvwUVBLrfkEOe6IFes6hfxOrrkPzSPv7SdHp4K/zsOoLk16aTP
xRgUgFY3gt1fgbnAd7V4NbaO9MOp8L+ZRN1q+QoeePVdGCMpuIVGys9tN27C2eF/
sIdRBpSC3r7tQ8UGtj81NYR7GhY1DMeGT4YDpGJK+FNtXsE2LWCAk6hjRTj0SHth
0zuDrV7SbEkSC1rN4w9+Eh2pkgfNEus8pqxU5xeeV8Zw7uYliJh6suAcILfLVwDz
96OP3J6p8s8Mc+8FWslxeo6/eR9bw9Qi9S7cyRVe1yu8iJaj+8S3YKLqwiF9X7sH
6z/PPcMh5bGSy6+laEx12n+Z1hKa7FD8gd2NZstBX7fHJc8CMSnlgug9iOGm3601
6aD4IfKPRazZeAJnR4RxHOuy02n2UToD2C1ZBJ8YbKid0lP+MVHmHz6ZFvIffuNp
Td39wgogXMxuaDI7NHhjFe1rFNUOGG/mDH+CSh6XLjvjqc3YIujmGVMWlDjY0eCf
+/cckeFdBFrqhOcd6FQwblc36ULq8aiE+v3ajilq1IfpGcvhreQCW8ooX0mv+0C4
Yxv2EB/RtYFg+ANg7gEYIRwNjnOvCrQkQn43HWk3Ig4RH7eD7EuWe0k+c/2NrEPV
uhal6ruZA7++adX2a3azRFnd82DE3P+nFTIolerg/RvbIidsrKk9e6G7T+SaK80d
OfIEcmRNOTFHy6bMZP44pP1IotTE/LUGZ7WrFFnxLfy6/62vWNgRWRZ4fsAv8coX
H2v/Sqhb8YQ0DHFzu3LARYanLBh7Z9WzUxosW0bEAPlLhNvUY7DTMoNeEc4dHBz+
U+vvCPofKeuttls/w3oCtayGL1yx9aTRL8rkB5w7nr85Yf7RIxaIrwUJN5sXmof0
/1IMC6M3TGdA41weK6qJ/3rhngcJZBDembpfHw4I8+1i5PEaLdQ4xEFZc9SPYtdX
e5t1qpqETQxJ5PUBKZqpTZCVpDQxTdZY+cAozaNNPLBtvdirSYX78utMuWe+LL9+
SMzzqatajoLqCTBpaw1AJJv2J8J4CKH3B24pyAsJzLYd6u9zI+MfgEGXiBmO7vXX
kMgxmm6AlGc4LZq/pXQOqK2J+cLnvBqvbqIBzE6fxi5kTx4uhKhysY7x/th5ntm5
iMnVjc0+9YiT9xK7GUnBfuITX35RPrejmiZmFqH7BRjkP6ehqbTrq52Wqq1yLcK4
V08frPVK2h2drDqJfTDSl90m1rhUfVkItQOhIUWH6Thr5OY8ja/DMQ6yfYCAv7hM
VfkUDjPK6w45iGaE8V81I9TB/ch0PAdqeu4IDdWLA4uyQwqVYgZYFE1XExhDEtNn
gcjLMhOA7VgoaEdhfdJHA/Q0LZIhU3S8kXSbj03p907QzczbvUE4qX6340FcDlRO
s7YlP/fvGK1/4uKlOkf6fFF4MPRKLAAhWQq4NoIIyTNIhZpR0FUzoRZ++PhoGyd9
Z5cdchHURiqfFRKNu15zq5eBmI8Mg8p63/jMHaAVTx21jslhIndC15KADfo/9HFn
jmHF2se5/+1zg8/0Jv0H/FNzBlmlJmwMAi7rL7kEibL23qJgxS6mlKAHBWzb7yn5
PnHUUhUlBADL90tYeKRxEbhZSi/P8fEaPW+xDzleHOcqz+WUSltFtwDzPFvT32T1
oYArIZ+kBlxLr0UTJMsnMmBtk2yP17KP5+bUjwnHscewAA6M54Rp/g28ULrv9ju5
6H8HeaYDnJ0UPz6llDpKxmrUUmUg+BO08Jn34qrSmlf81NJ/R0629ZocpIp+hnOl
z0YVAyPAWcabI1CZ5+7kAdx3Xc4Tr6Hu8m6SRjZPGDy8RFyxNir6mUWTh4lIn+Gm
Lssv+K7V6APL4JrENMfjRhuveRqzprAaiFAOOf1owJG6K1nQQURXXzoxixLj8KDT
zlBluuLiRcAnPW8J7EE4Sv3IkxYhyBwRqPC4VThaiPbcKmStWHSqoEH0n7JCUGZu
fcYe6ZmVwjG2VGSlD2UT+7vFQ5bh1sO8w5yKpW2ZE2R5PaXQeDnbTcuuWUl3h/Hi
xg6hSXDLOS4LRG2QbySc3G2cvk+qINa1FtnSoATo4I4TSY5d4GANfixyRf/wdHqR
zq1tSUgJykY3GgqBLuDBM8b4ynBIJD22SWmEyb9Jzw4O0nyonSk3//A/XYNQykKH
o4ELS27jsx4kxL5Nml3zWotDBVGclJTwDgn2Ljvei8PQshO8RsDAPjAdZV9PaLIY
/4gk7sko//Jv744AxLJdSzrgqnVyqzEd0VTQdmc9TOi/3muT3K/ApL91nHczuI4j
l0C80dYruRl17TL0X2DX3GTL/yKCADslr8I/ogQlBxf6cqv75TSiv8mUhBjBsGyh
cCO7dFCnN46njMWCXKzSJaANG2nCT8p0qW39FKB8NJeSAooAi8KpS/Y7Cqv0w4IW
73Sbt0RSSlxhTOf5IeJTTFw06VAaoObX+Z7SdQneLNCuMRZcaKHRnXIirRHRyz06
zBd7dzGM3CUTxNi+PrpxhtwNz/udcD6PSkXPABX74/o73+kcyBA9wIWAOv4RT8im
BiSN/nOaVONOPKNo8Ym3itZ5K1Xhl4fiRjoemEuCS5x1PLmIJ9a7R/UgTRx1bLIG
jR1LKlXUoFXIq0Dh1SpnoSUp73eBJJvEbO+JNgkA0fXo5HAt1oerUvr3xphwRD+U
jQ0QmXV03APEjRTalzf18uaqHEYMKJq4eDeXJv0wZmdW/vnoHiNpIjGuDCMK+uh+
0nxTJbr4FiHPEmeOeGNtyBNTCYG4+WH60zsoKKxZK6qj/TXg/AMhp6t0zubychbO
132OFE12ryG1VVNzj0YqsENX6pHXXhLwSa+z9JEyuL83wGdJhCKmVLjLCZFYYgDe
97ubnkOxGSC5XSdo+U3mtsudN+zTe+kTLrM9m2vcfr0Y4fv52reYLvttLPErcYZq
SsYsNaUa86BmCzEXMWeUKowEVX9Wtj7OZhQn696ZTnXTTLEIfISX9VDzHPSSm0qt
QmuQfC+gYh972sjh5BKyZ5ieVIFn4ybYyXf7UJKQ9t3seQIp+hmi3EWtodgeJ+Ul
sUiBHgcIt4zuBzJo72eqgwN/huNH7BBffQA1TP3y6uXmuYlraaFa6FY6uusMlW1a
iEomduCc9DzOh0+mbjrX+tMstSTxlnNsvBF4xU3RGOkV+cZZzsJW9JDiFQCHJ1uN
UgNML+DqG8TCgxGwBnJDmaP71oep4CQg9+zpwAPhablmzZrw9++elJaZMmHuGaD6
w910LZ6ycJMpTH0eCTTZ5wnTlrOLltcdstNhPnUEp+rlfEM4UOdrBuPtd5dHfUsr
6XKqM4tRHX3IbNCMvZ+7cUWHezeZ0mDVPnvSYFzUB9WUmKHNQKrhtDuphA3rWX9P
U2/Qa6ZV8R9/UNr+otKQiDHkj4tfUbVaexARLvr1+1h+VPqlBO/F/qcwfUHn9rxw
oBEdQFEDs2bFyfea5RmQ2cELwMa9o8OtlS26QLAPaOUxRQ2Ds30jMtXoLfNvq89W
x9Oqsb4iC+nqzILQw5lBajEZtYDIqi7oJNxNYWOGoBA8t4VEuC5iS7TDTU0zqFil
pL/eNX10geW7QxIzfpI4C1ukMTiX5kXqbMXsOv2tuMhhdkmmRMKl6z7I0WF8Z1T+
TJYnPNYu4PyxLZEC7jytq6N3z7O1PREz0+v/gVp7CtftUO2ASxFiklfjakzw3ev4
ILuxxx/ikR02n7/xEX4/sDghJx9GeuGqP3hDc3gBLBhhFRsbPbW9i9ihWKTXX7RK
LYlmMpZZOffWraNkD+ycHfsMOQm76I1na9p0YDTOzCAei9xELN/c2FbXsEW0ogS9
K59VKodyU4AfEjIHX0ugEAtCY1fZJPR0TkaRqaT9BTbMnPP6FwUFllwdvmEf0fzG
Uqe+3eokI9hsMuswulDSFScjv9CAMMEPReUvz62dkrkO/el82Ds624gJFB00iBRs
ySh8fIw9vbIiKrH5+inyZBmirhwNnmdfo+18ovMTREt0rMFN2nphi17A1t48xnT3
ewqckPG3L4O4zgS3suQjeltwGNuVQFlY4SkpXYZQ+HdGSJtz7ukTe1JfM8VH5iDj
AvneWiPh4ZqvGvxPq9Qhglp2V/kKoqEdlIhh7A5hhS1bu3u90TsBD7FFDJmw5TpW
AZV7+joIn8us1jtIz6hqQPc1YkzM/RUvomfq8oPXpulF2nFpNP+KiKAvP1Lblq7D
qMvFYMRJ1M9Zi/2+o5dXexGu4BlpyotZBFCo9ClgRakgF/eehrGgZ4eoIKIS8r1O
/mjiUIKRcEcc/9s5aOS+0J8QOYAQ1om7ybuOAC2AJDvB+SGb9NzGhF+Qz3AJbcXH
nKk//rZdvp42fm0R6dHr2nMh4yudovkeZKAOPhSKCJIMbedKqUFdlkm4GmLHwz0q
givP2dbAHTNbeI8TmhHT+0kSvVIgDFaxwU7sEOBg/S/rUrcrM7lX3dYT6O8g2H1x
9OtPc4YZOZRdC13GFR68ajrP+IrSPgntANVhzx1WOJxwcQUn7ZcRKoZH4/VclCJa
r+QhQir3BycbQKM5qv6D9uZxFkmAwUHCiAjJ+3VQJjPZhMWrPNd4tA2XzMx2gyA8
TSVPKw8eznbGgr531A4L63EEfYMe6TrR2Lm2GO2LOD4cZJI/pjwOMgQ4wT+CSEH2
i8atZaARDnMIqG9vwaAlFJ4Oykp3HG7JN2FbAJAtqbtXtjCE0AGgHbchRLQFtpZZ
wupjKYl1RemVcq+FlSu+BRArDwheUUTWDRhEKswYiMoz/VC21ZSXETRl9dwnESlT
YkLMWppoas7Fti5c/1YG9DOq5/gVXBO0fCUuRH3VyGK4ezR0ZQLevsuLa1gj4Ix9
Gtn8o1M35zUFrKoh78EMC5YmYsOorJ69ZcQ+xSxlT1xFqImkDVvNt+en7kaxeAsY
JR6r9gZcQjdrC/Pt3RVoxM6O0hBhF6lFC3D7dCT08RKnKoVXuLVXaLHsxq8WbyUX
4bYq049sS+m/wxHBpU6CBueZK7tpsm0qOwt1JdBX3bdcQZF2zMfw3DqoxxhyL5gH
DFvHNEeNDHdhUyqwOkzjdZ9YIvhgb9zzwx/qksgP96htiwaXkSzZYgikw0jC/Vbw
Qmet/8u1U0FgupI5BjXNIAEoex2bXlTFd58r3EVyPSDyakuudxjzrMzcXPDufDDH
NHzaLz3cJd+MOJO517DL38//6zHaBZwEZ/xdziN0RK8x7WS0fPoyFC7111tkHhnS
e8v9UAsi+eay0TMeUJLGPH3vi2bRGKy1wQ3ABUjc39co6Zn0MF90TDr8fCBM+LRI
pLZa0WL4Ty9BdvivMABe+aNjYp9bB/ZMZKLpuCzweqdYbl6NVBdbsY/2zabxIakm
TBR44DsK7WyLSLuainc7JtiI3A+/cVEpYDNqfD1W1xJAvTF5jENbfFyihQwaaYDs
HqrJM0JNxBFCs9LqwwB2V3WJrOIJfiNaraMWxXXK/xngcG+fqi7yjDbFrW49UgF8
OVxSaZWpaXhvW9qofvSNyBUquqkccJ2MVX340S16mj1DuGBNdl4MbUj4y6HMkZM4
Am+zXlRnTfpkXOKY0liDAEN5P4z5H/fkEoWRQ8GGgOVDfnEoTEkvtAhOqfRPzbdS
tiPtS/9rkMIh8+SFE5UIfHfdV4bz8a9OISfRAA9vRIUX/iQG9mRFLjKIBAG6c9mn
5IxIYvN9d3oT6itSRWIAdneRbrWzcG1Z1w6c4dD5RAvm5+3WoUDxuqc8dvqdIedQ
ab8xTBEahnkwSiGf6YPnGjUNvcybmitKCl4mfbiZrq6wyiT2vbNRXXs2iR4llGP+
QiHNIldyrWqtktKkyegTd2JlFJ9OmI1bkpeCqa3yt18KinU2Y2FMvgX3rWajgTEK
Sm7yZb+whEaAr6KeeuDMfKcrBS17hobqlooNznmdBSbgp6xtnvzooAIueVnrKfNp
M3ZGoRVXBgpABiDFrZxZ6RYh3vY9H2pbacrfWr3IDWGYNdkRDlG9Jgxo17um9lbM
VOobtFZvz849wZInVeIN4Yjtmv4cYN1Toex2V6j6W3FgK5GdaoHdBXl0h3Q8TOPl
NqyTgEpFYcGebmOeOqmGT7pactFJgevAXUVVYizpG4U1u4vDS2bU/OYdyDwpe0qK
hlIzDOfV3wf8Ebsfvh2WQi/UlVK8ARhUWG1wZ9ebvnNbyFT/rEOocpch0Gcxa206
I6G7THlKGaJZ2lB8nIHVzQ/kYhucIl5OnV8ERWpkNI25056Xb4yaWBMS1+MaT98E
oTuvyJF8WiauUZptVXwOGacQ3elH0xK+URr9SPdXtZ2N1pYc/KpP6GD3nGdsrrts
x7Jo08i+2GjI5YlcbAGX970r4Ld5kE9AZHmDibja2GzJm8zSZUYNLS1fz4i2nf85
GL1wOzpet+vMHeugO9srfh7aVvyh8dg1xUTkLA/1x8s2/zQPqGAmXSBc7C60OnDv
6AjeTs/OKLnFxNzPbGf9rBZc9rY5xL6n75HaenatLnMwsF8zrNJ11PYeJIXrOXYb
39IuebEYUyswIykMaGddLFqZFJjiFqH1qSpElZu3dh3VetRLGxLZBThduxRiFJOk
MYLTcpytiPtf9lA2JIw5qvq+WdDc68bMYtTYIOeD8+Uoyet3WLON75kLkjAF1sHA
RHUAxantS8ebKnihjXHgaOdkAFMPrGTmdYRiXNuK99q2ydxhq4IL6mq6lII3EjtA
mkPNKeQEldqbRtmesKz80NbKOPcO3Se0Yr1pg+vGjNxx/18sdWN3RsiRR8wIjg/l
DGwbdrkN68pVqV5VFTt5HHHDT9VDDPY4DpAtUxKvnTm7lYqDgbjjL5izcI1X2kGQ
KlgP54LBNhmf5hkrWfK+zRbKeqaz9HBFx+QDnoUUS0XvkWPL1fOAgGgrzcQyU6Sr
tE3RWJ9cea+2TExa2ARD2fN1pFub5gxH3wrp7S7DzA0eqq5Jo1+pnm9ngDYWVIW6
lFbZJ0JD9xDf656YaoNq/0+fY2fsWOH6wlutoG42uWz2ylzHj48z73PddqjoSbQS
DuTTqdTR26UhWfDes7mYpT+j5CdclT06YiZpIk9pmyJmvDPnBp3CoCLjcmLck3Bp
YCvxLiLW55bS01idoHjRBUTxSFAcNPKZDThXoQctx7jKfUPM1TBkcgtwjVgY60p2
cvy+SDu3v++pmh9XlbYNrduhU422M2ZxBiFYVv+PMlNb0nMzVw5b3AY4JVctcc7O
UW+x7EWa7hmI31z6GU33uxK9apS89PYM217SDAIG10HG548UjOAVTx7iS3TFW2L+
nQsB46fsfbsPsmc4zbwpA/qXsKBSU3CwEi7CAXgsJD8uJesg/NH1W3Z7ew+2Vd1g
2ngE/jn39Tv1/GU1STMHaq5RDNkf56oFImai9wZFEgUbZAIXrRsmM22D6wmHf4YU
aorM+dqrfRIhVr39az+PlIuxtsPOFQZGeVT0TB2R83QQpB9RaUXXPoJnobF7e7US
ax5jwdiSUXQ7QaK0vnnvDW6m73Az8NgC8H1etpZIpnQi8aj2+zRWIpqFDiOKTHPD
dfOy76rY4SVM3RjfzztR98oYjITt+E7kGvtWY0gnVuS8Thk7VlQPnMnJcInV1Oca
+XW0dlq3dlgcJpCJWuyggDRK9S9soS3b9aFRl8cSQm5RXfxjjBbEW0017Uz6BUkX
gT37Ii8N7FUyVBM2JGXl6VxhNkYIU4IucIt0NLzrxN0EWsLeZtwpwr3Vj16jjfGj
+03qABT2t3r0MY6Hr58JXOlTYmY5Gp9rrP8j7pWvvD/Ch86lvpqYyCESurMATrPI
GecXfL0JUrCBc7tPOa2c7Lc48TQ3QxJHlLKMHHve1gNlqaUATN7bmarAA3Q1YJ14
Rd2Mt2J67VP6uxoXHZzTAKKJ09zDkujiaggWdaraFX0yrwfhmQXciJ8a4M9lSVJf
Tl0c02+MHunsCVD+8hXYSl14yffimlj0NEQjAb9Yg1hio+ZBgAZLvzZLtw1TbvEO
e+rzcfFjigOuBLXJIzRRkzJf6QHkgIG5SxzMn44LZBL51/gVeN/ujKz+gSv8jLYP
/UUw7VWXSSLvrFDlHYm3mvbqzrpuhGE09HXMOWOJWO0m4sxQE3VmF7AzzvsgJm7j
fhsjmtJCN98grLOTGzcFK3WMtu+OCcjWKZkcC+2hrVXiKkrlNGMIIbvOH9uK+rMU
GbhXOr9NrUWqQ4XctkQAJ4vYw0DqyxS1PRYwNgWUZr2dyPqmvpNAtwS9CSckb2DT
1bRlF/Hw3J5Ac49mS0QiViqoWODKA++ay7JRilwdxYVNwQSmPPXx6P6qgdD1mgSw
i78Ac3F8L1ylPEyp1602Yj0lbhcH/CmPBBIkNJWcAH7LiWmtDf2do4m0IIMKjkbF
/bctDTnTb/d9tsFje511aciSkdAxODtVUAwkQMJ/Iwe08M5EAmSTD3bq389rQ6x7
BOp8HaFX4qQMIoRXG5BS8mEtkozEHkJAX7sNO7oRW98rgI/vdvosQYHeFJdxPyi7
+mdGNQyA7MnbytVd/tmiRlr9CalRaWHt6PtnhVyHtM8UEKHYrH4jjIHM15csJGtr
iVkWSu/ortCgyOGI4MWJ7/jEY+/cIcmFckt231MpBFK2RTOxjbtVtAx4KmHKVcUD
By1xcqFEBYOHl4dbhOn3RMfz+fcqIbnlRGHhPyiTS1ck4fh3WZPzp6HouZoAw7UZ
fZuYbJsCcMGUS/e/KJsCnMTXkCwr2TEMaUZTv1PzB9sMeEickX5BV4ZW1ohURRHE
2VYB5Entn9p4/500qYGiEBAZZXXYUiVjo5TnAsXzL11fWdDBTI7q0fnDmvynvLUO
9OS3ybqnkBgmTtfgklfMLZiIFZNJD6xmP4Lgl7kHMF+u45XvaUqchKzVhueQ5war
FrqlzKu2BMXOcyQW9kksoteEcC7B6cznX5wWXkIhVWUSljAgMZXHpJ/0H82bx77C
BLqS9ZOkFsLIpRg2Xt7gy2ljx5KD3fCPqc2eoTDCZQhB6S+S+7qQtmz6R3/bgza3
GyEkEjSnzFA+1UuDAZDVImRk6YPPVoR+rKysFdUuj21yCXGSIzvDNS8gd0Wc58w6
iE3z2Ym8tjPMf74uVTeTimH+u200+f+fIvS/K7pAAhur0W0Q15Tls6CsoJgS65cw
KuiQsdA3mqcDMzS+tXp3L7Slm0Vd7fPT/jbWsml2hUEELyZ6aLmPgbN9hi4yKgld
xWLj6Tvfdg4B1HRsv5WZX3CNzqEYCoB2eaUyvyoOnaU5lhHZF4KdK1bs7niWOiIH
M3kWcWG6K19AD2SAuJViGlObTCVcmV0osI2A57UtlQEP/pnDEloOJNuvZksez36j
IRjeU5qDPv11lgfLKctM6bb05fj+Uu6+IEv7GTFeLIg2r+WhT0eg8sLFl5vz5Fox
JEPOkq+82H1hmoFxdpTCtNtu0DIr8e2WVeWdqpBJ+oguLnbW78R8Yy4PahBrtFu4
boXCI3nGMkGQInS0baFg3HVqRykpaWeaURVewQmk7/DHxxrh6/e/dQaZKTVZAlTU
LTqLexyOGZP27FcmwPmLFya1c06jaRfsXgCFxTjYOvXGkOO5gRl/HOS5btg/3Ur2
CIKr/bFv34+CvScQLQkNbohPpVmuGsxbCwQI0H+/PIFWxzal4rxhFLJepdwAAV8Y
V/mykirhn+DjZh0muGGPRmnz7ZrkLXMhlpEb0v/U4epqkRMlt+x0vw4903JfEjg2
tcvfA2wjlXFsRvXV2HlDMyshmAAptv2NcWxGu6ogQslMTjlyBqegJHJRCjRi1tC/
zYyrakkDdONmanqL7xJ0vjgP0UxXs/JQU5yTH6hZ7WpMBGRew5z3CU8vo19kmXIX
QDBELRL64nbTWaYjbAdaZA4QFacnpRjHNZqMziRLPUs+hy3A6mP8oqHwmUj4Yrjx
uqpM6Sq5g5vw6DAugtPcwjcUhzDcOkrJrffgpi+AMQjX5askM8Hl9TQxL0CaPRwG
zGdUcuBTPnbWOSTIedb+AWujcWN5iQHZqxDbNWbse58gIWUuIcnMraJLI6myX0Cm
qqtNFGK3Zcj8qKIEKEwrHIqPn534Caifk04HRAz7pakmoof0nV8UHWUoS23PaXQe
9rUmqAIeldniMMGOOoTgvNw9tP4YUncMFZ6vFdiwwvGJ27QKIVDa67PGPSMMvzOw
415WsQFkbfNlCRGpZM2QsQzSOIKho7oZ7K7MZ5rVQUi1+Yh+3RZWhJLF/l5mZ4T1
hFZaboKP/7qPS+8ZZv8TuHjiRqh0ka3939C6qba1NliaTMgVnQEM+YmHToXuezZ/
exlOgFYsLQzSTB5jLo5Uh9JirM5/+dZY0BGSRdk4w01FpZhYMu4478TL/2X662/6
3Yra2KIFQCF6DVakhzU6aLw5GWH+mM+hxt3dPmUNlxgeTc1uEFtCXdUKJRa8Y2Ql
68nygiplOk+CLrtRTm2YtiyIMhowsQ4rIs7yrNdJj66M+mIcFOyqJgon9U7MQu3s
QnSVJH3xEhRtj0LTg5crLuuIWFeEESqOM3H0BwjqZpBPvHenbMh6Usx/hIulzHjY
HZnXO80VBi/xbHY2W11qDjB0vnS/rNszSGZEGEdao5nCPnDYWjsREnLRs/PyYDsn
uDDJTL4NqcRtzkpteKFUWAgK9FUo3EGrqonQquzKPPc0PFFOHlHgZ/wztpXKYtQn
e7TMhJ0xU0ngOJd9f9Fa1dRcLblpCiJSJKSM5a6sDURaccvOe7LI77Qzi8G5kcBq
SiaI9ncktMKCIsdE1G6IGKi5b9wVZhu35UvuMgcIz6VzbbOQabTYht0m1umbecpU
Vevx4DOUbURNDr0ReROE0BCvy0DCz61/WcIxenop+VANaTlDVHKcwuPgv6U46qUG
W7hEMEDSq0jkAyo38Z7bWUpgZRuLOVHbgLfw6hcNjO6+JP2W9Qlec+P7msf2Es4F
oFkyPKT4JK3eVb8looGIWD3DhflEF7GeQad9yA/X5D4SpFPnRCNLmcR7RQXotBmM
lQjk454qkyzHSQR+feTUWlqmxklGUpbt32pXU3shpo8qjdCiOIIS1o3uizl7NdJO
CZLbjquczN1G6FoAP3ISs76iFkBTSljy/nY+UtGVyz4/P6c1emz/gAFw+H/vSSgy
tytxURMzxCpIizJZgScQS4pfAFENcOGI9zIiysrr55vU6Sfow3/JlFbrkRjbJqN+
AdZUDB1M53JJxGnhE5Vgmh2Qg75HrQh4QHSyjUmrJXDwhl+w5Y3O5QQrhfX37o3s
S8elrhKwzjFHW6n2PRFuq15XhYSrktOv2j/4W9p/DIB1884s7ZWHQMy+jmlmSRqo
7tMICliAvaTUeWENoY1RWMBTUfXY0D7IXTFUorOXWtoGw2DPAwwBIi50Yeq9v3Je
BQy1gmN0EtklhSahAg3s1O3KYibw8T3r/kbqBR2qprXJX3KoaumFHDA9gVN4i/tN
Md0gNLSzAjWx/zeTOcxaRTBSWgaLkxQwb7Cl5Mfnlhslegm9KBRHKC8sw3SxsoVP
vc7NtmgT1DOmq+mOcnM0mE0K/AsMIE7k4+5B7Cr/nMT+R/aE2Li2ur3wUL10/oBO
E91AuNFbvT2CziW3JBDjKxoMThRvxZ+S7V8ozKM0X2BA9u8TAfi5/CPQ3mxuAEbL
YZFsjqpMHQbiN17CRMXthQC86ZqtuVJxlekExTZ5RjWxGcv/J7HCd7TaONoUXYs2
7rlnS25/qAHGcmhu6mmR0OH5fXXFOXqsYi/o2vEohCSAz7inhKLpHxmRoIbif6dV
8XCJPUiCcf4nuqS8v697hY1reKelmcy1mliyHqJrZnJ8q5zwGVNlc8THLsFKA9lA
1qpuCDFMhe0Ysi5fa5YSDFcfQOlExP8msDZs+wOS2/EH72EBmhczspsnBJBmHHXE
8u7uPcIiAm4s8sLbtlHW6SXc3sbltp3c0p8hGx5spGsMA0RI3LBcxG2GWUPBqDXL
BZDpbw1rmAp0bTzKjDKGCoEYsGVovZxmPYsc1ALAMlegU/lRBe7DfyvehvQIZpVU
4JX517JkeH/9HOE6GtifJycj3AVtkOdeTM7/WdzIiPXRTgJQAp9tNiHZBo+h6F4A
RGmjc2Ovt9JfFUqlONUd1iJSvMCxws7lDqqPdEXSDa5QXMhuxyXi4/zpdQ6OMC70
SIktst2k1gxSHYVEe2tBgfyol7U7l0G/FSsML5GTWDTKwROwUCsLedEWkNhdRfGI
4+lNrL9Kh1UKvsmxdpQxNaWVnP2cf2p4o/YZ0cpdx5WWxH28q88d7O8W3Jlf1duK
QZdvpJARAUWI/yNnPxrr2hPsGNC8bGfeKgLYzAtamO+2eSsewanuGtpgpytKW/T3
L2r5hheEJoGcXvOYXFx65DxQM61BCkRB3pV2f+UCLmpqpYKsDJLOq5TW6QoSidP8
oQuqkUUAej11crA9/jaZcDLY+R3Hv8xIDJy84t1z9R+OjRWrMRi41SqGHfA/TAPV
4hTAfc8E3CR76qzdAaVw8I0shA1K4pQXBMuzDTMV9xSdBOuHlF2PCjV5bsKGpC7S
rW6qsqoYxWGh5wSfIjyyDXkaK3HHs1kSuUW/pEozQfc5bX/fGoRJy1a5oRINBkDO
nUMaadMsWXhuXKf/gKVFG/Q5lsJ6/EOCeVtA6dJZylRU1OsApji+aVPVo6SpMUgD
SMAunZ1RCQJ/0qApniSapBIY3Py1Uwb39sJcLizl8R2+oWm0aG1Dc2QCJ5mWxlm5
aHc11Ri0XLPm5WIHP0BinG5x/XYatM6OOjVd4Lwb8gl/2+B47HinOD7ksdNEXvsF
RwSqUGVDn/6ky7Z/imResYBFN+qrwS9Je9ke0ogsVtc77UFeEtf2uyAQQh7G/f4y
vYQAZST150KLgH+9YphZOoCuogOxQf6ghdIg46CISyIunOgjNoQywFz6c+isxbzI
5M4oIw5G6h6YKAXxUzFvBExy5uNLsDFZzEaA2isj2IfFVGQMn1cXN2Jv8nlFM39P
31rCVRLu3mf+Uu0si3qewJAFzRBI9l6C/UO9/R32a0EmDAO2OkZebAIgauasHAFd
/kDAjpA+CKl9xQcGPMAVIv/bhFJnPOVjDjCuvDQuM6Mf/wGvIYZWnHN/XHOMsrF0
xca+S2IbjYlVxgSia8RQaOci2tG0YyMamdcjXZ+6kyIriUPQRz1D5J4OeMgM1yCw
AHmy2m0+Ms3Ub8feBjaWpnMvzjsTTDuEXyujRfSdbaMTdsyMBQSE0MM5in/9prjA
4r4ub9pUFvaTQYtjdZ4th5wpL1ZLYlUtwkUfFouf9dk6Dsiv+buX2BtvE3aJiT11
aqF6xlMUas64XrkiSBfG899e+kLB/BV92ZQhBMd6wWNC4FaPilQEJVruOmg3mX00
6MkpB95R6wTQkDDiv0PZKPeeTXeX1yeIxCl5iGfkKwZSIKqapbT3PnX6VdtqhqbB
traOjcJGnSkv77AvmEINrwV7uKHp5iw2kAWbJgimqcpMU3sOIO582aJQZfoUR8pk
baN+8QzrTQiAsLwzOsj1bWrThm+e67iSFJI5Ik/QkoSBSn19dctkw3i1MFMm2pcN
ZlU9+t4AhmO+mM55a6/jkhD2g7mxTXrdly4ddyHgphOI2g36dTIHNFJyWwoi6+t6
3ImFUby/gPvRCWVDG3E8sQHssnyaHNJcO1f8uRQp6LmrocjI5XyVxuaejWpDwQ90
TzEiGtPSetSrBmLLNOo+ZkjK6Kfh77RZMzrDU5Hm1TJl1LiVR2DEE6jtdE4FzsUj
a5JwW2478asREXpvTbUfwsIyLXRV9oLZ5B+s6VqAG78R/Ka3k9CYRrylUOC/Hlig
UiTaNxO+89H32lanziTSpSyN9a/Zm0aP8HBL32lZweh9+vQW9oJWi8gYFItgGHge
pmKjSokpnBy6cjADW4Q6D85ir7d98Kfi5oq4HJsLXKV9C0zeAy4YSsqJzXOtpGFF
WYnCOxBaoFKv0zrbK8ernNi7aKL3gt0/6U0bTkO/F8JnuicSZFDo7GQNhLYZk47p
7L1gpsVV3Hh4dKK4Wls8qudStc9xHHSGGEfNk6XZSkYYfHRtTJQwjm1roFATvIq/
Z76+OTtwU1nzwaFVFM2E/zI4n2hyZ2fhIXnwopWtUYtk1qfaztV3QySwCOBSXs+E
RKaUc0ESKbKH4M32ZqPndNt4VPBpRvsEfIlXVDGs+vCpxMZtKZHSrcKXBinz5O+x
05Tt829DtkA6OspMksJytDcBDPHIKlP8zkp0XUcjdeDCZ2qvjfLgmT1WMZCkguTn
QSUwVxQXTho0P6INhUg+nb2SptRlPuiDhlu/3Rfqrhoo0yoE1o4RWr7aUb8qCiWI
/bi2CeemYuDHzwRgOeevPqeyi31WxhrQ67J22EsPWDJIv9p8+L+nXxHYTQbzI+De
x4C+JZbpD/XN+hFsyuDbthsWGQYd2sTRl0yqtp+lUtqgSn5PdJ6dWJ2cVOE1Nvji
2+QssfD2mcL9lSESY1Q61ox5DKl0VS+Wg7Ubfc5chiyacT7phMPm3cr3LsDxDaBL
mGS+TxoQcgzgLBhlqPtVf6QbUVd9AKJOKOTjExNn+wwNLpP6H2ObUGc3GnhhUSag
cuY/YXvqEpiha2Fe3vH7Fy5UlPXp/+OZ5+WjMKssM7lIgi7X8YkZS7nOy0AzdIZm
qyrb3kPX1/wlZLX6utevNZYOuywN6KwODznWVNUZB+CXEF1a7g0cMRBpfhrQg82m
2V+lBs+E6hekgvRr1NvGuP4ngeiQaAvo/0QbgmdOmE1tjEHbT4bP0kT8MkeF0CMc
xBuSF+UKwQ4fYmA2UESQd8c7rSyBo5e/jR7uoKSp3JDqjoQ9OOPjihV84CdKY2wZ
sZtHE8mTgXfb/il5SLlGxEuQWOxih8YvbnARjUIriZP6CzJfDQyotUigqiiHV+tn
snn1xWpfqJ3+0sxZdBpZGc6JnhpDJfXwd+XylHf0HDySuHdu1yilb9TV/P/qvG+L
jJN5K70ObD7eX+bSKH+eUyVkEbSuhMn+7PSDJpzbpr0zEYHr1enVKBli9tgCjHuq
cpMXYjxpH/jss0jvSpmV84VciSaOhnuJ0EmtUx5HAzogjEs/FV8sNU97Ur3mpedV
IPi3l9mC8OPXNlBcC3nsqLY85qn4vSY1rP33ukCahehOPLZbp5eF3hLrpLlna+ob
nBv2DqSwnytOzEkMQBDuMGPyEk7BXGxyq+MrkL5ezuhWLzcafSnVaeZvFF66uZ47
enwLnbjRbWO7FVP3sN+5Hb+wnBVsLAk00A+FV8PQ7XwwXX/MRJydz0B3GBLZ4mFT
QFLJcor69mEL2LwKZb+Ylk3hu8nVEu+dY6fZILPnRHDy0uiH/0c4HSj9pkyW6jY1
u4iqWQRo/p4guJM8UC45ISeRg8bNMJf7TlD+5CA6JGdE4bbfWlyD8ONxySHXMYXm
lt2XtXVUYg4aO5kDy1MnfSkFTDmOVGf+lxMJ+mCJulH58cHBbYmKIFn9FNKXf/H7
OSTzrLYNfWYyeLFPJSXWLYR1vmDV4y/sHEWalcdVJiC8WRXWjNoAkoxkiaA3SSOq
FZXPUfuAJUZ3K0osmn9CcFwOvZGG19ixmB+awIecPheuxwySOLQdVqTTir3sNCM1
JHK4y1QrQPSohO0tOmuCmPasA7wwD790GkILPLj/MNeCJqpZYgNNqNGQ1TQUWXIz
hLT0Vv0S54QCjIxWcsjcQODIF6Jo7KaHaDycrEmWTbcUhPlpGSvpQyFbaxPjp9ae
ETMNetV7B/2P/DAiEsaf4KsfONx9uYNWhduE128K1W3SgN823KbA/1jw9WeB8VGe
+SNcKIiinxp428lt1Zx/w06XoTONzZ0vhSuTWWyQfeLkNmzQWOQ3yyJSkdwIrj1s
aDrpG1azpCMNCXQuGW0rWxB1nURbQcxKL2Xj+QKFnkjHWE5UFI/1wF86UaRyDnCx
f039pUq8E13aonNqaUP6SiZaX0EmNu0wc2UitEfXcsA4EoNpZoYH7Gl4Jcbo50/L
BWtNom0X4rsvYMh8bRmHit58ELBfymmvuIpBGMLiZjZ7+OipfJ2WC5EkD8cOpWEJ
Zpfa6LnCX8lhXCSUcn03+F//rivfuTF9i5eFgsxu8GdLOPl0XIXPVQK1YzgP9p3s
O65WbYhaV97rFkuEBA8BeOY+i9FmpjHQmptBBX0treuLI/gfushN2zTZ5DgcIjNC
YxqzLu7M9WXy7aRc+6Q/13eTj0SnMNzu+v4Z+7hyg+koiHtw+qGETzktpU65pie8
o8xE3axMRWki3ulxg1t3juwUX+3SMta/ZQKl3RU9OiAqmjpZ9KYRdPXK8yqcKSH2
AzlvZvd7fFP0a0vxr4tbwao7c4C9rLkxyOrEPYkkpmeqxJ7j7lJoXHSSFEdx7+tN
dMcAHezN/wB81jyiaNhX4H40nPzWjXlA+1QRgkcT+FDG+laImmMdiztHUK10kOIg
BTr08VjyrjNIamPN+TffAYd6EIPtDwfxB6mnTLlh47R7t1LesSwgCXimiioMxsOp
T4Z9kU+NCRNgWaitgsezgsW+kKwHW5JWtMldnanitdqx3dL7GSEVZECUWmvKBagC
wWe/ls8JAhY26JWTyPoTiDUXh6+qrQxNTKz5XY68yNmaehejrUYDPf1yrb7U9hh3
kSTD8lFwxNhOp4aEJgbn2H5O0xuTrJ//CdQDT5nITu9mNSQkdehI9Tnbp0yEE77O
OItHq8AH3eyCbV1ePX3D/6f/2FblWgJbqSueeQ5MVMzDevLOqudmJLydwCp0E87W
hDMOHue3bqe0IPwKgahJCiJNBgjm0njW3T5vHKL3jEBeodq+4W8ZUZiutC1HNEbk
yWFMwmRL1AjXig6kikTI9+wEqjJUh0C1y2/wO/G8TZ3jR0uMIkEjsD3SCdPmFHoP
klBLgaT/6l0fDpmLo5SXEKF7J2nICSsmNKwras+sAbmvar+/fvg+LeT3i9d8815x
DXGOs+AHHz67vOD7YQEQkVvTzu13bLmEQhAXEF4QO8oz4i6d361uBl2uccGvivRD
4zyw18YS61kyRPaHugAKxVmhNmKZSrjIhZP79OPc+cPu3ebbz2P7meflQe9QKE4c
wYdDmV+5RqHVfFBSepAP6SFu56KwaqwOwMOlLslcNbResaVUsLZ2iRwEOPOqbic1
Y04Zqmfaigp1h3VEJtHcWF48zXMPMLGDlyD6bKDc3+6U6jM6rGUA8jAZutiAiw9x
WNbdoHfya5NTwhYPRIrG5jwUe0d25TGFl0l/lTU/iqBiIbKbtHtLKG98kFzKlhaN
OYPm+Iuhhjc9JK/uFJCOF/cfnaqXbbI+fkNx2Rl8i5R9rGD2L64kVK2DGVZ2zBwq
2ttT+L9jGLrGrkdsVxPW5x1+rCIal2yRi319MGkkG5BJ29/rS5MuYUY8Ob/niXZ3
m8JMU9n7NOhGl12FfoMW5FD4TBp9kFX9MCxGn7giHASy9SdRICZ3Rq2E1Sxd+Sny
SSkrdrahV0TgEtTT9Wv7lCzut5/pgIV0UTrGkOKcAjbflPHMJyfbUh2JLTyUSXwI
0W63udh6aaej+OEKqRFxxrMjQj7VEe5e9c+8gRc7qIC+9t43vWWGEbcAix/xlYQZ
0JObBN69/0HYmnVQWuQziUdVcJpijRTISAwVnbRL1WS7S18OpmkgNMr1Y9XSsUlN
wtDzW4kHk6rADNPLZvAV6O4xpb1c2aGZF2wFQBUkRXYnvuM5jH7zF0RrukCUAjNv
PIcbYED4rFPMWscH+nyo0XfZJC8kHv7skDHT148PtryNVQr/2bzJOJSEgOX1TjrL
XXz3FwAdLJs5L1xT6A5puXb2dhRGddMafqMYxMIRuKVvggP9UIC5cm4gaVkl5E8Y
Ve1YFOwoZuPF/YLpGdCPjYY3auGH6LCT+3KlKj4y0P23Ktg7Tmc8K44BlmB7V4th
LlRJaTECDeB8yZCxZZ+6UoQ5/ZxMoTolG8VRmKXxqnFUjwsc+N6GY4OK4w2qeq8t
g8Cfw102XTdScYV42SdbBFKiQvHXJYTH1KJ93jO2YgrwcoNG0JFPjI9adPfPfHEF
h3+cjG49u6avza77DlR9GsUOHeOFX4IZCBPzNsW27/RfdJ28418dCdnzNXjEZ5VW
OXJdC6CGYH7xGOXuHqyUEl6QYQX0tyqpuT8B1/nq95a/ftV6ZfJ4gQ7TpIGU8Mfi
DcI1pUkn5RQlJrQbNd6UVQ1kVwEgMajfJqJI9ZfkIXXhckRcLAqvuanG3QlcP0ap
PDlgFZ8Ylao8nl9tpAilb+Xwc1BuWuyPBkPg1McwVMIMjp7uNgJajiMPS0VAG6EA
p2cdx7NO/0qtxzqfmL2n3vPBE7hSzx8pLeP6o94vc1oT42BzMLHJgJF0wIhgy+wL
HEvLJ/U1VY6SpaFbUsYTDccxzwDSR1D8axbuV6HhyFiRBzb+Y5kBzy9uDMJaFkbB
0rtKzpmxsBGkwrQBcR/8OJwPvTi1VZ9Swi3b0ZFAkT5PRt53sy5F2jX7UAyB1Ty/
ak/hRF3XWbPBgwb98PHl1irKoJOfd+ufWiVMIpM7A/tTB2uRco+IL89KxIGQ1+rt
64bYJziRlJi2MCCPC8ZJFeP3UT66lOs/llu/TFZyn2nrQQhF8LThMZ6TmThb5EVL
0QYH1xTVMdtcNiCtDtlPIRtINcnZU5NMymqustr77SfZLqeQ3hnc9ibEFCdMrAZY
ds4F/NX7DSFFDG/3hCd8+cQ4lW3cTjIQ4+1Nd+kaDg4jgoy9dRKjRmAqGvh9eerH
hwZml4E4wBetGz6MJAuu1/AT89iWIk9wYdxjtS5pArjE3SHP78i7euBiFRVe7Kw8
Oq0qKGmtscTTSxZD4FBPbKSJVcOZEWGHFsFnu4amnxeE617B3r0bytYqcLFVJRuW
57oAk8EsYUl4RX5wR758JfTQ60GsYkSn5w4K85uP0Vu7KWwRD5cUEN58qIqu5/TM
SDnbxbT6G22YG8rb0V43b2+vd+vW2P3xB0VXl6kug5mjvYpUgreebz6aX8GjoVXg
6ygJgxpNARfCEAglr/bQpiMT+MlkSQbpuhGTuxk1pSC4ZGUxEVKWBFB2KyxIfpbu
G3C9JBTMz57RlogcS8FzPD1SDdgg75F49pxBGoB87cUYk9/+LwAmlpnft7u0KQt5
WFqMrwLYDaCQSbZZLOydNONUQW6DrP4GuQxSXJm9jRvKC9tiuFplVVQa7s70HlKA
AfjPf4KWAEYuyWMEcsepP8F+a6P8K00pfJvz/49JZ4A+ij+Jxi/v+SA8LxnlBndb
NFnlQOTUcjgTkWiJzaXiQIDZIZWrqZ5EGYBGeBFytgJKvsW1opMnJR2WFpsuUZTX
G8OrjghUldDatP8qvlC7BECgNGdDwt7IJbF8nGD9OfXPZtj1zpuq1mX8cUTHesJQ
5m19r9T9co+6fDn2Gr7VnESYmpeYSoPZU7C+IMm5wOzjKSjpiiHgkXdlLEVsns5Q
sfEpFv6CyttR+gKfUhTDZy+vAgWPQ8oW2oJ05scULXz/tjMyQ2zajmknWm0PkqHV
T30tFImKmC7PBOkF5H+u/uzyeZbllBMQSHhORNtttx3XQVY7rkq68lRUg+sESdgG
aKC+fYZR2V4SQvOECgHaWWKCuj0OPwgmoZS64f3DD2BhTGK0BPCj58pramBpQU07
0KElgbzzTZy4R6mrL1nbCNS/H5SO0NxtpcbvtmkRUcfYeaO6BE75TWMEw5T6qH/l
E3F0Kr/SN7cYkw1XT3yI0nl9+E7TtT0YPwNs6FXPfAowhJCM3X3Wr9KBTose8Cw9
hc79HeSQadJTiM/N3VepeEqv7VgC7owgvSouF8ajXWJ6UmzylkD6SyHtfkOks2/a
/OUMCBrKSNsIycsMwS5AjE3Q8H8/XVaIUxv2NY0r1eTeDUTDV7lZ3VCfWPOz1QMI
XFDrWfpEPqAznV9h9iElsB3VlcA0KOltYr3iJmGxLkOa/YX2kx4Ojmnqq5ksTbcV
hTwLU5YgUzK/TyUCOFpIzTqjj/HkGGr4PoBEUfWL07l8RtUkMwgeG2MDrbjVjtbl
KVQZbIJ8SXTvAgquyjJmsZ5FaOwzQV/3GQabiv6SoxI7QAkZda9gbA6EmcV6KxOU
Y1b9+oVDROiMi5S3ciNLP0VBHF+EPpnxSjNvOGYi8VmCtCaxKZsFmxypguLKpeb4
YCKq6vuV/nC0dQiB0s6nOLmt304AS8U6i1PSxkGloFm1rFRDnkkVc4juJNjPMEjg
eMV1Y+Hxr+DVI+PeR9mNSrCHl6JlOs87SeE1DqvMkjvgBL3FwPTxv+ygvrWpvi7b
Lfyb/wr0FIbKyWyCawoNCDij17Bp2d6wWddnhME9Pf4rgsBtC+4dLql8mYqsNqKz
3mxt3qSkGyMX22ab15nJqmyW1OZxkJGy61R6nkorJZNm08IWgkqns4R4+vURRnxa
bepsZATHzFuKpLelJP23HQklURsINysjoAGweYOceA0ljT+R8QHK3Fh0+rkC+Ygh
TDyNA8v2tUHmwaPKOpbSgxyxQPktd9V9kl2FCNLagJNbKwkLXpnfpfBnFFYTsuZo
UMyTlJDU0BBQmudauoJqL496k8zA+01gYnFXKXnI50ieOSQwpIZ3AA/CbvPC0tti
GA8h1QvQhRbARXQSedl3U9Yxt+J3LN1NjxESRgRBiAgZIYsiJYKETM7AOXrelFoy
FUxl9eYpZICzSO0x9wry/FAz+GhajbXQKYf2lpXzvnnIjOdoyY3ySdzxvQ3Q2mFx
e6HMNPmAPp7QLYwEj4oYnRXym0ppaRMxhh49swt9kvzU6yr4OoMoj0ys3GkMj3R0
DjgZbPe536XeVCB9Q5rSIIvjcVgxYDpjpVS0q57s5+qu8I62Qw1MtKIJtxIsAC18
7uDuO+Rdq6jIynlWrQ4EXRn9DR5fVhWR4i5pkpx8Y3RX1UgrVIGdbE5dGgl52g7b
OoBzhk+3UN8bizrxmymWH/Wu+p7n5BlK5bCefn9JFmOnPsT/rx90gVsiik6DlaPQ
fDRaw3I/XOzPJPkbTuq0dBlPoAD+G6WP0cqGrR58kxP39YPakzeL2BlhNJoAFNAK
zbXvy36fKB/AF38KQENl7AfIQVOHPH3wMGffu557sIB3IdAnBk7lUs1vSk17olKf
/OTcKxDBWHSpXyKVwT0UPo6OIlDC4nkk9lb5iRuKaWBZedFFrqbXP9LWQXhTPQlU
QnFLeXhwli59w5zeNzMyfZPN3EoazH8QWoaI2Blj4xaycS7t28xatDKGpcT8oOup
hzMW36sD3bC64mvpiQzUIvVbqyGBLbNV5DA1QgH/ZN/a3F+5sN/HdVMFvocIaLVA
hD179p4U2O5ywG/VvO2JEDz6wa2RWxokmd8DNShi2UNTx1S/Lk4TaeBhP+OaBSCt
eFGZu9OJnh0hxEdihSfA0ejdOAbFKSl+fMtUdIOgh6WQdwLWgOT1RIyxb1wvYGp5
a8gMdGwFLANK2+1fzNt/zRShmW+iXsNUhMfqj8qFpoBpncUJ43dmqcILc5oH6F5R
heyneEZiXbjNow1eiG6rRzs7Wmax5NMXRn2rchcIOad6aUDpSw6+4Gi9ZWOLNsba
kj0K6Nxqiye92HBHXxGv4RqylXZNe8WMNL3zVx/hHRPyqzdlt+uT0CaaUtDrl5MT
pCgiafjRwErUw+Mi1OSXkYxw/cISZHMDj1R90oOKACeOsxO0oeInd3J5pA11CyOo
LRQdrkQf0UAR0AWsyiOqFswasrRxDlDf1RUT/ex83ZooweobK/tuUJTahGdIZzEX
VyTLKHMaNwdXHa69dS+cWddex38f3zOs3GUuGw1RECENpL7LM1gomV98oRnG8Pg7
lkIcgWPGoZjoI0jL9SdkVsRVJJG6pLhd493vdwYNlYMeLl1j3cFnM0Hd40KMQDj4
fiTcmveBwIyhaQ0MqEZs1f8otOnrcSn2eYusSW5XI19x33MI/pVKdp/aVgkTHixA
6Pxc8XEbxjeAqz2jS501LmbfubdWyl1VOCiSRVrACNJYsxWuBvRxMVm3m0Iw6oVL
zpJ0xP5UHF3yldUCdOawjM2J3mTUUrw0PgfjkpcRFmPg1/Wj564pjjb0Tid8m6vm
FJ7IS5B+USTsCvum75p63/Fp9hDjo97uwGaBLc2MKOOwvsqF/nb+5rRvFA3QNBHM
3WnqaTRFe915zrc0Cappk76LWJwQVfvb1qkOqweuujFq4RhumIB9hMzUb9zZ1ijX
vzdO+meZ8q/BDmL+Eviz1tIi8zNLOWUqqObi6AH8Mexdr8IKd7haMwZqOH/YOkO9
e56pEOIaeEmGpaOis/kOkKaiWUxxmUaow7Ld0lm0A4+4MAYk+AzLUV117IgKm9YC
3O8sotlw5uXpibGtvpGjLEKZ4geVu0BEq85XWzTzefb54+nhlRrkloP8LzwXAS3Q
W1nsvIWeo70g88XoC64CPErLLA1TJRb5cvBXpui5zw0da/uknLnPIBgKro2+XLmf
XuOEOmkwviOSJrN6nPsmyXA5T1iHhislv4E+DjmakZAapJ6K5WvaSI2U5xC3uvO0
sYJv+HppxJQMUMzOhCz7uYe0u6Jlqgjb8mroIBzsFaqVU7XmcnJMc0zrsRInHJMR
EnJweHJessiATGXmdTdCo2esM/qod/q7Upxq9B+S1KuWx1KSBTL2AeofV0degKp0
KU5G0Tz1iERC6T3lx0msUABS4Wyg643otscsh3WXmtQktq0Z/y4adF1cNpCth+/I
3OfQfR3dfgCNnHFueKn1WREBySikn9eKe3sMPYsZYo7jx1eoJgypCb/MpJ1hzXnf
uS0gBqOUefccmvQr/kY6lNV4+1Ifh1uYdyquYtfcyQRT73ZQO3R6wCc/zsU+9AFW
8QRpMP6BYQP3spi4/RgZWlQNWWWkE3nS8sMPFZxaHsNLnOH0wLkmOa8/MYX0IGmT
uRrzovxW0kgPUxqilPMvMsUl024jPsg/DUxS19+IdBGaZqbz9ZEyUP2gIdSddf8m
Wto9AYpTrKEK6JhMcgFeJxunvAJKdiKwVP2/eC4rQjNy0UPGfDaeQjFKY9IwfOqF
ajGSi3//uHsaPZcUT6kavfxopsXoqPNIz0KPp9Y3z31v1TdK/NBULkYUG7I/ZbbK
9/NIGyHChh1Kpzoie+8HinFLrXLB+xOP+7qAhFq6R01asG/1Ps3bN8GIK/V00/5V
PxVmswSFCebQ/zZcSfgWLEGAMnUeMmuGGp5dcJTIwXle54eXew2izEnTw4xuyNRl
g4V4d8Klupjlr0lzJdw4ujr7OJH5jceysoOYhAV+GsNX4U1Wpxytogdpt6IUwZz1
gl0mPHaRcsuwM4wig176TLG30LmEhlLCCy3zYjtWEFSh1tFH6W1YvJXIkyT8aWnt
34XYKNxGnusxjwg2MIxN71gSgitCuhomiIo18TKnQFsU6RfLii+qndTZxZYdf6ob
U1NPXCaDFXLXHRogSuxJNcneyaW4Y9UaPcs9mZaZB9JQv6jC+/uGJJ4JJhiG2emN
q8r25n01OoqYSRs9OZk7XlAFaVd5apYHm6HGFsu4Y+WwYVDhLJmikxIgA1WpsNo0
O8CZaoKU7Zf8vQ8OaDqDdElXdXKfGJRBcWopX9JOT8Vw9AGyqEB8eHqgLNBVdC6b
R30S2u/fmf4Bz4dfTPQ7wwLQCU1QN83dhBMoy661isruUZ12bNmBdT42bFSO6+66
5l+9HZ1W76Tspk4SFVD8f029st6tzCLGQe/wJT3v2nkTPOni9O5KfdAa/0U/Xy+3
0LmPUweO/Q712RUnKFOWyXEswoHXZ739f3h4e4Fl79o7HXrXk8LNJqmwQJ+0gQkY
fVYE9/Xd11v8JiBmAyVsa6jFuHKaSalrdUSkOoSkB+tabAzV5N1lCyj4UsauEX+U
m2lDdJcivIMqobUs97bFCgk/tD8r0V/PUHUIq7Nj0IUmYDkvE8gDxBE3p555fDio
EhxoeAWy2YkOlCjCvcD5s0w6wP0EjQuAhUGW9sXkOsggsXRQhiXaUyQ9XiMhRnQ6
LCSKUZLY3xwsdZEs++pUCFOvuI8XrBgxf1fUttaZgneio6lfA4sPgEC9yVgz9ocV
4WXKPRh1BXSygP3B4fcYy8wMowoK4/u151NV8n56v3BD2QWmSA2Idxsc3ZszkRdJ
4de6TTA5VFpXSOlvWovhQrJNdaVNZkSNnggV9Xn0/rnrUt2VEGkhop1kakJhP/La
t6Vlir4kVfJM8BOYL5Bqt2hzMbwnHPFA00r1YiQmMKf6w9SQw1i8CcE75+4wnbja
3bUDY8AdUIcn+imqfXrCTtAg75iVbGkFRv5i74lwuis6Hf2tUOZT1qKVNv99z+NS
a3LSkDzUtqsenxfcxWWU/+FGTVO3RJT41Web6KV7LlP/L6p/juj2XZGNJW0PLdSE
ZdSKI0todx5m7fI9RMqVX2O9pA8kogvdZ319aq777luxJzGMvP4HYXw8GDDs+QaI
ThkCtpGYV2Tjwy/BM3L1YmQPq01s3nQuw7r2BNFzdHfQndgXwbKlQsS5sjqplrXC
JZaZQGRIm6A83IjTHGoihCMauG7O3CS+lx2F0zasskhAYa3DDb2NGOkYxGviEfgc
cezZHkzaJPqp4y8eBmycPo3EAlfJYBrsgn4TR4qw696Tx5qg1LziJQVN6+1uL1e2
JVl+7txKDhhwknQid2GwouLEm2Z5DuuhySBzrsoKteiA7jlTtfpI8a3yuxwpZX3K
nThCZk3o5W+y2yMM8AID/dLUNNjMg5m8eJhJ/y9MHHJkvWnLvUniRkcIs/9bWK/H
NGGGdjlS2Cms2aBORRPs4UHvxtfqsLaukyr+URl3XBCgBXLxo7AGrVmaXR6uTcC5
l/6P8r9G05pq3KlmrkxKwC2I7GRfA/HCf7tbM952+BXi2d5RcAQGbI6PBzEYBPaD
kh/MV5ZRxQRPgnw+IVB+0QVuskOouj66fyjbOr+o0EMIHGWRl+P/ImelV7K+IIKY
zuM6gbexRSbHDK2lbn+SsA43xwTF9KN88qE9jaaVpRwGWIwOBk/IAyHP+uR0hOWP
loN7GX8Jp74LQ5ZfE2VplVUCNTbkXnzWqf/behlBsVFQfbcphrEgjt6/PeRM08mL
3Z9Bd5VzDfqFnrKB7Ujjncnp2v71kQLlM6kjSISZpZHgOcDqEoVgZnd2w3bh6lH0
81wmLnLBdyhXOVQy7BdQ2jF50Pz4vggAdXxyOPZXuIzEZdCKFmHyiAmccAk8Wt9r
lTkcVAG+zSbWfBdH+t0zP21SIn5FkIZVFFO+iUsUjVtiWR/gQhaVrT/aJeTGkztn
e4UJBndAAK4ht+2PAxeSZG2sm9GiZz3xPIA5WL9765rfEgqrHP1t2gYFZQdwyHxX
zUnHqD87kQX+mdhlVfGt7uXW9eOxGAql/nmZ47Sl8Lte2HraAJ2EKFUk4p1MvzW1
41Ar33nbm1od69+vyLE0tGeCn1d1GbsJHPvVp1sCY3xVmDUI0Z2UrOI168KpeWa4
kXIOr5Lz2+d5wht7BghoBcpiG8I5oDY2kAFy67/8CEZg9IQDquQlfA16dpoTFrp7
0d9cjbeiwr+EiZU44omsVuJJ1dglkC2aagr7CaG/0whUFwBf9HmpZdA1RrgVnxKf
LeL3ZMTtZBzBXYKb7pojhpOidfV2hYgCHnL0b4yzBkWfYAsM/RVFA8B0HcT3b4v/
iLksospIqesi4pdGhdkY42+3u3lsmz+V4lmCvftJtNl6WG67gweOxsyv3gwyY/zc
79b5NzuEXa7VjxdveVQ1/vHIoIwP4qlnb7nmg8hA3wAje3id24mM1VGRstVA2Bon
yThTD4BYDplMsn15FanubRc1si2HlXGP5H7NbAoMJdTJMO6lKR2PKf6xdkP0OFDx
FItV3K43KuYxnDfbSsgwz624qRX8EjRvecP3aXoFeCrIGntj+xTOXqQYAOTnA196
QjGZv8uRtabZTv+8SCSeE9R/X2GKYMhigIdoBLQwJnrtXHpn7kcZW9HJKOzX4WOW
TcuEx2N23Kag38j+H4oQ3jRxV7VuJvlAWg2ZYLyQuKAqroyNmoctZK416a7YRZIi
iD+1vLVt45hBDjYrZsMiqWKXPvS7CAB7nqP4a7bBZ40nz9C9vQZ8W/uRxsChFwu/
M9poQrtMYWg/WQ+tdJgXx9kxDVM/CvXH+RxpnMi7k+H9G6nEmXAqMItVEIDrV6OY
o7kWvsYz2uiPOCtM1+so6QREc86KXs9/1jArfkfzL7W+kC+0j2A/ioHPfdPCGcsL
jYnENPbDVv5gJbIv08lFE9Y2o2nFi/v+NmSpl47cwd5NknZfxZcSeeu3t7p29rM4
UlcPBv6OGdNQr7TO6lXh3KvQeA+Tcjti4duInVsy/mJEDH48DYaVDy1pXlpOiM7I
2trNPV8jwJ3mkYS8Qs+ENb+CUF6qyDLCzv1WWOQlvgo1Py7g7YPohDXmxP9v1t0l
GrOqu/sbsmntbfcVzG0vdnZ1KnjilL74qtFWDqJZ9lGxxcZZABNnUYR6n/yVbdjd
ibOH5ZCwFNho/sT5VtITfLQ7f9I50FK2kFCL5fcy2ZocPoI5lekcdyHuG9WpjZys
vZRDyW6uw6DAyj0LIbWe1Bal825BNM6QUdRymVK0SqCmOuKXNaIzf9jz11Jb1Tx7
V1rruvmSbi0NBlN5wuUz00/JStiIa5j2nv+i/FHKGjVX2R3b3iKkHERMxZHSNWOB
BbhQTO9CyzvOASNfC2lIuW0vzk372w9VF1kWTCIpCyLXdc06Egy0uyV+I4XVUezx
A7YDI5okupEcCW2wp3QHmM/xLb2DHA7LGbgPM3gRRYYM6J6gFB+hIIIqPebFAyPl
HWMJ3VbuNpzf+E3QyBq1NsiKM6lK9NKOfS9dHmSLFqcXhv8czLb+Z1kUwXp9VDFb
5ROzomdNt2MzXfO5GvW1CbOsIMr5V45cdh5mXF0xZk3875O8PNaJQ/9xB9pXux25
CfC9uPsotYPPBW3pUBdLxfS9/vTc7xnovvvxn3YYz+5Dv29l3kPU/pMBxwR8iOxi
seDqE0QQqfxfIAr7jF/jLN8PlLnPh5IzcIzUAGFwujz7xygm5oxtAlcD6QKdanys
J8/QAWHKp54cVQmkrEQB9c4CsEjK84ZiIr9GurkfANGD2OWHGGXaX0KpdLsw4qiD
Hj6eP7dP5JQCShcyNQyqhl3cee9DdXEdg202ARnX34sattieatrHBa41KSug8jLm
aiwBruwvoAdDb23v8PgU3Ev/hjVO5uKJlWsbHL28C/FIbKO+6RNoN83ozV5IcOVW
5sk3ZCiFv1t/hZnY4XkCdDQhk8a0E3LWcWHwcuYksjyQe1vUK6W4Vruq4iSiXVqG
xv2mM67s0pSZvvhB14aPr2GLIu55xCrDDY1fdtdQZ3lfRZ6gW8KcNp4hnFx0Gdlr
D3SewusFScQbzGVqMXP91OPxqdfJ/+wUFsTcUNehdLXFhhnzcDCppgTPLrQztPNP
UsSojg7k82mn7qIy/ZYZfO/BjgDtpvQmSmJTyn8dv9055Kb5EtVpwyDFVgQ0VdXS
fow5pENL5NuGy8L1Dm1ZNbmsxKkkh1zV74B55ul6Y9vtYbBxnnLCtF3p7xurTabf
0F4FCHqtqKEWdhnnWg+xq+6TdYNdRYD6Vzd4cI/Fpz1KUdvoI/I5nBHk8SYQVeoj
L4TkyE3KUUUufWROXEMVQE9KzF3uiRRjsOKgVqrwQAi6QeahbzBntmF47pEmrdiI
V7PqwWuEqUqoIxgl0GrUqDLfy22sW9DVzXiVkaZTFjssxwTIWjGtqMscAgWA7Jyo
8o/QDVlO9nDZg6WeC6wXtCaFuN1QNRwwz37MMTTk8ciuZyRbOYM25OwbOuHDEsAi
ytY8yWJJEsv1M94dyJPOVHauZNHCp2rELXurDsN2o0a0f67Xmo7qi8UXkj3pNXe8
OsDBjl25CXC38tyxEjU1HJsHC7QKtPALSzBM8E+uc780fKOjJnAfzFDn46i9V0pq
C5WwrbEcJKTBGFb76adkT8hbb68c47vYghONrP7bnTVfLe+MwWxIm7PcTbp9CyOI
KLzAbBLLlJ3rxddmzTW/+Idh3e4fiqpzXfUcB/4ipSRvMDyIZMRqet3Xd7DFci4U
+oR0PUm9a+1EBOn4WMdqcLRgXrMgfub+LnsaPmsR5t03XVBjenRgazpfn6O1Z43K
2TYEIP8vHqn1riS88uQJlZE1CGSyVi0SZ6XlOL6Xj+pbf1+C0vET/XLHuTIKd+Tc
H1nJk3Fhnyo6eH7V696iTPtwtvE608NSNr+B3FWPVhNqluY66ysAgvyjG+ku8m7Y
CraMOwmq8cPqFT3bwndglrq/sFFIQNnqypxweiAoo9YMKM5laX+dWcoPzTT8WGg9
cqIKv2CrfhiiNBvb4wERYPazwBLD4P11PBz2+p8twim+Ya13jJXQosoZwC3iId2R
W6YtIj12bwzgk1hmPT2n/Q/mPIarkhMbi65fOwDUsi72kq2c4OgCvRQ5KdCfS/eJ
2AAtG78Tq0p7l4Gk78JL9B2zrK2vWp5P6RSd9/DfhLlPrQRRfehSL4P5886CA6B/
7z9VOsLSyn9Cyi/AE3cYAVMM42rhyzX7cp0lP7kp1UkgModP7PMzxSVInhMTZ4mb
AvhKCutusZtLw+AldGbCreZw1oLmM2FbPdG9FZDgeTn0FeGmBWgIZRClPTePc/BD
59NJyPBDHszk6GmBLkWvfelwJVlHjhYTv7cPa5RCV+s2j9K5xb5l/lnAGhbL6y5y
AMxkZS4duP6zz6lJVL1K9bQelMqz2ksGewbYBG65A3QrQBLrOqTuX9pZZFJ9g0NE
hMgF983mZhA6vmNR9S6i1QND5uu68zNVQzOktWjDHaV9NDe2XeWpgTuyrjG+HPkg
VhYTdro3biCiprXyuQQkdOejZicwkQaLlY8s4IugG35BltadIwutsTTkPKaGVpcR
OBb3e7hTeQSsQx+UDm07oyYZT6EolgnrR3CEdZVhrN1frOIt+/C3nLQbX2l/Mmev
A4fTN7jVBeykK55MSb5dKos0ekkOs/auZr2tVzJR6VgEJrgUEqSAMyL2xxNmgrDr
ptmKEPIOiKYJvqYl7SOLBvKspdPZDWu/bmrW1qaXk23eoMnvvYVo26DETHwwBmOA
w2Lk800TTvY7ze8GZkIZr6xB1Y38SjrjYlgPnyauUFjgdxvJMS5suASmaXeOGUOo
iwmei7RoIO/+LEK4URF4R3LB1J61mcop0REuR2NWLF7g8MZuSIgb0HmU/UHM8X+h
72H4mrbLm/y6FOgHhJvuG5lyVmipi3LhEkhlQLjm/dawfh9cJyeWcgMjYznP2uol
WD7smjtRZayf5AMbH7RMIloIUu4qszGWGzxBUZZpAq3yhCYf3tmfV+mNGRwwdFVr
zAhgTuIxz2MvIKdb27AZyuAyjgXyWEePoii52OCKqMt2z2K4WZ9GytjU0QOC5K49
3PdGQywY3EREEYcZALnuQXZFDRW1MLySto+GHGl/NVIaWGF8TPSm8dzqQshhKIw+
zvzz8zqOup4dgpfVH7Pttf6ny87WK+NRPdFehYyzJB0F6ahQhyL62lg3u8FUV1jG
H8iUzxLPyp4RFa+ReY1YfSeCTI/7jWio9QqcbMT4WX8dHCvYXZT1ZGuV3xZX93gs
wBGBOteHev4Ej275BY4saC3xSLhOujUQW5CcRekEGJ6LwElRvdihGIOi9FjWjWa+
K6Tehb65g0NVg8QCvRMC9xrnQyqE9Pax/y4p94TVWBP+H3EdFJAWP4mFOfJitYd0
Y99Be6Zg/FFtOESmVKDC2vb7VX79TCk8Ey0hmgYuni2gnauulibsecdp0cIu1uOn
/p2FLby567qatQDiu0ion2jqnBiw2jVk6Oju4sRM4/fgnEK0obFTPxyrddo6ziyd
PRxPOjfQy2G4YeIGziFeHHMZu5IzNMAxEcayAsI/otFz4qyzhxOMd3DO9/fzEuB3
31XKgFWO8qUIHkxTsVVMoOzsVoMeLHiXrCaIoWasXLIMGvIZligddpn9ULKcqwCD
/M6/+LEsXtJUk40UIxLhRX4cCnQ3hJfLrrGIlkGR6p/PRhkua07JLVzLXRII1wlR
HqtpkQtaNutSZISmnmrKEWfVVWcDu6OwCAkikTiHV4XNhzDau8ofKnQJ8lumNdED
zJw0D2nHWJdQLhrlDOisHMvoOhtFzw1YT2cX7x+1M/l7RJssYfT1sOIKY13+amMy
4QHLuP4j/pC0CbW4/izLrviCaR49iodbYWIHO72bSWhjDI7KN74jyWi86BGDfCUw
2lUTBJj47Y3++CIyvGA6T3qiCD4Iz9B09yvK2U30z8b+C1ZMVI5hibFNm7d4cdbA
4VVKrd0mltuc017OJ69+3+ofF4OWvucdpWOIFgZEZ2KbaNaPyM23oZ+gen0gsiH1
7M5xGGoPXu5g3RMrIhuzsF4SKsAOmj5HWYYaCYxqC8LlHI363QnNnVxwVzFyo/Sf
k89/C+Wt/4R8bj5w2Z4Gvy0wcHs5k7fC+GMRmn/k4dG2+nxRiG4UC3jFy8wxxiJy
j8m+f4Nzzn8fpAS0CinfRKVV9QvYoH+wdXHs1QKNnkQgqUoHOARz1+c7xmAzRJKD
UjOSmRDmH/c9XCOP/m5bhf9KxO/tl27/QAh+72sjMbFazPbJEOscZENcFM4clj30
TzkOotH2PbIaAnY7v4MZgN5ZAl4AEF0xs5sNKHqQY1TUaWAWGu0a6KnbEY0DkWxV
pl2w8lG9vdAriTr/MivyVElZDZGnoxtq3shmLYuuCBVzJqytuW5IDF6+tzh9tVoC
YY8gchAB2g5/Pm1PM7RRH10PklYr9kaLugPL9sfRfDjegNqv/JMV6K9oRK43xq2t
I2OVIIJR+7n+EJ/lzygSkLutPhf/23NpUF3CmskpJfjnf50PzzZobKOWQDf2ES3P
ztH4ITYBjM2xhe0gRA3vAgBAqfhhi4wJ1S/zE6SkBHZcUeuJwNCVP2ZDf+ntXA7o
j7QRjdwWcA+AeV0EsEG70wTXMDc550w44RwWGQIHty6g+NmXhe02OFwQn8Qf3c4l
vue4XCiuRLfQ2z8p5XbOqF1jLtVHEiCpUPEFhklKwdWwp/gMVyXlvvVIMZKCaeRO
gXHKx2JyakRbeMWVULLfPmykbAEG9lWkNyrwGG1+AWoJnyRdMpzA+Iv7W6X1bbxW
K1hVbnMM7qWRq+GPMuuW+mUu+VksHUQYcwFee3Yve5UrBvAfw04MOCs/SX9Q61ju
n7LPn94HPgE7ZhYju5efKDkN4aNaBEtHxfhojcpgpnBDLSEhINu13BOCoK9PkIAv
MiTeff1jlxOSmx4x1wIVJtGfJJ5y3URQO+ziAXZGt0vNd8EHl516iSzDNlJp7zUC
PFerQ7qXy0mmlawBFJhkBc7Ynmt30yQa1uyb0gPTjgHJgngkaM9bqpv/PCH5aAru
jGwI+04o38PbvNkl7jNgEdnFZJJXE00RLVzL7XjklR3vjCfCFIjX+eDWzQmMKnbp
OW00qvIvVwRRZWjOjiuYnLU1pkFBNJr27di8JYEp+m+46U4hMLH/n/u7C95UiGzg
YydAYtOvzsL6irre5ve2Aqs3j7mmtiZ2LhjJWDXVw7hEnPk0viyXAePWMZzIRTJS
yuHg++p2qFyykvcLH8buh4fg1arh47r8M3sgsekNjWY3mGYB0kHKfpcfGKGRyYAB
UR7fg+iUq5Mxx/jn1i3xZwTMWjFsgTyOkoyJzSCKtypjbb6iA9BVIXOT0PIlyeeU
kWydJZN5lsNkI72fGfOBNRoxctk6hSZgQ4HTOYlaizcSMqlyraUwlUr0kLsT3x1X
hcwLd77/YM4l9WFmRVzYNKqGj4o2m88hzdQX4WWAz47SnIGvRD8KTPpLxU7IJB/4
/SqkxEShdncJKw7ZPX03Wk7MYX2BqAvV4yKXy6uZfz3oeAK0iLDgSxPcjAlIqcqs
tdoRU4fyK7MWw5YH/+y15w5iblVR8wZ0oMGA2KNjVSRXt6jXanpW0YLY6MB9MPgJ
pMCpOGhTQ1YplL9Ov6JOI1dOolzHxjt64tpPkafuRGoN641BlLrimach/dGBumCH
xfz1RP1vel8bF07OHwwbS15ZJ2nkGwiVWU9ykQFwmw1eg59tQsng6uOSWtPbmN3/
sWJPqGO9eac6oZ2GZvoN0QFOKzMw29hqMuJcq6T4XbajZRnCv9wySzsajN0MjBAk
/X5uQ086b7+iaJA+7BrjMTaO4A59PXRgafZJiObnk/mXqufBo5nqJ5Umzy3UzBhl
fHpa2kDdHvAHNadWJMEXlRJisQIJJFez1srCg5nvO8ATAYEykgVvAMrhLUeMCLXX
mEg9dXpXfeLCmQG65m8oMrTmacmQCQhJpTMi6WyPSwWYlajVA7+YYfvZnRS4/EBG
H7hjUJXwCa5v5T8yD7zBALzDdT/g6w1BdkoJzdgNMnxkxSf1yiItODfTdMK5TofJ
qYeQyVixQhhFgLviGTId2iBnyxFFy9Hyy1AZT5Uovd0pQVrjBMnfKf7dA2ZMZYkV
mixvXIttVueYmdDLTLFmk0XC6vUsf0nBO/Sa4gOtElQSr5cwblNezBCwCVQmBB7L
hlXGSWcrr4n5CQqql7avOb+WWuqMi/deznE/OK8r3j1lUdp/QeefRMp8KzfWjEz4
RBap5N/AoWjbGKcg8in8ysfbUkbyygX5SEhazZ+cKjKTiSTuRdISrBREjV/uZ2oX
hmPH6SvB5hfoPPN4lZttdl+U+KkGZL3peN/xmXhE7MOGSJbdQHOCLDhKLsibQjub
t9yZyBr3DlAyLMDhO6e+gk6WoDBe0xK+ykC1VlCV6sI8vCjkojxlreku2ewnyY3z
HnfC4nELPzdoNeHk91ceEOCJWdbtg50j3LNgctBE9Es317lmtlc6wnLfXxaDkmLX
zukNbBhWz1a74t1afkKXY2hF98eBXmDtwXTlgStz0kPPVd4s6FbdgpGyNv4s3A9v
cVL7VgC0JqepHyUCZYaa0wvMdMAEOXiaxdQo7MqkO8qhjWNoIdBumj6NphxBC1y8
jWfs4uxKsMj8LU1vq5ITvQfGeQNwtdaZKa5GIY3oH/85cERHgk83GDBfHFUoJm0a
b0FY4n9wEKbY1vDQbNAHAmailDTBDSv85NVDENeZvav1GXrVxGmAhPxGekqqPvRv
FpGRGoFnY7mFegmqItxxCKnKbjSmwCDaL7BKhfVRVySdDnDFUebwomllHUS3peZp
Pode42F8YVjXP8eJArLpotbKEHUGhuZXqjB5mQ+5/pWjBdlArwIeNKk3wAL2xnoc
idLk36k/veHNRgIdcq+P5SWOx0lYeEN7irN5OjQmshBZUYGxfDXmkN2Kr3xvZ7kT
A7yMTJi3pUUycupPiVuk6ItQZ+EpwVQ95AKzpeuRGDMTXO4MUoK7A6gDQ15QAPzd
opNfKJtlVaXw8W5t9lghaxV5sL8vMjz7eMxV6phJeGuB+LTXjyi4grXWY0LFNhNe
Htm3WTDTDUBAfc9BSbvmL52Fab67SBJZQybBrKFujw3Q9CRfoT9DM4tm37OTj3cW
MyxJvYgSKQJwM9FvYEo2nL++ZifoFxOMWSFv8Grlh3qqsfGta/CeUoAOUwYwYiZM
+5UgeIi24MhnDK1qUGpl2Wn1M7xqk8BbUr3GDA+6lzxFyrk/WMGQ1RkOBl8Lyc2m
ozE6JDs2YQOmjB/xGSYKNb0v9tGx8Ju/PpMWwkQ51ePrqBttxYy6ucscytFz5gtl
08CqBNUGFzA/5R+NLAVczaTmhGZLFShRqiZgFEianB1nkCzoj5Ta8v/6H2MDjTBz
fSEW71wCDzh4nf0laymwwEmQfkwSbvR6ZU+JERIquqpNCKvpz2Rppsc8sduY6g2p
Lsjnk+eWjLJ6zPqNGVVXep05/iGChR2yxYv1LhPLjdtOJoulm3Lwr8by1AdgnSuN
KW5Wpvjhejwq2w3jTER5ppDz98nmH7CKA9DfdsENhGUcWkKswqsPuTbzLNDxXzUz
EXFhMOKkeWp49s4Z5PX3lmR9wDOrU0SgBYPd00aaPsa2uYrP+4itI+ffI6hM5uje
NUg+TA8TLKQOQabOOdIlhzBPlh7wEXMe26XYEdIr+v6DHA/NB6KbNm+hANNxP63p
8M1LBjfYO5DBdecJPM/TJKSlrJq7ktxGgnfSPC0Wq2eAhA7QoAu3xaasWmYX6kDI
nZxygmkY/+vIUGG9ek+IZzZIR/ZeGjk1Qw66i/4JdqOvHBdP8aiYgVU/d0j3urfk
COIMWRNdqO1YLHRiSx4JZ9LRDv0GXpA4bnq2SGn3pGxxV9MWwRJGGSJxZHKiseA9
LsN7B2SLwTe8jyXBqYxaSP+yu6Hh1MDzRXb/ZTnm/O8UdkIDoutNsMAMrBMy9QGr
Q0xckDKtWAp38/fD2iGDhAMgVatlJOcEGCQjKGRqDTEAJhUWxgwULxmnHEBV9EG9
xE4b91yc+RfctnLJFRb2Be22v47XchQfzvnbKJBI1JIq+YBFEFJVVJDcquOsE3nq
bu5eOxBRP7rpnu2xH9NO819t+9zzG2iPqh4LTrUPvVX9glQMEmDHCxuHPmGmxkQI
zNsjnYfTkyyMj6OwzNCTcFQdq/aXNYfcF+YkLvdIrFI43wA/p4RR1dvyUgyTBQTi
vnMC1wVK8giDM5ao6Z0FtEHwXANuYydWGIpea8r+IHqyo96B1DbyIAh+qEvCDL4o
JnblT+DTUEBKK50R1Tm8FcPHGbB+vhCzh2w12HjqJd0aUMvWRMgK3v/Bs9KKWpfd
VpKiOGiUX6JEmUCJg1LATQR9y76zqsYBhpW4ZG9hlbQYBN3nOm/r9RARdrMbICCi
W5sO3gXNG2ETz2XmsXjFE6E1v4UA9O5043xUyiXy8lGVMXz+ewrb8lYWDboC8JQR
3GgaRkayihytP73nssxzpEao+e9WmlhS+p1uVDhZL3LPi9RMNC9OOZSWGRosucvB
96z5tarb4loIYRKVkQV4pVkQxCZspgJRNrtzSXeDlIBskk755z5m8aPDEFWRFxcJ
GWhLrn23zWJ46fXKuc0Azcf0+RX5Wk5Ww9FgEom2GIIcvT70UkFocRxRdJAO++j2
xSFkQ7HKA9YGiQB/8UP9ZzmSGk+6GVTSVuC0W5ceJIXeXY/Tlw1utZ6JOkqOSuYY
Gn2ei8nQYbRMoY65cpdLV7Q4b7FodXvw0Obos6ShrFIv4bRcJgQyP5IHSsa2cDRw
L0c/owUC7f10D3a0DwtzqWVWMXakKkwVSdpF1+Sw4b8Po2va2pOfMnwHdifzW0Cc
70B8XGqAHl0gx+OT2F2u8dJprkYo2AFfXm61YAe2sCbSULkjGclS9RfWdvRE0NTX
VP3qyn6+HmNAqsiqotBnoC06XcELnzUArqTLe3HK0e9fntZ0T8bvFMAcWNvAj5ek
Ru9noGlr0cXhDjwQvDmCLubH5MCoqedOmw8+Ue0m2CAgJImyBxChCHMluMyI4ah9
iqa5PXjg2ICNSCn6639h5L7I4m3jXIbKx1J3z7CSXeiplyZv0seL9ecewjk2YUGI
HioBQT46Q4vYrzZmDH57GyauxVt7Bwxdch223kE3qvH1jykCZlmM2Ti78aS/QL/J
ZESCu4GXHnxQCGL9QKv1dmmiPbXaI/xZ3y6SJnXfq8DYd6xSSNW7/Uyd+zu1SSBr
YznUcJHUxYXvoOlyjAgZllIUYOH//LkoBkfP3xTxxzDTRu37M+8kC98Oq9LThGIa
PHupBpj8zKAvgO0IiwiJzR1ME6QJDbA694TLmLj9t2biXM3BTPL3QpXEFjqkqf3g
kQVUIZNV8ozgz9O8/psERZZNAskVX6V0SaRnhfQG/q3uMMgGqr6vaCDwdCbDFLrT
HxHmPjPnH+5bWuPZPAPsxZa0MZ1crJWVNDjD6CaQBn3rXzVayf/nAzvx9n7NTb9k
/sg9Q/g2Jj8nZSfYBS72YUgpTMeI6u9LH9Pc4stNYmwMMJcqLNfLi/0LV7F5eDmh
+DzYbYEYA827r8WTd/HhSzXMAe68cZLrfjSImjQNjw2sDXYgIji3DPS6CUoNQv8w
6ClI1XDmyD2TzkK9SVS075R7V0WXYHaSsfis1MEkNMXCw6RjZ26LGZwG8AjoflfC
rYHKYnmYLynePelyJjuvOx/UkwHzZvMAGohr6lZewyOj14mChyueH3zJCieFoZY1
6YAWtQ9PUvqXizlOLBVClyc5eZwDdhwfpnJF4/U5ileBUwY1KAoCP6J7yri+TraO
OwM0ri7aYIx6VqfzryNptUULd20usmVxhE3J4JuZEgr1JdrC3K2uQoov+VkldKQn
IfMR51CdcrUI71SDTliOZG6sejwzKHNQBSgLOmY6Uwp+M/XY/kqg8vU9bIO+uFMh
Jkm5RtH2T7IE8e15nX9KBfvXechWNIegJJOU8pXt1MDc3DME2SfBJRkzGwlfZ9SA
LXB/YzP24q0/+RhGW4KW7RODEnBYZPPHbKkN12eXitAPlAfzSPLoJs6m8Yh/sccG
4Ug/8nS69QzNG3z1loDqj08bjJ0haF66n1oG5/pWvnB/9JudcUgj/UWy9Y+vUgPf
UlG1iYgBvOGbcvdASjL70MXbrVIS6sQ6yox+aC0xCTtdDZBsOr1R2ZrCn7v3t6VB
tycGasscDNYDwVCWkEr0lZh1zylkvR2xnbo6eNKxzoCLcUhz4ilmm5viK7QSNJmn
bMolOKAF8j6wXwMH/P6aX8BndZ6ap8uEzxQOs5TbGDlzJGNkze45s0OFNZ2RYAVv
GFMjPudrY0joGmP+H4A+3IR61EcYid9t0EilbaomB8lK7tS2L5iHRF3BUo4OyjGU
OJLHPgDA7y1+63eBaP6lVKlgq1uYSHxPJtsaAyroMiGjv4JDfas2M8T2JupLl3i5
Q+xlZ2xUUgpWkORQ9yvKNrQGfcL/KuCKAf/aOVr3L87I4YS6dMNluaTdmlephSiy
iLwB0d4l+kOiNvL0rciLJ2r3GgxYM+VXysg3PX5D9CsHPgtmFAONYb5WwWb2FI76
NgNjx5kn6LlM0zEy71Wfrzt/RGAZ4AU6QjUpkE2WiYjEOPOIXT4JaLKCOv85++UN
x0zFWZTU1o6UF0ZEu+IHKi5L4EOQb3Y0fWH/zLWyXpOcUg9ZZ1YAXUaYjP3KJt0o
xswp6FWhlqb0ylIvYNv4JxT9QACEinysdkt9l/qitmxcJfYSwj/xINHHmECjXHb8
Aqe68Kb00x25X2YFiNR2Jc3NhPpbLVby4UrP3K1sEp3q/s6F5AgGX9/3wNhmIH+E
m7/39BzgLJ6bGKxr+W4G+awBjb90ltwA7zpmVh4zUkQvRIWT7qekIPa31yMy0utV
uNx6oOsVrT1fmz8F6Lc4zzFCviD7qJ3C4GcPTLGk1irtc6Crsl3kO1O9BCc3ZHfI
TluIiMsKlnWVz90NfrEZshtgRyDfzW+tIWFMSTkPiGD1+1A8Z3qWJgiuGRIvngmz
JsSAGgt+2NaQvQMttw20/iWUP8LtC+nHvLcOBDHE4m1LYuWFZoW2KWYGsYrMfjs6
oLEGPZZTxsllklSvdbBJC5Ig+BJm4d2D25R1ltHaaiXVaU43tu/XBY+u43NQ2OoY
MYhojjVPfjtT4EnMsvGUKDI45j1ArcO0COLANFShS3eZapi5RIg0SXtj83gEGjrg
u0ULbfBss0n/yA/GPI7cHlY9GuGnMWkjvfGXkg7+rek7TYrRuKGHLL/wYukR3iZz
tlw8d5R2qoZymt+jFfD1VtPKswZOwKEewKWQXa+rVaHuZL9JbVmcruOkjdjNYw/j
8OE55tmKtSFGAfTn7V6+x67P2/fuTi4f8nk/oW2WpD3nnfnlOlF7d830l5zkdjmE
icw42kXr/jYS/4D603gdioZB7MpJidllfQNUk1qwFHfQ07its0hwDEbEHJtQcdrS
qcsn5Gb1Hy2QbBhGsG0xUJo47MlN01IA7gPNv3yIH4t8xqlFF1SC9oW+Rhgp4vSz
HsGFqQqJjfrj5BBSx9A8UTnrVvQ/7IsmjuIjvKexDmHnvDTNm1JbF+kKolpg6mTa
TtniLcJbzpSDfWJxA356uZc+Ve+aVZwMevecniJWvUnTSqKuZsJz7DCuQd7WYXhe
9OtGSIH2fujyOqm46mQMwToWFEKsXe2aIxLxtxLW/SzRHnUJ0V0ARA6lcLrPTuDz
4iVfcf6Z3nfZW9PHEpzp3kv6E8ApeRldo2BfZOy1U6yObDiMOFmPgWNaW3DhJHYm
8gj9MFb6sVCDzC5g2mzRW7dAr19wLgldGGW7xj4HRM9K/Reb/fdlQ5avtRH0oJqF
TufT9MXhwBeO8cSN3Wkg9HGZZDa6AXzmnfKDtXoMZUBjHthTQjCRKESTZ7VzI6+G
DQ9KWDC+D1gjHjGV7QESmd4T9T1r5RG8vk9Cv2btqZ90qraZQalU4DL6wui3bsTi
85sKAU+MJTOy0vxeMmZbtIVbaG5B3UlSL/YLScodCWTtwPes+4tKIu4xBFuiW0az
q6hvBi/7T7TtnPHGuQBLrAvOc4RxLR/4LhjfOoW4fqqvcGNheJ8WdU3zTQyNVGGb
HHa14kMC89clD60XxnDbCKUvtpVU93d+VldvjmmSPY4df9v9wyR2fd9aJb5UuUz8
aR9TtqrL444SIeGxNP+Lyc86ydfI3eX3Uzp0lB7YHAPfuP6Uw4Bgz0qU0vXyDW66
M8gcj0iIbvHXdymcnAKKC3yDjc9Hdtr6VtLCX2yyZj0OSYsmGj1Uo1atRi/1D1yt
/vyLGGpEJ7ez7MIar52IPIqSLEcNgyvmZui2ijN/uFRKaYSDhowI7oSgKEkzmZxg
OIVP18/DMmO7n88CbMvNVhJvpr8qPwQjUJ5faO99E2HGdGAMWhEkjTAGTrWEGSOz
L/82LLUkS5vBu34NMv87FVZ0WAMm4JqUImkNElMaalJEcWrJm/6WaG07qLJuFuoC
K39Oa/5JgNOWU4SbHMrnhGyfTQZxN/g87kaEXlwkhKy/fSY9uUmDMkmzeV6lyQdL
FHplFoml2+zDhriwAkBCStXUFeX5TswWrxHHK5xiRnXSd8s6T8hntfpJ7WxY73Dd
/Ary4Qd+GBKjzCd2fnej7qgKUdXeYrw2n3vLd+9sUB1p3AT7sDknfB9redy2cbge
ALOZTLV5159q7ghdiNiP74MwdCGm03PvWDtZ85uMudyLaJ+VL6zP8nV+g/9ChI4G
giPrwuvDd3a3Ij7J4q4b9nyzNJvstqSo9n+ReSqQIaFIKQ7ioctyTC2yUBbk30o9
68vs9W1bwoyPqAh/YxvcXGzQwRMBeoqZiX6QhXpVL6hqkzOtE7GtZd9WHztSDFnr
RutUvGeLY0yDHv1rw/Qn/Qr5Xn/oEPNw/tFON10TzHpdkvl69WbOk59Xhws3nMfF
sBcfwyro2bN1An19PaMYHNyJzPwknE/pg06JrijE/L9Vu5D5HPN29jIXWgi9t+V9
YVoRP8vPR2YJjD+IKlscHwM6YLeQpx1byadOovMGaXHvXj+YUW6LNiMxI4GrJzSC
8VvC0mfbO7wQxxMVY5n0AviNhl+SXn7HyTER4N9fIg9gaizkeCPTe68xF78atglI
WQ7SvdR/xtyUV5sBbRKMusTo52x+Us6jivGMbt8yvePbgJvS/6LV3oLFdBHScRHH
OsLf9Q0f8yFXR6vFanXU1XhLMPSDng01nmVOzxvXJaRU6s1CP76vUwmYRBO3uyA+
Pz6MPWQez80UIfymT6FuRbZqDqHBzOKJOI5W8l+xFDBrP/biflaBEDVGEvuvlIC/
NQKKRf3JE9JkRrpAeiJe7xDqTNNNlp0LDuPiRnpKAav3UnVTtjwiKz8bUFiaNSwN
AiBrO/CpJMYh794BCG/i2TbLdyhFR95CCPi790wAjMnO1An/I+QX5DLVqCvxXeB5
/o162zHrlZ7tlcbKHB326XOwSP/qvvWhAy4bqsm/JIKD71xzFZXAbGKbNmuN4sZV
jj8tg+ys/XtB7dFkj6HsNP3kNCBZQgROtltUhMK6LhCSknTZPb2bpzTE6Pzds+7V
6U/nCkllCvvTlgMM1/ejmKl1Em0wi3Q8i7OV4+2HuHWtNybwMGngIRBeM3ErlJhD
nx6iVGDjtGkTDxahN8BP5E3awSQzfgT9LQzS+fS/UB+VI467Rzv68U/dhHVVQ+hq
bTMbRwU6UxbzQywLTQaR9wf7tFopceJL2Mdm68dzAz4ZUPcvBU+NeEqJD8WcYvob
CFgeuOBSb+GhXEaTkWxRikTr54mQcc/iSMluEmLdDdyIflh/kf+Qijx3nU5Viuda
7U61Wo+tesspoAOzcOsakXLvNhnGxErXnGyG/vlYGHmOaoPOfe92T/IKKszzdJTz
oiFAjpeoB7fWlgs6ytp57uDCRo9QjElOImiUMXiQg9lqHcAzdfqH5+naQscvy23N
rWv5TJ4IpOLYcSyMNR41C/3/PT1v5ulUmZmbr8JthKgrWP9ojzmWb317vjxZwHnU
rCYYZxll0sMzAy4pTJe4PNFUHVpaa9LnXO12yYf6ctxVZyPXl3DQ5EIT7idl5Cf5
TDM02y4v/2d8h9CAT9VXXD0CvXxkcaEc+t1k9zkOkREU9Q4BOlfvWhn/jwYvIWkE
IVjx2rqoA+pYublsQaUaIIY15UAQF8k3iyi4pp7r9+ayJWlImmRuDrpfGnILmt11
rwoeLW0XVDbnsPfmoro7UjUMGTOlmzH19jg+5tQAx/Vi3bK4jAPE60Hsp0FLWE6x
TRq+mL5thTRS9b0Lbf84HinrUtUKKKINlIFww5soFuiFrNAu0KcPTVNeikN8U+tH
iQ0flfqlRYeHPjYXo4HX+rzKKUvBGJ84fmr32i0N6XaZ7FsHFRnoyDmjQ9sENIVq
qDj1pqMXuc9xqZ/gfSMNcz2i/d3tjUPYhr0zJXFxRsoSp+nlxGjaBWzimrwFzMXe
nLa9NX141MS3lClNIocZfXebOn794majQIAv6GDzliB9lzCmHgCEZAQO5106Ah2W
E4cpheddiJqmx4lA0ytfhh+EODU9LM8h955XV4D2ebIdSFVHm3rmPtb9nZh4TaZi
3jlGnhEWezlQpwg2yjx2SFcPQL8C2w1bJIlekFZRPmUq8w9CDMYhq7FHbjOuXxse
OhEMvkXQjGvROj84oy7oefVyMWr+PO6/gZvolZhQVzJCKYEm4DP1sjsxjHKSah8q
UugRvKusfjrVaqRZQP4a6wyDBHNhZi1pt5LA02i+DN0YN8Ri5d/cTdm/RjO8nhH5
ytYXAYyq/9ap/LkLOvKMgtLgWtmxorcf6R8oe1/pREhVEpmVd4ZARMzWZXyAVRXJ
9QI1iZrtjQRbEwZU4xcpFXPiJ3ikD9qcUykPocMTscPS+uydaRy7woC+p5Z+a+DO
lFxFUZDqWU5MoVYMUpLimw3qRo6Fd+2b/++9g+WOtsOhEInb9XB5+KHu8tKEyRwi
X0agazoLv30iJfZwk/asX0ygvMr3TcOsATo9Bzuj3ODadXzfVMMNpldKhrruMO01
uzp+e882RTbakpTAifYSrkE1HXTQRRtORwH3kWoiokVVKAm+oiNkwfgkPKZU8Quv
Jy+yR4E3ofFhOymWkGhZw4bsdJ8KICnWMkO9NNAGkhy33t4e/HJQGw9VTOl/4vF5
+meSjm7V4u00Q7YHuKD0/xBaencLBNhO233162sUQIqk5TJWsw0ZCY2Ri1CzBHo+
trsR2QYo0wv6W+sVgnne4ZxazZQC5qvAdwj5JPiYjelxp4nSi4ZVi02Dj1wHRwFd
qnEawzAWSaoWAxIiJFVhSMc5Pu6koKkD1ukDJM+A7r0IEKQmmSxC5EYOrZ2qPNv6
dqonR7uT7+LeH3DPIxDBLbeNIWgL36bOB3UhJoh7ugFk+4Pr0vVQy3uyO+TSruZo
/3Z2ExGfAAEztdSgG/ujHflmRYByVzTvrcWMYj6bAYNRxrU5pg1tKRbxtp1k9inp
40qQ+dWuMEGV+UY/rWZ6wWGJoNi2GLlp3m27CgiXmIsk5P/sWSNEkvWszin52xzd
gu7LDKjXUCgVuy8p516fSz1P6Od+MF2HMYfPB9nsda0EurpvBDiHd0VFoZjt+W9/
avhabdbqi/rhxqpfAxGxuwyLMjTew/KjOqm8u5Adu1U2aulMTESG7x8YbCSxFK7/
OGpATFphsaU9FsJCHFocqzeIjAT90ydBPFJhdGFnydMFrG3wZwmxXqCwbRvyHwS+
MLjXRGK3wAQr+bYUpLP38g7oCNTDkG40A2ypqwu1VSy0pdCRJkkn2hJ8nElbDq7e
Pqr3bkpi+GSuWxZDd2VYBlMD3eSGQc01GYlkjQy6x/MBhW6D0FhvqMqx3gcTYguK
m4jR/Akj0aHadoBfPvgCrmbRQMSOK7eVt71kYy+opjfdyXh1KBrd4jpwU2h3HoV8
nKz+BbzpSpepnb0zfKmmQ3pOEM+Os8kyBrPwDCQTeS9B0kXqeKjoVUkkgWk69qfe
GRU/5HZdP/VsbcHUJYMob0NPHk/NZNMgi5M6/0ZjrBA0/AYFv8sLoI/bReRdmmhT
tJ1MoZw330eo3SleElnVd9k4+YlRiRZ7dKJdHjGY/3imI1cUB7U9nqbZxzrYsNDZ
dagjdhXRiPmpHBVyD9BXbX6IngCEFOhIxJelj7YM75Xqfm4aeWBRdYWiQbZjEv3A
usTyLkMUtJ32RSfFcPd7evi4/1f2cquntFi27aKhecWKATHQ28dsDEbgspXGP8mS
CuZpsaBcxVjuFEdLMIX2Wy0U+Cy3cOZs9u2DeGtCf+iB4TqgwkC5QgepgDbPGWfn
ANGv/TDW1s26Wf+FVtZgpjUXF5FC7DNhhI3laOUq0edMi0xenAKENexBswX/aS14
j1pvdB+Pgcf7Hfi9JeZj02PoAG6E3sdY9yWBNHwuK74TVdcYrICPi/bS2x8c5JvJ
GwdKIyQNqqHsY85LNlvF/hLqAHtxsRa+WAUVcHtIv8LqvykbMlkhPpfc/MZOhzDn
XvtIWZgczRzhMKtZHoVJkmds1J5S/I+vGeqZ+9iG4zcfabSLmx3KZ6JJDv40ZQbE
Fm9xnZSZe4aR03B2s54EgGB4Fz6a/DYd8AauMJ5H4PWik3H2ZfgYLeHpthhAmG4+
5fHwWP+t3wSMWWaBKQasI6qSw1s+dfCKkXI7d/NyFAtnCrK3uCZ5vjX7VHhPrnws
JH8YDvijAD5JquKF33eZfNcw2eY48bmJFJzMOPOI8jET9csiFyyNqe5nW3qAYYHA
NlftLn+V68Y0o1w5VcI4M/FiPtyYWenQpt4XwMUaFY1NcmqheNLxvjwmfQjHLG6J
OcrYmY0QdxA+QAnmENO7ktrCurxxzWTPvQ18JAjipd8Andh/QTZ7JsU8AHgpWgQu
8NniH7dQAhrprKZEHffjQp/iHAsaKOZHDeUEmwrVmYWBxBCKn4cmzVXjXaJ3gc3r
5xq05ClF+1fVaF7zmcr/pgidY3w/UKWI9iPAFomhns5fhj4lDLk7p7MzaT2D+/h2
3z9YyuRO1sO6CDdAjLVseVJPKVgPRtHRYd/in98TcdSIp0lwuSNFkW7acQEcHj2i
rJfOaCo4C1yhhkZbQtQLIms7eFhRQIoSAg62u1/8Qw4o8VcWbGMQzH+CUzF3HSnz
bPlfELgL29815UXyr33Q4KDe/c1fdSjyg7/qf6OawXcseVWM8uug0nJ2/rwpYo5J
xnxg4yapSJ3uZZ3x9UJTsAsbrPhC3dESPl7CwsgvfBflpTQY96LXGD0fhHgiu90o
ENadusvR2nn/127/fD3DoY1igBD6INj2NTbgBiib/4yAer5niagPf45fG68CgCEO
6b3kcoPdKEkYyw2wFOGBxj17NZ6gRcJXiw/hYmddk8lm72+uyEKGTaTT5z4oZyum
PjS8u9lIpI2pcXJEuOonIaa/PnwyCFJ0gM/X4TGXLRGEa88VqifVNbFaDmwtsGby
LpxH5Nq8cj+POEHeP3fSg6YoY945GewIeHf3jkzS/dFX8J8iincJ0UnpAuzsEHKX
USdCkO+Qgsm9PEk0Dfx9UeS/urDWmoPe4vQQ+syuU8pIFnB6rfP1IyF9X2lBZwpK
ke7n2jZPmCqbthp3de675Wte/YnbMe4CHOsJI/GKACk1qSVecjlVo4Mx7LUmQPTK
PoXttfx8xcj6/7n4h1SMprqsQrCQjrZxeD/GYsVbVazYwIGYzpzemxGCh/reJBaf
5H95YrB9YllweD8ln+a4gjsMtOx0vjcDtdjVw0z5Z78E61EIyh6MlPoyCrUGpal1
2rFZS4YXJe50lhxwUTLS/eAoK70DvRp+J5eYH/Mh/f+j3N0thVJQfB/ETs0tsNWl
mmEQqJ4xEmw8YUF8pnLyBqmeANiiCsSrdlCpakhHws9DlRLtTcD9/rFWs6S6Vhdp
bvmpxjpJfmNmUnIMhNfph4rl0/VBN927kH7kr0Uh6qkAGHg771JDb2pBXl3+GeY8
V58ShBpCcLsbXX+qcytA7c61i3ptJmRJ61MpVJKpB6vUqEnxFBKRLlv99U9Dn+Aw
YmDZqG45TXyDyYGW4EwD/Xt1yGIarVcrvhTOm5ZXFk3wTl2RGj/86t3Pwyae4q/q
GEwAnjn0+PwrTi+r3bP0gIOif79W4egTLi3SfkrwfbhJRV32VKeXogxAThrNpAVu
95JaYKQRiIssXpjaUkCkEAQyg+VuCXKmorUN4LrUv7jIrg6OmqMmdYj0hgW2LpGH
EzwtQbKZ3JsaKt2r3HZ3SFh7xsWZUAZ88NZuP1PJg0THXJYKEd+Y4+V8CcT/LbgI
KkNaJ96TA7ZKAb5240AV3Z18yL5we98//p0CB0FkNMRWRfoMuYJXPMy0nR/RRB7v
6IOYE0iBZTEpA4eXGlS0DlTu5BXQD/RL5s1J3EbcKz2uODfZh+snnEagSkcHd3ym
3Pc0BBBVp5suKNqlp28qDXYp9JqrBAHeGwH3If7E5tLISbTUosc+dWBlfAr3GMbG
5HCT4ZITdizDdqZKXdAljm5akejegK0wwkSVWiYbEswHzw+qYJt4XKcflJHkx72M
6DBtz7Op0DBvhag2GLn92nO0xUbShJGRvFAy2IHEZJGnD9+sx0nDTYHu0QTJ52uW
N9yiA/L6ASoBjl1ICNzPexpPqFsMUhX/GwhKCaRbxFasYMkTE+Hn83DnLW2X8GMo
6r21my3Ao5r+IPB01dsoG7H2kDTSmu4a25OremFd0nuO6j0SeGIvyq8xYE6qj0P6
jNZr1nh3OF8CH+dP9nMkVhzwaYOJcxWYKn0+QFTOrTOiJ9/++gPVfdhTXWi0wRsj
0BziCk9W8zalAejNf85bwKb1pzhR1d56o4lf1+49MBalvNT/Q4FTh0ksWB3obfmm
vvJ4n1P1pfbDhH3iTnoWqvWPNC38alIlHvpxosUaJSbfZR9J+BrBF6ZQV9ZXT5bQ
I6bVtZ/0NcSjfmpAr8Amnzga5BBAomj1PRPYBIzNKnEqW9rtIlw78X6RhUPjamB2
uS/hMWAtHQcmWebLb9gTbktBzjB1psRKJ/r9AQLMRZ/ydO/LooFoCaFVyOE0OyCP
372TLCVXHUUBPC8xOVsiBt4D+uGKnJbLCkNBXP9NvgJAe63xYHs/DUnMAVIKFJwQ
j2di7hON5dqx9WGD3ZzYLYCzZZq1fAn+QSwvQY7pF5Zl4OD49/PgijMbhOScsQhk
MtypvYJa0qIUvrmBOUT27CkWLPAXa6X5yRvPZeXYYY2Ze22aiEX97JxeJ2T7YN/T
KKlERefDAYFf+/mvYYFx++e+jJXZSgw4i6XsUN+sWD4Zra/4xPZic40tb+JuHgCS
CE4HUoZHE8o6t26pWfl69aHjNZZSdj59zEHdcXv4oMapgDhoW/kYdnasa5mXRVUQ
ENGI7h7w/h5gTfUoP2aZRmPO9mRMcuhJ8i2k6uXWIgIXM7aJDxyUfo9/6N7mwceB
5CCeCKalIjoN36cMwmMm5RFet25jftzCpUFk91ccpcfdSY+N0Ca7dYdTFig6xwIY
vwC2CpNDigQiJsAuFGBN6GpXFwPSOMtXNzJTchMD+2SXS9Gd7fU0awnYi1c81lWB
ZKAFeFiXVaUEQzYq5+miVW/A38j8PaMiMMRzvijm5/eM+5hPQjMlCxBfnbnVyI3y
tE+UVvuQwn412R0XhZClPN5c1BznoF8gWZCX8o2iiQc+ZTG+btLJth9iw6KJ5ORu
d46+QoEwlQdD466t1HDqE7j9HUsXDoRPoG2fMd6PwAnqzHeor69PW7rl5zkS1wb6
lEVy6wSVUfV/ECyv0n9m3DcDM3KpYQyprkTZ7e6J6lJ4A1p0zSsRpfjIt6r4lZLu
DyAjjK+ptMiNNX5edd/AYM4iGo8eG1HwU46mS8HJrQ2jMJlcFz/QByH3PwQSDdSA
85U3Vh14aRVLKmmrOB9P3frajmXF3b/71DEW1508wpCZHNhQL0ge+PILkt4nu9Do
2/jf7mvCeeb6p9i7USaHqjVTklMYTkZ/8ZhDddoI+s/84WjP+bw+vvSLfQ3EHyP1
OkrYH5tpoie0Ecf1zRK9cWR9Y6eW+XnqMTmcYjkXrd42r4VCY/38hFsSFSd5FxKd
oECGBk1Ct8nDzLMaa6FJc27mykQFnVnpQNF4qhhxk++sCXAzH1ANkI+TKlgJalmP
pHZ5hw8EUWIjwqZDgRTbKRIEhLrk2kAY/Hl+rmQlXXDLCcqKuv3IQDFGZ/0VItav
aiwuzPIqRFde4tUwr6dLAbrLDX0q1eu9ZXW6Rotfk1Tic0KkaM57+lBgOKTKvvW+
SShrO7vwWIHsomqbY01/Te2hnXSqFm/VKHUq4YNHc/gnI2RnFAa0yNleiT87ePnt
3cT9FgaTbIRy0vR8HOly5IU6fqICsXt6hq0iBsSMK3qcSHsozmrt9Q0AecZG2H2A
+tFjyOQxxphO5xndnfYmGV2RMISpfKREm0BOLvUXmYXPalId8IK2vAakdxwvfYH8
Vc5BOZCPgMDAP1P+d3/x+7jKg4w1mk+cF91moD3xusG33klcYpM3sITUitvX7lE4
U6XX6yO/bmdMGdEcqTvtx6mZcSeCSdPC4I+x8DrO7ndV+71qXUfg/MNiq+Ue5Vp8
qCJ6itZS0pJgOm0V5dt3pwerEQgAUnjs2BvWE37RjaQelov3WpEWgKecixcY/dHQ
XomDEI+NkvJQfjZV4aGm/g67kdqHURzCtmHBghOeTt3tOgYOykkn2ESJoYLM1MWq
s+yfemMwcpU4JbsbZ1CKpS3Bx/vNECC1weh6nOfxjj6HZybcFTo5PYPmpnEkzRZk
wF5QBzKzJFMGdLnPFHbUeU6yI6aKzwWhV7Xzwa+HA8SU/tX9inM4J3Boy6mzFpwT
EmrIKXLZF6pvdTVpPi4HSM9THqoNy8Heoxhj05qGXrBkx91SL/O9TzzfVwtgIYS5
vthLy82PHV+pfvijHfEeiMLn30kCTJDHDBlvFL1qaDJGKjRVoBmRbiWRMBcU9xcP
CddEwq3Qvmm+ellrMT3U8ozNRRU0vFCPhagI7rd3SwqmXjZr9d/5QC6xIA6mOaGW
UFe2zi3CjjYWR7eGW9uNu7hLvC84AdOXvxCSr8fJ7sTQgJ1CnV5E9TAdZBwAlXaZ
CN/pD+b0F2G0PtkE0cIceLuLFJqxqpKGlVjtkibeED25Lmq0QvpxAszxSYUX0skc
OVpsgKYYFORaNKbX1dwtEGJ6fOYAj7qbCpmb/GM3XECw3e30oywKeCO4tfHSeVj8
uloeKYthlwnG7zXmbW/Gkre28Su91RioqbAjCHJpGqxPyPDnQOWyiKhPSUnJcPbf
QAE3/YOsz1ujMw+UVWVqEhEewk7uv5EeZK0Fr8LXhDlW5fiZoFaDOD7BOzopJC16
oNxiciiMXz3Blcde//CLpNaRvWOYD/OI1OtWmOgmS6JVp9GXQJUHJL27lnbv3gZa
wBtVS/S8i51nvbcSxdSFgk1ME9XPEMmKW17JQACaolc2Qgyi8xZjDvKx4z0iRB/o
yl+5qd1vbEaB7s8Vs5BeDCrIen/qdYjgtxZ7inAqHqUOcbuTeWDBD/HKYeGsCIx0
jxentSecG3jNZ+WTRDejVUhc03Jli7KdyyCXa9TfIl1Hv3hCCUOQOhtyevl03Wq4
AgyxgCirPPHl+qRb8hDvoUcNO4r3m3oH0dEFM+QZjV/MyPRpLB0r37cpZA8FQoAS
QQV27XelF9a1jQguLbrv6LceXvlgx78PQbo2YgZRvBaWwVOT6coQK6s0Wf9yhf7h
AmFrSmJU6br+H8A5HB7RgbUQYg3sv2kyU8NSFoPwFE69GjOlMuuhv+u7D+ZmiJiA
Y6r+FxxxWZY/nLlXRdIDZCbwH6iqBV++5HHiNT40CAXOrUrKJpcVOHU/Dq/EeLUY
kZU4wZ9jJFqDpO7QTfAiMWFhv9GP0LGet/KFglbaTCcrOzsiGvfMkKg7n711sP62
s2v6cHzMg0YKX20mlZepJA5sll6zxoawMIKR12zc9hTy1M5CAfhPZHqmcMR1T5+D
kDZcyNP05/dIpqsmI93KRwhjr6J7wyMogEvQfZL/YGloI1D1cdGMGDNH6ZUTV93d
RpPjpGMdpIOodMLqw48oznqVPZz1fpZBjNGPOQwjjrnB4vCaYoWSchV31lD/sXJb
BIzEzltp61e6AlxjP2yV717MT+lRcwdKidMZtoV3QpZS9Z+Zcim9bAozQM66Kxqs
qwjPqz6YKagnDz40ZzMBYe6HDkh4inmeBRPo+BNdgpBjFUE6cklqrDspjwpf78MN
EqbBXqvYg2EBVNhfG0ip5fCPlObGshzjHONbnl13nGoplnrb4gJtnJeSP/ljlP9i
espWq51dTyFmFI/afpImYfN8cbIabkhEZnxGnaE4coiuI8dzx2XzM+S9FhHTbftA
/JDScie41nqb6SqGHxYe7n0DXecGzbQgrFf3eWYg2h/AQQIndU3kB4PzAQsgUtLP
aEN8IKsemTxi9YUYQJfD3BiP/hDTL8Is6sAKZHa9ojcjeSSSns3x+IdPXI+GiPOx
28AUEGi8B4+lCicqh5LamyJxoguDFOOSbOIRXdsq9QsPH5b6mWnVSaDqRIyHuLRn
LkYftWzHU6fxIvfbx05UjjQwhbcCLNyNUQZj4Icq5ntqqW7qteVfEGjmoun7yAsD
Hjmv+mtUyNVu1H9u1LtMVtpjnuoTaTwuIU8WGaI75yhC2zjQ9SFvJhnPMEG6H3gz
FU6FYl8NzteK900Ttrr7XHTSAeEcJPPMz2pHaL9ueA36elDW5mveGKufEBJAib+K
hmozdku2wiO/FaCKtvFTtuJboNGsOdmkOOVZPlIODx5cn/M4NSM7WfDP5XHj+dfO
rOaWbblglwlLgF3owNK4s0lEOCyeLD4rOSRW704gAfEJeHArEHzsjlEBo48FT95P
0qXhUWvKgxQSW+9DLH+BTS/b5937iYD3rWfVlI2bv2qP2lKM0qwtoK9bXld1zuAk
gJzDT2rzzl5eCbL1y5STiql74HIjuDGsEhTtDUGU3DhUr2KHILAGEsXjI59uZNxm
kloL3ZS8vLAz2yPn0JBmlece3Mbfh8bcAQdpPvbfHtAwoOmPOQcH/XjfmiJe9qdp
eyRQjFXKyr43vlKRyZc5PtmC3+FU0YZ10xPsFJ4mrbm4yPTKYnB+H0RQVtf75pEw
wjNwuhaNKRBGAgJepR7q1UP+LWyAYhzTjpDmQCPNiIjt0xJEHBjfjRlgp5TCHzge
mQrsa5ZlAYZewdk0vSj6OQm+qfXP/z6tVZk3V7xcWUA068lMENxFzHL52G8vTosv
FYW5zWTBn27rQ7eCErgvYRUFTmKVC54DdcRYIoWdP4PjYf59TbBFCoClhTdwhp17
swl3QKoJa11YTWOF3gTqMNim6I4J951u8qdI9t8DhAFaxRxmj1N5Lccv8jb4YqTi
xN3SJA6sRyFFd0xk3X21TqBgLVwrUIFdtTdCuN44wJh7RDjN0DHrXEcfbleJ0hDm
DEtZhFoYosKbN5qF3c5FZUjQqQxkRRN/epQesSKqWPpC6YCmMmOwI4YA6gGTsSIc
i5Y2z1QqPtQpN0gJXIwKgJVuATzWN7+zUbxCqxCL/Yv9/4FiB/QsGyZV+XzGNKar
IBhAZRiB3DdFW2ReOb0SysP4Fp++F9NKkt8jLyPHX27S+8VD2dk175mAd6vimjg6
835mlf590BRKEaHdGVUFXfLz81aYLv7qf2N7kgnc4LIA1itRuRcl6O0jtuST24N7
4towIkoP+pETnb+eL6Tn0FNA2UbCCNqwnJ3d6AtURy73eFdl31w0y7bXgDvfttsT
7JmqCNCe0zpY+l/1wPR1dXMBxAv1D8Z3GFt+5E/bfaxNQAbI3T1UUtNAuHvi5dYx
53h3QDr7COgiXAEmSQsqfAwA+JCEImsLcFhPVBBL8vf/2WQZGVY5QZDxcCImPREl
fBUKrWOmQAmaUNNx/NTKe6ZIa2HQBa5QNYfJYzqZ92gTUMa4iRzYJg/LBqZ7IFmh
CwHV3CDQiZRh8BsNcmfpT8iz8RGqr/BrlGBOLBomcFVGiq7dheMbXIgRycOhh74A
zy/qqGR/BABfCyk1EkLXdso+xeY5bEa9DOBpjsKApjKPLcWj9JKEll8CIOYjd2aK
7/bjqM8SAsR0Fex0Y/mcm/9wMZg+9olp91m2HRM46MNIMi829sLHQAiWH7lNJ0A5
sF40EJzBxgxj0kE52GlOSflCZ2JVSrXfFROBR/doksRcZJZr/64J/RDXcJkjpPvg
jkybj4yVt2yqSWrsDpmcjfkfYHzLjPepcsjFYDw2QAwxoQaZS63g7288ElntVowM
iJrfx3CAutCrtmb7uXEAAcXdoc75PPzXQAg8sMD7Ec0hM1vvhpWS0DU1Vm1B7WD3
SuTk4Ptqpwt76GD6jx3l8DA7hQkTUB66XZu1HyYY6UHZMSGai6oYI1lr/BCkF8jZ
4DpSpVsE77qeTlbs9bxzfsooCmSVWW63pRnSc8epLcWq4ZIFjAkHLApOBfOGDte1
Q7MuQ54ypi7lSVuE4obR2F7ddsOz8LQhAUc5d37ubZ2oR6UwBkIRgbTyACMEKKi1
5wsNVH9WcwRsplOaknv+Zuar4jDZNZBrTAc0r85OZ6zWlMrULkJA3HH1ZyYlTwvh
tPgHRnSmzqB6RAwZyCNQ+aXz99mD/JrMKS+Na5RrVPwCROI0CqRalDJ+eOGBqGGV
U6zqKXel8hn/0SQfhYZkSY7ELbFLOIrMp5h+MGfBjeNeJLH4zMc7eKja26Zib77t
R+Iz6QJtR9LDSHeLW+eGXBRKEBLtK+NDutqegS97EBeQ1LEYF3ulL4TSkcmu9cEI
XIWU192roqVWeMBTkemzfRBqHL4vxuzoMqc392zg2u3TplMvj5zwoi0eUOCaYZKX
fsyxtDyQDBzJ1GCBakF1gaSU1b1zMqn93Hl7qtomGXI/rs4aqAaXfs5SrjsLr57+
uMTtAg7lyncrev9jktySjehRBusy57BLBp5ABUzNDytQ8ExqikXWmpoSw1Mx7cTB
NlsGCTSkQkjVg04os5hBNTzcwft1SrPrGCyyF5jHc/Bv+fMkze1p3IuqKhvxwqzA
CZ9es/g56fDpt9Sf7N3FudFwebygM/QgKvYcDFNqaeavrI+jHaSTVYtS5pHBvc/v
kfvIg7Zzt9zUTPbjIKyTHWxmke0Z/1ju2SBESdRDvtKCm+ZkDCl1uRuzk9s9Trrx
q9k4r5oE0QS1z11EOgW5vNoGXoyCwB5b3CJrMJs25HAQ6cZ7Nz/jW8sXoq+8DVU4
SUa/iRi1eKLYMchnk9Mwk+jdxkkcyrJCU1xUKE0m0BYfORM09IhsLIe8ZaOucrUF
oh4tbJLqjW5Qz7/+hZhOsvw16bn3Ll0w9eeTAe/FvfOzikvnedQP4W6Ck3RecuAz
0LwP7V/khtVo6yCa3FaYohMzLvWsZu0rYjmS+CKBi5UigAiT4fF2q5Pm4EumYEfD
S1Bm/P5iCSbCxzDAFlp32ThY/CzDlJ5KArj6NddjaBRNpJ8B7AfIwVyRhOj4EsUI
xU3fx47MRMx2OFFxtoKBL1yfFID/2DPVFuYWXg+VnrSO++eweMUgKoeGiPx8M6PC
pkvZNNAlZnij0e29byEH5w2baltqb8Yn/MkQOlWjA6IA9mukbs2dSuexKcoHkizP
hpqNUu9KqYgVHy6EBONvkwhmYnzYL9yRt5kB4b9PZ0D7IAoRlEjkAkDIiXS0czav
E2bvElny0cG35ihetotg4JbaeXsqiiPqgjJzsBX4OJLsOLRGXj00lKyRgzTlA4gT
rHvkS3TnfQrDF7Ses5pMvPcQlNdt/iR5/T527tpqSxK8QXRgKCywNdNIQ3gGewY2
lapfwEt8+craYmUImy1JrXzS9DqiEFrqDN4udCVrC9QI7RbQL2JBJprtWSX9lSc2
u5zujG0rB9070FGrvH/7ga3cF84N1tkGf6YhMN5+AllCB909+BfdYM/hQ4Ko7XK/
tHmJmLcO5B0846CWvyNO3ZN8MlflfpjJ0r8Ub9c25SYT6gFc4Zme8ViqRPr0WMnq
CurZ/ia/fp73T/xgODRCWelphWWBc+g18GlcYS+mvd3VPO2Z7MjzFePoalZWRkHX
yXsXLjvQRJH6jbulwY4uoSan5jvm6k33AMQrFVQM4PyUQoqpkB87nSdiqAIhPyuh
kBnSSJqGTpnnErSXQTr0+Yy/mEjczjhx2QHxA3hlzdrZ2/B4MQY+93E4dz98MPUt
OozwO4djNoSTFeknU36wkF1CHVHqrRP8/T42+pICydAHwaCvXmilv1D214dRknnA
XstkXIQXDGdqwzH6cWmVf1+qUZnAs/1SK4MEceQj2zWdSjadSv7Gfz4hufCNjfN5
74B4/cR7aDkB7shkltMAWTOM2HjEwF815aa1+ZE+4UWh6gRy9YOol71H5VfVcTj5
WA2KOfzUAuP9ruGam9op7kkbnX9d5Wtun7Xq9HkYOfGJ44P9NoorhASF3V7Fizvf
3fsBv4AEJP6HLoQyXsQRq3Uo44k7G2jxdq6bC5j5PUqzboa2p8ckf/EcEXBxethV
Jo2S/WQ+uBkmy2Xq5J+XZIEJMJqrVMG6hQ7rU697Y2nIeXX1pgm1CiSUKe1Who0N
nEcVGNlXTYt/F7ViOkw8JaL22NJr9FQ20lK9fv2QTTDvf5MHeCWnB8OSa71qmabj
TEht8gAl1VNMSlXv9lp+t7nlvTC64QdPgbQp/Ij1/VAWAJhqX1kwAPpERCbaRWZq
YLxgep3H+4YXzz3T0U32QWVQojOp1mX74OwYvD+Nz3zQQ/KEw6t1ZtAf/99BU/0m
jRSKjfwgAbcBtmwDE1HaqbrxSXr/GZjohz8/DOWNhVzD8B2LUOCALH6ii19bJj1w
xMvQD9PjNPeZBg4Zv4EpmEy9BqjWUMLE6v1usjqbDvvQMRnpdqA/inydVfIHcuWo
vgRqX/841mtP6JKQTIMmwJWWtHT23+eICaOII8ZzretfK9RWD2ClpvzT6R4Bnyfz
9O5rZncQmtwaKv/U1cKmCI+IUo/x8jUH3qlEG4kvgrEVEckGBW/MQrF1yATFChDm
jU+IVuc1wOC/ak/Rhq9H9G5IaLQHTFdD5v7MjpWs1bjbU6Cya0xWyr35GDcretqn
TOZcqeaiLSwq/SjIWg5NQEns/2NqRGsNL5Z49QziJlplB7bRLDf5m+BngEdwbelH
MTr9L/ufEVzNX9bpqE766zG7O/L4bbF3hJDC+Yn/CjJJTw5GTHZNx57kPsYqrr9S
N7q9WVRmJPmRv2dzM/ACYrLsqa/VNKRAGvuuBeUO85BgZ65QjZ+xXYn75dYWggJA
fhufHLoFepLuE4uDbU47CqwZmChq7RztkN2izujlNqLyyGdR+OejjDZlXJ8VGZW5
IB6fkZfEVvL375xuHmtJeWyUcNFnsW4rWi4uwplEBorIl10O7E+UTv09pCl3AyAC
T3Uxq6tjNLfvgsMpWXVCNWh2AXC8S3XWj1GLMmdRpmK3P9/sAnQ3ieil8Ej8wcTU
1xu13ztzI2j6kIKVzCy19/w5cSB1mhY9FH4Ewx1J2Ymozf5FWA6X3Ccs9Mr5icay
LOJdgdRX6dJXxiJvHOpi3RAp+wQ1OFMKRjL4xYdfAvugrrOo24jKNe7kmep8QmDx
mo/8Rb3MxWEYFh36r3U8e2lCJnNAsId52FwPWrIWA14yYimDI4uM6+2M4Q02viJR
jcHZ/j/ArqarvrB1XhS8Z45BOgiRsyDp9zfmndEAQ9BXevewiOUW+Hphx4i07C4R
O2PymtH7/A0Y+I9MwCw3x2AtM7j/EEcvSzPnGrIJ4e19/3MLsWVrmkCa1x9D72KR
xWeCmU3O7g1/6YxObTzB9RkLI914bLv53+HEZOJF5T7xu1lAbqPNIEEqYrmey41q
5m0kEDTu7B30/1jHkHNB2c0clr1Qf0T8mhFPQaqpGTDh07LcJDLKXeYygf61WcUD
tqnJBKCSwyyURhc08m+QNaFj0SHX0ibJvRk5ykQrZBACjJdJQtwby9G5MK6zLuln
cxz6JdXv0thfT+HbLJL98+VQaTZyt8d9vE4CbHLMHDPJQgNuqw3NCGySQb3Moano
higg6z3FyhGB2i368jGM1XJXh/5hNTxP3J1/+UFpkEvicfSDIBDItNPCQVQfKbsa
ydD8mEc2pUxk0+UHlbCZvKqFx3yCNYd9DyLqupeTO43ULTCAu1zjvD6tEXwu/dS2
lCo5Z4LW4IiPv88LO/D4A61MCxymNMAGr595ZmM3iWVwxT9POPY7LmnQ9AJ3yhuF
zqq/J3qKa4vrYMAzZmrwa8B5vs9iHlwFs8cHkqhXQ6AHgCjV7C94WIwjEClW3fYn
GVXQJTRDXiP3L+kFegko8Gvx30gdn8b2YD+wROlDA/tPNlWgS4b0C7SgZepCpLUr
awL8gADQT4SW9m0hZEyCyc3UWbE1p9wgdMe7lONyal85/MRxLkI0rVwmqIEWWnQw
QIhrnMZAbdAHZeF0V6Yofn9IFdYT+Ct0/ChEjEwO+icdUQMzgj1rxXYUjDq6H0wc
Gvw8XkUzv1VFmtebHDBlQdTMQhUhK7yfS9qFCrRCE23PIKEmUVUagpJnUP0P4T6H
pKMvVYqVmMq9ip+Hbl2zFFYv8ocD69t/F67UJZHtCsuxgYM4jUEfcI8Tt2Skz55/
IPrWhgW1h4ZQGzZydQ0EMCUU9QhJr3NC/klOb4D34jlWvJUaEuAJ8UNYaNnceT4R
0QrfU9KF3cLuxyS7k21dUQNbStJyiOKB9qGytTyRb4AQwKG4F2XN1E/VEnB0PtoG
EmAshg5sQyPvkVuxhSfJdpVZ8tY0AQ0l9yn1D54c4Wtg0mW1qDAzZVthKGR6jxnk
UXIRsjV866M/9c/9k+v5hKczbjIgjR+Er6sQTk3ZQm7HYu8xLusjAA996gRqUucK
/rlzol4J8+Kd1cZk4jx+RePNz2qZUadhSBXpxbi/dQSm0SxuRIUVOvG+qz3G+++g
8oT+RpV9PISmjRtj8nsROm9Hzeg9GmNrbqnGGxftsAd86c0QUZU2cc39b1izX92b
mq9YJ03PUQ4nM78o+ODLrHFO0xhrrlbf0ZDheWNY4aa2ul69ef7tZx1NKBDaKJnz
e+vUB4Rz/zwZLUThBEJZ0nthlv715QHqTePx2Wq0w4oYBM/ALworkh7PUryspgds
20LZnnikN0ker1phq9SD7JiSxS0c1Ueb0ir8r0/m+1Doa0fkBOA9zY4NdL556aPs
9m9gMOgQNwYFnyBKClfULNS8mKqeEIH9MLInc3HChx2iA8sa1leey2K4By0W/o8e
it6ueS9c0JyOfYIMy+6P0ayPsvvVb+mar/ckZYbEqW6JSPv0YQ8UnEK1XMqhqMeL
0bcBOTaUoIHkUR0pBFO4IR3/YSHhSTwwsOML4mkhSky098ySbWuHw+yAhFuqqmm0
mRhezyvaIVaIoCjjw5HiDifk9uBhXeiDQMGzU+6vXXRPGv2UH06leadN9mUkWnw4
yqvRcZ+vHvPLvZFzX/qxpdBYIYUuGthMGk0zI09Gfzp0V3q+xunSI2Yr+cZ2Li0O
0FIvB6bu3rwkbrrZ/eG45j6Oq6DQZkWECmTlgMNMyKPFCVK8XPTBHvPyQIW2EJ1a
tfq8pfq1HZCl42c4ayetv/o4qzqgmVL0uiSIeA0i44zxf45taJHIaeZL+vo0hzUS
V3fkj+PR+FM3HzkDI9IVdtC/Wr2qjFLYNni3YhJyXt+40Ef3m7NhBaJECmVTSPjk
ic1jAiErW3qBwqPBbce8yZ46eJRGuSojbcQWZs7UK2xhyOS3BlhiaPVIFcjJMgmC
MJCej7UYTgeniKODUnDEENYcck+Oiys3I3urGEea6nPmiwfCIr84SAxwJJ4OMYz3
7W2fwtzxzAy/nWxuknF0uTkoRZaAioJ+7F4p1xyOeatSQFJYxtLectYXWOf3nOE6
CCJo5Z2ARNG6cdhEtxrvM0dPLE7fNcnqm6RF16rd3d2c36D6N6kN+HdziexgNYrO
nCA4Askaxk+I+hNBZIsOZfrvIbiZW3+LNhrogNBlolct/28XksJubJLCEfTh+POQ
nTl1HLTsP1UiqkgyAyV5sjy8BNv/qhcYk+KzrTbsnwiP/RIFEE4VFmIjQMXWfgiE
3aUbObWnP/4MtF1aOGqXG7rCUI52igi7aY9r7ATHxJhKAPfbP8fqhrlqSAy6WDOJ
yqvYK/9Jq7NmsvcVQQBsxBw+3gb6H6RI6VfpUK4/URGkPlx1Bqs5qk4QjBfHsBGJ
fyzYkx14ui18Vf3np+XrAzT/2d5vK7SeGs6QBifVfg+hsUz4drNevtRIM7/jJUo8
t67LGIHnzFLbgP/nlPWSTErXqpBmwe+7IEor4XJtoLkKDP2b6nvd9YTQEh33hiUc
f0yh3lcUy6q/+Z48uFNzHqGNaGw6kRLnkNXgTeAFPW2N8fnMhLm2Qcge2bATKOP1
aCFsYn0TY957SsLNjfWsLVfVEoqnEFJMm7FyVfLUMtDbLR4OH9XCV6Fkeak7XsuB
dh87x8Tb06nxcyKwOsBBWSpyhaiU47KpEOZeucsSAZcpupAqfAvnO/5pUv9o64E+
U/SSJSxxaBrc2vErQGAU8+IW7lemlJh59IHbkxlvarryWJ2tfpITZZtGmMxK99BN
Va8ESGc2NAJiqAsvGJBVoSVuu5h5xIisf6o5BcXBuRKC0N7Rv4ipWDlARaZTU06h
S4R+lBWeB51MOXCA6cnQ1uB6lqoOV8xu06V5bt4lMq2/SomWlpGZF/OdgozoZsUv
K4tfxR9IleB3UetRXOqR1912ue/hc4TmwNXIXx7vRwi+pq/ivlYz1ZNzSHpwVPui
TmZmodeOsUA1s3zbUtYRnZHOXKZuvzo7c7w+4TdvtSQ5TF0pyqxt282khOq34+Fx
p1ee7qHL/B7Ctz0m5zQPy9DkQ4stIwjJ7T2w57pSyLWahDG54AuY0l4audjDjYds
HnAHoKm2RblyjLwjUJuyu2DDr5pKRYLc5NZkpBCGcQKQY+5EIarKaJCdOEV1kM8S
jBMhAoZNxuBBxuYlaTx3/1e3tYIhqaDGBQI70HiJdqni68VYkwNrtklw6LE0SpYd
0XgQNr+AtyOMT7szvPcyAPJvnwIapxZFkeiJe6KOK7Xu+pmxzAUO0PP56Zj/dfsj
div16gSYWy/SBzCJoTcqwkadhcUFbvEZrH+Qex4TtCxbWx9tDv/9kj3gYQKxIZdU
Vk844dhlCK6Bj+2AylIWRzgaAqmWkH19cAaJfU+prEW5tfX6zk5b4osNORe2q7/e
vuu1CETHwTv0UAg//6HCV2zebt9VXWnxM3VTXgzU8nG6/31dG/EWx8/U8IvkHgUS
dIOHCcP0mEwMtCwsxAIMTnec5ENAK8KV8dvU7UfUxnQiHcD5Ext+sgdmw9ZIX0X2
HXuS2KZ82O7gX1AraPiGmi40FoY3LqueGpeGJKMGLUQD2CSMxxCJaV62F+IQpw8h
DkDGMi7hl88bTlmsWxIT4sw46xqMmPAHF2TwwyXHC7VMgvT/iml1nNepS/YuYnqd
TQUL/UDXSBgGa2fSncBA8C187UvhaO6OUrbKOLnJWP1zvnJSCWwGWgI89mqDQQqG
Lh4tVZqD1Q6KstOgsOOWWZUVc5y0Uibke48tbR+5zrB5i9KEYvr4HPCcXFkAT5sA
jTOLtx7DEzcSGKrfqE8BcOc/DgTeiEyLJS4TTmJHsCh9/SznOvD3xYfTstTI5uA7
WMcC11E6L467FyUm97celIGvYSDdkWAbiKK7wxizKOmMfDLJj9ovA666b2h98BBy
dQXk76Y0syt63gTYHAmJhv7KMV5wA/FceKcPUl+q63xHxJ0EiUjjxNInw4Moxz+j
B7MW36gSvHrDnMtrorlIhu46FLNx2ejwadEjTkT5ujr8OYSZqXaHwS15um3o95y2
Ebqmxx7RBCT/sQlO/8bFlrfwbVFN8FOvnRs/mGIysLPRGIFaj7T3m+OvdzwdzsxS
VPrai7kz51lBYLBny0XLuPYdDTHXoZYSsnaOY5H9v9dOK4C9VZD6xAQLv5iHgDbl
aQBdNnV8R7CmbX1udz0AACRbZmC6eyIIYRQNaV/PfPilFdHHOiKdq5d8ubp8KIVi
CeuCXkeiRx1CFIW1iQ1wzMoYiy1AJ1FNwW63qfrgTx1e+1+A3WXtglH40nmBFEtV
yy8FDiw1FZK8Tx9DCY4F+5u4h8S2wnZkCIhqay5lHobSGEK+7WrGX985Ou1s68Fj
5oQ+FYSKD7W3yi5ArtaUte2sfPnt09/NP2q8FmaTGCZC14tmAEelT7OxKqVb5fBS
ne9GDAtnlszESuk2yuIKvlMM+WrCeh1VWd7/iDy98C/WpiVJrSmWllBC+4V0PSR2
YksC3pIro3my5bI3mLRsKWd5VzOAI3Rj37nglblVQ7e2iQFXcu2xpioD0C53P6jF
rI0nZqJUiaKXCBz7rY+UO0nH3bivcEz1n9M9mnup0ZruNpFRoIRbzlk02wA4RFf8
ojI5o2LUGeJLHLWtihNbkryVRIJOLqWQBt7ZjOfkXEUuHEayYo/x2/7CtdIoD6rt
zJ0UAMHHnIOvkdieH3Cutv6lH2PO5R6a/1Dv+k7+f690hqqzzoXY/gzysdoNpNog
8WDVo2zuE4cARs4GupGskOZZXgLuyMzQIWWoPlaIHrHKNsoL7oR3///M+0TsbN5i
HjP86dJKJjnS5IG3C8dcZXH+cq9RH8obM6r/0jzuej8FJfB6ziHQJWYMYEFpx3Dj
LbsgDmzAVqbLJ+qPGCIO/QbFrc4kcKckOh+66Dcu2b1wzWbnT+H+IZNG714vyae6
aZWiNn/3YIHWTlhuvJc4snh5/35CQdEMigBtdrawRJZQELLoM3T9vPySEP2iFdlr
7ke240SGaId0rmMd59GvKAy/KphLxR5vfYCkXIddhoI0hqoWz3j4OcYIlAvHtBAM
Y03fYCg3BmUlOYyWjUIUVv8iSIkxnjycW6gYWDJU27ALEPxZFWjQAklythzP9/Uu
UNJL+M1DtpukBQc0RpL8+/Txp7sJvzv2rwHRcPFfOgCEp03VcWsXblA8eZ49DFf4
UE5zpEbaYr+fC+oqBCmiw53LXYOuHbSHPMyP+iwVvoFTlXtPlwU3htHO4Mol3szD
XElUs0g9MNLQZJKimB4lti9pJxSb0+pav+7idpXsp0ysnOWwc2E7cHiMzJdVi1bo
BJ90Hf3vRwoPsJEX2N35utMig8p/aD2dhvT8aFp4wYq9ND2qTcNsLyhfHhGFvfud
V/GT8OLxFPy8BE2yqKgkiCntdlr2tnjAgV7yeMkCHC3yxL5NYhRQLIVId0nCBtoI
fumaEpHoHIQ4kWs7KlvCRlnQFAOnTuCk8neoz/RdnwhZriovYPiPV+z27lxq6OsJ
AkCarM+erZ98a/ZPz3y/V51Zmbrqc+6NEjruf29Euf5DoAVpZbiiYqsuUHT1yYMK
3XUX2D53KsIjxIqw7Dxgjs1oqUWpUuOXjWkkKvQPHwNhklwAhkNirtDAveE+Su9h
hu+2qxHiiFvFYW4aZ+dBA/0jVkKY/h9IaqGkhznsvGlqccfD902l9uMsoplEAJl5
MKeI+2sXLF79hQsfZmQymUIClDcAsXQJmREAiRDL6f/1dBEcRH8MHsY/MoqjbJHS
SBj198VnOLOUwgehvpI4odW3jfCOddhCmgczY3cRykv2JnXN4IdhEHK6GbW2+NkA
azs6QENu6os6zINcqtckE7TjRk6Ush+nV8KMFu1mJxZFVO/wcApxqk3s6t0lP1oY
9gM+3mejXYn7lW1z63vmc6sf+fXXruk0GdsSTkFU4HbIA03N6PNfGf3GgO6U4Ofl
8AAOhPULcsty6azkYxy5nuR3FcXF38yLzUGZLMsLX8Ex42FVNNBYQzqPpEWD8JRN
rdgr+dv3CvNX7JEcmb/EokD1brEh1GDr8LSVKX7PBStJ+6+Y2kmv7FQAIT/tI55e
PMJzrc/jrLPp0N5HcqxRByroYgbt1UHVjArORmZ7lXXS6HfJDN9r4xC/ncq2ilNF
Whvfa86ItN2wkyM9IIcpBsMcSblF2GKkjOa6r3lzaSKSXOtoYXUSCPC6k/Ry2S5d
orckDnya63RP2naut2urOI8MAJbihnfGBjNJRYdldtnjGaKTrFMwdIi5hJ4yMmug
2kELqAilOXStwBdlbGNSRDWo4fIzz4Xx8cgG5TMB1kbNtDEPfp7Z4Q7vhJTsDD5U
OKAuhq5Uz88loKqA9PU5oBLPo48n4OEyyEoC6CTLIN2eSeQrXE+KTalg7mOQseHV
xNjjw4gY07Nn4DCpn8l57tnCPCAIVcpO/zQvmZxLn8DzDApr/2+KyY9Pj2aUS/9+
Ii/Xl3728i0BvylJEzyWMJ8+zhP05w7Y5AXu6xmv+lwyPi9oT3CYNkMdKNtBqScZ
lqDG7BCSMgy+5Cju8CkPktxQAE9h0EsZzDgrW9Z+RKhZXmvaFWqRNA76dUROBP23
ZgZn2m2Vef6EPRmPBsbEVGFWS/5E1rbrzID8tLYzdog9VJpa1x6kjX9k6jMAdmoj
H1+mKEh9aMulH15H0UAl12k0ri/Ccwp9dqblhuHXzQOe4oMOOC37sQ7Ul3lTzgx/
MMG6NgbniFatEGNn41Qsh+mjsetXsUmoWtGQMLUwXrgimzzcw2P9fcG3PD1P+yD5
t4hilPmS2J5YvYle4I5DKjsR0tz6ySDuxY/M3vL+Yc7CYheNRf92oJl6HuQCISkY
t+uHdbOlCNAeAmlVi9iGfoFC4rNEQJ0sjMdnZbhS8ALXd5DwFrlYoZzeXweCn+zQ
iGzhR/VZV0tnn8WuF3x7ZMfSoeZuSkvpDfxWtcHA9yq1SQ5ltijTiIDj4xV1V7iM
6sRqYJJuzTpuidVJ0vbMaXHDVmRcN+LZQVRJcj1OhDYNnK5n7OAFoH2iKTCb+wBg
bLtL/hXHKOgpIW3QfoCKO+4iMONTDopVySlw4/QRuHfCbI1FAnyoQ4bqggbeGr4W
BbhJbufBrRFofwx1EOs7myZRdq0eJi5ZM95sXuPQJKtzVBLXakfiLk6O0gzQzQou
jCa//Inh9cTGujNy7HT5cZxDOiVTSycTNxh2Kiigo5H5nWgmQRU2HAL1g9LjvVxB
zwRunON3sAKuc67TLToSxzPh9zk8sMiBugpeifPzofyQviRMFAcS182UlV9pTM3W
UCtRiJpf7UDvhJyOuAZVOYc4lpMEIwkQj8KNCH9SxFuJxxrAMIo6XK5+Tb4Y+xRw
opBVXMqSySqOJPWiuFn0Gltc3YoqX2GpAdKEsueOv3wePrgJcEUBxJvny/nCZRF0
F7SwKqFb5malFwKSVVt9qNuAPcdiDkhZ83YrXtLtTsomudpRzF3ncecrIGM2NWBC
wWO/0nhN6dNvmMDf16dzwqQopK8f4ApjYRoZS7+1gGteIzsJq7F4sNAfu/CaxJyG
csUG/iX0UmgEhR1PKP1Y2ugPMbsB7PgLcnp0yNNQCplMVxpMI5t3rvDXorSN0jk1
TqyLOXm9KvkA36X6nJIltubySF3Kc3FNgFVO7vR4uN3fyEqBJE4YvMpl57UsCqcb
JUDo2T9oO5nue4sjRqbKnCosxsx+FJZVs3RdyHWCq5Q3VDve1BieblZse5XCxd5B
3F+wGzjUVzWKLHmleh/wIt2k8BFfBdp3mxR0IC9OaDriITVvS4ABcEFMlwgB17qb
Wz1FwXbkRK8RrW55C5QryzVMYB4mo+LEbHcjJftz2l3Oezo63wOOAZ6Wj6d2/Y2s
iyfzPBmcXsEOvb0C6HZ8p+AAdmtUs8FwDoId+RZEHFwne0skvdVeiDpK5ozXK7yA
MPr7ClMKwZ0V/1YLgNLaAXcjevJ8h3GxCEut0111yLIkfnAeDtGFQjnIIjPylXUZ
2HXmVJKaB3XWBkQZBQwWv0kAu+WuvofKVdW7JZ/OA1T0T1JgwjnrEyj1THkScaeQ
0pzhisJetGYihQwGo3AxSf3anWeuCPLg8ijICT0MV7Wqsi0AmGIziVIMB06Xvi5J
i+qx1c9q1tk/lUEMRtT++4S7sIXbq9CtKrAH/HuDLG7MTLcm+/Gpi8/kgoECCzd8
JhPEHRA7GA5+OEwl7fL9z8MLitqiIyVw8+BsPupgV1HA7RVcCAr0dqUdUXdiSq6L
pHNQxDG+cALVe136MVrdWUB2ymjHtsovHLmeHfl3U3y91yP/iPXMuoqI2SS2FQdI
LHy1Mo7NuQyArR/be2gqo48zqEKPmx/mTkDbSFpAmUZ71ArPiZ4vscF73Jvp++l4
hCoT8lGyOL/HYXxzvbszbI8gRR3l440m/OjogX0MQ7ZnrcW3tMfIQH+W+OOUIvpT
9qALWtIx5yPzEWU+i2p2WfifTjo+mo4cZwIiwwvN2na8HbUImlLmkypWOZZv837a
2OZ0TdtIR9EBeInBmOZ96aRF42+2zhqMI9jJl7Yzp1fXClJn+Axz6RiBbIT9q+NE
nXm35IaCJ/XQJWjWHBBSTEC1yuxeQi4pZwwTLD0z17OWEgk0RPerNIa0eVYeEUGr
VFX3b7dELBAmD00hbDISyc94nkhQNRL65o+6LYdnEZNfP2nsly7RrZdqYNQ4zO8K
B4ScuYJk9fS+DUc8IlkRfJadyMMRi3FrPeAoz2gkMJVRVzBVD4s3ixhGH3K08ban
a/D9ZEIeUgFq54GYZ6wTTKD/Nr1ke+Y7bN3R5AmuqCFidtKA01L94nqHClvNjhVp
4Svtxmp/JZEzepb/+xw5JvKl4hT6GgOlADCPwN5+MCQDNTWzg0ADV0PHtH14slm4
b94qS2R3EFNuTntcNabw0edY9b9fYsZnlvn9kFFHZCx8MrIaxQJlXn9Lg3ynyiOA
7n2kRsx5V/AoD/jMv+Vb3A/Bfe0PESHGVoNjqRcboH8hKp7Z2TJ8+GZup6TaqpxB
txLAi7jvx87ugvS+gWQd145/08U/pIU0gyJQzeJFPTcRCLZv/LJ1+83YtGX7P1Nr
BTceX/1Eeoi8du9QHNjFKvEI0ti10K3qQojJ8TdbLiydUApmtEFkKdk5TBxGoNSt
IqskOmfjDD7GXCB0AZ1AvSg+78ElVaf/9PoXhSW6D1ntBFevMczhaFJZ/I3SNvwC
3R1bMCq+C5Y4KqXmOJZ4RMspksHz4qzfcKF4DhXN3pxX6doRIf6+AM1t8WIkyVSm
lWh2DgxDuefNXFzJ+mu/196PUVshNLvnW93tntkRzXG9eYH3bF6UpgAXGRK0l0r+
4ouSQXazoPv3s7DH2q1HzvGTFwmmikRmbPKLwjmCKST67iuE9VZ705VtLf/2rmXF
SRRgkNy13IquONNxUnV/0015Ru/8AftrFCEVKWOp5eC8jg/Eqyhuo2jPsGiwKmNh
1GtsU0EUepeyVv/46W9hso2jXbbxAM9uY3gRtZig8XUt5pSwaqTqOYLDFfYMhMkV
ZAsJBdsD1MLPHONCOmTfU+h+lb877DnuAXTly+qkcqHly8a2/1KlkthLHYyZrr0S
Vzbr0j8iPM9sxb8NBLqMjGoyafpCmxjQOU6LQFKRyC76EzXtr6DLI1nQNvxvLbzC
E2A71zs0M+kbC0XX8l3VVNtBVUzneG86JWZ85pvOSap1FQtwN7iEJ6E9KlChyVCi
7IksjHthd1tQELpdzXWWVkjHL0JJk3SacTpmf3BJxeQCJEModzO4uSfba4SUyOYD
uLKSnZVy9wDDbIUhoovFqGdyVQhQXyazQplvOLgNOPEnDstOGQYcPO3qfpPXcyGv
5dkBxX8iDtMT/hkqJvWBcnZgF+erknIrV8nQjkQivfVvhdan84er2+TjuNB92MrH
F12ihXrndIOHwrB3qWmyj4Blzz+07CiJsMu7SVKPXT4o3kFazsUODpLi+Ki3nfgL
9xNKdlvfzDknY9Y2F0d5JgU9U0IiS97dAvgnanNh0NFQqfJzPQyunU4FDLFhV488
glwrG22d/yHTWZ+S99lWuiSunfOlKvLaSAhrX+ZJBfsXg5jbUcXBtdcvaw+cRw+2
l6g49u/LR9wpt11VaLp3/Z4aYjfLJIF1Z1GIE6nZEgYrQWFtSH0HZRgjCUd5Mfmj
Zv3bdL3fRZDjmk2ESe8GDS5Qb6xPjES9WnUKHG9ZYycFB/Rkqa1HcV5529Ahw81D
AejK1UO/Ro73/cDJirBvPskp9PImm4Bdp4d6v5Wdp3kLkOzMlXLPBNZCgUt1/VNW
f+lgak+Fixd6Wy0JrB/+FlEvau+rII23/q7bGJBeVbpTkUkB2JlEPOCb9OOU12/+
oBxVDMiyXHiVEXgtBPI5OlQ+eZl/satlQ0YLR/XB2OwOxmRib/JzC9wgkkP1DHDv
FLbf+K2afabbMUIPIc7a40Vl8JtQmeVMHpjX+1t/e8/mwOsU4OlKTuA2e5vmlZXg
T2iWW62jhzYj2K6VTAOnYFM98vtb2J3DRGDjyAQU6nK/6B1Ob/7nYB3DiKqSSn8K
96aexNp+ZLZUHMa8nyHBXTw4CjZJOVEkdWz0CmVXa6ZybFzS+KCuy4RVx2zW/VzX
+xaLrAePVdNPWMz7IOjJMJo+3pQXVqEcFp/tk08j0gOqCEgpJr2w1cOHSmz3613J
tKmpmzdGrWLPngmGroJtCj4Lar/sNx3B+JBHSZI4flJOK/fjrjlL6z7Z8MrUMwTP
dGKugtYehnPv/nSvT1MImZTi4fHW6+yc5gk5cCNbnKOVvyTLWeO3fC543UzQl8y8
Cx4Dumn8xdITk5Ps61jNgtWFRb/MfBu1dtGEjn6QURtMh6qMJMf6jJqJRnaSqQZW
+0X6srMzyi8eohtHGLqTvMkbthp0XUaz6W5m4klWgfOwduKdRlr0KzRLXtXlweZB
P18d698sxxdNwgxtKmGCGI6BLWeb2gUrgWNmUYSsr9fMgam8f5uXYAKB+Gz+ZnSR
zELG+bAk9sWvpGlyhkDv6awcLSUtc1yaz4aVYZarVgI2YCDPqKJzIC7lmUv0jUjR
bVtfulbJ3gE28H3e6nJAAdBcUS6FjUHrQRmamj9+Q6U5qS175dZdTgeVgYZUYLNe
r7A25RNPVZmoQLSEk7FQQuMBplXskz9T5GmgjZwSWNFwBOp9+qQcZzHrcVRCthRp
ubPqqexhOp3AJsXgmDnxl0m1rKWjQnIicSNU/LoBm9/znZXuRFZx3zYo+cahZJKD
GB/p8v4NmAcjwseaQqZiXkvr1P4cjZzTCWUWXEWDTWOjtiQ8WfFHJZLfs2vF7kpf
BPvK0c5BMP47ho/pCnRSCdCqsPRa8NaKuErjmKcswYLbsx3u8trH5mKPvf7JpDTt
00Fpo2AUubqnfY3CR+tuMgXATgFoTw5vN6LXxkdk2O8inzkWVCTOdZpkr2bUVJLF
xm/QFx5kJuGV5YszHcPThlXS6/YKCXPT4t0PYOhe63LLbKqgIk1Al5a6/f/MZukJ
Lb4KAS0QeoKqpwry2cYaZzbPcI0KuOnVR1fRPL/Akyxrow40Ds588htp3BWQh6S4
3i6qNPPOk2bmKaYgLYhzryj9BA3Bm24PsNLeItE5pXd4B6Q9k98XjKXjvGNWQsQI
ZgqiuAhOs+Eld//auA5YONnYiD4Finri3YfwUsc8m/lB+3GBzCORUfodoeAxK3Sw
SGq3odg4oXlebj5O8h62pb4XK82dPSUxcDW2cGyc8YNFj4oWa2zeLmV7kNqltetP
8hFx/tCr8dOBDqCw7tp51lg77zEQVqSBM8wkQUAUeZs1Gy0HVcnGy5yKFT9F0WV/
efXmmDtVokq1j5sQCyGSmdJmSzMw9xDyigqa6WYD4EH8P1qKshRYTVTBdwfuM1nt
fa8MA7iZPvQmZOZXDVwUhLKL6Hqt+hb5+qVqTNuB+Q47JGAbB0KUeRtPc6NxbCel
fIyddLn+nXNfzrw/XvMOP9tZqKbw+eluvSK93pRIORGMacQtSd/CbJcTL88XoSOm
uOCdMVS9Y9wK1+9l2ibtH15qtsHydoqGZ25j5l2p+NlQQH+WUqBBZQ69lUP24lap
UdhSvDPskRF8sYFCRIjgGEqfHOZS6UVBBGEAfoR//QyzHj6bbg8eyxgAWYg4LCDX
jjFyWfMkQWqeq05DPHiRgmcTGYsqnCWEsHTz35ghkkrxt85amil38Ch3F91pq+hq
Uh68V76yzjOm+BZbMmLGi9YvcqCUtNoFrkn26uwqNL8/oDVfQp8lXFn6wZtSBPgB
pkdhlWdgR6xJT6mdxH1GrY08i71XNbdtk0NdPNNX2cAVDjIS4GbE3L4f3VvyYwEO
b4Kw/CagFweWV+++iELJQzcXImhRZVaU/7N0entrGQsM5pvNFiU7f7F+B05N7QxX
duRdvI7TRm5CUxyor/y+dgcHu146FUc30+msSwpSnmDqFlXSXw5mNgz1NDgE8ohl
XEVTZedxyIXf9nQ6NCIiQ8ubcmP0BAbZXVYYmy8zG+16PbE/z+w3svBI3mnCpL+J
N/L1SDLqLmc4MPz2EJKLh+boGZgnjL7uaQ+HF9oLkA1gn1n5NVp3P0LDLbi+6Q8k
3Yplpplk+yviwXNqOzTUBLPDOzWyojXoSSR8Elk5AI9TgaFDF3urX5b15CeBoN9y
zW3r4wawDROny1J0R4QlrV2UJLHap/zCFWi594m9LoUprQl6zuDjOi2w7tnZeWDk
pb/Q/Luw7tVWFMP6418NNeoq3hmC5e1/SLF4NSqovTFMFogNXqd/Y/gTUNZsgsHM
gd+cG8/yAvTfzfTXkfWf2sTHtubUH0tWQ1UxIa7pQrm5rUjNjqbbwFh33eviU5Zg
2ft7+uMf5TnMvRVgdJFZ3Pzd8urHQRQMpADY/vgi6tXCJJ+aE2qpZRMT+05bvJQo
Xqo0UZ5rGdBo3pv+y9TYJeSwcOB3XTH0m/WJr36DG0p9eQ2y+OkH43Lgsj0MukjH
ZqvCa8XGdl721Xt3B8/ovEWXhqj0upjAACRHrnh7qA1uiU7Br+YW9t9+tTRARVDZ
syXw9/uNjdJTRSFv1zMeIneifWcmURXhohAuUHQRyp3yulT8dGbx3VoJZtZd3UO+
d/dWdvThAmU+YVKNzQ2gG6y7rQhV2YAKc9IXMUuDJkYBZaY6JNCauQHC7surgVCS
4Ktsn1vZcA+IATmhtioQt0BZ333jQFRxWHHRQ0FyzxTHIsxtEiQ13bCGmq01v1lc
fz0uYVsyilrYGcApK0YfI4AoMwIY0cH7KkzQn9FsUtyvnPxsoKSPJndGDoGxs/6i
2PL+5md7Rbbnkuok8J6auhuqiw1jix3scgRssZ+yhoersY8AXMxxmIIbaR2ZZ1XE
ajJx7dMkpGzz1Zsnh6fK9zinoDRuB6mzEuvYIcRpIVjEaqyoiAO+kbKytQXR3d+i
mLXeYDde4yCz9uLNoiHXHFTXGb63ZkDsVQobpsKGAEOrqmFM+WaA2mfo45KAZBoI
k/obB6nGbHsu2131pSU7WtDi8LX0z26rHU5tzVvQfd/VscxVpu94O8CfAznLs2EE
hHJIu8uZS9DhGCC6AjJsqt3r+9xbfzaBk5WySfr7VAgdIOluwWDW2UkHo4rbW9Cx
/wY+Zygm0++6dxNQgKw4KXLD8+yTVPNmnyEi+eIfLA6mnIxohhTN9GW4KQr7Q6RR
nRd2A5AclZHsPaT96XJLymCghxF0S+XyXhqdY8Jf04muUoKWwV+2VdjhxkkE/WGC
QTn5tqUPAtZ5vjAfgtF48NrWmvqaQzvRYoksY+oJ51cT0MeXImlH6pnggoLqsOyn
9TRvGr6Hx+CRuxtyqlFCTOucJqXtZEUz0njjZ4GT6AdZn5rayEz78/TY7tWjyVZC
daYOmaxZUFqtLStStmFksMAeJgHkEvBIMNTDjgPEUNbXr2qNKUal2mVakT+unDLS
rWAsRuLkm8NfIAL4dKG2O8l31OnWr2L13gbw7kBdOy2Km2j8gNZ00zyP6eLcuD85
0Wq2Rjosy6sljiAF3s9+hPW5rSt7lmSISyInxv8Z2cEweLP1/t4PBOCPG7OwZF2F
+OCxrBg7nuaVpX20ejbohlFrTXKL68Hhj5wh5xk2Cs0X3AK4n33pzicZVWabs87S
RDNrrHoic1lNWTlMZrGiSYW3QoMSVAxHbvg0wU1pbJXti/Mz3Z61iUtPqtBG2NjO
jsQ6zcL59l//dMh6ZQ3agVFbSgzEDQNH6hx8uFxE8DV0zF0R3jMGuib+XwQVMU1V
FBBM8R/jZYVPryKtP5qKOCBP/OCcLunzobPzGmGd31qVv1hhECxsqHL2qNZLlYqi
9MkSnjDqkXiN6thAFzbsKKfKsR8XG10Z/ymwRoL2+/O1OI/mryzO8Haj4x7YTuvT
Q1pq6A3FdQXBnaOovJKa242hDe8971VLGK/7iggsuyA5HSEVjFCVlSJL9rZ7cl26
Bqx3zCfLw2ta8PA8okgJtATcnO/GahX/F/oqP92sCTOj1znxrrlMe3OtP3PH70m0
xTlVvRN1Ly/ymZcpJEKi9746S9u9n4qVVQoLlRgNNdTuHhLgj6kiGiZ1OLdR1vVJ
hgP+AYU5es0OSopgkVrdAZX8tQVqLZVqzNSM6R19F5iwD+QeQBnLaQ+mC/scNRZp
NqTWzN6gAf8395qjO68lJtR5td0QwB25u48rzAnkafI0hS14FuGLO6kCrjANGVd1
DrLgVwG/BTrZkrIKZh50yoh6pZOqVjeFbVd+Jf5KfBnP+fa/W41Q5p43DbhOhHpC
+IDf8kJhV5qFzbnd3f0wDg6pojrFn42LV9ETiSAbK5o2ab2ZRRXXaTLqefs9sjdf
yRfIEwE0Mr6PjR7Zo5DzjSuLnoPMu2jzwuxFrRP0XSfvaIyj94F8k/fyj1sOnRnN
tJeIutimDxSXIP1XnslzA9CnsbCX4l1x0fg++MDGrRNsrOo+G6huT+iw+k5lNOqg
HtyCmm5O5MqT2bFm1oAiwS+rHi3x8jbjhQs0ceBPAPV0FS5ff0/uKXcmwflX5Y0N
Zqfa1KNzyvB0dpLSi3rnO8LVhhWZWqKTaaLEN8uINIuuidvRXE7HUxucBlyX/D22
RfD9uQoOaxor+pHDk1QdpaFWQUKAhCJG2B/7LKAGpKVrwnmkU7eZUEnGt2+WnKxR
askjRWS6a1L+5OG8n070cO63uDx7R/tBGn7SK7NK3HQbIttfF0nTapzZhyNnnaUC
ePLD6lo2GiJ7Ufb+A9tGbPKsEGxsR27bqhzx7nUxHuOgyF/YOOke9qIcMZCMrz6c
XakwY01muuZVk89BFgAIsjA/FBxlaPvSBWzfdUet12nPL1gnxiR/nBmQrMqEEvzk
vf2Q/As0fp5OnnLAKMDqnOrSOaH/q97bYDYabRV54cxdZqIdRTKYYqpg2WbzYDKy
m0RgHOWyTDvhXsipu7wiOi3b6s5pTq78pxOJ1wWlDGx/jU7Ji/GYNLiVVmBTeAwZ
LDYLW8nhEyg9jMVuqp9DuAXCUMIm7IKxVkk1/9j1/tkoZGdt85n3Lpga3zYTOiic
XPa4jZKfEcBFw/QYs93Xze/6TejB1dYHc9JODMhbBkqCs14oMO7bJQm+STExWtpF
KS3aiVQY3C7hIZSZ/+Zr1yxGvv9uAo3Q16J8LwkR8jODtuR5DtU1Nh5LtrI1rpg+
TnEYbB4zDHZqA2UYk6BByXYNqgXa3N4RSwzO9KfJgXhxriQ/uDfnM+zyBcvQernA
3XBaQWTcqbbmwRBvHNf0v/WSdDeAQ1yCQ46nwgrD3/ijqkybj+xq5pYGJsVDx5uf
mRG1o26LcAhzYJZ2O/R/KjfFAM9O7CpyOgcZVAsvO+giCfO5vrvmv4iZ6ZRdTkoZ
L32lfArJ61fekdoI+Vr3W+2tCPbdSIZaXnxLIGk3w++FIU1z8mygEhYOks+YUYMM
qoTEfL5XiXPY2mfnkb5tYQmezFAtVNPeJTr23hvuF+J4r5a6fUTKWx3VTFLLCP2v
PljuGHpCjcwsuPP9bk7fDGfWnodo2p1Op8yCOtQJfeg5f9XWIafAxtTLnfZtSL2F
/subuZIUfyGn267zJz27i1f1iWDYPoXh6rSfR/ZRnnyO3p7OuC0vGg0l9s72+GaU
o0C6LHh2wE8NPVw6c40TsxQFb5DMQExauNcMwR2VKBN1CmUETmcGgS2Ny9riiSpq
ieDPxPsRRD0QWr7NMqFVRHIZyppNOwP2Ga1C0ubbt1zPoy8RltXKYtiX/C7wUGD0
9yEWtH91b4Bx3rPE5kkxUud0Na+1VYuq96sxZOxi6k8uha6wStH5NN6nspYLdHd+
QpwSnQ50hkijJ5SKm75e/xfBwgg0NwnACXki1moaV0hXw0Rdl0IJcUB6+4QYm2vi
/W8UsRV3Ovg4qtUlSKyvcnjWZetwtNSX9CkaanG059964iG7fIlHLIYMi/v6RA4O
485SCWpUVpyPquQ5rRFkzOUr/i3USVzmQTPvNMsG3KO7bqwrnziaQLKvtEvdPOG7
5P71sMO3vxUQbiPn9o3fVp3FzurawAF0cSYJodwwEG997h0I5AC9FDI0gFCNDTHy
2VHiAcfmadkIR3XRxtNVemRBSNubF3DyDt9XjzEIDqkzm/0Of6tzHXRBZb9LYMqI
kroZJLdfX70UJ81kLJH9QC+B28Xc9OwTOtn1zrxpXRNcq4dMZT8+d20zxfphzjQ7
TOQBuFrncysRCWw9vyTPNVBXhN5YtFmVGTlQoOI8ednTrlyVM1UDuIF3Hh4GCC6G
CgXxg09EVxbxd1gGTdDftybOzaXP6FNFaJaMhB/ycrgpaT2bFKVVD9oecxV6NSAp
y5UKTw7XbRSCDdJIBsNnIN5F7aBSJB7QHc+Q+joWowCf2Zzn27PgvgivnIFC5b66
pdQglCQad1I/HjExB+PIi1RZtBXhpKcvCkum5cM86VOOgqEbgrdHa/G6/Yz2FhS8
zl69rdARFxo15ij4XdjbcMOeFP/8c90Igc28lXQEIrwSNeBrCtjOkVk2bc+gRVbu
uKcW/kzgsLK0cqD9Fo9U4d001I2PGLucPJ9rNwP26t4a9hnwfIVcvHoSvuGEeUGo
8ga4IFExm2PrZoM9X3yFOUl7Xe6aHMKig3UuwPZEeXvDXXSQ3gPJ8ZKL+8KzxHaj
5CagJs0wufc9MBx8lQeW3DG1A5sdxiquB2MfnnHg8p5D4i2Pz1hOkg/7mFRHWjVA
i2fhJTzpKbZ/ZmOIPJfrL4iLE1LAphE0SXqV2ULtVhzxdYE58RM+3RIKkQogF4+7
+rbDRZ+K9sR5z0X+RGloG6o4RZM+JzYe5btvhqBDb6hTNwI7iM2KlOUEHZ7k2gGG
0b6bROVP9I2r6I/AAbIPvr+KEMgtm9rDkMqRaVVJwE2ZDiVxOthqOXJlpf6NQDKq
q2X32hMES+rWSFejZntcCzst06enAvfrvKs7lf5yUe5CnKqauQJ/WSlgXf6hAHzb
7NQmBqYijZbRILzW9Ku07WHbxyItu4XWbWfh0y3LLahz+m2s6sBlb4l362xU2J24
EChyqeO5x8pxm4XglGJvaUBZ8NE8cZIY2GGV4jMIiy1uleNsdkPW9H9OYYr4B41x
R/Pi3n6pGvN2b0gkH2zQeUFUxAUigZUTMBIVcOm0jQTahCHmxR5CW2zR3ifdssAW
WWSuEv6ZV0ZqcpV74/CvHDgLNtmnk7VGr764HrLrQf+fj51cLfnlsiXaEIUoYzVc
k9loeFMB5BaF77B3T0wE5JYqlomLLp7FJ5VOFB/JXXuMBgn7qizrqaB/Af1oozuP
9DmenasAyFbydk2Xgi865gaAfWjP2Oi+uitk45qslJ2BSw/F6EVyMXdUJr9kl1Zk
DODIhgylXnG3sZRqCKl6PYLSM0zIU54vd1B8PLea3Ro84H6Dp3ndIv+I/e4TmdoP
iDhYxZdTWmKqqdi4OLtkPcyVJWhhCegN6Wrs0r3X2Pq817K5UOHzBXJtANzZAnlM
iJx+ZZYM0QzdeLMFHqr8UdCmckcYwRwo1gi+5dzSsThOfZii9o9JmuDR/eN3YKSL
KbYyq5nGzL1LtzvL5SZqsLggYDCU28hiH+29d9Li1A+9aSonx253MvNQVz9A+N5O
0xfepjEHSygAorrCMJJhQCJ1PPy5N03dRInP7ub7V5co5ffkE57U1VjHqUKBmkjt
hoZvsC79MQpgF36xpDQb40T+sDHYjsQIIvOgc9vzbwOMAxq91FsuidSAKJDwV+9Q
5f9PHXO6tQDLQfWYu1N6fP1b3r9luotR0QNOPAZ0Vk/T7LkLBqIyYY30QUpBXhxr
73PahODH+TPcjQSzqvelb6nXlwEjKw6WtsyO2Kt2VyaXWhWjO/jVBJ0WDKnfVohF
CPnMd4jhQeVsWXVZuO8Jrql+w91sARTpFigRewPtMUAyLsNPqdA5CmbHXGXkLp7V
3fNm9zVPydMulbcRbMh1psnDYXYsvs1kDOAOO39gLMMlGJrDRByZXPpDcZwfcq7J
ZxVvzIml6Jlk1qEO6LUuJYg5vC5tdGFzmNWjQpIm9PQLD+x8hN+dCcz/x+bMvamY
EotzKDhttlMVe+ckr+Yh54DJmyNFJ0bpPILhLQQOKOsgaijaYIO4nulAVoa2vc66
nH8wzwskb5SQmCzkpI1bsorYPntExUdlr8xq2NZut9Xp7o+G+Rp8+wWIh2srV01O
9LRGcSjfw5+ZLESzV5/p+KwuS4h8qIVLDrtKcLGfk+aB3EX+8zL1BAoSfNSReCOx
1HnQp9Hn1DOXwGxeBDO8CDwSgNHU8dbnOhjVHZfp8gv4T4TKWdE8N/pHbbUv9d2I
KJ3CiQbiawct/qdR+av8XjdaQPG3zIK8IynHDeKI7AAp2wlrz4qna+ElQ9FuZrXi
ayrYp6woTcs3fBjP005Z8B0YusAP74GS5tmFVawz27Wka6Udg3UdeZRdKelqN5Jk
5B8C1gy8Jt0xONuVxTf9oJNEkHZKrIUvXnBU7FDDIKo5JNkHmyHkfMgTitQOesL7
eLO+j1M4DPG35pBzdhP4KW6ISHtkhdleD37hdxNM5mRTQ4D60MX+8toG8nEPjrx3
thf3bG0DxWfYqQ5h9nsM5hl5UEZ/ktNZLjHsP2LjncANhyThIHdgp8rJc9qkhBgV
RCof/ffkcHdbk6PGJW2O+kqgDusUOq21Mzcg/MDgNarjDs2jx3Lfe3LDLZ3o+awQ
YnniU9ygaSBTTwZ6y7nrRaElakyT5lPU7BIqHsVgQieHJyLp3tbj6ghIYfTm9HOW
fzpnHtAX7X8DuZnGQQkE9gh/vKLOXSiIH+uELMJqHh47fOKwsyhFLOcH0YJ6o03F
jyFxyKWYF4LvxkGGejQoZn11+559i0eRn91sXTJGVrzhxrTJxE7wibRzfkjt7Zs8
AweJXCH8wfMH/QWWgA4KajU0woIcQ+EOAAonUdL2VCaMNqRY1KIDNGOdjzGrrsCZ
Nio5t4D1YtrgKvIIE2VX2DGXR5zFIZjgfDCBAQJs0I36JsJyIevY2Ink1GaXVW4/
HRhsyrNCAYheR1Nz6Wqt7B2RTy3vB2TiLe+HFFOJ/4wmrBonXUC5EVU1otONRp6O
q4g9r1VHOq65bsyLd1IaZavtUKTJ32n4nuQxIfjzRVWFI119on+rxFXuLAyisoR+
AoLWKBhxryRgF7M1p2J7UUAo+zvAUC2Yla8a9t9i8l8o9m2H0pYF8/KgD8MHiD3r
Vw6YZpmlQZqU15RjtkAVf9m9IlS8n8rajthZkSzgX1GOMlbEbABc00+9uFOQd72B
kZuytaCT9pQaiMXAWMSkXuBJirAnigwf+39MyX04jJPTiHLgpILwTGmU5+zP/H0f
pBpdIYuj0nnyxXHW2+IoFb+aOY/h4VJrM6DMeQhOKiUr6u+CtkLHbiLYoSNMToTF
J6yjPAI4pR/57QiCLbAV13gW8YW6ldTZl1KtPBNmUtB5QoDyOdqjm77XCbhlN4K8
5HCg2OD8xsF1XmYqXSgLkFCBTmCtdLU0SgkWc2tQo2rV/NvIHpTcubDvRU/YjGiX
2t2yZGe5dMiq6zIQnqW2npRlDJh82TfhX0rmxXQP3XMLTgT60E0UwqxkiCHCbVVV
KLAOkWOW7tNl6Y0celO+IxSpzi9PeIJmrABo3Fyl7bF5gEA5i4Wf8zsScmR40DSu
C16nC+8T7j5zEWIahfSS348uhobLH7DgD9jjHzHZJwYdZSGf8Bt3n3rvnLF4fLHN
ZaG5TEf1UvNVwzO1MdBA9NrI9BFYYJrhicYqIME2lCKFudN6Zyzd0/3PTsSF8GmC
6fdLD6Wtc/gkZshAujHhyX7sLr5HgWWDfzwxslKunV7Gym8OQpgujtYzoDsRXS5H
74HjRrdU6ZIcWAOgFiv8nUwFgRqtMw0dqPFpHc5OSh/hF6pWwoOyHjxgMOLQn4Cb
1sMtayJKTvZkn16c21MVEuI4BbmblIhKovFj0dwQTgx9vZbOgl3lavR6MzOvD2XR
x8uwm3MJhbhUar/JCqIUCSbSVPFlwMozcp4mfFwulhTdhPRcjeyRXh5vsGgaMBv8
iA9sqV36ODovLGge3/tJpkTBdUQkPej4Ci9SGWT9dZ6GQyOzkroylV7Wmti1lYsG
zSzbdKP+514kRmy1IEaCMUbsP6jWFNm0bDHc9GT5Owcs8SIfQIDzPIAHV7kaPbLm
fXWdLnsl0xdd/jF52UQdGCLxy/dfwX8xFchPKx8XQGRG/T2qV1JzdSrJPGlGu7r4
ozXqUttugaeZtDsKJnlw/uXdxP/ljW3InkXeabWwjWTDL65/Qjx35JJyQBm9rBPY
xzlli1cIJ0TbrO7E4nZoZfM/8mQVBsr9XGRAXAo96Jfmu5icLred7mbk1gsGurt6
XPbok7qKe+UgvwdoP/gSGN7hXGhDe9yafOW6JfsLCVXXFdaTJDf/3b7yIHzglMgt
QMtyZeMIJUBF+q543M7KsblFnUJuLyPXNwUrDn25vsiv24DTeNYXB29EtLuIiNgI
kaE+zYgxt1ATkL+yUefqw7OXLFik5wl/0sVJSp3aXf7DhGXkNKnJOB2vv6c5+If+
3l4imjBnf8KKQW1dpzElkr52T0CVFbhqGQzXVT+cFh8uCwmbWFHJbtUjMh0kCCTf
BaPE31XTEeqxXz0ZQpsReKO+HyiT17MSIYTaxJMNsdp3bbvKZe54/adFVMCZsnnZ
ZquIhCE9y2cu1FKgSAIZtl8H49EaSsw/+m87ewSs7397eIEjT30Htu0G2ddKtpFg
qT+RA9C3EQjMW2/EqkFeR+l9KyfsO3l5zsK+SxJnhRTvVSigCt6JBJrGBTpOFn21
+5EeuLdwWwAZC2JHMiTTU39of9mmkgPRcoiupUMmJV45zn1DsakpWLeISWaeGIAZ
DORofgBwvl7q12rVcbnfzu81RT93nMcupRPlYxbLcbhwVJQw1+OREWECjbti95SE
v1oU+dUd/V9qkMFJxDMAfLxIthbI2Ird2uzJhihnFBuCDqzWk4ovQBEhHX+XSL9o
wyzmQRMTPkgg68ci0OMafbfvwBJh61K/YVV9L6qYykRH9g1IfyHGUyv0Oxos5Sc4
7kxIdoJhRHdiuZVTIweUW6ZqUGtmgxr3/CvgtiRbJvLLu4wyrjUWy27LXs/UibOB
eG1ph8gVoGr02Ip4rydPgwm0uGBFhLw0FKeN7R/a4hmUcAc20NAwQfucdVIhwkL6
tFY4nPc8J8h1aY0/QAcyHGc809BCt/cJaEKn3wNw0PLat/D0PqQXiETBaP92zHI0
ekWcqdzdZhCfq5NSbHeDXOLxUvwAKhsSyQcopxbpb/F958e8MrFwEBWmSYD9Ldyf
fJNgvz4oJAxwSq21B8W8+Efk7MaXCtTtK74kFgcsC7AMfgl6VNKWoVw3pobjVD97
VTtyya49dEqOF1DLpd4b47jSHPzyuQlAg5BhP6yYeyKQP0SI5cE1M1xti2Hbb0y1
RQIwjitnPXNXrrHfdheC7op0mJFhZrqQTvtYya8F/gTE1e1bB1VYqqkjnvXwYriU
MIqFjC5X4q3vhs1mwidlU4F8F7ZhOz77CdDkPi4QxlUIISEoRv8iwOnLuDQmMlKS
TyAsP4pRK+3gefvhrsyvluDwcvQlPDx1t4ROkKTVK3ZKP/t7O+E5go/EEVDVqn0d
D8jjPJJNT15x0oENZIc2+d/IFlaSp/iEHpu6K7JeIQKJdAfnGlmIu8KRwJAvfZ8m
e8UjstQQRIhSfqnrW+c1Q4En8Zre0NQVQhVHQWjRgAANnw/H8Umgg3vPk1hjTbtq
b5cKQ9Ds+eD64/QR53a2IV4KnTxtfMRkmxR7kGQ1kQtwwHF6sGiE6aKXJQJa2wJd
uFxB9qadPK/pLjEgC1mlaO3ZdpmpXTFsO/c7tqk4I71DE+qCeozSslVxlOXKijFo
bHFl6TJ6QKdUWamfaUOoG1d7wrCxQoPz/gj4obAwR96EjiBZJiPPj0d3fvoQlcIf
5STl07gRS/zPA9MoBI+mZNdpvQSP/zrX5Xp31NRnN+riHdPAtzw2oE7niWLkM6Wa
n4Nt2jtQ5NSKV0o9upB/SkzDCea0mYLcIWw3A8dSOKk5ByWIDZVR6xndtJ6+/hUV
eGjznTccRR+r5cSnJej9LapB5VDI9Ua+xeW2DSAtbjsEvXyJPnmI8aDjzonvOs26
hJfn9PekCFSHy5Ct88qzBiFUJxYaBeIfJuGuJdFtG0W6tufvMf2WklSNeaQwKHOs
hbpdGjrhmCvoRPcS5D8ym6SA2de1tG1WOF/c62s5o1c0eYlgTraTlm875JXo3c0S
wEXLmOL/APrJh79bGhRtjTCplvfhTbV/OgwvVOmUhJ9We4TYsvolXRwZ6djAdo4+
LIojzq4i652wl0kqyQ7xmmsFAY7CODfxGEobHQqjA89vGHSiyQUGrkIMMOCIXwGC
bGUxqitBvs2UsRdMFRExxmrGh7Jds5FhwMw2zmIdPS9soVSs7DQ86upUGQFPinPA
nMGdcJf+TCSxt6rKqbvb7u9HDUVLDcGt/9nDCQE+e61iN2QaQUO3yviRlzXRzsNz
cT5RFCZ+Ncmx2VhSLRsTz2/XCYsUK2cw3iFvYVQZXZ9MZN3DMPGPxguNsC8Hz4+a
MzgVmv/FRsyL83HZJvurYriMZ4F1rGd0YY8kwV9HgvgpxuZOZLzoAoyPXbJrFepW
klm4zg9b5zJtD88dGCbl+wHy5AIk6mIMWaVKHiXder4n4hlIcnKo3T+cWHG4yied
RnN2Sys+MKzlBqEim4pxdZvH0MVr5MFrJoMcDtw7dTBRAAuj8QGSpobDB4w/NISp
aDLc04gCJWA5hZiruk+Vtaq2iKRLWwtNpl45dIvIHcYrjwVTEHCGySVGjCKifilu
zZ9CU6ZtHE/OKmMNkDMTVQsNt1eYRniaNFi/sM/Ykk5FaOX+zGxGQJ2lhIEzLnET
WyWS6dwoGVhDCQF5lcLG2N/CcpOiR9t7Z6Rl276QrBrmyPbA/cNxMGC5OrgCxiop
ZK3LeimI4UgjtU+LPFbymY2TcU+2a2117BtaCx3rcWxhBvDW7LpyC/2itwBpUkHv
69jTOA1dqdIGM292mlwyPnlgZAJGdRU0578m5GMD3Doy0bwFqN/ehhZlbziD5Djn
CCIxRmovK4WABuXN8txkBSlULAZohwKvbnyg1AOEjgh6+XvbECkjMgKwm3L43oo7
ZkhBaHM7QctO7N2pzdIbOyOYHyh08JvfDL1/gJjj07hJooX0Ho0k2+vlTox6uofA
gdqbYaQ1ersv302OYV95rok/YBnwBrNGCHqwrYbuModKazuAvb7IlLi9+yz29uFp
aBtDR9cdee0uQeRTalUSWHbRdRD4lRZUEXzBnHfmk2VvuZlVNlRea/PDzfoLcG+5
Hea0X4fvo+Xi4wsph4I/40IWj7X4Irc/iHU9k2Ra6jy0VTA/5ecIaC8gfl+n9Hnv
oIcErKP8apiQAVdDE6JY2GxlHH0sDDnURk0a5rXcRKtjKtdJ2BkS5thfLXUF8qct
z+FNrSc5ESdBLKgxNF80Tj9DzksfBgbFao3y2wdrYdC8rWzpgazOrGNhbILo5qd6
2HgJqGSggYyBbi2WKLu1+dApuFgj3Rtbs5lavlYYhUKAfMyqljTsQ+QtivbV9Ffl
IVUqN0f7w4Q2K+5Q7nS9DryTWPL8wbk+4CsgySjLfGyE0gkNkPjXXroP2eT7cl9H
7yDVg5Z/Rk/UxobJtmXCT4BJEbrc3xyYi0jFgbGxwPukkbz811W5aWqNslIQpoUd
pSTkOSPdT068MCWug/EqxYTtCLkAkU8B8RWc37McFMqyNU2k3TL6tHUXxSEkElAu
9FaIYbKj56ZFanaFpLgALgQbDrU4M5IvqisKG3e5P+ry29GH/wof9ND0oMbKlIm0
yB+fJvXEokD1VdUOhclv9bUgyEKnCXTRjBDr2VM7VY4lr1/zptqb3qg473SI0ehV
6AVPexr45AUtIWqAER27F5XBHNAZGiKrD4XPQUrwB9LogYbnGEVDIMsj4i6DZ5hU
BL7pzbbEY5wwD8WaiVvG96RKbG08j5rHbK7fFr+L60+s1T3qKC4Fnw1jkYhl0npC
8BPsKmByPr/Dzp3n6U+BocNwA2KJKHSkrHumXKA9lbWCFSVLy5Uh4Jsc0CEI/2td
92iJVrXWNjREzzFFSaBSZN+/N4zMUL4O1c4hmoML5o49fBJD6LUEH6ifaqs4MLfM
njqr2vhYNsji6tLspYuu1iwSW7dyVRZrKBg3+NI8BBaA5/T+Pj+/odozhtVDeewj
dGfVGlHHOTHKhzzJ6utZGk4iR8jQF19yqAPRbBlvlrZ5HcyAPqoeshfC6yaq6PuN
Cl1vdMQFU38AOikw9g2iOAxxlu4wzuhzTCZ0PYdGwYEWp3gXTljk/yriHOXOrXU/
lKSEty1xWFS8dzlpEWOk0QitoONsvlOfANZbL3GEyAXCgg6/b9pUN7wqBTU+syeZ
wH/gBDjHnX+hJW1KKG0hK1oN+bK31pb62drqHAMl+fUOULg3XxpWOfbgBrx9QOdr
Nib7LUTEFa0fXNshHOSZniEEBXa4o22nsmQj0lLw3TLN3PrZwBXutInO8NJCfc3w
c0MDGM233SXEQKcrAzOQhU2Pmk1n5NlLNlLz7jkwv3idIDTxMtjApbhQKCroraBu
160egtjYhqy6nqPcQN4Us9XqARrriJ2VFXj+fPfgJlt1N0cbfM0JpAoba2QXWcoz
oD+8W1fvWaE5g0MLnzD3GIcuubMft8pyIFxoAZXoMGgmbG8qfPqSEMtt/HwgKti2
19BSQSpC1pouL9rtfX0e70oHbihkFpqo06dgOrK/EwLOvr8rcqTLSoTHtRYlHByN
78eQVyqJl737w0AZNJ3wb8ms2K8VUgjGne1ibw8j+C9iuukddFxMxH/FIHVeKXiT
fuL4KpLJkm3U9S13G44/juwE/84nmhLOCINXe7DqEkDyZXKjSnvoAae6gyh14bbA
VhmVNhUWOfo0tR1T99Fr5OD+xVwYYqcgJloInNfSC97hnCvdnx98RJ8bDogRT/rK
k/0x2HTtsbUx2S6u8XQQiys9b2ibODxeNMN2sLqmPdcYLqsqTyHTiTa2h62sr1kN
9MutOYm1M8ScyIief4ERQq8R/hXoHNfSyE4E1kh5Qjye6smQsk2PJwULMuzDDYXq
qKla+s4bGjxuzP+7QJm9RzFwR0ils2R4MehGQw0LVfH/6MCe723GLy/RoLDZ2WVF
h1pEC+bnGwnUWxhU1ckNuALkJYoZltggL+cQlB49TnQkSi1zEMmO6btiladZs9NE
wCDGl6hv0Hsm8xUndSBxFV4WYqj8H85L1+sTpuw9hEvgSpsnZib+/M8CROqLzuns
w/SG4T4W/XNorZg9eqijK/YE7IIJc6ooMi9boYzhVaktlPwKhNHSNDwzxZ+fwpRg
WK9m9Mj4xQ3oJMVuml+kznvMratq/xTgBMoY9JohRmThsvql5JKBoT7kW6uioN+x
OKg1I4v2V3je/nPbpD/Dn5hFPMMexkmA6OLWigNzH3Q1xR6gVKVE+xvKMb/3phkm
rsZY0APr9+Hrr60O6mAIRh/WJl+cJuu6ABFVZTOC+MM/I4cPN/x99iE6GnalCrmT
dv1Ken/nieURTKEkC65GR5u3x26BSFvgbj5Mf52+xmyxp76obCZP1y3HhCNUeV44
hX2Udcz3/ZiWBk4au3T+D2LXWpOpjSbGhpy02qXBXtKmFyS9lqb3BUJsIAS6JZ06
HysHLTfb7dgYyWNJxHSl1jmaexgAvwVjb3Qhqu+IsfKxM1HjKMl6BMEEymXOmYLM
mzhjVj76/z5BoIiRajHClE2cIpBr7WBvJB/egrQjWrfoOPsZe8M8Gv/hLXCh+lgj
89WjgBeqJ+kDmaimXvgBY6dXFxpXndr1YQd1tnRhefOxb0a8p9z48hbt4AIioFHS
BJy33Ee1+If50/NbzuIfewFNyygjKq5qPfPLEizF2djZHIOwgEQ8CPgJz9QANElz
5UXRE30SEEH/CYjm+/1O/ZP4WHwWDizle4YKkRHYlFVlqdFNobceW61Bop9ld/rp
0ds1OTjA+6cxcocJ7JMyJyLK2b0Ti6mX5DAHZX7pn0/bJk1CgXZugIb6+ZmVVbjg
QzNsB9q0o1MEDjgUQrQCYD2wxeGs7lS/jq//VSDu0c1L5U/j7ttSAvrI73x1qYbr
8h4s3y4sq1JJPAv5p+iVymzXinHjS++YcRY+b9eTxHa/b040mTN8J3zQJprp3QjN
QWSVpfJEsPkapdR8lKCa04iUuZm34j+UHB/uH4EN4/OEpO185qe1JtoxhGit8mdR
GGZN1OHfzp/wWIDR1nA9mqQ5VSy3sgGcKuQQFcMGEH+QhrSXVVq0a24BiN4henG/
tjhea6E936q58nwqkET5XXUl6O09VsF10yTqybQzPnos1KYhRqYiAfGeWe65D5BO
5yzluKpWPTxDQ8E5uQ8yTf1j8/9gtNoOz/IDlUpxCd24+aexJtRfhgvQylQrLYh9
W6x6wp3jd+nFNzfr2L93ohAoVmptX3r1xCvKWa8vDl3SP+iepqAbCKjhUGjsBvQy
OEPFa9/PMlMXXVyFYdNCNVU2/+lwT0qyCYuyB2US832vDRNEBTpmj+7w9Q8p/Hnu
hCbWM02Yx64KM8OhuaGtOQxIDHxRHVbJ75lMdOexISH4ZO6poqGrBLf+sTbLO33u
8ICeTXMO7ub7at4DDezGMXsvv7TcEC84XIV+b5Re6pxGul1jBdISyE9LGshf1quY
bcyfgk1qvQHhsaCEd4ePQ2QrF5m1rHbw8kv3rITVxMTJC2g3rZLxApJZNUktm3NF
RrMkyik7ngq3Y+jq48APxeflu93jA7af7Q9O60RWkRTvlPUsOQSz1ZpFDqP9h6Ja
NsvwdAKbxG8F1IJC5QfuaHpFXfQZ9587IMqHjx/98Ybi3CmuFHFlRFGvEzPfQnFk
KUe2f8RB2Tad6G9yUDDVDGVsns3zxFBYS55j7rkDf8YcZEHdI3CxjxG4NPJY18r1
XlcYWprnIUlquzDBb5g1eRUIa42KVwAjAUMRkhWudErUUvofQ3xMRQTC4fvQF3cY
SQVASV4hA6Rgdfx+ZJqaVYK8gOEaHSBcK2Yc36jvUJW36be4iIk3h1d70SwBILuZ
3qds7+LetRKZaZB7hkcOD4SOUap9LoPUv1TjyYGhZZQ086jx/E8sgeUNFRr+ADQP
5TFzLCFVOCY/fIIdHzV9F4AP4b+9ChSUeYYiC1Kkw4ihnb1R9hG9ntM+a+vNu6+A
NstxiKk0+FMyajkTty1hy3xjQ1Tnt6dlJGmgpa0b+9rdZx6DqD8OXIVsuBqt3wPh
wID9mB5VIh0W/9JqlHgqOvLiG85Mw7rN9hONCdNA0v6rxnd3udyZvAax74xv7MZW
he8yRvduvubDCrtn1HvyFkEtCE+t6Z2HGFmj3ds9C6rOptA+KwvyQ0Kum5RA+Xg8
r5cOaeHiGFeoa5uUbVvFRhEYTuioYOhoztMixHREBkXH3U+wSY+DEm+hN2bQUKSk
BrnlPmq8AXis3Q7Fgdjh7twjunzTxNeCq84p4CSp2Rn9PMP2/Uk87Y56rT0iOerZ
IQYrdcSKMzia4fcvU31iX5zaEJqR4/FRwPqumhwzIvo9zYZJ5HPhu+nORUWGJJ3S
Az4R9lLQWnLYnNPUVgZwJLr5Gr0SuoSef9MtYfqCpYMlHjyaRY/I6tiYOsz1C3NW
C3RimOpxPnwsl4JrvPc6oG0l9iIyWramXz5NL/VXZftg6UL9PcXkwDtGgf+pLFJZ
loTj+dds3+2aPfc+DwLB5e7elaNqAtCIShNlB1QgZV/+fC6RR8wpFmPBBxWa6xGF
MgahtpdD8LCAJI0rcGjFYIQJyBtlmzfYzMEZzMtTO1W+8hf2MSRBf5H8B/mS/Te6
m2HoXySyR/+PD74M+baej9mZvS3copgghVPhZIGy6IK8t6e1hBOxdZZI2N3i0L+A
5HkVKW2i9NF0G5mMlThYa9vHAJZA2/JDoDJ5e1S/+UajFYa4jEAH0vrjuqIdllJW
xh9KJdaVK+CjPf1aMKY+yxz/Xt2lgo4kDo0KB1yyCc2XtFIVuywz5I88J1SoVYPW
wL06/pKTCZh5Q9WcxkCJZyji8GwxaY0TBvNwiPJK/UPaFRkbZo6tSGNj8idPCNE6
SxxXFIl2UHwZQCqya6r48/YIlcrEfGdtw0FRoVNVDfP/0RL+0eDYDhGaL5OP9jWv
D2reo5qEpB96qqTMSfz20rnP2IVQmBygQNDB8MEepC17Tb6brO4OyXZ2usct/syf
/Lby8cVDlGuDoEO/Rrl8erewDIACKKPyPFTFF5ULb64qSe7fRabuB9pH1J1+rv0x
lWSzEQDMrqX64WIawxsk5MsXiPUHik07WQKFJmRM5kpHGWyDUk4oNAfvLEfCvcPy
1plv6wzAYN/jrX5DragTsH+D36vFdhao4fFsfN4G5dL7Z13PYXNVHQg5RLeSTkzz
uYkg5dd05YapDRMxeqiBu8utqDy41FEw+2gMzB1M/0dyzbMTbz+NPzy6IpgY4ygn
vsT5o4a9RHtabgQIarRCk5+0ztP9crIzFFAzAdWe/agwhd6l72WsShxqat18GcDU
xZLxHMWmnuFy4qT2BqKhdt4E+a1LZJPhDvTJ0kfSD+zuBuPYWYaanwIRnXw/grWr
93+LD0+KZNA4B9afVWJbKGHuWSjgE4iCRvWKbu4hYG3n72iFJfanCjW7n9BTJ/dy
MxJH67EFLszKXt2MfzWH/vdwOTNj1jsrUGhoEv/ebBuXo9i5KqAGJ4AwXllSrwdz
oZOwkoOr0FVN2/eh0WCyeXPwWDz0Kkvc1Cc/fnDpXGSjBz3/F+stgJRW8h74expS
ggBLOwruTjtFA7T2deADNq+cZU9HEAKDnl5dnnkf60RbgpvgEXpNYF2VkyyqKqkN
vRCUxaib/dDc06DriAA49jFyW6swml7LHzFTJXd2yTdbH9u4psU1PgkvuEShwGFO
PajP4jT4I9Pjmr94LpYpIWK24FKRrdVvi3MqRmjFb6YoQ81UHa9L4Dyee9o8KZrJ
UYCTPZexHdxnKze43UT3z+vOD4ajOTRgVfYpdNfJryGLp0zpfNeZONiaq6m6YULE
0kG8AeJpOfC/xCyuivq5d2Jq1o5CfFCXDBLF3MY59+Y69AFv7YTRPJ2NdliHnVMR
6FCz2TXOeEJx9hWN3kgpNFxlHdhwd2vrxfnuA9e+jDXOK0Tla/kxtnugQYZ/IFOA
35g+ZuzC5TKgGqV/wmOWfy1Ph1hzd94XQzJg+XRhv5zvSI4n2rkWyYaZYhdGH3AJ
FubcazmrRDC/KvqW8XM/+PfJXm7CskoTJgPAn5MdX4T1wgzcilVKG1Ay5VhvYmnh
ekcnfbRz6ym9TX/za8vuDe4s1H2qqzD6Wfl9jqpbFVmrA8jab/q82xL6JkdDSNTS
Onwv4Dm/IZWpVsoj+gTlVLuyfzUGt4PmhjnDwDhYFK7ieAmv4NY4RK5xA5SCmoMl
L1SM8cf03n+f8vhYK3qtIYz4wiXg45t6iEXogXnOENxhk/IcyHPwGCX+U63l5BfC
H6RROJk6a61argMygX/wxcqniTd3Oe2oeKud8N+UIPX2+pyWeELMiiHNgB6bY1bN
NWYQdoSlvy88Tr79ipzi9ZKoq6bzWNqpacGBC4rxo+SxaNKVU2yxrUoic6RYvc8+
K123TCQpSB7PF3Jk6k0V3frc7ceKJEZxTDtIv57STCbho99DzXofY76efJcROp8c
A99Jzsoniydh1Vt3F4zgIOE9bGAKzNY1IfJ6RMEXyCMn3w8ghoK+Z2erNX6EuATe
sWm9f9YYsJbu0ZbvXDg/fEECOf7TTXGupC1j2dqeXcSn1HNkX/aL11q5bWMCIb+6
ul/NhEaZTn6z3aleZl18AE5HsHR6dHrPdLoCN3cnuU//Lx8nkdqXI/FoAUXvSF7c
BzciuyUej7pUOSXUcUucWWmOulKbGxGmMWcbDR2ZoCm3sHqIVpqZJL/mtlOt9EVY
33I6w/FQEzy9vFVDJIJCfTf3TaCBUYTkhU0k//Zqnk1L9zEsQeG7dlJh6fV2sJkj
YV2tHZBzOa8icNlSct8beG8t8epn6CclHUj0kmqCnf3FeMssvem0YP43+E/Jdt34
piZ3qy2N545PcCjo8Qyo9veKTcmjFhplhGz9AS7laN2Sx0RWrmpMiuEhMoNCAeAV
7Zo8uagbuLGUoBqA+yWJK9T3kZJhIPsTR37OUyxHPyDXkH2Bf7fOEYzkEGs3eWLd
8o7KeRhpzv2EEP2yvQZnWB/eSbr/MFDU2vuz74DPWeVqWy9c7fjU/nyRDWGmtKCp
ePnLVljCnWIycs25KjisAVWP/45n91hE9GYRbV9iCxVw/uIGG2tPPqSoLUg7IV0P
/ZKUzn3hF2ttDVPKvLG8FUOvvPGZlrxVNvD9EHAAv8qYnS7j5HlgMZ2ZY20NrTWq
oR0Z9E85yHzTrjzatcufkjk5SEGwC1uTr9LutjAO+HsThyZbCk/V1OIO0LnGsh5V
O7wDh7XusBVFtEELwocb4B755GgoMOMYogygekD9ovBKsrMSX5/l6X7q+Wra7+WU
Ld+Ac9vzMfv1x9fs8+PkvISuBGpq3ja3NzsLIMxRtixs5lf21CgJyuoQvyUL/5RH
vdSVou68O9jKcXSsv/62g/2h/+mjXeP/WgQpyllY0oVtQtxYXUdJbXnmGD0sKmYp
phDUte5xfKLZSXCzhpzzPhf5dY58jqhQMc/Rr7VHf3+wxxaDlbA9sE5Qm6W6MSjs
gIMmXyVik//jQDgtBcNJKH2ulCFf9S6E+N4Rgk6DXQI/Lv62XRp3FywyOpxmXD/X
Csp0mcVJ+D65XooDnUUX5ncqlIWCczxImPKq+0Y6YEdZyaii7kyYWJGXtSxDotNk
M0iJXwjBY2lTcBH6IJLpRXn1nNSZFLC3IbBdllUpA9KOSzC0GQz5iva69WOPHfMi
YDPt09T6VDn36WImBfrDoN9s07APWzse9apAzzOofUEDpiLSdP+9uRBeGx+UEWwI
OBKJtMqV+oubczmGePPwMdzKcfCNpndNikC5miF8s9ytLyYXwwqwYoVEdS3UdoFF
uxLNYcaMVdVR61ULzdm6Cv+R1+FIO7yjqDIdjCJOTDyY6fhd2Skp53TmzzJ2BKm4
N23fSuwBsdME996ZvgBa6v0+OdP324l9O+UMfnI05Hf3sVk/qs63O3kfJvOYyaNX
H7G0H7aRxgo2qm2rSdsnIyEKmt0+YYocP4sYEcuVUh2iRx/uJHHrcnO49JGM0X/p
5+q4F+HHP6xqoSUheAAr7Ii/8J6fnC4UZo2/9n6D+vWR6wauVskuRuWQg4i47bPX
vwVy0cWJh3OZCKJKPs/D89NkAVYqNzBG2NtDGwDalQrYAaF59abU3sJGxlbHYsXr
UWc69iaGMrhjRDLc0QhuoMgRdhKRp/dnK8ZPfxRa2AsZr7GXYWo/JUij7QurwLqH
PFMMbNOEriEttkWbJUrTMsyd7J6xCNIfVI2bFM4wGyMYZrvawIBJGJxojBouO8En
QV+9wqQtD/MpJ0PryC7c8q2GK7TTfJ/sMtoZp3uhxe6wXYbWfQsM4uD6FyXlu8Qe
a0Yai8SZ6f4l1gVH1hwH1pNN06CoD6sGEXJh6mBGiyw+KNrb1m+uXFqNM0r6dWf5
8NQ+tt1JiXbMWTl0scz+OdYudlJWYqTITqjslRPIMwyCHsOEFbLx1tFX3jB0kbnm
ACi5rewBBB3L0GF9XjDterg58w7vfqNO7qs7BovAb5S+IkzSJGLRzIEFrQYaiwvV
a3D52m7oTB78PXyumsJustqNlhJ5ZtGfEBdU02IM5mCpxtjG5QcHKLDIA3MEmRjT
1rLhMsSgwXFePb74eWRwXtC1ChrKO4M14m/yNOwTM80PBVbWXZoAfUDGNAj5LptW
nOydsPfXOWl/OCbkqJGLapx66xn7v7gr0FRUD1oEXsqrZ2374bvxbJFn8v/mjqKa
iNBdjjK1KVaST5uCjBtxFDXxuwmoHsBmxIh4chXEyimqiDqgZpfmoA2AWjmSyizw
0NjR44ewgGBjP9NI99hL7BuovN4lpOCg2YvENmJesF6GKaSWAwp7UB2fA6Cce52L
t4vcSQ9y6c9vhrT7lc3jkjxQHEaf7tMUVjVzgdAuuPs+8GV9fHUhu6OmCieyS36+
ms7DtZfYUJeGnMZV91Wx/C6inssODK6mD7qPf3sbHQTsVlO6PW+/bT8/IBp8S822
Wqgrv1ckJR/mdWGDTCZaF7/S1TwJtnCLfxum3Eo+7jQjTcgH9DP3Y2RAK7C+VBYo
GDoz5bTi5nrL751B1+IoqYkDXk2Z5oOcnVomfDpbgJf95xFRpDSD7ijYUDTMWVdQ
R3yrgd/8V9wIBxBaA6oH9TSPS0d+l7G1MH4hBsjyvzSal3nvk/p1hVg5DUDB3nTL
UiS/DFTjLvDPy1muN4DdjqlWP6MnYk0yRAsqTu5L3E9dI1PcxtCkm62VT3zsMVEO
pmI8lOwk75NTkCtvEnBd85YdVakdHshH1LGZoVTrUCpNHxBmvMoTaZTIKL93CxqL
VGzcM2FJVFWuln00AxF/Gpm06IRboESo9AfJicvvJnFQWVkR2OpVYJ5bee+lU8ev
bk4BHZ5ebQ2sV6YOLYJKZCIlqZ22w1l5P//CjVYER0CDuRsMOMCoqdaudRD35Hv3
Cel4k82nf0wB5EeT1rO5L1vsItVKTmwSCIqUAE6g0hpxqUdKsq0ow0/3qaHXxjLq
6C7T4nkHwvTqUg+jsKbc/Ue02I/wm3v97JuKBILuxuvAxV/1Kzoj2sY6H91TPPxk
l/TtgMrw2rseThj1Foq5m7wjckLNF39FDnUjiHRwu30nHc9R1Rn8bbT3boX2DR8l
upw9nJuruqsaovskEfwH7PdYXmQPC+X/wamMXI4gz86VRuutEp6pijtDTALqgxV+
N6lFy1rHe6d+mIl+8ZQ5y5zCFLnM7Rcv9dZ7jKObExzFkBeleWrUx7mrYFw5ku7+
2Hp9e18B6cZr+DuGaEHj550T1bpoCA4yBvUYTpJfsEOFEy8jmpxBXESrxb+KzUgx
hPo2pLtJWU+0KgpnAiEi7cg9f0XZTvffjoCkeMS+eM+msAPf7V9zAS/gcOnLC7Ji
dili8is0Hz4jvtK3dTFoaACBC3PLdXoH5xTGgZWj8rw4vz7a/6ykNBnIEt0Exbcb
XWJYy8NwDYIrjYIXcg7tF1Soj2lk2+evscWOiVgkIT0tH+iz/G2Z3m7874M6eMch
PqIMcw8XB24eH2jMQ/TY0+Epi16tNCPfTblfWrOcjNawDwkuemA9NUOMql6iydH4
Biot+1mZlk/3R2hgll69NCKBmFfzPnRjYoL567xIQdtLi+LM69bNe2dpDwZ07bhD
4dRyji6efJdMsxTVR2rFBBb4/zPM8f+6Yy46FXUzVBCfV4qsJ/w6k1b8V3UxZziZ
iWtqOzbenfMvuNq8pEdCJjly98qRaX7Vo4fjBko4YxpKMSI2ZMbAbQZiE1yfNNCc
sHTb+dEr0kVcHkUjzk1m3OxRBLLjxlBWNQ7S+GnTrePmZk0awNjmBqLbBqbsFkmH
en/C7+S8RVXZP8lk6gjc2XTkFiLK2/tvg4Iaq+CNSPYRvuej5AGL4qo+YNDb5RZX
1n1cDm0adndX76jARQNCQx2k9xdsJwo9qRRRq2NXtiNugzzMcFAjvA4/XEy8iSMB
bnmxX6P7Ahy97Uv0ZcUc6HfUvz8/EEFEXZ36C3wWQbUppD2EX4/7fZ5h5q34rEn8
kIQauwwQeD0iI+YyJzgDvbW0AoglbUODmpdQwcD4dIHzTJvKcMqM+O07XyojPbFr
ythJvQBGezdKWJ0IMm8rztNadEG2SYYKtqv2dhyl+ASs4GuwA+s8TJOkSHkw24Is
Lk9pS0+UdwQLMOgBtLWMiPSEKgyVFxhkCYsIAJJPZHuXdY4j+dOj5ThS2l7MfkVa
5wSO+r4QirTxQ5aTIZRx/LAQ6NAmU78cM3FuyS8A3gL9mgHxoDzxW1CMGm/9lgp6
Qf4BUMfTfgWT8i5+OUFJRWRoq3aeXHFaIKLqbIAsrcq3MrDN4m6mjsBJmUir5oTq
+x9zgxjM6T74ShRXhsIqx466jBVUTaI69KjQwrm1nRtir7/Ut2+STWRAbBH8cpJ2
hIBYeYYSBM2TZ7oJ1S30gDJSW0pBbAvUkx10hwfwautU5TAik/a0gxcIpPJshjEs
Hohh3/wOOPwXEe0rRIbu8TVZEebi8OkrCNcS6v4TDIwLWiz9UcvpGyqAbdS5kK6I
cXucZuRkqP/LrlK6pIU5SceV47mInxakcUG9dV1cQ42cszkFwlKeWck/b2oADeM5
FRSUDEXpWBVpF8QVz8jYJglMZxUqpNkPhPkhFZYwyMWPd0hvo8avgcOg+1lpEUMJ
y2h+KFLIBG1XOJbKFE5qnUlhUS5Peo3h0bpEDabVSopDg64PKsDQdIoT/2Ot3f1c
kHTbKe2LOipH4MG3SHemCETMIX4s3XRCsIBvySYKMiUtMOwLuFTz65mGUS/Pj3LD
1YxZge0W5wOt4zioOMuIfmfAJLfUgL3Y38mqqJjy/Dil8u1LoF0HvrepbB2W9wPS
87KIHQgfWXBqVgb4ePNQXjyFoKoYSqSmgX1yewegwT/Ck+9X9E1kBh/ZJpaIX4av
P9dyefERcuYlostuljuGIwn6qbwXi9NXS3lET5718yZyaRD6BKw67fAnOBmU//XK
6quMYQx/kwDSOkP5wKRV6+di18tkaNTvSfpa6QbK3AMqWaGMIFmVrvMXcwYmuCXm
x8G7/qJglRlTBzyD4Wtb0zl7aDMenIdNTYfqJVQ6fpII2HUKxFRxdFp5vhL51Kv+
HBrbwVDrBnNaK69ShonaNwagpeH4i/AA1U078gJB7j+5BZNbhrnss2gX/8TC0pzx
5iGBgJuOVvexH9VCrfPYYPcKuSBnPnPN3IEEPLcOVrrpFrVUUOkqC5/9KqXWEgbM
3rJ69QiBJUjkOD9WG9ctIQqVrmNiLMqqa+hqMFQomnCoEWCBNRiJcMOQ1Ju4gWY1
vKVv9mbgxsb/Jyv7s7vxkjTVs6X2Hx7qSckEv57C6L0YLNq3nWyaBZuiv1NSBTd5
+LZdJC2+d8RV3eye6kfBMELaiWCmHN/bGpTqKGAIBoo5OkfGKeNFEXKNF6LaOBEt
/Qj4oFvmyXiSc5NPgS40WRkXuTrJ9Pkk2mulxqWX3EYC/Y55GIU4qDvVI96GdBdb
jJ+XORxFA1MVLAlPAUt2vmf0B2vRYRUKpMdc7dgAcPjxAd7RBQYB7RctMHWeQD7i
4KVQ1WJSx2MA5ZWV4SGZUBnRuaN8GdAyBKY6i+9JrkUph1mi7IUG73VYT04fy0xe
GXyKGyDw8W4O66AuoZPpVKPfQcaMIF6d/5ZP88SUCfzn83FbAjd7B9m2VJGwU0Ig
+WiCZlnNond4Nm6EUQ9fS81Kndtuju9hVTjIOY3GvrLoQxxsqq7SdBW3INdfTazQ
V4EsOWQnMHNKZsDaI0ILVf9ler9Jayf/f8jXWRvhE+tB+r41L+P0LE19DfQVjE3g
mCOeNJ+t7cUojfc6TvKxNQ8xoA05VrxRXiER9R/NsCDvMRtKDGYfbz/jFnV27iuV
Olr5SiDBtIU9EIGD9gd4cvuDO9vxoXIgcTjLIEHcLaHzOTp7jJeYbQKKJwvGATcK
Rh6mHu4F2/NLwVOCH9OuTGguFD+82JYY3dVqZmEIbkQs3g+/nap2J23wSvXfeZiL
eaTP9mqRqTsGVeMsv9Hq0KSxidnhs7qNFGjs2O75bycmuumzzs+1Ot6b5VYJMfd/
gg9UpaoDat+zMTpfCnlrSP9nfio6d892grfwHcMGCu7fpnUYEjux7Xw9nqfXRHEK
aNxeDNIDs7B9TAEqRM8BbJN+ADEPd7H/rOURS6YKabBIzsVJxKA04q4Mrd0WHkxC
1ivWblSl7qaroNGUAJvGpQDhPGHRu81TFr3EOne6ZlY5ciiR9ohtt7ndFkiN8wRv
i3KXT/WUTyDvm/EmO2HN+WUwo1QplMDEz67juV2VF9PEe61Kh+IukROLfa+LzOSI
at3nsm5inbhdenZEGlkvWvTvA8MGcNNkFGQ/6a1zhbNfm4mZY2fp6JulUCtfFYtM
c/FelviK4yRGuR1iTINvVoCbpODU2qeYzqnjX3bXygG1+oPohxSHmBN655St2PlU
9dLdcBkVPM7Hw+NrglzVL2iuTxGYlqqTL5z72PAF6yv2ulyqQ1wipe/qd+cf/knO
AL3/C1HwToWhgiLfMOM7vBiUwcsUJMXI5NJIELMC0A2k7iffG42UEC4/WjwNQX8q
D0wcs3zVRgch07FPC/4Zkt0jdJpeYMZAAQceyMMwmBAaUFbUmpRKbMuNXxPy8Ibb
gOvqJaKid12PLMNaQphYLoiEVXXRc1jjjCapydeQqg5/ykLSLg1354QGxdJWu9vJ
TqeRirbQmHAZBfDrqKMIJrc3KuH18P9zEhqSkteu6cLkEBa/IjSgO7k3e11hWfqr
hQUlyap9SOJR+5ImKPLbuBqM3arNP4zK5ZdR02T0xrfSwddnrCXHvU9T+jxeTjnJ
kk86H3PmkRY/yb2ORNi11OFqq/7ZNUt1GlsIKU/SwBpjmtwrVzI2TA6Z2OFmFake
2+7rORV4HuPivEZw2xXJIzUQZkKLixkJ4lOS/Hu5LiwNWHBOmcAB/K6rAZ08zQC3
QdsDtZBkkYpO1i3TLRiTi/QyH5DmT2ZLgTPc3grbYonF5T9qVE8kzdzOKzylJwEy
tKkpqE/ln1sNM40HaGptNIKesCTaYIr22pT/TRIB7VQeku5sSE6KVFqZZbOELSRy
GR5It9Ak2H3YwRmA1Y5mhmueYoYoPLWzzHJ1f7ChtMi8CAMtNte74fMPdmZpAHGU
pyPgJZx1erncVNEt+87KsKEKtzZJLPRzmoqi/5JuOOUE7uUNyR2quwr9jVn4afeC
idyYWK6ZphmpkNQsZYSVwQEk/sEmVmgpQCkvvBNe141UMK97oKi1xhi1BkPWIelQ
J6mgXmKm6Qqef0PT8Lm/UGiYX8U0ckpPs7wSObj+133ZVIt+dk8OOC9iFlkQ2YyL
Gv8Mh1O6cTWwy6OwQvnLOi4GNJJctwHcCxJTOJvQt3h8W/9aFG30a3RTHcj4C6K9
G0aO6AarfRKjGBUXMWkh5tVNVAMEWNltTAMd+qG4BQyQThR+CH+2kul4j8JAXZes
WrLFusoGEJmEwWbznwyVSDm8G4180gFkarLIJTSUbS3UWhFDJYF2f52c16efQcIe
06kBolYBAUi905cD30d6K6DR706n9BBbYZsbWbQbbilboh90pL8swYVNPQuCcGBt
dFRrHPprClH2elWtDdPEbWw5U2/TToiY2aKmhpDKmIJYMNcF9Q3By0wIjOjsrNlB
z+ssh6yCSmLhJRX5yvyM0IJmqU/difZjgOMrCgVI7/uLlMuF2lAAuGF1hebP/m+X
waGkt/BRrgad13SHSwqXjazrgfTzJnBdRns0ltk723KYm5IjEgnjqEpwXlpSzxcL
0uU+L2vfQmr7bf8IfGVUy9jbTS2XLCXzU6i+etXBu7JEAQhrwczR18P/bPtfuogo
hfRMgt+a+HC8rwx7vjmSyHlCX9rFhQjmrmYZ5mKg34RsaytZTNH2iCcUS0xjhl/y
GXngTfy7nYSnt8WczqAr2ARQlQyVnCJXlmpkTCMZ9+aHl1YRgnTjw12wHibM2aCD
Aknm8FV7fwH9Td6vIDkLQJE1n0R8ydLZgfNr2VGssolJ4zid1kB5Pq5dxFwhOzk3
DGEzpwsy9O7LxTTo/ZhZBPONPHyODS1PZ5A1Nejs67mn9MJHfvz2u+YwkNB52kAl
z8Ejb+zxk6cUjv2xOPeT8t6kikf0mrxZFycOmuSXj9o8Lx3zEBfDI7pGZljBW9vf
MTdOq/KIgsTlPXJrMOQdFRxPJPMzbG74Tk7Xwh1PthKut4xIp71ARY3iGVZ1v4ED
VdiFT9x1zXRJBW+8c+szLBGf88vuKoQAk2bGTIsuc7QTpT/VZ8UElDVy7bHAFpry
Xh462TbzTLEpUqjKtXUfxm/fWE+dkOO2W7XiFyXTSlXF3+7O6UH1m+DpKXSgFdk2
wa/0GF4tnaueQtipuzzcmAS53TTokFd7BW9jiJNDBVZ9VmLZCyBqBxPWLFX6P5gO
ouzkvzb4iL+5eSeXo1tUfG92IqD/TrnEdIbknm+6tHXAJlWPvDvL2VIiPP98Uojz
QuML8ecMczBScBlKZTIy4akmW+kGFaJQ3OaVZCF4WyRPtnIcEwpx0pfX3Kh9qSqp
qORkpb86v0ceg3YgBaIC0LJqNmIrtyk6b1PMDVv9EibOe4vpkHi1LO1Ht+EwMYL+
btgaEEzBboZaCmBWZK/Yph2mhFGUs9odKDmakAAbAujR3d46iULexY8m1tc5YtnN
VAtynyvJbvzOs4eU7KuCu/LHl7bVyZ/kAux0ZV1sHDNZQNS17CloBdzpxgwdxKqr
LVlTDr0dNZl9zXB7gBYaXf9Ggl5Rp8PawaHc9oAzxniUmAE21x1ewEUKP+xd5WOT
vdZ8O+cKgSx0+zzLTHRPqJPbxkotzTZTqCBblrz2QoYD9dWUxg50b0jKkITorGKL
iP34frnbUpEFv/kY048Oe9bodessEvBR/zJUqPNrw02FkcEdBHOE1lJAsbtm+bSe
Bp0GF+KMDOG372U2XHu2nluC93FE03A4VzvLsmJYHI+ZxNpv6Sd4nymj/t41PkfS
+dRInQtfe1fGExHydND2Z+aRyF0xy9TcNMcU5dOQ8+KqHsmHE4slTJ8HdqawTvbV
xjSwvfsHqeUtcrgvRi1e+fcfH+aouK3rn18lo6YNp8UqWF4tgxhhenJcmdb/3KMY
X3wlaVk7a1K8Yb40yP4Vw4bcQVQcqDGguqzbWktpbS1cLHm1zX/JsWxk/gO76XB+
KU9iX0x9qMeh/W1a5B0dBLlTW0+G19NOXEP4xaWpeZHE2JoPoxvpZV5AIrajpWlU
nAlceCEGTVHZIkOcWwVlS7YY+q520aOXXTXqnPiAaQIPUjdE9qvxBb0xcpz1eAxy
iwdEKsp2Yn2iKOcl8r8LMr5KD2KKqnvQyR6ZgsH20SSLevHvGoQLuOBy2C5kFY8L
XakZ4kklOPbRFMrkAdAOCv5X1GhDzUbehf6N7GboZUdKeB44JJNZoPRcPX6n99oh
e3MUQRj+K2Od4Uv3bF1p+jIiHWJJ49GjC5Efw4JcFNmzznEt+6rYlFTgWIv5HeT2
T+ukwwRviNXJ6r5JKr2A249sw1Fcek28xgh3oIWxn0NQU5EImO1bRSC/XB0CgztG
StG6IJ0j22Tnhq0HC2ScK8QrF+hlYMbux4qjqnyjc+9xngbYbdiO5povms6gfiJx
zQRNZJlvwkbcC3ywC8O03JEHZsKnudeLAYCs/O3CsbkCbiNlWHS9wPwErIWCrY8J
5n8odr3lcuhzRbwfzf/jzURg3+RltvgM+753et6BnW+mTah6e5zH3X838kR7BEOC
6WI7fQept6lMUlHs8JWeckCHn6hH/SyHT7qCF8wb2nEnhLKXkUTwNHkWbGfmEusP
ei2cpX8BL8BeWDepspF6/WRnktAFYw6MGFn90DV7dj1BXfJ6BWuynQUFM41rHJ9D
S+oWwh17HwXrQa3HUC6SURCUZPQtBPQRnYQD+YTsG0T4dPy17w2AzRByKQwYjUCt
BbIyz5CQkvvXAuJwO5+n9Bc+t+EZ9u492gX74xhpOW2rEmbGo8uZsGkVQT3UTHYm
bU/XLRzWy4ERbsUbCbuMT6ZCym6kqOhuucvgVWG5hEsbonX0zu72ze05oXUMAoN9
7gsTjvV/PaJ+U7XrJb06n/yVSLnB3doiohIEQXhOQjXOg3u0S40+8gMv7tmMC/0o
q2/HoStCLh5Y2Wzmnf9JbrdR5wtvgbX3T/+CQuFxiMro1jbisOqZy406Z0jwf7/r
pM2nCK7+udIBNDlCxNJpaR8UuakV9RK10PVUnSx17QKdbDFYOlZj9yjcdWralhIR
Px0TycJWPOtascIvNv3N7Z9Rv5mCED6fYdqQFUK5/HSOmgrNcbJ/BBEe2hF+EY5C
hpoS2xnWd1BKtx9+RhCE51jxS0zcjGciuGYNXHkszya9QX0Sjl+v+tyH8Mfq5Bno
cZlgvFlO3ipCb1xJIXimXu8swFA7PczL/oN05weKrAGqv9ho3PcFqZcONeHzfDz1
CBuSEspKDbIQhsQ7xKJXmF/yT7LZL5mPgpwOuhFzF9YLamipoovuwF0yRxhXmXr/
bc+04I1kWTA8JAoEwpDSP5LTZh5kIFebaLvBk1T4MB1vcvYdlM4l7tgZiu90RlxC
vEQg3HBeQRcqOKhqc8x7uFQx1XBl8cvw5+91Nh1jMhF83czAJUZ+IWZEnMQ2Tgit
P6lxE6ZH44pk5CeKpLzg24+y/c76Rb18tIzyH5whJ/uyF6b4oqMnVtUIcCG99qtg
3u6FK5c+ZB6fbh+xmf7wviWhCImEL2RbXekYgJau5LFu0dmw0CccgspV7xa5EZJx
BM+4SUoZAI+sq+JJLKfzxKxDK2nuHkWNQyjRHEImVNNF7ASKOhlCoTKLsBFIIDe2
XnCU8glgWDGjXRVspjRyoQWB+J0oatz0gfRXNFIb5eQ8/12dqZ98AfgEsDZtUkDV
j0c2LY4IkHv50FZv1mgnbZYxzbm2CYvoyakJjioQXP2iAWzXLdCybcb2ObZGWyXj
L/D/q7V/Ia/pRc6ttpfXYLmIGN0vizNwKjADR+B0z8UT6Di+O7nRhpE3yVvrdDDg
WQ3vot2BpG3CF6ID+R/ymvJqiW8fqIx8S+ZwEJczCajavz1DykJwj+KKKSmuJL+/
1XrNDmA+xrKg2MrJbwvkqV3AdbffSAe76u+fogUyvvPEGWFb/is9NCd4GwjJ0VkV
Mg8BBQQB5xZCinOF126TzR7ZJYRTW8RGpFEpxp4MjCXr2lEiK9YwN0vINarJZ3RE
IfNvkY57ifAmqymkEQ9BDUKJsM1s4C2pc2NVQ93m44aNe2pPdhkaw8VjLVxMc3HP
AqiFKkk4/r7XfKUXacmX2Vwpq5OZRhaLHrb1TDsmzEo6E7zEyB+27VyAJqsY3ZsO
w56v+3yz9t9PFEWCdbXvmMaWxon5aRcoWit2+AqktQuGn1tG1ArxK0D5x89tn0x/
vFYvA7JHxL7n4yYpXo+ysMdzr6Wqw0PjwvTE4pOLXaPIPV62f5E0rOcCGrK1LZxD
ceyBhWdjXVlLe8qaCWFpbKNjSWLElFWrFnFHAxHB/Q1pt+4EzjGf+vSf8kZs1udD
wxJ0fxt+X57KnHBCJlNPnTw5vpylCYLrwXN+mOOF1gaC0kogvRSTQgcYC0jnyQxw
/d+00JC76e8Ts7hdorWKUbz4z9A4DFp2LZcpJodIm34QbNKYtM9s0jFVPOqUA4yP
lw/ld2Cq5M+SLK/BU9goTVaU1kbAPp7E0gvsogBsjho9MXG2WyFMyGWYtk67w+53
zuCqKBUUcM/VwTiXhVhh6uSdhoyfeBaVNhIoZsIlMyPodOxI5Kh6bqrdlnoBudQZ
qbN9/WGFZs1/+KVWojywfK4iO0AWNBEvr4SgmUpd0EzCsHH8oP0D99tptW0DV/AO
uJG2laFbsz1/ZN4flMf9/J7+u72JAJQuzxeTejXXiwWLUqJyoTrgk88dSKHleI68
bIY1EiUKj6tDhBaI4UKskP3grOJA//oHO1BKyvCWFd1HGM8Hb74O4J9iypE5/8mP
YCOjCZDZ2S0AHWCTu+BHe0PepbWOtB+GltM22wtRulwOhN6B2U5T8fy0E1eAPh/A
s43gbON0Vhfur8KIxq5jKAjtBblRONg/iHEdilc8vZIHDEyGQqr6+rdES6Aww66S
eYftrfnYbS/U+X0Y4jxf+TCTC92h+mcfo0ald1LkaaoSbksmEg1gBhnrWQbEBD1e
RxCbN8GmS7zJ0RpZXIYJe7jMmwDHGXaaC0RV1JDsnbR8sX5U+hcvWfcKCtbgJjyE
rLGIsoB5613JKAaEVKF+BocgYvXuu1lLG1ogsLORCvApQkNWx0WN+0mpJgnP0/on
WSKoN+Fnf1l1zJZlP4j4ib5BUEGhWaVUeoA9yDmCfIL0wEpSlDvcJUZxvFKSz4nM
369NoVJkMLveazfhl5oQs005YTpW/lKarS9FFf6Uq1zYbk38SdPQg5NclkZHJQSk
px3PTZhuCfhzAgwki9xVPWKNVJNHli6OWE0BWKNqK8ckhsySPdl9A0s6Ar7mHW/L
Z6lK21KIJIxpRYX5eKx09Z4JjYSYLyBDJLnW6nGL8K56i0Pi60ykngUni48gZUEm
DvMFAb3sJCydsPFyaHA5onJd0IO235e9dsoGQiUtpnsHBV6+Kbqv20ME6pHv2i1y
S9vhgRLwgaM/Pgtu1yR74ZeK/KunxCYM1TY8ckjDcU+prNT17YmwTQTuLBWL/MFf
kRzJmD7pm5t/MVrjvDogzSxiLhGnmQGHL0CT2izLVOhaUW5N19avxT6wz9jVIk9E
/H2vwy+bmflGJBYxywWrj3WwaRuIfoalLDuIHJpJuenOaewpnL3pnWuMEkf9Qw46
YYidsEEnB/Jo5H/XJelUMoCffo+bz+duoHyYqA1GGWMuawMRKKDFTi0x2JTCV4HF
Kq307BWmPoe6t8fomTscYnxJC0QkyBDxlEkaNJ8owJkoxtjz0CjH8X8JMEavrZHl
DGjHa+Uf4DjyHzhk3w/6u52cTHlp/vuqPP08yAnGojeXH7abQYrLjx1zub5/Qa7j
yX5qvBDH0XayFiKlnXIT26s+54NTDOMejdrl04RfXjMIvUzkAKTmv1x54nUYgTwC
RqX8o6oNw/O31Y2A8os+oqedsr2SCpGNng4Isvclir6AWbXlPYILo5ZuekSi7j5t
BC0xWhPmdK4sI0IBcOfv87kL00OABXj+0HcAkT0UyKnlDr3evlBfglt+yn3KdHs5
1uZoViqA9028pcizozutSForBjM+hG6L+v8l/Me4cNnNUbpnU0ln0D1wbaDkNV8p
lRrU3K/Q/p+ArSFALOeUATloF9FnA6rsT70YT3PiyGE2q0T8obUCgA1r3sOBC18X
KIksiDOnm8PClko3QE4eP9W7w0WFyEiSGoXxTduxg8P1bcpH32V+ROfuG9S6LpeV
aleiDqkdbdnlDhADX1Nr2hQOyiRfWnZ7QQnqhR7K1zvr9ye0rCXNu4CsV+crdaJC
tQdpGEupRpB1G/+LYopCVZDU0533gELLUo9p2AJFzJiOaGBu8eudarNLrjO+HV1d
oFcn4UEv2zgVXdWxNOukvrGg46tCtEUdW2Sur9gZNOPjdDX7k/izyW9k2C/VGWJ4
s+16Pf1Srv3FykCaxoa09c7i01vGXGO+h7zGFDO+ajeCiKa7X7bdldswE68S5j+U
/lu21/RdEaVZJXJ70juqs4vpixebhEDnSdMhCqX4AHgrmskgQwfVwe7zAhgHmt79
7qv2WtJUvD5W/qQCkTt8CbTIZvJyWY/NAwlyECWNqzjnuGcEFJf4lwlbq3uNlGp3
QcNnEmNsmeN297NHKMqJh9f1RRpMqbpDXtspDalQlrBhb/4oaO4lc2TdmBEmp6Dl
rDzC9jbC8zL8LM4NXFxXsqYoYzL9TtKnJdrcDOgbVIJHF5sHRCtdGoVIcMOpsPF5
RvMrRDFTmxSISv/DasYaAg65UUKgsBrJfySdGfeAgbP8sywzhwaikyZ2IlHi1T6G
w06bd7J4YFKI6alVdGBNlHNZh2tK+2sDlYSLcPGSjVApA3tDEsMIzWdHZeTJzO0Z
Nuc96pI+qdqCGpvOUexVNqF+9olph6gGRZiEM9dGJEeVyDV9VzRT4pNSXmTN0zKv
NBRSKUU4OHLeocN8UxyJIDzP7TLzkRzPrxJsg+KdugdpGK06LnhUpookS4eMc44C
sujnhMlm31Oi9zcEmaXYwr+yrrLZFVeubvRSKGQ1qSxeFns2YU47ih4Gm4gD4RBN
HWjPI55Uc9HvjHIZ2Afcv2Pf2Uzyj7XXwmRJaMBmGbLAkUnM/paMXNGbhDhwQdTu
U5iANtbKVrlATnkzYGBq/MHyYzuvkw12bAIH7SKOC4FWdu4yz58Um6Iv7nvg9O4Q
Nr0TQbgiJJ7pYOdXD5Y7mhHA/XPUFddAEAcTov5AdbDcKB+bXnRELISreP+WKNlF
U7aa16TWRRLAIN7zQTnb2wBLthfyJw3qGxP7lrf7SFi9vgG9Fmk3OG3cwq2R1R6x
3+cZZ5AGqI0NAWEBG2dV7+hqtqsp1u5Bp/3hyV2LTEp1LYmSi9pOZDTKaGL6K0/B
uRPLVqAWHE0Q9Pnbbuj61GDVX763UEp4Wb2Q0oujpGie+5Oy7SERAZb+nk1O5Id9
5BaUgWXHHExPOUTn3f5Pd/dLr9n8oHmrm1G+5wXOHThMyKxg/m8GhKytk9AdnFyv
sHw7UxNHtHschob3z9PrZKx1NFIPQBd0sXEmZn6grBC2A3W+TntGQQxAipiA/h+7
cIcxmtEuWPKAE7EnBvLGOpdxrmPWFdVg0veWv+YLi3b+yMOmozxivt9/02SMdNYW
cznZrbWW7BfL2OUiRG/nz1rWC3uCYAdI/u22l8iF3KlQJ67JtNbym1F1bKoiuJNU
RLrTY/PUwnNBLFnW3FmOLj/1GlFu8No3jg6pcyC2fB4QlwBZmZLQ781QOBGdcV+9
b6+8iuDsLdspj6QS/ebW/bRz2gI/nRQ7FxSokXXdYofauxwpp5Qwgu6Fy9v8g1Rn
BUASLy40SbER+dZbedKjUxJAKIjVIOZ02oYZ5/ih6o2ztdDN2aHwFh70/JoTLI1c
VG4L5BtkbXEdhY+Hz0MkvvAsfPvsjTBJJAi5w3ofDQUfZK4RrHQs34i3mRpRvT4U
nFKvaS0NgamiodYNgQd8g4IPSoxZ9MnSW7XC4mMnZpdvfOvNt+51EA9AMFoMD4iL
HzIINoSgy5jQyWWBjXno592/Q9JnTq+QjNe+CHSMvmNmbJ4Kq0vFk+iUwmtG0IIM
FrqO6zbxX5Iqv1hMOHVrUEG3gOT0LKoX8O03xe8QlgaH+lAk08I9nwJk/p/rML/X
J7r3GUL5BopmbnXb8fLoJBW3BnnVH/n8uHnZdhaBL4WVvpf2zJrO9h5mGRjG8mX2
bqMI+kI8ibdwboWTR7cPlzS6VmrOwWT67Nl8oJryaLKypy3he5LMLjhalelHoK4s
SrujiMmJU20XIRqrTs72Lrv4oQe4lXO/PS8d/xnV7nQAbeVTJvtIP58qpFdzPYdh
WikzjehjM3IRXlGr8h8O11UYyxo0GDUaakF5SHiOIJmPWJGyYPCpIjGSE0cSqTK2
94HLOjcpck0d0IAvTVLXrIgqXY1wr2XdHi7hSOtoZ47DGRcbNUjBAo4YllNemEQm
8PjDtXKoSMx0Y/2jecov1g5VczeP01FXENJjanRbgpPNjKioLcQ2MDZ968vRTD/y
/QqqAllN0S0twO4A3Rg4flh02y+wklL3zNdQDw+oRmKIxC1YXyUb7GkjuxRCJR1S
uNuW+0uft9L11i0y1C9z2fuIfQBSgx7gdMiCo+uMFwTaB0fh5sZmhZ7hCrmODy5C
J4FxR/UjwCtyf6U2dn706NzJ02Yyxd5YFuexRAEOlHjGfb9DmuyVPLMxvS8tyEkj
BBu61libMyCpEOd1K87Cmye1CuX6wHKwiL3YcKc7ER/di/zKuQ9f2ufHhXWlOqPT
N8oKRcZYr9dHej12EnAA3IKyKb3wleA2uxNNVDCI//XnH8g9Tmyp6Y60Cw13sBQ6
LnF4trs2If5QSdNbrxSuq+GRguMZMaAuMi3hdyMOCp4rjDEbGPjXLOIsYyK/ILT4
L0hnv5EYmmO1Nyl8CYS5NM5u4XkVqm6JyLdXgIcwTyv0qf0IJzpQHkB1nakZwArC
IFf+P6Ylplxe/0ugwdwbv7A1FWxhrxtXT/SpjEznBXPbeLZb9b/Ee8pt7KoYhSFQ
XPSASrrnvgCFhwoRCDNnuuUENph0ZWkpgTywAw1adnHy95cNN0ebbZUiEN0Kpdqm
hZeTY3OjRwf/bQUYlwUnL0Ep0BlB8/2noJzb8ullhERqIpHOwqngzzSa/mmEBKYd
UJqOkRop6pFCHjdONNxRNYzQB8QpyEzQtaHTIOTKj6Uk4ZcWvj5Qj0YIF9zYYD5F
MaJIoLTyKnf9F2I3zLdRPZPTHjW/+omHwc+X88xRShaChkmQ2kylMaHOoUdEz79a
EHGdoLa+BLabIBCAXJFgFXYXi0c0qjh8EdQONzPAmVnfYFuSGWumQcR6/w8EBLbJ
jSdnfsxglrDHTBWXATj5M4Ulmsw363QOz81N1wUtqJwGr4DVx94wstRYbh4UdAdv
F3tEyfcCXzRpE4P15V54GvU5mi5lx8z1xZ2fXDOIma5yQE6PgUjQvnUcUkOllLwY
fdHcuC2jHYPVYTXs5sf4zPrPWDLgVsW/pffR93Qlz+eJ25v04KAzNp3q1klY4wED
fPkb9BnAOZM6Y4A06quZFQspe5VUr0uMayn+m/kbWvn7NPKbYevxO6Z7SeFFcNMZ
AXPYnC6hnTUT/m5l7iiYuKw3ArlYHcxa9znD6akyj1mA3+rIP1Awob+wXUPpQK5h
lmHU+lvHdexJeKI8jfwEXg4zFLX1m88DTpsjvzSPlFojm8BRJaiK59EiOWDB+Fdf
eLjzGWyDvkdi7cU8kdmZGeB4nPimnC7MrRjGzxPVVnW0Bu9HfvTuV8T4Oym/ISBF
q/NODjy2AEusSIOtJPYv+S/mNlmgHa0DhzfVtsgNhqVoSjpOM3jWL4zpidHaGJwH
r/YGvFvnpgJorPc6DzXg4G42OXvx5DWEdIPoCLLD+DIU74B0aXiX9ZlPrDE5uejX
E+HaKXRvNLiRFZGD22qZt8VlpeTjg/jyTGbbNMJJ7Y3QnVJhHYWVMzrGBK5PBkxT
8ITvK4rZTmM8Rq4BqwUxpiTtfiQ7MLWN58WmG4QTnFoJGyk9aLF1Q0Fhx3RJPtQg
S5keNcckzJdxStFxw/2QUIL+zklv1B76LSGcqet2wGOEc3t7SRWhhwIJAoMfCq9T
OJgN1wqeHke9f75MXuzjS1vYzQnU5NoYSo6YVQ1Di3SReAPyFAxIIM+6Sm1jxAbT
PwHTxpWvX6WPeVSY02lR8Jt31Ii3A03zXE+zkCA4CWYaFXVlSsOfCJaivm7y0CQP
xsJ1rNogAK7/opmkcNd8bULJU8VNW6Rl1eE8R6EOPd265bsN3dCTLloAkbS9P53H
8jQjDEMrdjXSe8IS9aYQ28kRopw8X1IJoH4SYwDnlV5OSv2CCnfOjHNvEMVsRISf
vGWHdRpXNJ7XAYIp6QI8OobfiyDmcmhMc2VhM/lRYDezC2Oj/L9wSR90ssJKUHNY
0z/MHPpXXOfxv7Pu/LdlIZ1wkn1p+fAUMUJXpjVrWh3yjP1QsnZS8BobaNSM/vWX
4QaiFRl/iSn+zUTs57KPEjORyJTpoisRm/C7D3dcubDd1cGfe+IGQDV4PJZLe3bb
Ij+x/p8opGHi7zCkLwkI90w61Dird2XcfXxQ9LSbQv8yLQ8o2lXQUoPiijLxgrgc
x5MG7yHUa9SBBUq9ZitzpjX6NC1WOYfN8uUeibX9eIJZYwq9Aw+9oN8iSbwnnmKL
5SlLZtFFM4Mjz+q59Zsiovh5DV3hLH4MQwqPWNwdXOyBLLS3DiIxGuu7YKzbSYby
Ytlk1Y42lPBor6swHFBWe4q4Sv5Tpyz1DXIwhF3G4m3KZj/z/mee+hNRtvyfcKse
Blsw3Y/UBsY00gtvzBllx62KQ2DABHGjD3BU+oQxo1N6p/SfRyUFVRfJTflGwABU
DxgGkPUIc0+bYTCLprOT6u/BPjPe8uQyCrb228UcAEcuzB5mGssGnRgY19x6/oza
SuSY3mAvi0U+pSqTi/8vdoeUzNBHINWouJw7clKUQFuwal1NvJ0Kl+j+hV3Rodvr
wzxtKUkCddSIAWzgvsGXApd2EZdLRC1ZJ/tmny1VzArxGB19px+OAu+CHy6wV1Lh
f9nuYNs+f2xLCLKpRFHdzoSbow9fK9hzv3yWcM2tvwIUUyEby0nOrbN1H1x0kWV+
UJjG2YcjvnKjQU3mcXhtxTfPCbdzY63vLMt/Txmm4OQwbHWHQT0onkEGmO833d+H
irRO+An4Ok+Vmr2RvrKDNUuv1iSo/Ah4TogKK8QRKF9cj82XllqBu5ZesZAClbAV
T4mLZtLPC8tzslZJlNeSB3BHQdTekvng3a2cUvu5hCaT486A8sEyueNn/ABlbze7
mM+ixuiAVssNRAVBevFnWRAVDYnW233R2E5vU8XIsInCtFVnsfLj57mZPeLBPp7C
KSM5akjrAADKimRbAJ0XAh46UMDDEmSBFyB4ZQmCKqRwkTPJWFU0k9R1i88tLebh
goJTHiRMVergVqUgNXd+5uYvVaijY8eTmM5XjLnLhsSUUe+cFoCdk2iqnnwcgP10
sVrzkxO7Pi0zM8tQAy5grBER3VlsR94dBnnhLu2I5i9kz/VXLQW4SGKmvC/TC2pc
c6e4zJhikjs/neY45Q6+Jeeafw2PzoJz5tiidBuNzV/gMOsYNJ6so3s9w/FWPc96
+SX2RTUFjDvrsphYc/ILHomP/yY6EOS6CI5H8OVZhiAFwq/WgIv3CjMvuz/qJ/Fa
6JK6n4sOQ0zui8rHwUzIfYAX1EdgXR2u3fBapniUGptllPPTnPLTT+orrPAqELAk
9qNlWS3jnUG4lVwuQUGylmwvEF+pQXbD4T1/yhQ0P/J7Sj95o3YtjXMyO8uFAXGF
Z69EW++n9wlvnNzGwJpEnB6o/m22xUjUOnwmL/Td8Fmk3k46nzX9htmWU+p824G2
tvZ2bI8F8sQTqhUk8nEBiS4AfbDu0xtT7E74i+TG1WyF84luaJEuCVf0/6OBBHxD
Q8EGCOQrnRhLLT2Iz+bZRZwcAAQNdeTbI6Q4vD4Q2Zv7prxqiO9XbT6cZGreEny2
ZHK+R2xrQ7hKulEuLv1Z+QXoHtDBjF/K3FjnbMWGDtNFN2wl09u1LtMXLTnZqv4h
a0ron7d23eJ5NMg54JHd2PzP/N1KTM41+z0aoBttY7TqjgrbD04Y8MdqtTJZ36ZM
gFzHDdNiUxgC+lIZ7I/Kuqx61AHnjoxZk6YnsF/ct0WyG6/EnPwmQBoRx0ZOcIcV
nb/fpWo7pIFpbS4rZHXZ0fqpyd8iqDwAsnQ7Z+A5GAi5/ckSH3ddp9YAgPsyzn/P
5Lu+qJlsLGgDKZ7TK9uOEQELuK+DSViphhP8z7/hWP4Au10OSXDmBb/HczBU2JG6
S8GwDDwFLPsAYS5vi26DEsNx6TBba2emFhj4bUTIiubRnCA/H86uGZTyW0SA5Bf2
oCRjyrcT+P9FUNo/hoVRKAFjUULmJu9sjJPt60ya1I3nY/YiwxuGsoCVeErdqY4J
6Y9tfNYgTUrQ95wy86siHgWyoUG6ojr0EEtHB7iCMtN3Rt2R8FeCSMMr+qaLy9PU
7cPZowAQk3n2zyvaRBcU5n9ioLdN09DeKB+zRcg8K1jogUHnQJKyPeY2291ysZDl
xvWFflQrxSczK8E1rZAFWQhrW1OmABKj/h89ICnLGtqg7JTY28IzYDpeaiLDLxri
Z2DadDKfEnkYju915qaaGNhTbOMlpozLADtVk+yfxjv24v6sMCSGz+a0l5gDD8OX
eNMxW2FelOSyCNn1XnHIxtTR6ykw4/ph6v3kI/OwlvdCLhZCMTwK1a0zqO04UDUm
/HFFKyhmaKBSDrqvozCJSZ4z/ETqtq4LYO4lU2k8Yj0Sap42uD2gQlctK4S4jfnu
29Nl4qixQaVDeKuoGhXkace4aWqQFp1tTfZi2UNFym6uug0IMfMtijSLomoKPGJs
3WQKQK1qTzpwKjXVUEOETiSiZdp7f3xo44CAQ+EbzRKrYdIgmi+gP9kD9VBFztOa
C2Gc5PtR9TlHTLzd+FonjC/7u5GQPLwj0SlH1tEq/p6s+LScyGKtZ0bh1ct8qDri
UFcYIlXfJnIBk2acFpiyL94K+eQcRnx5EPfjRaC/IPVTd/E6Uha6rhha7+zBqlm5
hsH444lsAFcrxx16e/+BhnKV8K59sZCQfHtABa71gbZRvUcXpTI34uASdaYA+nT9
IBnSqritpRzERUcEvW15gNV/9VwpwdH6RFME23cQX0AV3y0oce1GCDokB96GeBcF
41dm1ZzPF02vpddT1LW/BtgfLQ9lkwsJzkZVUgQMGX9DmeQXoA8GXeK5dO7sdNvR
9XeyodVgAorWX6UtoI7PsYvVnk4961+OLC53/LRwOVn3bu95SlhgSY2eIMoezku2
KHQKqDc3Kk+OmR45J5ZARTFgQZMpSl568dyej5a1cluw4rzdAw+Sgxp5uKkn8uD9
Zt0ObLkHucl+cYpzq5jqOlMJsxFl5Lm48HR7xsOrEQEb+GyRZL/YI2oLlmq9cxiV
mMbHKzuNzOdeHRFqwEPlAisLIiqkKXzPe9vvlF9Dupd+dLzLjd2MEZ9/+2s8spLA
H1YDTRxHfSKEqXmQb9uWLqWQO9uGyEHZy5Juo9Sn4fIG4ARdH8TBPR1jxe41GBHo
CiAWZq5YSqBY8dS2dgnQm8fuVaWSkVXi3HIJuA741QZIg0dL8rycKAw0Uhq27sdU
TaWqvLyUeQv2SLf62V9QrADp9JpKa5zhDddwHbw2CtVq5lAS9eLnGUF0JErhLE0c
OnuxHLUReHXqxcEUs8hzgMwozxpcpFtefsaAOFzqALUT61o5f3TFt4WBp5rr2uih
dKKZUD+lWgh9IxLU/Fj/6yaH4JqEbqKXWt/NeY2B32Y+jl/hSkBwsUcyVl1itggl
alPDjNNAbMRSJWSCXj3m0Q+F6hySeH0iguo1JAus2Os3Ip8HaPSQDXSIMMOs9d91
Sav21LvPzpr64DPBgd9jifCrU4n3+CPp/a6xiEv+4F8w4oDOZjJloHe6UZDHrYWM
7Ur0ptJC71VdX3OVRGU6hyauM9AZtsyaVsdgPVuwKtsp4SKWjRoG9lUsl0JEE61t
yDXFzjgeQvTRbC9PuPyXx9QTGE33HSRC+G3CSUMnmhFxh3Qru05thrnIJO/l0b7z
s5hFn2wjC2Kt3lymJofObkCaVms/gwTWc+q6Bd6uhErw9xP1ZGMS7C54LalMt3if
92q83Tk2VJTbGfpLTDfxmT8OYiyE8Mr5DscAgRKB6xKq2fYGLgC72xLAO3XiMrbt
F13mAg1zFqoiySc1ZH4zM295YegUfdGyvWy3CusmIx8SUhh7UncGIOxG+NLKJTNR
w4ExAVTYBBrfu2v4bAObIeVSWWCi2Gv2tf9HML98K/rVT2HydPfk+2S52nQY64qc
uOZQ+BMfT+t0M+7JQU6/RTcbsHO7oigkNeLqn5XQgGCVbdXq6uY6FLE+TMcaINKL
YHMRuJRly++B1JpQGoW6aBNG5n2SsPJTo7fAUIaikiX6w0EI9lDdzKAnCwUyi3sV
1D4GQ5+1J8jOuSQKvB3gUDYi56kkPLNYXCbeJ6VyxoWK8YGf1wd/bAbtbyLGNe76
trBUPxhIxRerWwKXljHpVc0iHcSEo2DTouzCI/GbmDmN/3ztHPpbejLyx0X6LqFo
D+HrLUNwM1hfi56pI/M67vUOGwE8O0PKtJO1ZhdlfyouF5cv9URaLUgvVfJ9KPzY
0RbeofvQtCOjfosp932TntT3SH9cMk/F7IdeLQsKjolJn3Jepn0/9FI+qe7bDeWF
F4uK71GRthhXy3x5hxzzJpDYvKiOX9Al8Z8sUjME8kmgdQWD9wFm3Rw++GQeoFUq
dMOdVKG3fv7LSjhdrekWmiXRLn4tR0k2U+BE0pCwH6HNjfuCYzNae/usTqC0d1w9
7/c9SUipH5sUBvDiv8dYrx8Kq2/+2MGjEhZFxaeVyV4HyatwUEeo9BSwG2GJcgQw
Zee1v6m0KMrsz1eLQ6Ud2GSx8nN33yLSESuVuCfWqfM4RH5V+Ry3cPvVSl3vHdzt
rnDqBJXY5xPYixEi/2juKrB+bD6p7ij4SmHBY0n09nDWVTxsg1MUhl/QJu7OGL5c
82oMbB8HrsEfqk9r55eEczToEipmWySqrP1b9uobtNg8gbhfE70tYmAUqEH9NP9Z
W0rahm1DTOhV+DkhXLOJkB+W4pjLKOAU4WjGOusXcpc+FCtDg9DT9PAO0nc+Ky44
ak0B5V8LJ7zK5RjVZFD79ZeesqBh07wK4YiVlxNmST5yXTl04JvSYCcNNUal08tO
Ig0Yypo4bigY1pekzZYGZkmIiLjxfId2B/W31d36D832EHCQp7a7YDRJQJXfVzaX
jSfmion+D0ij0W0MdrrXGhXQafz0ONX3PCdcz/FUu1u6UQoA3y5iGLFT6u1pk0rU
ZnhqFYFE0Fp0v1hMHru8rWUf/9QovOjiyE9txCfC/8rcGob9oYKpSPBbGxloaOtr
V7FJ5Y1vu4kICIxOyFIQBhpTZZolD194OKTTPphiPGcIlqCWVLYj+z8cfoBuFicM
GwdmRl/oJD53MrW3yYpR3IRr4nD17mTOMKK8RUK7+a15p0haTQY6J1UNhx/MlIAp
d9jsX3nhth+tz1DzNJVHMIkV7ryDjpUIv4MdWe2adWegZ/YNKNfY/R9eokGzyz8v
OCooPaLH4ZZ9N4mXB+4vJ4C9uigu6180zgvwosUjpEK073Wl1d8lwd+F7sWTe3BS
in1eQCcG92rSX7wAlEMlFpPp6L/UDknGVWudMzq1LRmMQymgXu+OHhW1K7iNKeQV
d0qk9Nlq7DTPfvyUJdLSH9094l/QReT05gncsSqs37yfMWgM+u+Srst6iUelw8kG
d2+RwwtUsPhGv/uRmm0A5OsV+sXmA8gJ965/nnFavmXSXZwgZPS1NlKW1sGcCIt/
eOt3AqD7fLL2qeL3ZJSM5qxG8fNKkcLF+fnpvnpORwighaEzLtfmOIjeoOxb2Xg8
tz2owRQrpVV8U8TZF3drKAhM7aSQ+e0w7chrbqV50HOotCZbzxRrx40BBApxoFXK
BEl6oSK5ZPqIzD5qq8lwEXFMbWE8KHp5WprV3TvtoeQdWtDoaNALjOAbzdZAnLb1
Bb5CwDGiVw/oA7D2NPQ33z/yqVBMb5J54H1A71R5gNXH0Pkuspo+0yKTQjMBZoe2
9P3gA99+oMC7GnfctLRYO17N+/wGZia7iTRriCu91f6c5Svy3fijt1nlsQTkmr9D
qq8IlRuzxz9+DKD0SsdVi4CivqMjTH3bvqWfUoouzhvq2Z7vq1MZmNni95ZSQiRV
aYPmNLvgll27d752jLbkOzE+ZZ2YIvfKi7A3SkWcrVFTmmC9uCLRWYndmiIBm5Zi
ev3RsrFuTfINlSzcNUlleeKMovyNctmmyPBpYxD2UeRjvwJTSsCyEK0GRdh8DE1+
CTzsDyiQPTFwm/ZTsQrSxECZ6F86ufTnzlPY6hYiC4KXoiu3CIPrToUxm+TYw7SD
CU/+JrqbS0/oDf+yrYJfKMxlZdFv+zrz/Ve1COxuuXF9Nq8ZaJHzFYqmvUCXyq8C
Old2ez3ar4dzieY22WQtwURN66RL8yGiK4S7JsThtJklGDlHBP6jGBw51PrsP6So
XP17LoRnTdN/vLkWG12qJFKpTZMfyrphxndq7AJzLbD47X9a7mYANtRPwOf9dyGP
7Xpt7reXOY9HF1jPubl7k31Ji7mP+Z3oQ+5Fc5NEsJzQ72A1jyoKbPc5bXkfpXJy
XT6AdHfGvRC+HWtUpfEkqCAm95xqQ3gpLVxuG+SPANrxRMRpUZKgKmhRrWcHur07
Z7wp9cCUBUq014kuaYxvZTP15Dcn4W/ZtXSRjyqAlp5NTmM9WBUsgU2Axqp+J45c
MGD2ELBsTQc6Y1DW/S4TnqjGUTlUD2c/hUF6SobLCjA7ywVQHBH82FJnXVzemtjv
iKm6k2/3iTp4wPtqLmyaEZf9C8A7sTL6uyB2EzKBBdSvitUWeU33aqr/96tM9980
tLKKH6ZD+oKhlq790zj7WSlGZ7WtayGMEcPd/3lIreJBfbn6JJ9vRAe5NpigHzYS
24CvFzKjEhquOKbgPrMbGJp2JOrMKVNyKHaE6CRz4pRHy43E48YcpsdxciO1c2Fq
j2rixlzxoOTNBMgEREvnl3x18rRCkO2Te/A9UatuQi/r4shfy1zqa9l93k7UNSB5
Wj7TBgN7yYBHoqoW06m51ITh+pRZnX7xCcWI5uTp+vaTbnkKjld/LF/UobQzMyXI
FrYffeOIRIWZqJPw/KMEGdCmnHme0+w5NXubYrPP2mW3g7mcpi8d3caMI37fpGUQ
hYbJ/bqxE1qDRsgrNiS1s0ZxvWkJBL+b1h5iEZW9xfhl9jU3uhQOASHsYliEH2oI
nbPXPc4RGNxt9+EVQ9ZiKAd/zfo+80Rgg6c7+FmxgCe8acny/wdPsnZjVE+qLolZ
Nb4JhUEN0bIRVY3RY5UXVFTMKqSIuxSWke3dyZbTTS2d323XRKwKrEWezMb2/u5r
HQfbhRgpwtcJvFrps/Bin+0tF7vpBuHRsZ0AUQsKxaorQSomE0jWFLS88cl8ut4A
o4G2c1Q0xzlRCPceDEACfRdEpcDwOWBE6dLBVjbOlCLHps7o04WL6WEhdUKyfCK9
XPwlToDoJ7Oq8++xDuLdvmb2Tjc/mM9fE7tNWm4RAy/m/j9OiL1EzpFxUiiwf5DL
hXoM/bQffBqWxmgMcqcTi20wA1NTSNGS85299SgGDgc6NBLYbxJOoCmfYqay9Gpu
6jz08SjWOQ9C3EvUHmF3z5W3ogTrwThkNmH/3IWjrUuIO0eddi9FslgpSY2yyxAr
ALkMh+ptfkVuJyHKZkPaiZ51zG2GyG13K4E3jGbVstCTEnHMz1ynEju20m5cshmG
dQG+SuoSACTQ6xlCQ8nFbI15uqMMkhVYwDnQInt2r1pvoOo5K5rwYxQwcBc2kOq7
tQbyqocFN0PQlZX9rmxuDdHSYEVB1d6H0d/FHODCkmJZOcT92hTd44zRRGIi763E
mQ5ICxswYcwnGLtDtlUg8f/PlxjYfxuWpDmbudUkc0ppcS4omje16sG+WRHkqXfC
XCHwKRr4r8ZbT1s+qGp3JG+g8Oe1HjrsXmvPikzOyxRNif/T4Y7WmmG3qeBYc7qB
ehDnT4pyPcq+Axf4t4VApM6NFqwJQVKyyJgydvdGL71948b/deDVhtpxUQAeJZri
gJTgRHdDbeYs4MM0nhXLUMeh9+30WA5g8gy1cW+SwpVVnWcbxknlaziArSz4gOlU
0n7+GcTEk7YRBlhkmQrVTPJ/Bob2Z9MODR+YBHwnrJMY22yqThvSbGTMfs16Rdtj
JqOA2jGdri0ekQMS0CtOMRn/5pbaqpHJC2RHS04yzZYhLOyyr501NmGVQoG2RUim
miKCJPe1lriKRHMK29MQQ8DD1jhus1Yak7xqVluRh2YZqcovWyYLsrMNvC20UlaO
D1ksJJXKEBVLRd8pgvhHa7Tny6DwU5ME66M7tgcFAAYAhg7h79V5XC4rqiaKIBXt
EEWt7RdxpudKSuYP+RMyyhdycSfcZnqywSiuOsaLjcncYZ6mJ4lbJ7TWvSwrNl/X
myAfELa5sUwHhla0gQM+H8F6FVByRKC9H9TFTVMeTlfNKRo2ykDmH8373ar37o3O
ePoqWgTcrU1kvKTGrD49WBlchMZBGeN+Ve0E6nVeEGZUMD3g9EPueQkxJhOMia7r
v+zgTozaBeaXqzWIWFFYe9jKa3BDwdpbEJveiTnNybfLjkPdiSVgpac+eJlAvaBN
2G7M2OqwPQp+EYBC4yM6ww7O5lsMvjuumt+tdo0nPfz1fuLEWPMhGrD5TPWT2uY5
3L4QtsZPpjPIChj/y4aP//dBlT02VGew2EacO53FtgLIKU9HGbOqJXH6s+gSbGoB
iewi+Tqn0r2CRVmmWVy6M+4EFMY4JQPl8sp3XX43kN8XtCoHdGv7IDmKyUm60ZjE
fK/P5e5m7gGDRxx8FPZ4XoANyu1vctlVZN+ZNrHqmuN/KpQCadnqsFogXIi+CpPj
E1DgXwPxJYl+KibIoSGAiphXLgpBN10JSHxULVBg3cmfJ9ZECz3kj/VjFsFREC2w
1zPCKwTanpszId/wYf95s5ch+TTX8AQDyx82sbbyedo39diBtFbr7aCDrsaRtzNe
xxFLZN4tMAw1RqUHPTVLIGtFYB1znx8m0BJNQwF/pwZifhFFjs+q9vlfqAMn+/IY
2TYGNft2XH7LefMyF76AvBcQ3qp0Cfd3alz+6KUgq/1lKe4RgfABmju5Q4UaIfR3
/wSoKpg5NPM57BDRJXr2DcPATcyMcVcsonQtaIVix4DqeHKWTUG3Sv/JajzB48wj
/SH9LaS4wdXP1ENAjc3XpDXUExTc36lsZSbAUb0/srMJjwo83zFJVAmr4HNvYj9s
Rk1ra8mSdumiVbv1ehtxg66fEqCUoXUQZI/QTJtZlNgCBwRrP143i21w7IE/Xvi3
C7u+m2TcKlbzRJyODebREGSWC7ugdUhnsxvacExK7H4+YkEMQKvx5V2OMg25Sd3W
j35OwSnPtmVlGFjhxNzrGBeybW7+x3dxScv9vHqxasBnxsqbkfUUtgiPk8Rme5SJ
u+xn6MeeLoj0CvxCbghKa5kGVFlF/tc4ZaK5PobAwo+RkBL9PtQ+gB/taQxXQzQs
686jdf/PopKUmimZN1KUrt4n7RZd2iatUHztFX7dMbt3c01IZjDQQsZXHLDcPph5
dmxho+k78JFRJM7sBu9SrCXiBpyCsW9WmP3S/A9x754MVpiA8AIRKbFjhZYjq/3F
YWzystP2qg/eZ6y7/UGDUSRETmzp4fTOsTKUr+aJNGMTImCFc3YKJAvfjaoJ2CnY
76BupNgnTZ7CfTRaPAQIJNXiFZe0fCecnZ9/+s7VNYzK31TxDhZWfxmBhauNZND2
pKYY8y5kAg/bUkZLdAKz7lQp9pmwUOToB6OA8l+cdtnnPx3lvsDUsKWKUHjg3NuG
XkeLqt8Vb2uU5ivK2JtpTqmQSIivH8nUpAENBqDhpOmCump/dxNkWZuaxqW3mlp+
5UTR7BB7IAoSEyuYnHNL3ckm56Th6QHNF++IniEVujVS58ZzI0Rgj6IlpldfoTOy
k2Q8yomrflY+UNL7mrXsvdCyFmXSrEPu4oRVEs6o8VB+NdYZ8w5le6AEwtdIO44/
M9zcvEccaPzZpuCB+eul/WpiD3MW4mAGFd7mF+WHYz/jl+K/jmiRt1uOA0LNdnRv
eTTaj1I42JecS08pultqPBj8rTJNVwQfdyYV9O1IOj7TMy0m1uK+8Wy1rl4uBfjr
DY0+OUOG6yvvSixHkwt1O7Jp1aRvGO4fo3k6J1p45RuRsHPyNujxSJeSsH9cE823
wqws/DAQdX2LLWUF3+ssSo0uZ8rU7acfwv4mxyJYnbq/QvknKqZcaIZc0KdSdEfZ
GmWfzhm1cVWjhjetkFfGS1nTzXLTg7nnEOHTL/cw4/T/ciNRri5mumy4/rNz/aCD
Xs1VsiC7l45SyH+VW+gYnCCNJINaK5DEAkKjw9dd+i+q+kqluHvINVqYCOHvEK4H
BrZ+KlUKplmEo+KIG0fpZ9DBzLuUJJs5CxcB+KKnuJUlqcYXTtjJPi/lFr+PtSpN
g8sep5suJ0FJuDOOVgXg+k4AvNk6a7pde7i0PrA2BvCQ8svyzw2ClQKj7OIrIQoU
Kx0hVbH/w/Wvd01nMuTTkUulndGq1RSeowbN+P5Utt2awp6Ed4+et0pd8w1M2vvy
UI1wu+6rn+tO36/00sa/FYAil2jeEVYh62BPHE+FIk2/YFx9mIEaldu04cUxf222
8LmQmYdRKnCGzO56u5LIoxElQF7jdOZnW37e0j+35mJ2v8THKCnxTMmSZJ/kTKM0
82TUEJQKb4OTuOnKLIUWmJPzUqn+2DgibpFFJnPvgi6ak27/jBg0869M0Qe1C2xE
k6U/8a3jotsi11DNG6ecMaWI6wEpM/aE2Ylxl+lMhG+LWTseXLYvJHoVyT11snrn
C8OcbuuxBI0wH70EgMVRcWSaEEJWnLOEEKLXFZ8JDWNZT9/uGwo3dg0fofdEMPSS
qEEHhbrtdAuymnhtHjILdjw5M8UfCBoMXr/wrWmgt76R029jk3gVYVC6rMq9jtLO
RKnPTxcPZdnxwKsDg9HbYE0OkORXNfnzy5DWnMgzwRP/tK1ZXf3UtmlFPQU41gFO
Yh+EYecJJbjEqwFsnemnQyUdIWHshKOYqg2nejUBjD99ic6pdkcQIjd7uOkSRBnm
8l9zrLk6s1TEcW0pm44SzTW3lFOvL4PSzqv4IT29p5cr0YA9szu4lM7dhEIH40La
dyY2ShGe57qWOgH3LIZ/zvT3CJpYK1eHSmRPosg4JuwN0hUH7OBz4L+kso5qLozY
pKpuHDY1gxV6L2+OwdGch0qfvoyxUBxDVHZN4ZlOlOb63fCIuevmOkPx194ZYH7h
31QFtP3KgMkaZXXfRDqfCXqQTB+KFjsk1ZfAjF26KtLEGQ6v1PF2FxrVll3C6Rap
npTEA9QLyN8ITGvjRKMhBuYn6f3R0Zh0LtK+Ar7t3SMyhF2143IVixX5jZqdJnjR
hJDLZr2ky1coXEv8zszN3sBgVs5Md5KYTCyyN8LwcK664BVqhVaj1ZluwRzLjIRW
kbutrwrpmDPmGnOp1h7a0+h0V3TezFKqD9KfuOIp+OtQjVWQpfFywcu9bmLrnAEX
uUftJaWglGBqq3fMFyCoLA9JeosFGyB4hHd6P//A/Ir/ppuSYZrNNIIlPX0KCPJI
QkIdv5WTG2iqWWJDlZgIi/SCAVqfc6wsaDxqBHwAnw4UswPLpHpbBW+heRoctXTd
yti/XbB2Tfon8uadgJxSecQki6MjuKnvdo9xb1Takxi5Vm7pqJg3//lK3AJdEfuI
2FDoWaZqNTPUVuJy2vOYHU7EudLnm6vUVOx+8HrKnWFHnsYIBywOA/ay9/9Lr65l
we6xAdUIMjRz0t/Q3qWDTcx6PmXEMMMKKdnNQbhVIUnEdreytxiZTtHcUo3D4y1Z
DEaQeKa5TwvYXTbZ1gOzY4cTE6sYhLT2cO7ChCNuayhgUNZZtju4NkAWdd41iRCC
6gyxGX1XpXciBPnmsAYSfh1vyT80GfqlH4sP0fseFJcePXpteFDjXu24IkSRcJGW
u/wzqOnD/3RXkhdDFS50dwUF6o39YyH0yxP3iIX1fgFbqtt52FN+VqH41x0H7/8w
F6Vq5RuQ8UITyXjdkr7wosZXl3LHXYUmQlda50nK2aSzTuD1vfBLWH7sMjXvl/fb
3Uejq0Cz9oCPAZDEsSFlX5HM68VAjcva1iDgE90xmsDUNxL5/99f5qal4N8/M9cX
LAXzqKIG5kif8GouYOvUSIU1XejhMTnsGxZdxCzaqMTpdvYC8uzbQx+FIIH9xAiP
yx6lbJiKP2HTTvTu17z/2Up5VHdB3MXR+hnfDGxWlac1OrGC3KtP82JPBoyQCC2z
NIpfTIhemTHwOTJf6aWw7FaTbIXyYj8GnvBKeyVryXem7aTjbQqJWOGmOro7GTd+
y6kMqjriwHk57C2DTOxhz1MXQBMaSmwMfrVi7oBFdIGE2MfQEEaR2IXnae4nyV67
bvzc8HC+30VPSWNJo4DbeE4UXGZ+BYp8199iFWrY9b7r15UnaAxhGvld5nkc5WZJ
N1BSQtqQLDSA2EP9JG2zlDdQqQZjwGvelam8jeyhwBfhX3sSA0eENnoFkP6U3Q5U
JwWPH/9fD6SE21dBcl9RsbLD4Msj8U6fHIRXH6gi4f16RKVvhD5oS8TOq2I31ofe
+x4aO0D06k/ESc51p0W6bBvhUssCO9LYk6t6MrV1eaSIBGNs9wWUop0UHVWI+uyQ
YWsN/ejDThH+76v66/1onmifV+ekoNv/JzunkmWVfkKbYl6homq8wSOdeoM+kn34
0xhY2i3L4ke1q4xP9q6dsw2W5yb4WvH43JZbcp51BaGKWu0NUdkojZh0zF/Cx3yx
hgi2TsucOXcj3oFbOtVaEiMYSOKLcsxDhHSFW4mKgXUaNuUh1K4jOFxVU7sG5zJJ
GJJqguUWMhcl6p/cJzGMXaS5V2LKhpM4ifrTqVYodhi5CZKQaTtWFNVRB259OTGo
rSrzN7Iqp4A6ezuis6s+NIdzsOW/2bAOUnEoEUdUxEku0k610A/bRpb3E8qstbuG
OpuftJy32fXpcuzwVFG5Qy/Ya3rybHij8GUn/YYypfHkVbp3YNs1NWVGHPin9iKc
b5A4OdDoOB/lIPscwEIW6/x+6UGbVoUB7FyxdGs74VeoJyR6YrUP2pB6Jh6R6KSO
BPx9lfqfAvb8PEVwsecaZ0gIVPsRBv5aCTVA1/pGU9MQQULkiP3uEHgIRFsyrQG+
JVGNxF3N1LcI+n0BQ9JWNts4/TRU+Qc/7TPGYH7cNjyp9a/UXnTwAZ54wNd0kDve
tRnkIDYsQv6GnxpZHC1/7rRMeW8E4OtJVsKgdk0nrkEJ/MhaDhJ9cCUnPRvPmL3b
AAcD4xyce6IYWMY2U32bYNIM/pLf4KPOEuF1gTxpCG1EhCg02RoaZNwBYO9FBORj
4u7KXEkfnVcm8LcIiEJKxH/ofcQV4EuHVEJo7zoK4naCub3ohRz1wQ2+rvwgEHO9
hDYbNakC0AuKtJ4QoiT29wv2aZQhiTYlxkcDCPWbFt7yDA9UYgJysrJyjSTVyksa
cTZr16kbxvjk+naqx7HllRTJC0CuZv55YHK4HeUlGa30rRnb+EBdyhWAYDCujCsx
10L0nqtNgLIjsyo0c6Rsi6V9XM8pIBUNBtVNTMMwNLgnsvUpldQDhJYHKaZ3YAKa
dglcY7pygZcq9jnphvZnupSbunVW+05lXGq/aB6Rg9cnswuSw1g9CwlNCmVmLccK
mD4/AnXslHA0KbAA9hlCLFAVsnkZ9LVIA8qmC+lsZmlD+8dCuufnQgOsa/hxkGpW
LUzYOSbyofOTZEtawGvF55LGiXL04k8evlB7pTPKJ00svEDweg8Tj8fIkulf0n3H
wp1TtkywkmdRpdXzNTZh3eBrVwhDeO9U+UZeeWefw8IMl1pYCh9MAW68YJMJRXhD
zRRV/YNZxpwegWg8yPPs5vQUBfaJfpIJm4xAydqkkixbXOCCvhEfZ0MkZJP5sKtf
Sh+aSSL/SxUSExvg2I8tW4GXN+d3KzofGoOCI+uJUJgrlkoK/e5U+0qA0wH1fwwu
gZLb8MDCCEaQ21EciWheZls/X2XAnH6kUdvS5vjoJwIqLnewrhodIVDPtyy7Nz1m
IqYC2TPV4PJ5QMAaby/QZEPd6dPaiBAFd6730sz32d3kjXHqE2mR+nu8E5fZ5A1L
b9+d1KouxqtpmE18fzgaadUFWx10pRep+zQMYYI8Z3h1ZT8vzJTrFtjgupS2ElEi
evqXjmKMHQtIDXRtCt8WJgxt/ZwTnQAzMMr5URuTDgrOyObcEfIq03AW8JbrGUdq
d4ETfLPCpRVx/n3H+lmnXuCspzdydFZHgw7v+NjyXyogtckBl9dYECut9K0JmUNT
kNoHDlUAjKiT8iawwymUzxQDyqIWwSmsJ8WeoNEokbUaDOdtH1GOkM5XzYQ/ZlZ1
/ALHBvBpj6IoOOld0OshhpdnPyTCN46itbUn/wLgNJ7TKRsenxIvs/BvsfTW/sKS
KRWntzk9LTohMECQuNg4fk+UonpJ4Ub7ZHxrZlekL0h9AaMEQop4/DlfWn9oA7kQ
DI5OUejHyutmhZlMzIXX6FZRoOWJ690qK7ZISknQe0Ab+sfyiLxr2MEjTjOMw3Mi
+fG3EYUKaU0V4Xk8Mf6tistoCHzHy6pnnHC+dLBc5rjnOnKIz4ExQ6dHYSz9ilfd
XX3xqPNB4WQOmV98/1iCh6Qw2mRoJn//me26Etvl+EPfjaj+MoYtAB05bWyrsq9d
MFy5XFtDtkL6B+37xXFAJJqEgy5gJatRtvXikQxAZJzOPqnpVu4/nGTOD9bBhU2K
+URajLdinZEdy4p/xFPewE5as8i82Sugp3GVKzy2izCLYf8DKa8uxp68JFOB+BU7
NQtoXyt8L314ajDictd5PwnVCdDjch9K1jsfLeUWjlHiuENfGgzQh79Bz8+sT3hP
LB24JbhTqf79x5WC0ZdTgTySETNKy6WtOcq+dfTRI3Urjw39ZsIggh2CyYhyZ45P
g+o2gP/+PTbsZj+5CARQA4v5NI6f71sj15SHchrB1Q7Om3VwEbJ2HKCOU5XyGvXH
2tJOAJgoHKPPojTnfDT02Glf9GRqp/u3xtWUefsqQUk0SON8huqc7hXsUzKzoyWZ
F8UM5uVxRAXUif5VBYTU4Psx6K1IRQqcSDzuwccltXjcqMVqwun2sf4PnAFxfsX4
3qeG2hykRvDu96PzS4oPFU/P75CQwvMdrvrJnZHu8BJfVJw9kb8EUvheveutY/qe
BNCNI8VWeVHezshpFCLQaPOs2nmPa0mfFLgV7+aAUqIF11Tc+L/xdZnnvC1edpg3
P+95+VP16XDNpZmk/JnKYHmsMl+mGvnKaxRpQE+KkrerS9fncb0DJu5o1I1l2I/7
dyWnvTLL7mA7LjXERPc4UGmcbOL3N6cuN6uuKpkEIZLH5UMdJAE3CxJotCctR2zT
BDJ2v6OqBSa0uNE1/sntkRhQmMBRBswi0W1Mwl9TZPtwzZvQBsSORJYwu2fE0UnL
e/hDH0emQ2Kt1wijMLyHZOWUozoQHec0Q68xNnqy0MDaIjLj/LH0uDOBPlqbsBOa
Wg7qio/ANzbgVUqBYbJ9x2gDhMRNHizALYXBU2dSLV+em2P4Lg7cgNkrB2Z4lW5o
xpv+CkCmjVgNUQWAPhyX3qP+d5I8rNPQz9dcz5pYleXEKSHGYWPLOkUykOhw+hLk
qp0BqAQgIBPbTc5r2MVAQNL6Oj68ukYdd7H8moCeAUNpjW5LHLNdNdfwNXDJHO/h
Ha5CNUNCrEo4NwMsmXYIkNULRiUKj11wgswwsLszV2SGHpPMjugtk3I9WrzWXM75
pZne9gZtpkIkhvfYka5zjjl85O4vFA2dadem+zdSlcMNH/fvwYUrKtAGDHjZr1dc
59czz7Bxx0SnU1uiY8ClgtpX9GwKjM/e263QXIpOfeL1x9jQkUDejGPxNTHHbdU+
U4czsht5UF9Qsmiqa8mfpSZZo7SJeuJatwr7QVaf84Q/I0TtYSm6/XsaZh3l9O/6
NbjKxJugZU89q/FfspqnUmnnNTymFq2DZtupcPHc9QCd4i1SbGi3zlfesuGrHO/H
DLGKbMhjhofa8sG/g5rGOJ2YBk5dZf0b6WF4kHa9F2+/AFq8J7SwYXnW5JKG9Ngi
gS+aHsqihT2ZfWMyFYQkrYnDJvA/WU9YAdfP4QQ2jR9KiYGj7HuyMDWn+0ttvWaY
d2LYZEwAfa6bUBPSNALPi8goo2lJpnMfst7MzMXOtbCGMcgr8IdLuEzd7fTx+MQC
Vp33HRkN35XPUXCy2Xx25pGAs1JLO/gjo5sd7E/9GzEicSlaCu5fRRGwVd7rcLQB
k1w9K/PNyHPQBD2bBkqHJxsXTl6V5nLd/WHrttYFESZZ1ZgmbrmxUws55fm3dw2U
GZNBAtQLRCvnhSqTH6uGbPQ9qZks33i6LPGXNzICPIt6D8h5CJ6oCLwyBgndK4Va
5i6sWcG/HgJ3SnGjMu9L02ASr8Y9GWdWJt9JOYSVbl/KtxDzq4hlySdjOcqfBGGr
yB+eFYz9a79A/v54o0GGD65tozCJVXAk4FXP4R0XKSbFPk8emU3w23kyjTdbMdTu
v/R0qK7yAktZSrMDwJc4OK6cjHwpQtT1QhzLZcRzvWa0pfyoQ7Vs4YQT/3vzOFMy
Kgqldo1aJ3tEnDAVnVjWIqhE+uV4+soAndnO4HHFiUHQGl7IUespKh0mvhnFM583
KFJTiLSCE4vkRX1wF7CAvMkrtKNZLPc2bg4xOlcq6lKzmZa84y+1jwUZKRcW1j4n
i4F/57h6v7zqQ/Bl28gqf5lRCbHjfjb4lwgEbXIl0ISYxEdg7DrvHlX7mvfrR8ue
SRTUOpPy2JyhfHwH+iattcQP0urS1x+Xm2D1SPhQp7oQhXIXj9EaYA/TQQjQe0Ms
x+0u86LWZ+D+gNhyAF6YUKOH5vLF2tZOGMvT6c0lfwraxnGDLAfIyt4NRNoXdDfK
pzf0MnsEdrmboT5LFmZPk6dsznjtm+EJr3Jffw8fZl9s0KylF58Z9cgFtowduw8Y
HfryWNfn38lKjne6N01UYdXZS316LS3tSvTxMoREjPW/RUtuYOiMNNKbMbwOuDNp
kRD6wvn326rUkRUOBIqdX/QQ5oo0PDYKNDeXUwIRgPEHV/aKwf5w5xIT5JNRk+Pw
EQIR4nKEt9yV1JsBfTiuoEwISoskuDLN1L98iEgMtePIWMTyAQ6jbFfLP/lACW/m
42tCBlrtvvKTtlBf5LbhfxJc4cpWD/Cnvxeg1mTVzl5ID6gPmROBZ95I3g/UjTlg
3X7NutfOFQ4cLM3wky3rDXlsOYXShzYNi/8qfiu5FxYA/THhCmUrDvIdLn+lWMZa
p+hicFkHFZsqgB3gtj/NRQcVP6XjooQjNnHBDNSpx1X54CayFlNOU6dsoPsr3EIk
8a71BNsZFQaokB+g7121TBYqvFIHAEQtGJmNRejoqGG0kC/FWRYx+2VXb7rtS2p3
NfMhJvgKSGo5+lFmAsa0KX77sQ7l4vPE+9azKoGrfJUPvXNPJp8DJYxl+4WNwszP
rxQnjYTFI7YVVV0oAIEFXcMdGICdH4Y/vMBQL9r4JIl6LQ4FHd1bekou3bpaNbFl
FDFSvmIZJ4J0cy6moSoaXQlDKrh2OvDQ+TBhW2JY8YwSD0SfTqtAnlA/qJSlAL6T
lm6SD8sEigs982/VC3W3ZWI4qJKtrAo7Fzkar4kayxaF+IEDHAcW4NGpoMllKOz2
GYcu/dhaeI9cIZ6wp6Gp3F0avXO8eKt2PyI5geOG2Unvx6jmF5mENmJY5ED4KnYt
rtStSW86yPThlhG5w43VhMEGghn+d4AW6VeLlXOs0iz6gaplfZ4uLhed4vG47ttE
XeP55TGni3ZVgjP298QIU6PI+AxRVoFyKF2mrGoNNDDtsIHuIW4277TFrAMreyll
Vc0lCWBEvQzcRGSGvqoxdxP+ufhwfb8MVyn2btMARv+NeCmlJiGvzNRfox0zi134
YC8iCa60eHCxTsLXxaAUX+gZhXtU/MHN915vvcKoMOz35I7KnQhSDd1T/LKyqHkf
uMjVEk3l5dAxnCrggqv1bxRoM+ILvKUCx7LETwiyKZtlkrH82AnUc5mjuuziOMLa
j/25wRdRt+6podBZVN7rsTbG2kD9aG7w9tqOTWlnOA2QgGLG8mEr5vigaU+dH2om
xB2AgRxmQ7m6pDarYjy/3I3Cppji+tgx99bf1nlFr9HWZ2rTrO8SWijLvAf5cQna
aPxIQLoQLlkIsXqa/M4buAFUtwKtjvJrN54FJHGzF1B+VKGjpzjEoAg+9FQk8BIx
+x1v5vteuBK2Po0BqYgXny6H5eufJ8nHm49MlS0RN/AXMFT9QkD50R8JBpvPO/1r
bWEyZ1bBCsgQIuuor+XzOAPjP5G0sTycvtWj5WCsbU3XdLXoBkVRf7cWtDNOv+Vt
XuedclqVLOOrcZMsI6Td58uoqKZGDWCG2XErSE+Im5c0ohu88iveR8gkSGdyILfT
yK18YvpOF7wL2h7GNttkA9LRkmwnnaOhNI2bPwJwKduaZVeHK10XvWAF21aA8Wsy
irxOJXD4tf33NPV4qL+JqfZ9zIiv/Zzxx/h+HOTN9WEASuFBUAJRGJJ4halHooxb
2X17X8r97aAq9IrW/nwULII+VZaSLRBOvbBEF/Cd7OcIxp8VTBFq14z3lSCvh2Gb
IXACcBl2Kb8HPZ7fVkQ6qB0JFYDrjYNESmgweHBACSBAfcGSRrOp6EdOSkxONqeb
+tUw1TOHZWZkayKWwU6Evkl476C2WNFG00fdrYxpDe4e9RTtK1OTmYU08+q8XB18
OBJ95I7EwU2toNm6g1bopFFtnQLpdjedjHMGp6pxd3fQkEyl3Q/+2NJg1tdkZSBu
WUmzROHre9rdi0LczeLoQ0b5pjYwrvZVdfbsuQnSDsn2+ATe2hPXu2LZbUpTrzCu
1Hi7l1KMwjTSyzwUQA73L6UmXPerTzKoLItnlsgbuargVqCncyUw59DGC7EYlY5r
IyBZROa1N5CSsS9d7Vxc/wVwI0mfDDdI9ey05FzEa2J++0pRg6LL1OvzPHa3ApKo
CxL0rT454RCXpQdJiGrsLaTj5ELT5hNWNyFo09om9YXq62tOyTKmE9TZK2rUvMAC
XM/tJA7xY6XQJx+W55pLvSjdVmBaUCBs24mgO7dCQsm6taB+XHCZ7a/AO+njJyUL
GylZEHC7vrSVkc1i14QRP8Rk53W9TCkTkNT4Yg5C2WK0TameLnaerFGNgKaxUx33
cpqGNodRv/k3fPpv0sdbF4VLfNUIYivuLXD7y7nj8cggEG8+8g4d2Yfzwu8dh+v/
XwjLR2X3UKPeYmNNj18Vg/DYzg3x0+xtnsAbUgwBODSKA1V+XzUyJdhEbNw3cZEw
4YK4a6M27UM3SZAuO073rAALXXDCbcPAWGAh03i9GLNP0MgQx9nWwJf6pwujKn/5
YS9O3sAmuvcC0wvf/q3hZRoOvffj/BeujA9FHsDme/i0U09wjNX9K6A62dmFqe9h
WH9/j1MyM8y8qsz6Vw47v408b26kbo4Mnj3S3ZVL+XviCNrle+kQJzihlnG+7Wdi
qpNj62Ys6wuYf8p3OPBjeKaVCZ4isWh0abAqtiwF61fPW595Gu3M3GcSpqrtSZSE
uhbzEQP0ERzlM6z96jXU/MmdAvcRn+FG3sv4ahReaDhwToP/O3fTMC8HpCG+QCEk
OBFdd0QeHMvmX4Gc65cJ0GRmv5S7pYoBiiO6Zz2yJMgytp7IKRcQt1E1xvgCNu4t
r3LVtIQeieiC5Lv71qcdo33dmx0KiVGCe0kJXxIzsQkKzJ87a7haxI14cBHhxHWA
/V2M44Mm1p4gtOSlFH7FsWKmA1RHsR2A3byDatBc1jhclmh9OAHamnR9MKPCeqDA
IjcI/Wg8mmcGwrKAZaaVAgeKlHiPbNmOAvQV8vhv7Q4vgmqb+CaOUKRPB/xS++rR
DOIInJTsRQSTzZuOgtz+72EcCiT7+adyONzq7kQ3Vzgm3nHhqXxMt6DeuBJwC4HB
2Worl9/jsE3edbSS2EosWupZoEXDDiLCkvK1kvYNF2tuLqZn+N1asOHAR86QnVst
W99/O+IKLSgzf63c56hwgeYZrCyFrsb4pEyctkyPDXZ1/2tthnsEB27fVL5o1J4T
1+Oh1euWxkwA0uT8dCl8/KoxMiDi/M9V2kaPwUuhDemjEZTwy2xmO5f7rVYIvTfZ
f/0FQkK7/zmv34B7++PJxZLVpC0O19AJfl68jilhLefUUZZe8e+e+GXqtEr/Saxf
8u4lKQS4IWYBddKEN6U9Z9ic/rFdYdqJWnCw3xALcWUoXkcQQ0hZQiJN2C00SAex
uCHC6vQRfRf+GLv9hS/LYtYfF6LwQyjUmWMwm69IZ09cWt67Il+rvR5zUNb2vMVj
XkHQ7/dniCOGy2YiFrln3L6v3vnt8E8hlAcPE1+NZxaYoYT3irEtniHjaAHnfJjs
eOzNe9vTPLqDsVUzIdE2slu6BVqVsNwYDvayP7MQt5IB6ksiD0Hu73dRKoOtP4Qo
Ogjy12dpmbaOAZp4KdpPpEUKktbB4zo0Uu292/X+7lOgzEXAof252bzNQ1Zgzwty
z+NzsTnFfJM6JUIT+h50nollfZZbmsjRbJdddae0Dw1WtqJV6+K+zVcytvs1W1ct
9cbQ+70OuzTSdOcTQWql/DPhnkeR0EMtn+XLBB9PD5pLTcWUOdqrbQ3E/AfDVwjS
6zY3Tmw3FTm1eODsZMSYyunteNeA0a1c03cfDPxnCvQ6aTQCHRy5JQxtkBGMH93f
TCK3ZTYpdcBge4NjE6ZTgfHD21kHB8xP0XdV7HA0VQr2Scplzpc7454tFJZXGXE5
zPobWrHqnuTdhgM7N57Qq6m32u2ODPYOJG3DdR6F0dSIGgcAEDpUdyRMHyy1+cf7
gc6y6Pc8TDghoixhJRmV+dYeuPppQtH/iGw6zVCOewivWEPCkn6Pi7PY9eTZ35CF
jA5zzHKyvPgoh/Hdq+M1NXd1jaI+Dblb9B1DXHrRpxxEMaUNdq9Kwi3j+/fFNHpi
8sO3cgFV/6X4cbOz7hzDvE+8v83AN5CcVtthm05nOIheg2e53LKt3egMRFIWz+Ku
dN/jpqYq/ZKf6W+27707/+JN22N6GyRY52Re+sqMmkUe585kkNue9M92F/o3c9Wr
WF95pPh6ApFpQ2pq9amAmvIw0lH/9ZZB7dcxRidCUaU6WX0lFoXIdl41oRgJuNtj
ipt+3vqyxGBujbbCpQlJBNpycW5B8/nXNLsNiEKA9dpyu3Imio1Ku8LlHKmqFcHt
ARNSeaUEblpXeY+YKS/U5AZ4Jvt5POY7W7Ko6b2NoR8IbrGE7c7SFPnG4LDaKsGN
gdbgolGoMnQ4/Q4MQHUMEog+QhaGBz/wxFUX0DT7vq2dXiwoFxY23EZuT6+FwT7K
1/NLtKYmZzKBj7+vHMlKA6JAYyUcTnupxz/viusyEU6sM3+ayhTAOvhnflawcuC0
9j+FDG0NjYQtCq6VHysmu0WgGG8w0GCN7dpjIUIgOfLDINBl22TFZ2QSbi6YHPXu
cc6boQDRCxTv86kfwjy5pdKEkNpaJ5Pb4GmPf9t1NZdkMr3JgsulH8owc/5aPhDD
br/sCrxOL6KpcwZs/eK9eUFfdkNySKy73WSyRvEz2EQ2Z5PEB2pwFACiM8FkooWd
3uULwiv0tVAXYKO9OrvTbzp5uuwGQiMxLoEYj2vxy9SU7hpFnCdTYf8Or6R1gDAl
Xi7ZkChIuPLjagtJwv20sGvDo0nZ9/vlYBToPibrZcpqoQbGs/Kfb2rE3OyJpBH6
TvwPw66/J4HFQhkDgzKb5mYON2GRvd8f25uMN/ZxIxXo83l9+aHuIW32Fn7qzrTV
IH0Fhpjku1504lKyPEPSFkyTyq5wn8HS9hI8a5iTN3C/Fi1xYzyAAyMs2NKZDWSF
ncnfnl9WCEmE1z6J33Bb/NEBaBkSBlaM6cKK7G8Gq/1uM5h83O+QXWAyo6rqsts8
44kVDwnIMH5Fe/q5tXN1mJdcjFWpFP13nng6imbgMEQkc4uY77PbLOBnHKeYa6Sr
QcKBrpHY1lDLi0VCBkoxe8x/bLjnPGEUrhFy+SGYzw36kxBbFisCjr0c3m+zwJC4
IrStg8SWdLOU2A59oBl/UvSG1D308jb+ThMtFpAvQOqgFwyO8tfKN62jeO0pa+rQ
lQi5EkxIE/RhAKdOwdW+/YJDY64n3OpjbtZw12GQlM6Q9x1Euqg3O97lNH9JTqnT
HQgrIbNNe2QwmgmltGXyPw1Vx41x0SndYcR17DHjykYNh+Czo9pvYINNRBVdDp3U
WpB/rIRnmRQjeCS6kzT/3kuA+PKhIU+T/p2EVWfGF99ganWkCoPiTS3OaxRDcPUl
gRcXzbhfMobeo3OttjLvCTq//VstKD9vEXym9NlhNGsk+DreedlyZ0rt1Q7KHs7j
B3nvK0jSPQETq9kXoxvoadDAnz2tJJL3X/ijT9GQleWhB3cvx174zWKPGGCWDdUm
4LxFzGERGjB9q77iRrQYf7cAnxR2tXfDxGUffp8D5qNYyht8ekfGBGGOv8LlWLhi
VULsLfFyWA6b22w933UbTtNEhL3aMYAWbEyZcv8Yap8pKb8Rn86N7RdtBp/VAv8z
keGacphuuKu3dTmyjQ+RiU0MiEQ3QIXvbR8o5RVdzOdXUawAJMYyEzfx85H0lLwz
9RqwhIBD1PLYxBtnJdLYjhqPLcNlq63IKpSXI3GRPepF4Q2rqtULe1aKokk5LNDr
Kldq4w43Bmb7V6behBO6llUgtDABvfNdf37Sw1iUnAHcFSzuwLW1HVK2B1vpl3ji
uo7xY5KaUZIPR8BYrszK3X8+WD451pnj4pHhkZ/UlVilPUVSrP9W5gLolE7anK7O
SEpKbWJI00EWdcSa6j+37dIvIzzEO0PJySg7jFn9sp3RYRnZpXgPIAahrSHqc2gC
mp3GxMUVCT+yFubXvIOAR9foSI+UNs4NZnUrE22E4fKiEoLsO++SY9xmbx05npZz
Gl0pvqn/3iafsu3jHxbSZL8E7LS3hPmiiDA32PgR/1rR2l86sihbQHEoTCFcKEs4
mDqi4DiteNFQMoaLSVTEZDawTCnNOWlm2FIc/qLJ+pxNObKy/3BEUiaSGlfj9T0q
VyYi6GstFVmRTsAScpCleeL+VKtXLOm7q0IDblGPVPegG160A3+4HApc5RPt2iJS
GlSmdXWWmtKNO9gFfs0gG8htiXsDYQA41Vm94FO4z7Vmu8CO07IeB+ly8biimSS2
u7suZ2MM1AHcap8Vn3Xd3WPwFpTlYQKTyaWDnFzzq6cQkRPbAzA6sD+wvslo8LY6
95XQudTH1sXRZ4Bw6VHjbc5M4ystNu9H2K6gchrF24ly+CiaB8edP8Xzies4ILib
7GTcXDmIeIfvKSivoEO+K+NhGKDH8C0lWqo/FSd6O8PuAOee27OUdhW1I1DWkyRC
YEFQz49SjSTVS7l+YCNsQvrf6UT9Dgv0eD9PbC/LQLyPb2aKy4DrxXyrRvD4zE8G
pvXObawoiKWOpStE1uSkki6RFr0dTZh3/ZpaTlwBq/oomPhB3qzfJqLogpX/GNWX
b3qkmwHlqZP9ZQO3wPzXwBC3h4j/qEZiaUZFOL+YXjgDIH8wjzn6RWjdNAcvLObH
YBZ9glQ4lQY+1khbwU27iwkpn9CRmq9pxMpTkSxCOvA1t+yfvwiYqpfAuRBeh8ds
slBwDzYgY+s41vOKez2j3hbX9YXqieTLreiCeGOeOedihoqjhVwvmcK0zq1NLsvD
Y6jH34A1b9SwQLFr3id2bb0IC8xhY1z8uXLMa2ZHDOwpXV6s9+h6/ohJkEHRiIS6
DwFttkb0aEpXjvA8uQhm+cfOzt5jzWdzobtDPIvEVwr6yIwI9t5gKOXQzJCtt3P9
Mjpd0kCcJWkG1L1G4+jLrYEoRNDkw+lHRidBkI/WnrziB2jpNh30S73fibELqnbD
oICsrYH7YpRuxoc1OEAD8CCcRu5BLAk7XSY/6XikkSdqjkdLe8Gu+AYkOAY+9MRD
5HcvwqCNLfrIPsm3DCn6p3F2hqX11YqtgoEgPLBO+Ss/R9aA6Kr3EaPiSFbDVBQi
gmQNRgxf7IW+HNnqDRCM0lIhhhiOQ/LUzMU1XL+Us/1KBTQQO50xlf7oJp40vhc1
yuiLneCX8RJEje5baZ3zpjSd8JfySq9DjDHh9/qe8P7icMunb8e3pxVuvazY33z1
7yJ+xmakOoHHG//TxQhooaAr9/KdwCpfaHGRlaY+FEOaVXB3w4y6SOO/NxQ4SthK
Y52TB12ZBYAXNILnIh1WWmUXhEVbCChTDPdmIiX2wk23Jp6vH4Q35xgA3tFGca2j
KdaLN2h6Vh8JoPhypubTlRJiiVzn8eXHOljzXSU3f8qiMfwlGe++C2mvk0DYvV5g
8fZR6wk8HYWqIw1F5cC3/dsajtDf74JXJTAjSCw3K14ZCRINbgzZC239g4RvFBLF
4TM+ZG+0gI0WrLBROkjEfvsNawwl/Dcc8XZtuBrjWNErou1tQcncbkpz5s9ec4up
1HOeDMmpPJ0aIiGYJ7fe8enq4f/j1blN79M67IJcoDpnGIX9eobYHS4fnJDvR60S
gpwGMvhrSjV+apxMQkmVhprutmoWqdUxYKy8XSOn1rhNZS559dJwlH/lxOnRDQRL
oFogWz+6sePR/3t1wlPfL2KvHwF1HHn8XApg5Y9D6XU7bUqFV4GicLzJf/GnvQz/
QoMcUoYuYXRdFgWjS10HyRqjxS76ekKNll/aaEXTWG20XqvwZs3vzFhNxP0DcBhZ
WHebazShDcuVO2rLCt2ONthTa3J3DfmLelK3IAT2F6m3F1H1ULpDQX0omlXDPAjW
JWCn1EkH3KAwb9Pk3tp1UqysuC9M6J5pdHYmb8VytG+UB/qMA91QPr2icuPseEHn
QQqvADChpTUdsZC1xSGe1wfgluLUNu34c0YhhYdEcAvt9g/zTEeUhwLaKmA7Qvqx
A2rz8wVyBq8Lp7EGA0g3h4xqmUcIbZGKNkD6Mdd63ffsDQOSS57cXgzKcJHyi6rd
lCvNB5KIFFO1uU0F3h+7vBXg4op4Vqu9FrZbKjpCjeKnpcyyma5AvrRvKRkQuy0v
sTJw1uFk3gs7yXRutTPHZgd61Q15z8qN//v/og9S2RxqpWN0xx/NwkUOVXRD9tVo
25MlyiLjLvbkLC8pKOHEDXso7GExkJsh7FbA/ksHyZ6KlnJOdk6ft63/0jcdzGNF
YiStpOSTwYX2N1XnzG86rtoBzmkF89DbqzhOnjGu0n4tri8vsP2oSKq/JeyLV4Zb
Z8AWRPJIlJIJXmq+ptE5NN+fCjsESoSUAz1CIZGsqWRdfra8XBdkq0GmOGloSYYl
i4hM1JvazPqdiDa56Obn2lYgbuwxLGa7GgjVsOro3wn92spjavgfPANOgpPWgu+5
Z0B8ZTk0ogj+5xLiQVbg5hjrbBRVSCuJyAOQY8K+GmLyTabuJtpRlOPl4kkbZoTr
db6Z7VY051IvQJc0dmVMEEwXhHR0NeK05uRRP5uRIKEc2Sk6k0Hu606OlpWvfan1
HpwNHcDh0pnYzc9qRAcCxWTucwcsF1a0qjcDhm/uS1lB4VhGE0qgRfAmf/PSGIP7
ynHlI2gWWJ1hjh8yHQurn+q4OHgn6zN3j82lU0vrlE/NIUXXgcHHtuUNFZFWCTjT
NZ5hPnDKQ9VvM3X5v0Us3VqMEnW0wxCkyp3XncGfocCVQpDah1dczVJUB2vX32zv
zin+V1fUYqfRRgj+k4LMLg7GzIUIlES9HK48m//qgIBEHEKUPDQEpT7GAMTJGv2F
yrpPHdVSKl9BbjRhsWAFRt7vZCQxoc9WmPS3uB7AaEkBao2N3NiW2BLZk1wQErtI
5uut/eBGW0WctKjFgwRm82Th+Ttl9YgjI2SYz2Bakm5fWueK5pxL417rPqBijpbA
rxNajIHNgoGQ+bLYhj5qkO9eEfhF+HSFDfax60uSdrmOwqhojtcw9R/ndYr+gNSq
0Y3vEviB/kMEF0mjlOCKXsn1MrDc1RvLZjMJ5UoYZe7AlfHO6+R8i4SRWCjARfUo
fIhjpJxt5hFvMfna8zSWpjx4uQYFHE44vb/geX6rNNM5tRrRxGfMvmscu9mtzF2Z
bKfpw71hINUyxjLGeLmsNppVF4Y8kh1T29rkBheRcJkhSRu5wQo3ghNcQSokAwqp
bTeCJmCC0NBxkQ0I07ZNvkrTq8VicrYmBuuN+cOdbxV4WZU1k46HOUzSfp8Xy41l
IHDva69XsYaew6Re52TMRsKREYzdi5ri+U5eToLQQ7PgiysXQN5Dv1cSyAeVij+j
v6R6aRvtimUPgPjZn1OsB0VAGnZ57AcQZ0/IoVMLWy7sk+2oxAY6a5TPKnzplYz1
OVDYlXW29XWuu3cchDrD/NxhyeF9+ch1NHG0lK5givLiIrMC52b4nibtYB7h+Q2x
ozeCKM9uFDGDs0aYIIF0qA4VJKL0Is+VE3FEzk6HCiGmg1N7gvKOvLp4rs2eNODc
N2HZPyTYk8x9GePkffOmcFasdKAJlbt25/ZuA5NOm6SEVLirC4zUTSIZs6DQK+nt
axd9nF0RvoFUG+a6MThg+dqBiWnJd36ksYYosK1ySiHZbiaJVMfvOXjJygJ3WrnT
vSBd34et9Qinmda1u220Jrddmx6TjIHgtV3P1bNJhMi7wiJsWe+KHAXqb75H5615
E9n3HiswLlNVaCQU6k1DQyfc8a9xm6tb+ocopqsKyJHsxoPpXN6OS9QIy9D0Tm76
IYVrUOeD3SUwM7T68Bz5Bg3Z8p/m7YmTayVarFckisXDz3sG3aSs7Y0S8aS2nj8z
zSJDQvwGgUfh575EOhr79HoF80Q/NqxOBBo8jtCAjsjSIVc1h6+NtP9U+sNZ0kBE
GpI7o49mtI4mM9bgYHf9fZseFmdOUwcVgHUuePXAaEM6JnNWfqwgpyoFo0+VYh3n
N0nV/kPIDjyOlUa5nGI/+w3TddWAoKOIYQTzVrT3qYbjsehPCqkqfbt5OLZp6yv3
vdJ1nSCkkpNHsn5VoMqzv5GNMqkwRUC9eQfEnMUbirl8+pscw7A/csGmcOSBPdIK
V0U0Epgh2xzaYghot5pxklQ8+Kerit50r+gcln3iEqJ4oO/iszV4hQEepHtc1/jn
AiIujJuI33ZEH+JsdTmaaO1KTh3VSsHN6sWKMVEXBLJIKrgBN/hqKYU829XbmceT
Lmd7H+irn3gN3/LV4reewCp/QNQNR3I/2kjRhivbNWVDOF8vMUCxkRj8jWbpo9Vw
5SJspY1eGMhC4qv+B7pMpCgHjkr8pyg1iHNZr1gpVY3kytiCb+z711i3SgI0gdX0
rdlyVCWMg/UF7prEZAfFVT9mM8Wt4dTELIQIj8o9GQZ1D/GmzzTdd1e9/EaBSDSB
dtrmJepamONN8qi61gM/91moq55PZPnAE+ckrg5FHZJz37vgj56ZdRNYsGObuu+c
cvUYKSh65WiVdeVJSRDt+7/D5iKv7UeKMEW6QELJbwZZdbwzwsn6Kxa0s+28KJ5s
8uRCnQfmfxRsjNy1tJfe6yHS6bw3gL5WyPqx0l0jEm35FkY1Y7pNzy2v+n54EzGp
LIhDb0Zuh1BIZrRrgECAhzW6u8BjhjE3t8C2zmHwFx53BAtoHt5JFj+W/l6zdDg2
VDoICnQwZxL1agzRaLP7nyWFyKn4RqtqRZEtPDfGYc2kPTEWDtlOsGqgwUxcvLSv
x5vxLNOqxEk9JlAkHY9eqSmCQiWx69R2eQFTlQPSaJh/vDFNLXkjh99FvQrHEmFD
3j39GbF1LUDxFeySq34p6FlthpQXV6pn8tUzW9ygatme83uxRW8SJCzugD+5SdTW
Dozg2Ajmzdc/J1+Vs09qeDpymnPLvryVY7oOT+oY8tLWYYf5gEf2QPwD00PauxQ5
o4FwMoynjAvQobnNdb+bvsLm2U4Zk22L+jWdm+2vnafFyPB6c9+QDy3Gij6xekjz
p8tvG+2CehdgbCC4k28t5M+2iXGWnNKG43m1DF7HSh7G8pJFwUNrre2qL9DBMLD8
WuwV4eqWCi/1jyophkVa/xHqbHIDc/0HuL6f+JyLJnPex1m5F0opcwvgU7CP4F+m
Yv/mdwyAo8Aw5xImaV5EIfTN6r1PwCU13ss2zMyZIYkaLYoFsGsevl5yQdv5nPcm
EEwAE0i7f+2CPgXGPMHY1Oyx//vw0z3nIB5spD3CpHGV8IFuFZTEEr7VAMnPwxSr
/QzywuAIz0HU4kfikbQYBSGjuHPt02kIxI0JUJYToBTRSSdep9VTbjmllCpnJBYz
md9y9w34D43y8g04oaNm+eKoT+nzyQ+v2VfIskgMMjQ10z3J9x8L1DI4pTXHDY8u
b8FQXe9RVEJmcrpDUK47XC9GCyMs3SxXkZO9ucAExok/hxmpKj8/xt3yflxzwyjU
ddgbPxrmE5Jx1VnmMP7fYkUBJAbhGOqm6MqCig47XqhClF8Bnmxax9HxBoQDUYO+
xbShVwwnnBiAomwU/27YkiTHHFrLRZBBAY7ONUCYyfqOxTveWMaZHw2LjqaIYQQ9
T9E0nTMH8i5i5AYy8A5syVzptGfsvXzkxy3COD+gsqySsiHf8JqTnr019MvBNULd
2kLRfKA//xIN1e3IUfPbUAcfEym4xCMBbHGbG1gyZXk+vxJSWZj0B42bFzOIWg1H
MbApOgAYxrEo6gsRSunCidadWjeK7DVbd0TdoPsHnnoY2WPFKaEmACqOfkxc5Ly8
wlah3MytOjURHPCEs1yQaWJ8OujDgRnbOCqoNpjwsqbCa9T9O3yA9YF6Pnu7xo08
kg1kiivp2YsSF3H9us/3NimHCx1oH/pv1BxmNVQfM7B85/ZzCGk8lol6Kcc7ZdyA
iRPfqXCd7hNy7+XDhJrcAAv7i9DZGVZGT3GxgYeG72coFgONwa/I915cfOz85Q84
mtQ4MuD20a5LroMSwOUW1sRJ4GQoCRbMqav9kp63RqowNjaeNQNoFgQf5iUePTQW
wWMjrBfdToyutK6pTWoda7V71x0DIIAp8iu0LnVkLhsmxF5ohpM7eKrPRb8ODo8E
wC7wM3Wcr9DJ5WS95tUZSqIcRTBq1eJONVW9tBSyoXwlbFFD71SvK1E6uEI65+t1
Up95gxWZkFUM4YnmnEWB9pM1oLKwSPYjC/5gtkNnZx5SxCe9wsh+1Ep81eCtVqTW
f6RJjSmKxXCQeKSV5qp8J5Zy1kKuFMpBcvVApX/1cB99VfmEYhWCvr7UFp963KzG
JPgGKU8+megaBd0+YFqUMcu4IWiquxgkKxHwnrJHIb9Jg+NUs5Pe397M8E+glgZG
C/BIsgVYaXuB3YtDTTDBUMRT29o0JkRqeC0GgF92ahGaC2xlvY6QYwPcBrm0/R1Y
ajoOEHz0u92hLxJdixLpjELOOJkrr9RZEOgH7pLydMScspK4X0Mk4T+Q0VW4JCDy
abbMkzOZcXqgy1nxU9DGu2qaCalzr4eRXm2RahioEZiNyEJUKTviM3qk0AO3L/zw
dS2VZwHhtCMwb0oQ2oSJwhRAWpKiYaWN+ZwYBIPEuyl/chEAk9lop0kXSxfXAyc3
mntd4h4XnPOxexdc9WpGncG+mSqE5ZCReeabPhgptwy3HyIqF/K+cuV8nscBF4pR
jqbnLLcZ8e6GNHBOrN+yxRtE4vA8+wdYbDwNrb0pNlD4AEDTS4tCwAn9cAIfv3jg
GJMZUE2CEpchJpzYl/qKWO4epvwf/aU+5CYsRqVwMvaAj5AtgxD8SVV6ZfF61UqQ
gzsvWz4lal4UCIuNThjNFeeZA5Z/BwElzQdXJPq7Gk0dC9le7JOhL9seZLnwjp6g
oUFvTOCaDnlkckkhgwyQ9mHiZzR1uU/SsurTahT9yz4waKQLKU/cR8ODf6RikekD
ScYef/Y6yv8+uzcsR0/VpXOuPKn4LsdK5s3k4HsDuvCm6+ZB6XsYHIeeAFnNTZB9
Racsnn1cnb/F7uTR9O+C4v2vYRQLvpv+A6imXA6FHR1AIKqIcGO8d+gUngCYf35g
E1f/G00jYqRDSZz4tHD/KEAGe+KWvoPGEplRb9LEF8WOrGh9CpUimbT8yJWVObvC
Mjlkxyxyi3oFxaLzECylxdgvmCwL6LYUyA2+B5+vn7LT97JyUNsRIB/aiWTaNpII
efTWIkuaBMXNd5jpg//AIUtuERyvQjiAXlELVFPC1v9uGpDaUPcsnswkDdTuO32r
0fQhxZgYIxn6ZpmPYwjhlpyLYReyz3O+Ib6Fx4F+nJJagu/urGQMgRzVX+ZVQaob
w0wDdu0OQLPgutSmLyPSv1xRIfwOfciG7SzpwYkzZ+3Sb19ZjjXtH7wL4wOZ7cRB
6CrGxNpTGG8gTQ/F48Ktd7Wv+HHnIzm5a+HU9xmjjWOWKWl60X9WcE3gPN2hvecT
gNcee1XAnRXLPwZKmt3fN2UBs3uqJGobR0PP97O8lx9TQJWz+NrJHqujtupvb+6d
OGahW7nICTX5icUYDR68DgqEN/aN/5u+YTFqaJnGqA8UOEYqlx6NV4tAiMukjA8s
ui0oZWEydRgiKO/RIsLMhqpzFgGq/NfnxjPgOOPzFhOrtS8jkouGcvrZ4/HS8a5e
pBYke/R3MiR6vP228iqpra9rbGEOohZ50NQ28J1J94iQG4jVq7L9ncWtigiHfc1Z
7hkuAuIWsN6U7STBsolH1EcJLGmvlPZxSimmie2qyO6J+49Sfi2pISdRwigEAjHs
jbUYVYVMSmtfeYeT7D065r+ZHEohavALvW0MGZdXUACiCXUuc02a46c/RLsXGOzL
cUW8V8bvhoof2ZJwNWoO3NxXfzJ7oP3c1NVXh0vGAjfcrXB9KG9QPrr10LIq7pg8
zJo28UnTM9DEZ/qlt1RG1NRsTHixGghr4z5kSsQYQ3zYr40Vm4wSpAmfwrqwaEOl
lv88/Ol5QjOdCMhbFSBR5akVkNZChfn9Dc55CsezQfbBjn/AdH2w6oydMzUtNxRZ
JvIj6dfl/lRtwxaXG7kGMIezpVrtlivoBevJOD9djDhytEtyO8K+cdu6nu8bavEo
/hF8QW3Md2FlNCyu/EBii0tGpFIdskVjKxxjM2O7sIOw7i/+E9eONuNzxdGakClX
j2rIJcomRZ+xWOz2MMohI77Kn0xzmB5F1V3Ch2JFH1IRUUyRCX4bfldGFxddI8Jp
ZYvJeGKl5zmK84wqFNyD9JorUTQ0VhRNtCaO21jcEIY9ufwHdpfFKB9UUOCR0xYy
WwJz0Q21zndbXaDEWABpPn97h0l7zb+569a8tnMstkIgyaBy9BmQ+PA11JJU6QRy
buVXZoh0ZRSRTFG2y/LeAGkea7vf58FpB4l6J98CkCoIlsU9c8bPz0QDShUHyJFa
9MWfn2qt4WlpeW8h+FQyta/Q1KxMzUvyDd5RJu95wk5UNRBGxvGFWPfQxzizbPJW
15LL93cKEhAqGnLpHRTgelzKdDc8sjOnjWVqbq63eq9lzCveR+3Mq6MK5/6dXt6X
9ogv0pECMdEVHv9PXsfblp+gRcFkzxNeTRoL+ie0JK4lpmJXJUpxI7w6gTFamUtu
wri8M3WiDDRdvLw0fxpEAudjWBsYaHi/2pGXsndr6Ne0dcnZaRNfT5XdUNiXLup1
ehzft4fRRLCM8tmhtzy1xLyy2UzPixfGLEoAHZJXNEMeNJblFpdYDI+PnZ7GBU0Y
TeDvwbCswBHJqTO83pcg28X6x4tFVuwe+INLf7vCUVgfC4DbgqQK+SIrfHBhyXBr
QM3Ci194Cg7kwx8iy61L0zLIX5LQSKSmsn2AFrZUmZlvcn9+B1PJa3aBz6Qbglmv
mGVIlVFEdguvm0egaLcl8j5p4R7iu+GQ64yAyJxwSQPnYlQytFeXjAF3isItZ7Eq
RJTC3hbcXp17cruwPE6j2KSCEkX1VR3PVMrLCItAzKWZ9DFSGu72GFsUZBXS00s6
bjT5bOJvNyJUfjU2tlWluUZJ4LGn4sBcW4lLfhbtNamPxT3fhttXXCvwbfhk/5l5
k3LIFrE+97Z1ly8r+xK2Trboc0QuatalnPlQ/G17QRgJ3cS3hNaWaUCzncHNra0c
NlLeVA9ZaTZhE1gYiqLR+chrqD5HY/6/BYOlQqBMjfeF4kK+mPA/2FFSRAgkskFB
MU51aemHIBsueOVSaSYqhibC0ACLFQ8BJMgz/UznZV9VdqlInVqSdRR8NqjJJb0r
0RsG9zkP5o31m88ni1xE9MpsCopTyvko8fko3FAu8K9sAWFrLXG7u6acZvnL9DP3
JvI7mXqv3fwM29GddAhvqvfBD2OMkF0DYZ7Z0+yyYfuCGUdXuMfGhq1JJFVjnI0O
qiPWSSXrhowadVv73FH8k4TI65HaBILpCXBMEz9M5MN1FDAV/+xXjUXkhrfD+hDm
V0uWl5YA/DpqXGlO6fouxz7UDwAU4bUPfCuPdUFzl4o3eMsDbd0R7PYlnOII8pP4
JiSFs46ZFG2tkeXqJb6pzPfql2nLfIO25SY8+Apig0d+f/K3X2wa3qPvll2tdfCS
9tLWC+4ZpcgNFtK/5mcODlEbhrWw1xBDR/aR61Vyw8vqDjFvPSoYUKd29BQwb2IN
Tr3Iv7eS5WEp31LxOYTKBFibcdtTZV3voAWZPU+d5PMwJ89LVRgF+d2PYAWSOkAO
5Soxy07mOvvgMY04DM9CYocn7yPdCrDtdyGEERtL04jqXGHGmPPoswxEupeAN9LK
zg3BeaWwmjkvV68Ci/k9AfoHl49cBlqTB48pew/1fPCS3t2fihO+6lcC3l3BSIve
kxQH+jgLSbll5feoM2J3s10J7krqTnKY4BE2ex3Vegb02Oufy1zyKxhdy3KhVXMD
L55/D0e241fR6Yh2osEP0uJxZzOO3wIhsezsUq5QCfVTrPNBPKq1zks5k3A5SrZn
8noySCOD0CmwnphvuCK/D+GWJFjJmzUzfHvExm5jG0AJ9T3/aIUSbsjt/Dx/pNfD
SwdxesnN9NvZOpIrmXWSSKeeTeDXg+C5muBHByTt6v2F7FchO13opTfGAQu40dLG
GS4iplcnIgJI2l5KmDIwGRfSBYGgG9XcUXrcUHRIX/e7hpOqb+Qpvbq4/NYk6DeC
RklgaMexpNEImts6eepUNoIK7E+MN2RtchHLsLAE29bPHTWh44im+lHqA/35trN5
nSusMHkrcY1pFzv/TwUvxFNLzqGG6EWezlHFzesVV/My0/+Nlr6XEy7pTyjVWAEV
B2oPpsqMH3QxhftkikYyVXTinuCaQrr4r2L8SX3Aw6wK2vP/pmsmttH4yb007JFf
33fbzQqlIfIm+jlpWjP6AAjIVO54XPC/mIm/L7gB6ccOSwYB4djGUoZaBHJm+pqI
7YWaLbvWL5EmwBM0KfJ6CLGfhjjwWzXHudb5o1HZoJx/HnCJ4hiAk9lpHrxJHaTC
fpewbReKRjyNYb2jMMZrpDXdHKQBUsBlZD1NkJdGmeXI8Hi5xJ3Ju4ebSILbvbI/
4y3DjrdeY0FzfJTwdnVONyVpLFO8Ue0Vnowvm5XshBwP18Nz1QBxlZi3+7Jy2mps
a8aDKc1kakV4zokVrT2q2Y884Ga4cb+sE4RpwH/eJh+q1fBStltejS7Ke1LqR9pA
TMzEQhkIZtoL3sI2/ADbWQA4WL9jgDRssGHYtKCP2QQLCJPJE7hoB67jly+gAvcz
qjDXIfCrM9nWl2hfuKa4FvOXNmZYJojvBTXPEDurU1oEKXi5qso85H5gOgl3LOur
yyUhr+ZGmu1KB+U65jyvijgDZ6CzwltehKJ5H+TI2AjH+FPWYFa5rvTxQiz3zDs0
OVC8E2TBriVhC9duZZmPPfaXOrdLP78xFAkakp1oEOMTIiJDDr6Mo19V16YKlx5I
TNUdNMzvRnNzlFsSwALuUAXfTdC0c8TXudScGuAGtJQKNsvUBHbhavd9/e5H1sLH
YXjnRWIj0D0n0TRPTSGg2w2LgfLMUb3OrFGXnbhnv2y6QkcDwgr6Q0kUI/mMm0SV
jbdcTz10CI1m5AN/a179T/oq9HdtJqyAY8vw+HZFyKfJM2P6yxaFWlceknEAdAzp
i5n5RYP1U6tO3iEeL8a285QImKUohorZdQ+0KkZkFyUJ4/A8sKyUKgVo0bYLfvwN
Vuw7xSr8dK0UdZ18EcajQZI7WaC9IaOxIc0XV3V5Y2Cqh4sWkUF+yYDPoTo5Otz9
jguGu5LGziisw9YcgZYXF9y9bJu7XxekDhnoG+uOrV8CEz0QqWq1rJ4D1Xlc80oP
Xo/EJJ1tQETnz9bc2VthhGIO+SbvfcWyGKLqkH9UFQq83J/6sjIdlAWTK/z9kkyM
3IG2YImF/NygpaXAiAoF3wsJ2cqHhOgwE8zI5+uO8pDFWvV+H4EYF1huNPbnV2fQ
1d+IfF2tdWP2xmU6EuoTpwwVaz5BK/N9ejMGnqj2N8IXe5BXCYVNlEyOxyZ31D9I
POCUJa+xaVAioLRaMiqaLXRaiY8lN5ycqtp72Da79RmjpHWwKEvy9MviylUHnKVI
Dt26gX0Js8AivsLu2G89/zSWyeJG9Yyx2Eet0y57XrqhBhrsnl0DblXE+gDzioZd
mS+0rPgnNDYNmog9gaJYxJ7Rvae/hCWZl1zJpz/QjO3qWGsRJ5KTqaGbjDDGUQcB
eRd6bh3ol5ek8W9sxzuE+NtR5WtyN8fZznx7DdtwpGV4vAQ4DHTNHkigOCkKlOLC
gDgJ7Ff/KUxVD7avP+vTVqjg9QMkDQH35FNRFbSO+7MST8hU/ukxwAMrxSbfyLo2
qP+bmAlz27dJlneTfFIYrN4zsUt/n0yFy2bAHbE3Fy0gL2Mvi7mAnPGZSIlLr3/e
ujGGQDpm/szNr90Z/XsqqJX61QB1CBh8de9hzYfjqjdsSJbvNSEpAdzW8KOmVKVR
JMOjA/RgeipRU7+KKECJ2DLVx602GnaNWHuOGiWbvm9jEwgYNZkVApC+JxnriOvk
Qhgj+ogKo+xo8Q2rySYGZWOBN4Ojzyp3sTd91YJbN7blzpue8nr5Yv7rBa2CDlHt
kP1BLQmlKTm0Gbdm111imp5fkAQRqdFBdJI6zm4ajwOCD4auhvinTwyScSqO3HnR
rBxzAvCzSwz/gT02/gnFTH26hCrGtY9mVAitNJKoQUS8q5AyhhkokRgl/CCALn0O
hwL0w7+5bpy0y/F9XdS76ENNLqInD2LCksoYp84lTRprR9XJkr2JnVOAWyscRzbj
4A0n460x5UimdxH664Tq44DAzXPrVzlb3h58A1ZHhgb7hu5HCv50+V0xH1hPoK6s
IAX+3TaJiTV+LjCTz98dFTconEL75DGHY9VZ3nflKZyRtcpTsCf5YGeQ9EW7vSUo
xMX/XPi3341o9BgwCjaCq+vumZ1r3gi1LY9FNR/V+HG3nUuqNdkfUFHbAOGOL1jp
lh6UGZ+jqMLLTzgpDKYdCaxpqewSUV6y7BfxXfuG43LuoS743p96HbgzxsQU/AWP
Fcpkzdeh9JXGzUWosiYH85mDwerjMkQvgEhy9EvvD9F8ZbuhpQcw5qVL4ws33V4O
GQP9WuO4nnZdmHvtyFAFexbSQN58+FWLt2wPFDSxcqqWxrVnY0slDN7zq8MgXTf4
UhAygXnxjmEHkkn2bQs4lQ9dUpaddSaPMFdbC7gF0MaBdmlZTIWowX+7uCFDxrUX
wpeZrU5BQAzV0dQfmV6XBcuDHXLLi4QJYoFIZA+zc61BxP0XnQPo9VWuU/OP/ZpP
GOonUZlY+jQJ5teonR/+OScnl+N9oDxKV+ems0vYiFmUpunPY3UV1VSnxA6GLL6X
sFXIZxqQmw5dz/fkJnlIkNrhDJ/Nz86wQcr9Cmy08Y6K5k9JT6KU/9tlQYofYmxf
fF0Rf07AGnP/1jpAzlvfIgEuwROvIo5dskNO05Zp1tq81Pk8YpwBBb1HZtfeF91Y
EpXK8dl0eZWZFyDNp131C3r7vylI8c9/UC1mTOfG73WoP4WKh9YUUeifb8zBottX
k/LT+yLNSNFLwzo0zbqd5y5GzojYxvPhVphc2ae/lNtHg9jttmETM8Z3Ke/7tymr
9GQnnwaWYExQlbqAct/Xa9mQv7//J8jp8yAI75/JRUP3w9rWToAfUjCpMM5dV2pk
MPY6iO8BdGd8Z2Y+A23zEJxtrJcnQN8UpIWnfZXjL/E/encoP+WLro9Ng1NeQW0S
b+ZS7sdqdzQ+pPW3g3mfz7K3SQq6QsE2fr66QFdHyhM/AhueUqRxzE9vLrx33kvT
BNT9yV+QeZRVnZfw0nSz7pOQFKkvhSb7Lr/d4EpIuICYo3oiZvl0KoCwAI2YzX33
tQ0whI4eL1i8ds2i8TcEsOyHh0e9VS6AUv0uQLJeetSxiS+EQxFYV6ykedndgXpK
qAvp+gErLn3WDQ1evo3Wi8zmE5a7nz/aAtRtt6jMeef82zTaocK0o50OjKOxEkQV
FPTIcXX5FklYSQJQf7fA6XJjOT2D68Um7e134QAqUPiYao3SQNN+JmUu3+SVoYeO
TyB0aYWt6W2Cd7e2auIwpBqAFKJ2aw44jjypklki0C38gfkV6nplfecDMiShGcHF
cq6ECA1yIHQslG3wjD2ks9ufXUQx/aGD6CuHTmHO8QAF9iZoZvOp48CAMxRG+Tq4
WAiaipu2Yrov0itvUpOeN4HMgQxInTMxoPZKb+foa1v25y9uKPb+iE7OGe+bmAmJ
u8UGXKqjj8o1O1m3HfB/mEmg0o+flYs265YxjzADBiqSOcMRAEMKac5jDeB8vEoP
BFNiFSHpyWlQOKebawop2GB9Bx8/htgowOhvmWAE85O6ulRRMrCH5sYFIjoBCMhk
6sQJC76QBZdZAu1bPdw5AB32f6o6t+koe40Z1gGLQT6FTOA6Uxv6vQQHCTEkN7K5
sTKm5yBRuyTHd2Ug8h+w9zN326rzyu+oGtyop6dcBBCAd+gXpInEi5868i7UDgBq
4/VNfXzCGGg80zDlme5j9qs3ewhnqCIVNXLcKYpQjO5AmplA7FGGLCO8AtTG59kW
olfa7YITEjt3KbM0MJrYi/x5JOp9LVVwQ+5U9v0qMNbrf1Fhq1xiV7Imxxk31ICH
3Lsj6UfhNfkvD5f0s4w0csEu1//2trzXHHRxd5b8GVUOWW3tUQemoKH/yox+wGzM
jzL63tnoQQpCMZZiaBUN/JgUbyvZ9a0ilCH6E1TNvK4JpvkHhNUZ/Do2crHjfeeK
o7y9hcYTRQs0LGIn/rQB5cyHVSWsy/RMcB2Mv9l0cFdozrUv+IclzF2vr1kAcC9F
d2XFCt3L+hklcaiGBN2yZWCxp+ckpZPMTagU0CgULLVzr2DTMTdNvq4lsCVWOmqd
pNO5q5P+st4wkagc5D/EHfIFCiKEIvmqjZSXkghCEIoiUYkEOkOzPmAXpIFHsv0G
1UldqxLQA79r0OYshfWDd+ucXbVbPy15ClQQnAm0FHCygzXEei46M1SvW2C6D6TT
Dp/g0EFbcCe5dLb0BhK5hBzH/croyNJ8mqkiL6RdA0h941qdftboVlZW36k0Gfwv
Tg5DN0jMvLFGGQMo1mgJL77K9REsgJd4Be3gbOrdYR/rQaWF2dEcma4UZIsLyKgV
rX76KcYO6nMaTEl08XmmmljBkjbXKMNe8ckc6sBkaBZfV7RWDWwXJwFQOxibn/7t
028mScujQFby37IvLWbvOXm/Hc181o+YWCVUvQnpiqxN3P0g13EFcmmECsKh0g8j
illSrnQy/ThFpIeY8FaAh4ZJiqqLzVHliBONaetVThsWG/h6CZJ6EAI3vR/ZpUY5
6FKEFuxN4bXRd6JVWVyHaxLQh07ILdO7wpzZA/Cvx7/Ut5LOOX04Yq8CIroghmuW
xU7Byr4tKcY35wOif+TLzMCK40YIg4v2AKfx+qQXDchiEaKYYGpxIIs/NMNqQ4wn
Wohc+GwjblPILctn0PSerhbHP4ngk+3zoSP/IVNooUaFQKQTCFqBczdYztS+Twdm
dBTXZIuo+s9lwqKcnC93ifzmfPAKSI33Le1BEEcpYHjHIythTz9dBbBz3xQmAUVP
DG/6caW2gmL4HSkgSfKPQrUY/jR/480nKeMjnJ7G7uby7YHMfuGknXQibv2RoHmC
dFd3l4cJcEpY9USdsiUqZrRoRTLxJ/uXuOo5jkKvfUxIc2LwVXVOtPBy88UQDO+I
OZtoYCzPZsdmXZQKfJGB8aGpa1+Xgj754KS9AhXxz2IAd2G8xvBKW3a4GA+hUnWE
hAEXLmm3uFsNcLFD0yyWbFHXDnBVFtj8MCUz/bo1FuLHkYbwekwTY2o16YNv34VP
ZjxnYVsmnXbNWj7kn/G3+lNxDCkbylMctkhFS908815VIir42kiMP25SpvaUKGXg
GuKN3upFA7QYT5Hk70P2IVL/JSH8S8xBDusBMRrDG2pSKEfmU5N6y9845MrLhyY3
/0db8tClH9QNf/ovEGaZhIIsnWRlmHFpLgiEXOVwMmRFomlz8lYbXTBQ1tL/5LBg
D26itkB8yaRCotl/bmG3IAjFY5A8pzdtMQNE62ssJEilRX3X+7I/sgSJ2ekLCB5B
9vfmcLgF/HNP3eplFAGO9T/D1gVJ99cb0WPvQq1HiNbg018ZOx/S5sUR0r5WkoG2
iA4nEFWKslm/lm/udQaF6vovg8ZwIfLvqwQa+40V+EXx9joKlTTFo/PdkvZI+Jxr
4yMlZIwfbo2rMXFE4URUXOS8aBNEdSiR+G/uHMccVGphW2MSvKxOlKcvbJUl8LTe
2VTJ9PdtH5Ulmhkf6aEWi9XAYdQH3WpndR4oxB0QQZOonQfNxrC4gHZrUCowOv53
ejg7cvEy7zqHwxgx+3NH0HokP3lim1DUOFXxENiKaLNms4nwm0aA79Ecmkbp6q/2
b1aazWOsEwHYpXmbm9vFVOBfcs4RFyB0v6ENxmBggeMnLhYTFDN//UJOViumopAc
RQAPLeP21xdifEec292TWTmqShS8sBdxKDe/a9WRmnenOrE0aXeeF5ZvJ5+cpf7l
qSVawN807HjnY8497ZdRZ46/3vTr9579JiiLq5flDobCGYU9GbZwpKiV36+BzpFp
XBtBLHLPjtov0WCz9q5g+cUI981gLKg3GrtjJnHT7SthF3ucVCOo1YDMs0bgxykj
FpO1ODHFEcKxrfIqaekn2RQR40l7CdDPeXMWlHE2z8wFtKU5dR3qBeyKRDHqBH7s
/F5DW++hiwn/MmO4bIBmLqClrPH7qV0o6LnUE6uhY2WYDq7DJKBKxd/JEiWYMTlT
Xr3lQOUJedJijRf8PvnpSEXfmGTpsivyMPZfbzgshd0SLB8FyE72QWs78zOy59xu
cys8lgNnHUB7fhnhqqnCT1v5I2tSRoxEdlqj7h537bEU5WjO3smxWmRlNxyO3lM5
ydV7JXIBZEduGPIxGb/HtBYCJeUsLLg1ZgoA/8gvL+q8VrDKKlBOsf/Wl7aWBqcB
sPnFKO631rI89ap4UZ1aG3KBZB/1Wb67aDFe5hXbqZLYi+s1G5GnSsbAwCAgukGZ
T55t6//4+9f3zwAM9TX362H0S9xud3yIRMaBC63zLBIoQO4VMUdprHb4j4zvl/61
2GxDDtxwVBv9SmMtVWyBIVDXeFrgyTzWcMYez3mOeE2AnQBiVCSrgX+dG+2ZjKbt
bctzqPbJDlNivZ6HOgG9bG/vp3adEgmJL8ebQDEegGWel44w/U7CMwbsJLvWgvpm
nvpMEH5N29OnZEStF7IlJH4Wl4EH5bieOP9+faqoox5p6X7K9fp1v8SFDLj+p7VK
wiZBxiZR9ne5U3oH3tVIz9OJ5i17rAcuTJLHIfKmxoheu8fO6KdDfjwd9v8Z2hOS
A+tuQKpRWw3I6LS4LqCG1TsZIOegITtGY5HBHHvKU5hKmpV7ve9DOCgY8iRm3ssJ
S9G1Rpa+/7wqaF7/NDL/KH9znM4rhTu6CAMa7icZbVPghwP3Kj/Jfl/OeAmhwiYm
Aa4Ah1u4iJkfkYPBr6At1bLYe16aUPreGNCo7akIe1Gs/gKFVKRdQ3QC79vgagCZ
gOv8PvRS/E69pOSHta9KhKXeJIZpgK93HkAdynp+rqiZlDJ/opbMF0L93XjT2EU5
hjqmI/aASl7qF/6ONLWxaT7xx/4bRjAK9vvNq25MzubrYQK5L1rnBOsb/dsEJ6t5
iPw2syRz9D/RNPI7c+3CvgiZEpJHiyrJL0X5Q2Sbkj7aQQ8enBRA4QO6zUtMb+Xw
DyZSCYLM08OhAQP5Okdqee7VIxY92gpsuucOFLDHcETjHox2ajdR0cDxl2T9P627
qPK2pXEjKIRY3y0EVUuLtvkXA1o7c0yfFXVUOTasam0Z7WoS/+wtqp2x6B5HW9yd
CU7RCkw4EjkdBV77xumaEmTw7QxRo5n3qrii19CJE9gdrNVJwuxb6/WHEb1UcW7x
IXBoMr9RmAwH6crt6x3TfDozslsGsVeA1G2bsDyHGzgke2/61A5yzJ9HqhSIq2Jf
YIUoc/rrDjJpN66PHBFVLqZPTAJNxWzs7esWxA/qdZ/okNUg+GFVr+dBZsjDDZCr
oKDfhh/8Ddcm04gFMYrqhSNnigd+3pL2OffeqvUzGkAlNoFrjRwh9SBOWIk4vIXN
cM2uIhBgDoOwMB7AO3wfdQkKLyEnxmhVHNngnhNBbXlBUNkxYk8V/enlZOeUD61j
UAyAIqu/O+/wZtimpgfZLTe1lsMUudXkix+ZrKg3N2VeYtg9qIfRBoBmJmQNGcZ5
tMu/JWn8kSQY674Qi0KoBr1UnMZPUOt+VrRH8DyySapL06qBMeIX7rMVe9jtzW13
BZOImkS9LgFB+Stpt4zmiygLP6nuwm9kkDGSSOuzr86y1308LCIU5xroKyxj9XIk
lv50owefXeAcR1YbnCqzjXi6vGnznHIQgXxCUF2IMtlITWsfI3v+LAM+OygfSXMS
GY78jjVhfHrSPPNRaKlt4nGkBhW1umQE9DHCLPDXSWJL6RgXKAMj7tSD6dEGMNGO
GkMGy/YxDCo+z+k68omlWA5RnEkn/E2OIOYY3um+jtHcURSFh3iTa4594f1FpdZg
eRmTLpyy/nrD3JBPIpw2ElvgV86o+Zh4YuGinoQdwsGu/dFNSmHewguLks1CPGGC
hLK1Db93dLjgQRMtncqpQuhm1ygLfn+OPdjtvPJq4//ESR7fKkTMTiXy1E9Cg9zy
LQ3PCr+F93fRt5OQW5XM9ocIY6J1laU34rqM+8KcMpR2HBkdqSgprMsDVfggYfxv
+x5Yh/u2E/yWIKEfOvEOtJFaudJDrLZqW9+KPx+T3lFRiEQAOZqh7YkAFdkHT6Wg
V3jBbabupb5Ijw4LWacPZkTfrtCOeKId6UJQ/Nhib9SjzFyF8aL9tZbjPXbUq5K/
FQlU/qSiBQAdaujJGg8nDO41/r1xv+WRyQbWoywqSlVj7Lfn3RsAQGqE7bTLGv6O
Zipo1g3ssqIaU6Xj0HQXARgqPQx2cKTUWH2olfTC/S/Hwrl+BBuTonn/zZCGVz1f
KQTqntmlQ9KdFUVYQBQQXYqrm2dJxcZQZV+jcZ9GzrDYM15ZrkOji3nLraH47p53
buzgFlSgsWBl5O3lukgk+/Ug7wbmdklWhwURF5XcscAQG/UnNybR7FEKDo1Pt31b
22ps+XfN6J56K5tnYVZEXB85VIiFji+Jj8lhqjlBbtP05S6b2kxJ9tE6VDYjNGgp
PlfgUQPWG+wYPZvMzBVN2mMHnjd5044C6GGn+0sok+IyerSi6C1Clu3e8WDuiYXI
+f53a7MqJOyt0nIYTaacFDAFEwCnTOK0y3qZ+wIqCg57vMX2kDoUM1uHVWYYMQG0
NA0t3+p+oo4ofWdjboivRf29CE5s39ag6PPYODu9+Bv7kmG+brpJBzEHKQsWUWMt
cquqlreA+527kIJrDGC6Hq6JNKmGagMWuRrtmrSqA7Rj81VJAuJg9Rz4x3J3VFcm
uYzHdVWJQvJ5ykbCxEw3wkPvOg5xFWBTmrbxJQ8/Z98JIPhs5K6g3TeqtT9VRT2Q
5SKD5npWpbscpn0Y60pEKX/t5S6CRPx9g/7o3gnJbyF4OUClqa3t1qsC777KEanK
TuZis/n1r+Hb3MTBrSOtMTttANOEITElVpZ8lynJrsT8So2FZE3R+h6l0/fUBQo/
PcyiGXYdp6jICGjoaYBlQyjxq4JerrbOuliKaiRf3eUIIGvkE8EUtitlGXIbPJAe
PPdecVuqUldVIOaKjJbtYjWPRKF+kZShM9AYlv2+7oQSzw2yHfLm2VhUTvzG6Fro
1Ek1rn6KeplO1UMI7mvdgFjZ1wjO97l1SHAJT9un55/BSAAwtWLSZfY7jO00d824
6K+GkZtExlr4CBG3Uic9+bGupsMIdchIEKm+PxrvdsvXFhi9vujemAMwXHAvODkA
sLwoauwzSs+FbRg+UjnxKggG/bWRYBR4aBxXDvhi4sD/eQbntmSqZxFzZvJARdGY
9N7U0W0kS+LSDaPiYJNNXWdLEd0i5jOrR9bFfxJHrXvHxCnOJSo6idZCvrRWpzkn
HuEFURrHhe8/njhUTOCj1IKDFYMlgQs4vUoXK+xuKGGgce1fOzk9d6zuLwx4Ug86
0tRzf45B9o3nVI0yYXCU1J/PObXHHjXaBjaTL4KViy2xugsuOl7DTMv+ff5QDQak
2YekSwsyfhXFvCG2vKo/O+jNRVRXddp0II3KUv0eM4mx5ZX5tH01l2kMC854axH7
P+O053hDVLeeSncn6WhCM8gwR9ucFytAMytyLvpZr2LFGZOGC35mWSRA5Pb/Uh8J
2f2TKT2YDTFrKa7NOLMCl3gqFE8u9g9yBQPToP5vwo4SSopSFALtDFnt8WXzhEG7
Q71wjAcp7owFwtMit75QXOziJU/E5n5V2IN9Z0dG61wNQNIafpO00IGmiS+aZMPK
AY5ey1zoRD3s1dOHW35tU1K7OolWy67kj3GhDh5c7W4PWRvxBl/ApawwInLLWfdw
lbWVc5idaeoVvD0a5/qEQN9eWUMfcfpuT1fERSqlgMviP0Y2k8ZhzWDbWLXX0gcH
XAfiznIYilYHQxZDf0/oi7l86lG1BJgJgtDxycJK9h9cJSmPsngX6tZnZpcMd3bB
zFbF3MXKhW4v68fV0fwjDsQmr2jJQR512UlwN7l2qSiAXOmeYW8U2F8MTEvofOKT
/II+szP9KPLbIPpAA6QA1vioKpxytVOV1eJ86mnFkpcf4sPXRVWvdGwf1GTBl0K8
jhJxejrR8jwmqq0EvnfvE7jkrgHxe4kKxcfoHgpfGKB7hXhotNDHu8rbOg4YUenZ
fMlD+Xs4nOU9+d6X0upi11tw/cy7cF70F+9iXlvW6U3MMsSxwBlMK5u002hi8PNq
FYsNhwk8mMunXYiKR3RLCETB6jDersuKHKtP8sLfIAyNCcALS/l1pKaXnTsrfHRb
1btIzLF83ecOHJ6sXklVfGyNqLmiRCfP9ZVLaicKYvbrzJ+Icfbong8wyizMrXdO
1Agqkb/0tVowhr47RsKKtdH5HNUSPwsE39GVte40ZFj/XEkJJS1ttWlJKz7QoBhy
7+1Y1G6lAxprcZG8s2bp48gINtA+nRKxIqGahnCLBbn51XknxKqitpakXss+YPWE
6O59JYxEqg7VNQ2/YR05kWiyYgKXPhCFqTd6eHMzib8PvncOQiMAwXTy6hj8kU1+
T+RA//867K/80S1qU9uLo7w6xg06hId8hLKi9k9p1g6gjPzzGUOTPEhc9CZqryWe
F2RSKThwuNG8s4R98ExSwFh14ua7UTDebkbix1tDJT0D9N912t1mZNSZV0OaZG5D
4PArHKD+5wleIOI5FkyG8n7Y5LSxm2nzrQsi2xaDXEesvkgA00r/ix8cvBWXFwlf
On6HqU4zJOEuNX08RglfoX+dQ7rsKC8ZQ0fcve/U9MNbmbiziSGAPOlN4uOxSXBM
zf1S9vhM4nFRW3zp69MSEydtKqWGDlm/7V3jY2saotW2YO3roC0aPPDzot8lFi+S
JRxQiJuiTx3hPOS1Am3R7CrTMPVgMidxOZYa3oz+7MS/jZFeQkJHNZpvR/wtpNe7
WQ86TMgnRHAcoNbeIX0Vrj9m0G/bMAGIDBIoxQRsGEiOh1XYudF6X5pxD12PpVCg
9IsGWEVfuUUA4w0ePw91RGmuA/tcLs/+81p7H93+mI9Oig/f3UHKBWwAqkb388xZ
lrNN76Dyxk3EeCEheVnCakepEzJrQ05OeiWivmuprQa/bj1EO+7jnv01kp2NeOeW
5ssrRGC5LOX9HV6Expsvr19qJH+kdZpDmynty0eGg8Pj3KoIbsLyqRAK00PDLG2D
y85LYhTl7rTaxf6PzaHuZf7wxy/mhsJyXzBEc01yOhkkereldqqWZKi7dybuufsX
DCkyasg5hpzGMM/YA+D8bAJRePrygEorgXUWzK41oTnloNVh63smUMpPP8TpX+kT
6JBLq8oTgymkvYeWUkH1a8f9QVmmQ96v4DhidA4CskWLkKNs1Emlaxf33KOD0NAm
84pSXf1DapR4QHLyKBMEcelWrI7PtVvbf/CtiBLOqFi9nonuB0RtA9Ec88LSQvZG
8t7CLNnhYGjaqWm2EOa6QdJMEBLrM9bOuy3iG10XVajkTuasmGuY2WA8jyNVuahy
9SE7ezN58WgyV1e3ACJVan8+OkmWF7TKJnzDafkk2vv53OyWyXiWnvTKc2F50yDW
CYWihLE2l6t4TctjR9iKmysZK+hon2bF0bYKbaEgSVRan7YAvP9XimL0zIsazcAj
Wtc8V41FVmtT3X0J0CQqnUO66teelp66XiqSgn2m7nKFF8fLLHomufndrLjuj11s
nWjrnMeZtDEPWrRPXFPtIpNRgNo25fXApsGSwZ4j7wnEcbEULlnZIA282xJ/xD6y
+c1kRoZEzyE3gmsHWSC72CVBWX/f38p22YY47AQAlaiaHFXSIOXTnnbXf2IIHzy0
/GMkNzdjcnfV3vyHT9aXdu4LtCLh4Nurs+GnzBORHaL3JE+tdG1zxxCiDuDp6MYU
7klTGP2ZhBaFbwnjm4v+xBt3ZRPvXF4X9TliH4zPgMoYweE1hsaxYGlTnpdY0v4g
8AXQZWHRDsxVIgLHgcnyg0AETx7+zxsFemTOX8v+3sFNXkGu3pXG3ZLW7R7wLFli
WJPGvdNsLw1GR8e65siln7Gvh0ck4RW421xMz0ZQkEPargfyLySU9nHvt+0hkCqH
t4u0GOns+wb8enUOUu3L1lInPkV/RPDDT4bCc+NQw09dy7CxfVvTaq2LCBUYxF4Q
Tz37qZPZq8UurJZvMNnDAl/DdKAJGxuD5ryOru3t4NDkkjPXUkb+gBJVPfXBH0Nl
fUFR9ibo3rUV3YZi65++9XlunHf+1W0txuTWqtADlsS720ipfbKdSc34aWmpCmDv
XyEFSPq1yQbd/Dm/EtycM0roddR8w+ZbaolIY4wEUqGWuE/qDLnTiVQgD7h+HnsP
exbGrh5yKE67FGzZk+XTxqMLVvDSjJFiLrGVH8XLCgRp439Sk5Me8p+HPNDM9Iym
7HnAvNVV6c85cZbi3BITuX95LBgHSqYwYGEjrMGVqcnGoIG3H3CcCaP4JjHTze4f
jcAKx5w74dzH7EzrFNQfksi539adXgP6xQQbSc0NdQSMYh+frqxtJs4egO93oy3s
PhMnkSrg7Icvuhawj+9L5P6X6FtoXujymAPb6J9gCA6IWxv2DTp0DRFTEtZEmzhU
ES8PniQdiZ/YisPuPjJ/5HOu5mWCeGRHMtc+OieMj93izLYUgrWWbviY9Y7STDwu
JrfltFFQqenI4pplYxiZUWuScCJ8uXQvTpUS97g9ExW9sYv8Q9Qiv5lZjDCe6lK8
45cAoq/3cgeJ8Y3Q3t87LQXdgsbFNlGVg4zm7DP8jcPoNZWvb+G0gq4qBWC/NEBs
Vl/mg+VS/gudTH5kn5PkVyHTajUO6x05BgKTOK6GXmhpE7FLFnxlaecXFtB1G5Qd
IqE34hN7JroiqZQbBZhrihjAGyHDtg6Lp2h19bYlkjaqaMltoASYP3TJfxhxDSHY
382POKq7ipzXkEn55FTouc/DXtGQMr1GTWDO1FlkLmCZzMv1c1wDqFkwpCmXHKhi
sktV0PDdDYSJwZ/Qb56+idsfvF2JeDQBBNg+dr+WLMtdsM+xK2crQtqW7grgRXNW
eUAC18uYy4daamBURZA9jNGzLfjbjX9+rA+kuV0jgG3XuSJwcfM9e11sQj/mXZIJ
MQWECXrxb8RRykn6+b58lUPlrejyfUEvbUd0MFWrOWJRZ5Isokg43NJsFOLnYM0l
PE9codfVq6aaCxRQF439oh/n/PZpGH3QxiwfJvQjOlfAOFhIc0qLXzB1LOlBqdrb
c7SCcMvVW6blklqXBr4ADL+hHh2fG+l0mykWgvEJIcqipylOP1kdCzF/QrOQy6ee
hapP/+Wa9F4wM7zazl9jGEl83lJnYyge8v4goaSf5Qrbbsg3EU2hiIJQuuHZlCCX
pOgk4Nxdy8oYlh+Bks0lTTy76DK+aoZ9bX3Ol/6rU9apEiV9DXCmuErm546odsmS
fmMCEqT4bWxulp9GFdwaRAc2g4rjaXEZmQEBIEnQ82/FTaK76D6JFHhDKVrj/J7u
n6Ywtj1RyePyaP5KKaOIxPyyj4xK0XNJHsELzNEbRZhJ2TjT4eP//ELlFfo7F2bB
kpnRXTF3eegoi61MaG1CIdjD3oUKSMocvFoSv0jWu0C5w7hqUTMt6ejtdJvVf6EV
Qh/v4cB1oQlif0ouNVJmdHiI7eOpmPYY1mktwhSzkmPVKAP35fsCMMYv2SlZ6QUy
o5FJh4JDqCHdaAQ8aGV19nxvPc9xbxy7e/1PPwJTeHbkU//FCdGoeY5aMuAdjc9J
LTdGq0lwWMya+r2M5AnoScICoVvVXqXaZO72IVRPTJT/4AM0T0mZhtIBWNMKOiUV
p4baJKdAgd+X/X53pVWz9es7sI/dcVaoPvybULWSrTPb+mOWakJ4Hisfy5hMRN8b
19Rmcl26heW/S/3DwdU88Dd5MxhB83uVujYsqyCVjpfBngNKvjjIL5aGuW7kkGWf
QAVm6QScEpoWHjWG5G7enaGh1piTN3PPOhZjn7Mb0O8e7Ki6RF5uT/IVFx3eP8zC
YYLfVO5PyVY/XE/t6Pu32DrTm4L0U/XVVogldz0gwVUFNTpChcBu2cpd/JL+Uyt5
lDGXB/kGRXvMYePIiopyhrgex8H4ne3b/ED1BClQelgmj3M+SG8pnKWfR0cP94Rw
FWUZjCVYKPRfUFT2TK2R4gkmuAl7Qor6mklVdg7Hois04Rk6NQ5UneSMKMD71s7x
dr8Pp/67CnHbKXjGusuakrVbsBo4ynLV1ugU2iQ8EPIGvAxHd13zAha5XXX0pLGT
vPumv96RfnQ61MVTCtNRUUP/dGKeoLGtAMgYP1s6L94nSzt0q1ooxIFSMLwSgQzt
IlEu9RaMwYr0k/lTPqoWvaCc61EEnQHnWGznAktXdco88AHTJ+PKDK0XWAvuqjyz
VAXt0qumIi6ftkwJYWiSEO2NwRyTFhRjSHgbBMenRg/JHOgNyaixdKbgrI1aDH39
kyWKSa4TRiqodyxZ9E+q9ZjNzXYAOb51548ZYwvPACW8s3PeHy4B/ARnOdYnLKFr
8uhEiyAWCBjHJta8AD/CyCM3NopTeAL6p3fYrbDCJU/lhjORTuMd4mQBvs5w42s9
71YSTE410b/xJ+9Mzc0s3SxB66EMgQMXmUN0LQXLM7VKAntmw0aUWJ8Cy7tW6a8I
V5qkGo+lpV6m87qSVZgW6SChYKAnPegCCH0twhQ/YbBy4S2+ifceiTbSmq2G7hWS
MQzcWNj0i9RBuv3HMGU4fnzUyr9Arbmcl3pY/ZhrtR9xAGycqIMd52IjpFBlAeqZ
auB4H6J7lw+z0XT0dECabUklLOyoXZbC6eriJ4kv6LeLx6bEWGOz04UxEDu2l3SQ
2CwhvmIoNBQoKtdFaYr5Y4DdPRC/6R8nHrPO87DeDOa1IblLK/tHZPVJkc2XwXk1
6jJTky7bK1gBfE96tSItUlka9mgRjPg48iBKwD0Va6V6ibf/Qql1JFC5AGNWFj0G
MU3S3DmlNcjs7Y/7QbG30rIn+eEpeQ9eqwKrIWgXnu56NxVDUpWXPx8RzL2s6wKr
cZzKH4xp7afsvECs9zJAvsWlk/bDxOJTV6Eg1qqZQJ//tgfPZWfKnJvBN2n7UFBx
ivLppQkhtd8xuwChk5N5Pu1I8SoJfGQRzgsXS6eC0noR3Ow1uN5khc2Lz+0Auux/
Y3ifnbyWPyV4i0ySQKXHsvIlH44SvQ0Ddkjc8x4wk2EQbE9kUQ7H8pJATJdi0eWF
3k+rhCo+1jbUW64HztY7B50C3Z0YwRlILB4Ze2FL1BRPdVPlg6w3XMAv5lnyM4d7
q2NdZLRp6dA1MLUZbjSL5ZSCyKsu9Ew5q6iIyVK7A3YiamSFuZjJwj2XcQIljMSW
euwGHx4b8sDbUKy/tTskq9WCVQqdcyDtrRhmHeHhcRQXVscJErweXxPpv9u0ClKh
MFki3lEPeohoQgQGt7ynil03wVGmGlcBzek1mQjJrW9/ztprwrpzdEkU+mDDP3GN
8OiYQ79iUjadFkpE3DrN8/og4ycBL4WyGXZkA2pv0KGSm6kOwxWIPgL2DOc5CoKz
hyMuQaqd2+3PXQ7a5Oq+9YXiYa+HbWZ9UqcoO1EBLhDB2StB7ExI4NGjxP35gOUn
JUCpHqJENkt5RL2KayBiGDxCQAxwdaG7ZFVDcklewJE3kMEhp+X8sZjFI/ZYvjr4
ah6H4XtH5y0Z7p/0q51FWGCtHms4zVV2AKuwlAc28Upax9RmI0VVXvvARU5dEZN2
S1DqpPMgoXLIcEVwZeVm2gRCRJnzEArKwg/Kc+VvvZGev/asYsegF6OyKVna7Dy/
6+m8U4NZCDcIKr+Y+4yggqZQFJGsZcJ1VT/xFfPhOppGDfE1XapzOiToQ+4zG4ZB
EOCJ+JLuJKzDJiEzRwyLxtrVbYCHeQoqt8BabRepGRVdFnFcTGObMHVM7hXbgoK3
/v6gBzOGBjqFoqgjUAahosnvzZHARxxqhMCnkLbZAdZWEyTvTH3ZKDxQGU+QbsyF
uU6wxMCDL2wgA9gA7SPd/IrjbQG4GvcqhAFDUx7MVASH2YkAkTHtdA2uL2SNnAdJ
W2oS0ZlEA5XVYVObnmU0t8zMeo9tYg6aOP/DBBWtDQzdynTHrsGbxDg4Vb/zK1Wn
UFickq0XQ8mg/YPz93bisbwIVmx8EgYT2Oh2UpTpuGd+e3P7aocKMm6ZSSWL4ooS
6/08CHea9XRwR40vgH3DBGO2aKc/yoojli2kdxGUpbZ+J1FIm6WZ3Vn4UsuMpxmu
UBqJTCQbBp3HyzspIAVo5QbYTX2bkgNO7u+1cGiK3Ag0y+EOLX1SIDe2/8vK3bHj
2Mlfii5OaUyE9lXZtqYLSgPoxk7B07g53OofN5zz4Vzonn8TA79dT0aBCnbuQc9y
kZ97GbcIyBFG7iRZymVEQwAywBR/jyceTG3EhBb6t2PfikJhRG7tZ1qA1TyXoVwb
4E1CHuu2kf0cm3CGKEuN8lbRap/XEX0Gfy0IUEC4J2rPmbq0eJNvLnBcbg8lH5j8
37cdvAnlYL6Sdo6dfXgJfpDrHL/q+UNRJ4R7vuxW6BCkjbGqR6V3LO7VskTisgqx
+B1THy630lolwE84n5N7M76ibRKflVJAngYsQ65jiaYbl1/JgB9paBzfoM/Z7QgI
BDI8et6exwmXlHX5Vn0HEnYCiDU/XsCG2hERlv0Z+Srztaf69YFGiyTFaew4TVa3
K/z2uRoHK2Q9sh7vdHAYr7v6cCmc39jXYQrEuUwLpBzfXrE97pv5Nm0UjR1KAnDZ
+m3v8ZSp7qIQIUD9ZDCwCuN/dTaV8alFcTi11doRclpkrcnk6z6trSOeaLpMkDxD
pSPfgCmcYQagmQK02S2rKPNMTQVs4cEJ4PTwWMxrvKAfxjXkk+PnBwzxNvgOSp5q
iSOJuSbcgmZX1GKiRJ4l+OsB3nBHwgExmvShhfsKjFaaY2RNOnJSBqOifBw9W2QC
3zp8xuOYkwE+Nus9etq58EL4srGQdstKHgF4XEjRIaJIGzhaGfHpzpw4nPaRQnMG
ffauc/PI0oHil3mZajb7joJR4QE9h3DI55TxKd0gWD7pNBBQnl7A95D+7Su+9/hv
Krn7phFNA1+rtYth1qClE74IkuUVNZbYD7W2vCAb4o0VN24R0hZ6ITKaV+nh04XE
xpyXSz2me78dy2Pel0AOt4O0d2saN8j5XCYN3pGUf6JxYYq9pUAo+qi7GCHSYHhu
UFsEZTbCw6U+Wsh5neWwivVYmfeDVn2GICnfN48i4XB0ky+/qKl/bXRu5nm2ttcS
hiIu5BsgCHhQQzzZnxbI0v4w8F9PkVMB2NEW0NTlMhdWGQjY6Ke0Uy3P0NkWRZhl
OYEqMZK37RGga4+chUvYlHPg2hig+JxT5ei2o2doaAxf47Q2EQO0bvFZ1HWDGyHh
k9DQYpCCIbWWvicLDCy39Odzblw6EzWMcyPj9mHjTIiKb59rr9NKHQ72G6Nn/6V+
0IISaWySc0iYgTp24XXUSrj2TwRqHCCiKWWDJdwAwuSBJPACTnj26C3At/rXw0K8
7L6ynDLBC9t0aeoKbwLsZZr+koOQlQnCmpcif2HhoaghJCAl9xyslX1WRE3vlP81
StFTmeovhWhKtR7f9H/rVFXJ6lmSV9V6BZskIv2bJqhudBjDQi02ym1n+nBIEJ5+
H9NDpGZ37gP0q8iNPXZf1cXSRQlmdqbXUnSt2ri4+tsMvkNP6PEQww2wFB3qYLDd
hl4qIjWyRoVaT5fBO15t/pG7S2Ja+vtUbZbnzREENNZdmNnRRwoN+1ktcmeww47d
NkrcOLGvFONFxWM4n5clFueFowVcwZJ1NYm+4ms7yO0dp4wlRIpI9sobKJK1hjMP
QetRyrqh35B/gxXg8Hapl2TefLUyY2ceuj7wTHF0yXLKuXOo8Bg97b9xyV9oOK9/
9n0Z3tzh4GxFFbKFBseL/ExLXsGtN5PitgJAo/Gv5o/IdR+PqtzXX+tPRKI0+hE+
jyKgWF4VboENaKnpnaWNHtpJA6i4mPKgNpD8lthOYe1E34aTYd6ykP8SA8lcs/mN
LCaTtYwvzFbsTycMx1eI4GlMQSK8i+7naaGVr7nN6Y4D0ecA86jgavkeI26Am6Q8
3+TxXQshpTWFa5QYfCV0+k5X6smtwODOCq3qjwQPo2PMjSsrmxK0tivHT+0gZzXH
4P20D0cMcmo3djKn7/9tE2c1mWH6sMAo+I+0hpA3zC8m+heaCBBLgpFZVMfZiQ97
j+adR07StDcEJdmFPERs9GLDAm0UUWoLLPM76ZyJnyL2s4LyfkrPQ1nTWKsApj7Y
R8K5wTWTCU4KvpOB8trvxgETXbzODH+SinuDu/pafYT0jqPavTbfwuQCOMVdy5aM
C9oqxQXTBnIW1ikQrVIffZyOIhXEYRaWyqKNKRjeOYghdWze/Z8Hm9NSSRo8nrRR
2XT95ZAudxfPTkiGzbRNTQ/H+vVKIqaONTGJuWyPAwhvCQSbpwsPFh2wSeKkbFhs
3oIvi1q/n5bUpU4VTZaesyPcg5DFgfRl2u9EZXUAODi1JaSY4FzSdE2/Axnhp+y2
N19S2FNYQhs+Yyw9WBh+hY7IKip/T24x+Q4jvTF8SUl26s1XoGVRT3PuawrKzg9T
wGlX7A2KH8O6bepFvpbi/O1ZhM8Uha+eJKuuzBvLBnhUOYQ3SGajtiI7oftzpzQY
dgVj0obcp4P0vwiuDnydw34dwdqh+8jLN8BWGzS72aJLBHlouIeqUGQbjMKz+Qu3
cfIV6xgZmu2sSFQMz4bxERItj52G6pvniqLjy0pulxWAJ197kaaNiVH65IlkxUqd
mT45KtURpTA0BD8dSCqBC1bua4+pVnzf91kYVEBfCi5b/Lmj1451iu1cMFtBy0RS
AeBYgUEwigSVlKZeVUDsUJFQVxcwR20Dqs/fNJ2i4EwvF6Bb/NsF849ZejK5MO2S
h1QKCmm9rcstvGMo+edvDKDhuDo7dX7ItCWN/LhLTcX29PNwgCQN+AT5VMrIlK9d
gynzhzN39+HD+I+68Wm/bfetPEG3Kas2rZPUCCW9+lnUCf55LVCh8hm/a5hovi/A
GBJ0ngNBMirQayz60iK4ec2oTU0wgbmHb5RSOBgJC7MnKirVVHUX9ruKHjWUO/Gk
brIJETwJUwjXwldDtkcTbIEnwYSL6fLv5ETw7RLebg1mIWntGrZmUlDoWlKMJNJx
FsvQOtU7jdDTb52LcyV4J4JbXmjrGGLvTaFog/tibdzwhvpQRTxi2sTYjrhAkwnW
1CiY2VcrP4lbOaLxF14Ae9LYLauu95KfUHOZyuzGobV5ct/LgMyYDby8IyiyEMma
q3Qr2S0NdoTe68OUqOvbr8+x0eFc4eU8TXCeeWxb8LicIv0qlZ9XPiTgb7WpJgHE
jCFcHplWoStMAcYK4Ql+ZyE2zZ0Q29mL26fnv2dRkZQas0G3Ke42UyKh8tm4w1eO
G2CRLzIShzy9XU+Z66LtaFe6c7d5A8b/vusHvj5XLLZJMAZXEd3T3CeCU9AFOcMZ
GxN9goD+L1XIj2LLDhWrbBKe1fFn+EunxK1bZZL2crAX9IomPk7bFmmo1VllV43U
QNJOoYDgqi3+Zr9BmBfyju67f6eiYqGgGglZiUaVeED2GGPt8uR5Nb7tr1HWBPiv
GpoFtbBsnzwNjyx43H48LMTnBy+o0VFFSd2mqjD08K3QW/gx0BOhCBIvnTsUe0ab
2KF7LxbLVB7hS7U3JSYdR2zExPO49HkkrnDn4HGkwjX+siixbiXjqJ/kVy8n7Rak
Um8K2UEPtSnSDbwUwKrv0lz8dkUWhJKgw/r20MRIiHmHV7GWdFMUdLY+B4KGwy6x
yUxr7yHXHrEetTMN52U/sNN004mGQ/DQA7B5WQ7K0GuITvbnu/bT/EWlR4xcLYSa
JHnOv5Gd4NHJWyWv8uLRaPgvqHl5b6Gz72L7R7eKLmBBDrxVQHjTxYV/kaWcGh+4
+d1ddUvl1EjflyJ9nj/d7Ry9/MSdKpav5kZC23JWwFvrVV3aqQrjDla5j62spqBT
Im29I5Hzfh8UpbQZvWhmAJhxuiNJz6W1OlKx2Wu30Q6DnA3CfgS1nRWoDYv9TyAs
qATjHmZKCTkiJ7peuywJmLb0cRSI3EsRaIVlrIgFtyZ0puDJ/kUpVb2ZtiSJOMyi
PrlmAUrmFVa4u6x7CRfePGz10eXTuqUmbH4DytQJBR1372u6CBuQJyXdOfQmQyxE
LA51DeALLcf5tTFtim5/BBdD7v8+C3sFLSdAQCEOrdBkje7Lj72bV9VRR3LvMxRj
1r6tRjPPJ3gEJTAbTUo8Sn39y/XvVllx+1k0syectGpoyzDmfJ72YJ6sF+DEtXS7
SS/5TQtXiIeYZoP3kinR1ZOKEVJox02Ubql6zJ/Pry8xsES8FWSwJeMyQhTjyfxR
DOQbFKaD0g9hjREEAvJf6lAv1YNXiLoTLnZfA/DFHO84IjNX3nUbiu5s9RBUThEI
ofV6pWxYepRU6zErEnzXV9iTgG48iaDe+/LiEkOScj4BYQyjpX8kuOSA6BThc4T0
VjgToR/s+tuqmRnU3yztNkmF+RCMWMaaLzfICy7RVOJw0u4UEXQlrS30h8rzye7C
Q/Q14TmEt9bmT5/QQ3RIhNIb2dDTI+bAmnzgW5kuuF5XJnP5CGcz7PzANoAWQgPa
FTxT+VtmfGbrp0Io5z+QT7a4bh12beOjgu+2G19vnddgvgf+iWP3klZ7FGENxGsp
ry3fdtp8VyflH9t7FlywObVdE2k0XjHx+bq1EJlcdbWOseuUtGLCsOPYLpIdsfbv
vyQvYHZA3daHFgzZC+BWgpXwvu5Vl6lYuV+U6gaLCle1cPrUr7DavKJ8nA6G1UCz
4LQis2Z48XlOgrL/6RNaZf85C754cx+DNx70NuH3TP33U8YryXMfMYNzqkudYBxS
sHPWi2ZwJ0isK2R3Jbl084Gb1I0xUVcwHZvyQCOan3HJ8/I7mwlxpAfnpETirl6+
EHPmixs6iyqRdeB3vejSE3hnodNjQUjOjDVvv/zzLU9gr+YE0ve5f2mX4DbzSS6M
lwgbShtfsag0vBBhf1EZAii5IGfFOlCaiXDrkVlb4SpYh+G2NIswlS2IRVAEb1BO
UiE3//e1LYPm66var9U+kQMVW4udrHX2RkCooyyc+QCxKEeBaQ/9gAyRZoXM9526
bZ/S6ctlyzK1VIvNoTJTCf00Wce8J4yFrzoNdMujqyNho4QbPheya5d7+z/CLfpQ
Hue8rl5IKRoYhyei5z8vh9Lr5AiX2jqjP52FGHq5PIYFr3XcT+cUbhNVdjzXSKg3
IRiIQzeU68Cfl2OiN6inoIWfQP3nQE/75uEoj1LtlPoBlkq6Cy/Qubcv8vaAcaHz
uFmMJpGBtlIR7ZlPCs2fbm3yCOygcdqR7fsFVgLJiZO0KB3VO9Hvr080EJEGRyhM
tDJCI8PRlnJj3K9pBu4hzvZh7/YKrbYhaKV4KZt2nvVmUXzAg/GmdmLWJrMpUU2a
wh5v0UhwmXl8zd2KImlYmGQ/I8GyAiMNOTgFKelCfD29qMMb7dfoMO41odalfaIy
heRFRswXDMiI6WgAxiGZSbV/TNW9wIwG5JHdcnIyrIO33VcSUcGEFZbO0YPVd+go
3uJCu9nfr6vsqK2Wps93qx56SlryUX+pv7t7j0Z4cHDZW5yVCeOwoq9XcSYLI54N
jD+Q0oAcgrf2W++I6Li0q04I2WuH3vVR25cj2+q6291pWWDJALmU9ZvPQCHomBuK
kMCQiJTZrdd/QuNC2/TBJPLGxjOBUl531TBiq6vCSqWHWxhahVsLxJF54HS4qCNh
N7p/8YvPTCktFGYCZ/3LKYxNoVa8isd7slDzvdaNxk5RCHh5TO213xvpwF6LlpE4
0c4ddz7DukY0uY3y01Psai59LMLjB15k7KTFyJgyV5eG9vZ6ezmP+tBTLBvlBucz
VHV9ukxIwpU6SXkxIbSWEXtcgBB+/fotSfSJIk0Y80By/575dhKFy7xH1bNL/isv
ZKN+Y2ovrd1uEs4JqajwtyqxCuu4J5LbTMFqcG9sYCxqjuqKLAL2UGhleZG4xZCg
SSdcaP8/A/y9rxI/AOLn5i199hK8vqkhtfDWqatHv4uzkQGdMXInbx65aDbIzCkt
xBvDaGNiQZLLebv1+CRofq31XKEK6T3ExNR2bziLBet39nQc0xf18KeENU6KNBlv
I4IKvwAT3RFTW2P36+nnOVUA12Sw1wVHfmjPFZT5HmbMRin1BryaNzrBv02mHJhS
zqpORokQOswhwJDaPaAucPJWUJKjBXkIdpaGMekPQ5EDFWoPfateW6t1Rv8XkomO
zFPmED7rA5h1GKrQEGLq2c7OCnK1TZ5YRuf7g9iTDHLXU7dP+/EAHLdoEdXZpCcT
JnqUuV22TBQqA+HfaUSaZj3ddD7DTOM93UokH4mS5F91glUDkYXCnAH56zFy1Rpd
wm49bcmL9OaQCWlcn6Rlfbmkldkp0F/Qq4A9QRYktEpNxzspgPxjzOmfvj3CaZ0j
viDijZwtosMOsjFwXxgIFT0hzofWZ0bUT+/c18P4K+yrSlSgNrUXYkCVc68Wkir8
r1fV5NcorRHc/pjw4eN8rjR6UnDKn5TO9bjybMKmTpnroWk1t7HdKuyOuBbiaKCg
lMY3diQyJEVyx5TShn2WLSNmX1ANChxKzD7ELeCH6qNsOboE9qb++h/B6LEAlXrM
rbMDGCpuqT4APFeKzKSMbjW4pc8yw9GG2iPoA+RNQdJqqb07znqIKmr/uif/VBvw
KRLPXd/HxEebR3vgKH8t04MngiLBW9LxVBUNd59FDRHPxKGwtDtv5pinRCRzlcf6
DhLyTgxyraBt1Rgnw1EsVbp4a9UdDD9bSY/9iT+GBbCGrMOEN3T1i3OYDcFgQjwz
3B3V5iUsrgxe8K6aFcWidRME3vHJMJgmxktHUOb7WsG41QabeKAfLEdGEmg1owIy
Hrm5bIJWWFEcjof5BJbp5IvWlWimHLWA6gdRAt+/PZxy+mkt4GFFxnWOD/n0KWFz
IpCRbA1+NkymaNOywdtxxnHIOa3RksS4/cNuJxbFV9UxUSaW3xYoJIGtyzeV3sh9
8l4p4YT2flDhyrtg1sawofxcCd4s1F9ogxIwZK0q9dlxqqSFPalDIKuLz059JrQp
8zVLk4tcio3Y8fjMGNmFCiQmGKe+ScA8G68hyD6JTdYYuMscUbaPUcp4JSWrFUTB
ei/uOJ2BOCYamb+ES/NmcCKydNgBI5IB9jo8mlmjcHoeRa8xXtRJmtw4viKiO50U
fGHcmKJr/jIdGMy2A+1q6XNIAmbqLkuD+8NtbRw0qjUyZNeVFNA9Wqcfzuy+VXQ/
VjCNhAERikmA688ds5G6anuhJ7wdRnF5d6ZXG4LX3sX7OVPvai3bRn49hi/a85nD
dTuRHeiDehvmnhfd4vlXPkNdOPh+ZCwD05+19nV8YuTcCbp4Xqul3HCbPSiaQan/
JmYQD/Dfo4tdilt7X/L4Su85X/6ikibSzzNbrPMnurYzOnmvgMGX1y1cdNfDpuSu
cFdc29XOiocEtSknmYYPHHLOe9VlIdCtFa4KGvm6Ch9hvLNdwj4xsYk+1OptvUOJ
4ohsJtRIlbiah+qGpMH0xbx5DDdEDT71ZM4brRnxxrPkgpsjYfiEGcQ0GTDdfuMN
+lhxlQ3WFerWMkaECDKZhE/TZW+9MBf1COGstRu/QcK1J+o84R5Dvj2oT3GCMovb
cGG2hkuPy3qm+RbLwZInkZN5YK7zxarVt6seFBIUpHOGxzMfMyt671QdcNGktMzD
2kYAR0guXbbPsMvuW5+Sw9qxqYJV/fFsWHuzN++RW8NGBDHQkipettQ5WPbbm1QK
s4YfZ1Utq+MeSb15ClE04uN0OZR0iA90dTcyETxpVmaXZzUXGwiKy9T1RH24UnHk
FCxC2xCrMf/Z0TUoQ1LHpydJs3RgZtvxT4SkW6iRd6oRJZWn9gKrIi0d5Y5jU/Tm
v5WwcvA825DxMIVpjP05KtQ/dV/AIdIDn6mMbpid66T8JSOQUcDgwsZFZQvca+Mn
q5EZJTXunqWiLX5ms4afUOcbWhNA756AxX5HQ4fZ/knElapRu7Jn1fRooFI4XCxe
JjTcelyVGYn5FQhzpOaE0D+R4GfsEd5D+DXWgVB3VFf+f79sIy4VM1uQn049BUtx
bVXKSjgTG4kYYO2oZLWHYZ9+eSSGQNH+NnBGFL8e1Y+Kn1yIRPL1o7NYuu3UvuSg
kbOD85Fx+KmBXYtL2G15Cto7nMRjw7ha9yjP2QuT3YxGIUH0jMK4I7SWfisYf4uK
xK3KDXfh87AvuTvvuPmpKJFk/giQf5mXgZZC6lIycybMwcX8zRThqwb7bwjyTMa8
OKyfy99TXvpBu5LGYCxObBbMRiCpCLmxAebTlGVnFF0p18HGDb48owNhBrp9Tu8y
6/aNpxQUyAl0gk/VDd505ajs86JfpHKaLN3GWr+6VA1c5GEvO10fOX6Gi9ktG0vI
13O1XnghOORoF1y4L1UwuikmLvDSC/aJldw8trHMmnTg+GKDxjwvJNm0J5tubPXM
cf+Y6cLdHuq4CcwMrit9cKjStGgXi0iQhZSkZcWtbZPMN1YYjpjAdWLV8yxgFF/F
cIvqtgBcCNmgMrdEtGKdq9+ObNdclcy6u/LT5hdilOltJ4owYxnQSjUmRwzxKmcr
BpG9yYZhE8xeuHuu9CQCRI66a3qVa//ltUu+ca0tQGlKazBr1T9J/geVNrMniX+V
N8autgsL9YmfOmRU9hHxYT4bv3Xrt+S8FADZ7hLiw3q6NhomK7cHLYGvQSyIxhZl
3L4i/LBfY1DuVwMVENu2tXd7fFXtNvEwH1PAoxqtXU8dFO3qDKsHSA5/LUu7MJkO
2+/8Bpivqalvd4gLJd6FpbohWUBM85kcuue2VpwHsSJTNEiSX0wHc/sxFzeBiepx
SV1I7nAi3fiblB2owcUZV03xUlM1DpF4XnpgNURXViUjgqPtsTpggC/q1bbmmtVa
9YPRaD/g0vfFWdlS3c6yOLSIToj4ua/c0ZH9F9immPxpNKUaXvAlecEEt5f9Fz7q
OpBTONf+rdikGsGcS/dVK4UDFR057aHcHkNbNUW4896OxxF66AT0dMOesoiUySuv
djj8etEBQzE1Rvw3bNY5XIwU1REbyCgJTFuFA/uWtyIF3DShDQEJMdFkcpVsoYs5
xTq+pXohvB5UdxTrFgACLHuXwL0w3WnvMQzQykcU46RffYSlhaLC7kBn0Ife/Moi
XWgtzT+QxvSViumX0HjxiHjQFLbdYKDHVqAVy4qnjCbMfSr2+lR+9VAjJTZQ714o
U+/8YUExSL4VuwzcOWpu5kY7JXIaOGLBuvAYjUZXreuV99lkqs79E83Hi9Vymje1
usVd9eqx2n8gyGuRD3nqB/VjUOeMhyl7SQt39gv7qx/U2qPRU0lxEg7BJoH/IP31
74lJBIhEQxk61f1Fry8dr8L72LTqQMUsPQjXf5xEvpwV2QPJhz5r6GZNogH8lWpk
jz5M4hj5T+UGHAjTaKM3Y7niAhG1Chnieic00QbBOQuSi4vIilnttYZvy22+kQJB
oYc5kwmwXSjm1X2EgekD3MZT1uetmOUrunAGcJWcSD6pagxhbZDL5H58pHJyEJ2n
B3+5eTY9BZ2ut5iDtRpiglpN/gkaztSRkARWPsoWsdR/1sB79rtTHCIBRgs7Fq27
1jQZdNEOTv9GqZdaK5SHLDRhESXE1cBPSwi5AuZjrTnTYr6+hvLi9BKERnMswhUo
DaxbuUuq3t2Xm+nBfVzmD/pKrmhdoyv0DRRJqguu2rhWEH9zb4DrGLzWzA6sumeY
BCqnuTU7oxsEDkvWqv+udJL1xgHjfS2OzE2kZs0L7JH0Ee6Dm3VWfzORjaiq3GMz
dUz5F7SiiGclmYNXcZrGhJ1Ec/vNgp5OW0OFq9PIdTWn4TNe0G6tLtPQSEmmX9pW
sJRFjD+AwX9HUy/YrlhFc54ZvHktZ52UKx4VH4zw4G3LVk8EKqrprs43pJ/RLnIp
CaX+7EKfRMo/BbHYGs4JbzriB9BphY949UHReI03VqmUpFi1cIPz0IshrZeMNCVw
3SJp83jtU6+15Iw74EEjxgyn0g4jW/GgBr+QgvT2rDEpx0Aq1n94oRXyf35tTWhN
pq27ko1Kfz8lGXmzlssXnnn1q66XUkWYD3BhQ/L06O2trcumWTBdpTGWmkIFx5BL
jJN4azcPo2DEm4pFyhpV1aj0XkJJiSEm3AVI09OCJu0P3Y24Y7EwQcygRVzciH3m
h9lJumqqYgLNOX7GaP7v9CObLe3AaW5Pi2BhCDkNji08wgD04UdrnD4SST1AuOeJ
tS0uB2G3PjkiNHMazpOB29oPp+flivLf+ysRWbXCI+IR4PHOpqclIpx+qHBvEtM1
MvBrorZXIbeEJJLLNReSu4zQ7o6kxqCvPbRt91ya+SJvulsoTZjgk327Oo+2hLZZ
BGgaArM189fvy85mQjeq2WxLJpOgT7ITvYNE6zRGu/PeeCwDDgV5kZPz53mgm03i
GDoOjYQxYNRSYmvtJfxxY0HF9pZoUCnWCZcb+u+VwSH6Td5h4VsDcW4/P8sAxWP0
cDAjcQkCW/ibQRHPPTrvSHY6GCVq+VNswGcHoEfFgTpZte2+L4sUdGhIR5WFRyc2
6MUlSjgYSeXvIraaidDMazbYrZtS8woB8VCwzteJNIE9nIejLQe6qB9CKWL25akm
2e5guQwGRVS2YLTaeOYLxETZCyn37ISAZjXYgclW3zmhUb4459hH0jmr7dlia5R9
bzJH6tyrKFrzlM8CaNvPpDpahmgxDRNJ9XeDGkIUThAWFUtWZcjslDyCyUaKW9AB
R07esH2q0QZ4nuMEXxU+95S85JuxldaIaEuCKn043BEIw2kRfjfdF0hzmV5AUnIk
Ao+Z6x729f2uFcru/B704++L8Hhka7aaPEbe8OYLWBkziTpYnLYE7rtmFvrlckSN
1+vIzXn/eI+yLlNgIK6zag8fcYj9FtEH45bR6ZAsezBvqTYvA4/vsoNDtV5UYUHT
b+lNiSEuvc79IvFMTJlFV8Ipzze5mgqtsB0TcwdxZBuJaiERjyELIQ6xdBNwPyuC
uBpeYgqQL9dZGSJLCSf0+RwpTJBlatPS+w8MKF4Gf5CnNvtRSU4rLimkugKYn8AA
dvCFdIyfNTMhZDaCymCJ74FWg5ZXDtkRD5NJETW6yss54i/sqruEI44ZK7kR9i0U
oECpItSBH17MxBwtxTwsAbQSEQqepJD600fqtE3KafJDCEm38AXP8cn4BlFeZQLD
p/ZXY/E9IYua8KotOpzPSY42WjxHmqNNTzF1EWAqxwSjCd8cLtjgUjDWkNtkFUMf
dIBxdzxouGCbsB6XujIJCJRlw2pFBW8bLR7RHULfGsfnrqXqMLubquc4HrRlDQbZ
oWcVgrbTB2T2RS3fYfuj2cAYzagh3bNrN/ju1tHWTFJNQvwhIC3vNihPLPHLBubp
4gBuWk59s/K7/WRP8xRQyGSd0wMAO7wobAPYsSBS2BjPF4Ja0rPt1ew6bllb0wUL
IGsZOFdUm4njbuV6Spye+kL8mcL9XS6IzX2hrnfuSLYChO5tp+QYt+xZgECRQtxO
RT3vKW3LBoBnViF5Th0OFAZwN1VpgiF9ZK9pAiiVwdUTtmzv2ZS+YPKx9Ti6/ii9
GI1fI+tMfykbsEL39WEP2A4EsvgT1z4pJ+tqaAyXIjNP+JpJGznZRKWlR/UZsL5V
Vx2Dzeu2L+a3HAvajvxrI6LhEgKoYU/LSDjfOoXEhEJ2JJfn6l4wwrRwStL7m9o4
HODbllqSod+QBl5XGqAn1idSs5QT6agUlKf045+tYzzY5usESogZOe2l8NR2mCBN
reoi9dHO9HaSygwGDAulJQRmYDA1KPGKQTWjKX3K/dOnMxbL0UD7QkxDE1n5mwCy
QkQtseioIQTGkjQ6XHOTmdTmgPIKFs8gWWNADLgBEAbRTLZDPzZqpoWsJPBBjVra
7HxOpFR0C2JcVwTQFk5iDVp0QAs5NVAdFt8XPHgVjHMUANH/wXAQi/lq0dssfJuF
LvHvVCJlOqrrVLmYrU12waPOynC/G6URQxojgzw7FEVI3rbusJprci3gEW7Mtphy
vecPSc4FEFlhUObwreOidQwgXIMOAsLY0PIE4fd0H46QzuDvf1ZH9MJqIFXq6g3g
JhdVkYkrTmqlS1DvGboRzkDhPu00TEuT6AoIaz81iZYe/E+FLFpfZ+RgBoS7sA6I
fDJ0lGyrj37zzn89tcOcP9PIeWdpXd4hpn3CJzcLA+/tJTYR/oUxIgm/5fDKFd3m
VeUlP18Cr9J/XA8nDev/5j7XZx/5uDD8SZ8BHTmzeJvrzYx564YUWToT22m5D5hT
QuhbXM3XOlrEDiTki9jjlAW3pzo2ss9rdR4XYrm3/2TWb+6YHcYAkDGmAQt6nfGN
lbKLV19mc8YdZP8erPI/UhAZY3o3Xn/AtcNGUz2cZWA/BzOdwJrR3EwCy+xGuB2O
KcjXNAkbTD9hMOGISN2lIK8n9dfLsDr/zQY40FMz+/sBEHNyxTXVZDB2vow+vXbC
NaixSbdaYKLqjiEdTrLA9pcwztPfZALCifcRpUmi3F1Mj6LO+8lfsNLpAx7OzQ+H
kLY7rivbL4UKbDb/HKMYeXy56VQDbY9N3CN1Y8Tk85iVCNxV0f1qDAFcRnLStJp1
Tam3jZlrjykOGoGElOKE8GytjIk3SrPqBnAaVhkJeGWZRMw0JC/jlm2ze75V0t8i
xhGbRvZcq5VhTQi3CltBa0ua0zjnPlrJ9v+Efl0y8prNSI354MdGWB14TlPzhEw0
iVk0R8LluwgyPBMQPDZaImsdBQFFczeUvjDXTOXZWb0FrsYZ2KYkoj1WxkReZ+6F
Ajg0HClqx44VFMtPcxL9k+PoDYNJcL7ssaVDGfqwpokEvLbfrgN63czuZngKfPhs
ycf02kD6yVy8Vzq1dYdf7KA1wj6hxKIz935by6m0mktaE/GyxH2JmClADSTQimN4
Mnr8sg6k2VNgEMgXjilfBxbOnevBbD7uEkZ5gWUd7dIpyvsFHoYOKkbJs/s+cVlQ
vzHjMYWROEgLwCsZH3orTrshhxiqzuPqQjfASZHeYTLg0owAvpKMoMiZw8FbvMb5
ng5Ogp1l+i38+V2IYmgADvodsCFD0QCmkAbJ9sgLw4pTf0f9LdkJR9xtk4Bv8ZJx
H3iEht5Jatb+XieEZ3ATpJ08RDTmZSJTkxIQ9li7ii7QidSOLqOWM1xZNA9xmQTb
fvCXxVlCQ522xLvYqTxm2OAzpK7S0llEfBlbsFgk8OQ4JNbVHVMxBQ1obQosSBP/
dpQlmF67vK0b1u3Nxkcu6n8b7O9PTeHlK/QGNpI3LYuW+Yj4LwWIUDhpTxRUKqCG
C28MCf2J6NA4Bj+nBLQdGKulCIgt00pg9PhQoQ2Cyey9S1OG600TkI22++dwShPP
GwDzyjdx77ui1OUIACW0aWX2w9hKRYkKOeSjVDjoStZc5ZspmmDhLSIjMhKP1hVs
XiCiXoyHH/LN2LCD14SghRg9bItTqhBT/fVHAHgF7yPGwjeBcoBmDb+XaVB8Jh81
eUvvUirjWanZ0jaViTdZyhyoLz+uKizc1n1DvSYtX8rUumpDIJ4V8t1Bo4//Zgpu
VylG7+F3bF7QsKAt4WjDy5ubJlf2ba+cFWCQSCtYrHCdEp2w1JVFfAtjj4cwgNAH
KqktToYyYFkzk4/ApHdP2UdizJQbCWQu9Z/pPdheJG/8DNOaa+gU7rSodwCb2X8y
0v+6lyFlWkpwV77eYE7sGs7EuYXVYwC6nMZs+lusDhDmmxjzzqzhdk4IRx6z9W4/
dBprh3WfANpW6omCvQktALCC64nGiIypBwKS7C5PMIu7XcgtBcdYAclpFncGV9IZ
KolDFPCPUp6dSDwoKvP1ZJcLLrkRILclmgfTooXeO/NTtRd9BREtMftqFc+ebEM5
NDk3F6IKPHcNii58mqhKJpoueUoy8IFiESi2wal33QudBHxn69gXk/yBpAvrAhMA
UX1dwqrwOvASDSfj7mlrS+2yIcccD9qhY6clLpj/m3FZ9ej1TECCdLu2E0rjbj/2
V37pEpprf3QNI4rkM4nOMgLAUBaRd+xHc1uGYtmJd7rK6NMk8Rop8lpU6yvvFIOj
kX9kzC1vob2ClXjTw2Ru6uaY3/zrJJLKQh98llgI2kxhB3z2ya0I2H9/f9zQhL/w
4SWUvUIB7KZezPM7CryUkGJSkulBPNF5QXHhZwyOyyH/gt3WrPl4DVcwEjkUlTXs
JA9CDKt0KrTPBMaHANAqDELOa70a+caoLEHbHYwOpAvdbwr454VtROiwknNM5V1X
IGZrO+hiFd8o9iCNTdjR9Pis/ufWRJGViAadkz2Bm9b165KF4E0T4n93h2PIpibv
54sd7PUA8OiaHYW/f/nT7GU3k7Mc26+dfoeiYfBmpK/p0mmnChmFmmWUiMih4rLa
h1tChBIqj8iqVL+BE/3IkPloZU/rD3LJxSPRDUEJS70dcVdNL/RqZw6wHm+QJ5yb
oDvQffrcmZyzF8mSm4CWZxtz52f464UEYBUX31/qeobnR+fb4+Cnq7oRsEQVPaoh
DxpbOTJndg6lqeJJ6VrX4Mc7jqwxEPawTVA9Zt5MS2gjRl5i/ruql151CnfnInJ8
pil+5s/hnkgoELRxR7UwLTtYvoBdvklNYfq1Xq98j1rTcNUAys8cpZotNfeHUGUV
tpemZcRV7QmrOMXi+hzvmJVHR0LM3y2gUbUIurmzJSSrICOeTVGKTQ75zxTGU6nE
AXy3NwupAfEs68+P8l10szQzQCq6Otko7pRVT4TjSqCsPGD8hrN6YgX9uynJJFtm
zKU4ltUtEhjMrvqc6lpEg01tsAGWLk79t6+jSw8Hoy0reo2Fczw7BxmV+vgjyUue
iRbSYtYHQlGSJpLfNNFVSY44h3F1bvOlWR4sLgAW77RukUfJj/K7AoE89brF+VYW
ho0CFeGDv0EzRbcKgBpsc8Nm/GmqSo16emnL8DKhh2M475sTNHKpOaZYDMX6SbWN
USuJWv1Y53u+2xPKF6xnaYK9/sOgnB7xmTbKnXndImGLTt7Yap9fbtzePUKtMgDc
ubt1akEXDBF1ljudAVswt6HNdpec8J5v57s3RXTTL8HnhqgsUVrNNuH1qWeAcpaI
I/dQSFMlitnmtxMcENNmYFwERWZMdyP5WUQRd3w9Awgut4ZZ/5pc+5WvFqcuco/b
oIQczvKlZUMWgN71BLO2D/5EB4jZ9PM195zmA7dnN/zw+PFRYJzpt/gPB4+Iba4I
04m3xvQ5MX+6KJAnFfoSglhWCm0kiTvYzKCCHyhI39Utq3QXTGWhW52qYUVgOj0W
a3EBDLHJG6XeIjUzK9zq64zRlOw5AE7p78T7GBQyKzdBUghyGk80kWjQ1YGY+6AL
EFkkMR/ns9MZoC1knBBxFr4dL7GGNXZG6aCEmijLBqb67E+L65ajm2XFr0LSidCl
FHhVvJ3O4Qm1sFM/gP6Ulz5H5yslpoSQTze8iNEbs6fUxmr8twVmReKrXwr/Nc32
XU6h/NwYbVIF7Ty6+NI+GYM3He5BR/GwLOZHj/H1smuCNfiamYduWacSkurRAy/0
cwDEC25z3fucHp1MIj3sbPdKmF9uC+gZRs/TvwE5oSs6EXWJZ93TMQsunTM7X/pF
uiqs5NnjRMhl8S+FqRQ1z20rpbJS3Myaon6lLHgQtQvEtEQtMEwkQnY/P84PqpCg
V/aILPUE5stkh4BjL5PjVg1dWNjkK+XvJqKmtsv2vo20Vv8DeQ6dFUwcjBdHl3Ls
Nk1Ik4npy00kPo15U+h20n1XdVz51mKZJLcjI01bFpH65CowMs721HAKy+11WU7R
NQGIDGODK/Qew4cxMX5Lh0P4DxgADpoS8mLvCvEKzUMJ79UXEgUZXlZpz+VPQPqh
rrZ/2UgKT4c25Uf7yoTtAmqkkqh4ahimvV2xpGnCX+Xj5rxeBRn7E9I3GjK/M968
jKqm/fnnZ2IAEV7gpPZWL5i+bg8K4g8pQ0CMrQhXB+OeW65YfnKx3bfGhS3oDxH3
J5W++hlMhjlj5vae60ZLChzv/ul2fDkTZ1DcAsZPDHWp1CBz1DTiWVY4mtAs7PTx
3+GrMr5WGx5LNsve0qnR8Hd5b22ZVNUqFvhgzLs0MsvWsK/k0qhSUVdSpR7dvtpX
Qx1htjjs55ki+ASkCLp+vVLP1NICZluD+B7qKddsJwq6kC28JHdwX3RylXkJsNi/
Cwju9PVIkyfKE7UNt1Ohl4oDyn4DVt9AMGTE3QFhzLIXcFuI5v1qqS0pgtiKDLyX
iXStvJDY/jYC0TxZ2TaEQpvmXJfqGb3Cs03QClZU9g0bqj89u1aG/eN/hDwlMikB
TyFrnww5Lk1w1erBaCIqgILMtot9weyKos4AHEYC6ePZ5unwnpAu3yD1acaGIeUo
cuoUy8XITLG+f6GjLAD4+GaI0X5tSb8jbEQ27f324gf0H7YRUspGcb813Ku/aQ0E
7uXHUe/j7rnA3WcC70LpNt0gao3loT6uFqlyZR36s7fGIQxUsh4DtNpQJt/4ZUUs
2e+EhljS8OX5+Eh9rpyYiAJe+pEccH3OT5+uLMJ+suMQUhM2zmSp4d1bwq3K99He
f/oiB8+3BYeaq6MuhaAaTZWoVb0Cw3HxpNzwqkzJFdPiSC3pWtJAm8q3/YZ0qKdq
5XpfJ4C4vBwWLPpQlj1Xb8v8j9nzcXHq7+5DWZW2PoGptfXQYQzUsu9xX1zclGBM
+uxtofzCPpezZin17sH8Z/z7hq5oSaUvYGIyUjqk6kUwLHtDVglc3wEWaqy43jna
7pmfYI8hpW+if/YSlAvbdpvIIxLdJ8JHK4r0UoC6+ARn8BO5faTiXuVsZFcEVr73
bFkko0vLM3AVjFMW86Mytou2QJI61oMsHZ7FB+Z7HER5f4AO4fPlYtPqGub8LWYy
CjkGJhOc8s11QougzP1NqqEp1jCDrBF54lV3o4U8Dy7pJhScKS1fypMHjo7DxPVO
Gyu+NQgzzd6Lfo91v/aF3d6rO9JSkhrQGn7y+pK7vbyG033b6rmLg9iYpJzbuBlp
pAF6d4s0DGoM61xTM9CwByTRPq0JcM7A7ZiZOsn5QjRd/UGYLFseaUVJt+B8u1aE
VCkIvV0yDkaW4EJJNHcFtXIHz2yOMOt8iU9QnJzEEEZyTsKEy34rHTdD5lf+7Wef
xO9x2DXZMjWPVS9s550ZNgApKsNc0P08RiJ7Sgw2MsZzNAPk01Tye80zOZnJ+Mt8
KTUqXmquGD6FM5AZ91R4wGLrK8Ff36JhiibYdIg04q3X1OE5VYpGSag335t6BwV2
WOdHhcKZiSl4lG4tyI95hVQoVb1pXXGCSKmAyKkiKpklN81LaqoiYdH/Ixm89S7Z
zateXWhjix30006ycSMbIWDuOL/Xp092jKvfFkEHv+nq3YFFF2aGkjDYuJSM7mcY
4GLhroeGo+o98YBalOey3e4XdjeZUStfehAmkUhdOO9E3ZCqBSLYV8Oa4QY6+gYr
ubCicO9JT3GRekqRlYmS7OmT96seRJLir+Qk7qoAyRypDeDrHKQ15dotb9cC/XTs
2Xqewc9znNZ5SNBOyPgQ2wkFVGFY3jdIRtu1NWBohtPleKjEY0IMDlBfolqwfDgN
ly4Qr80xuDdMIUenQKkVIe0Q3vJQYg5hpir8gxkPoCeEIMMjZtyIQRdO6ude5G2Z
8mQVVQN/Qffsvdxjv1qf+2PqxYo8RitgnH3fsibXQelLG5nLqkuVIm1lEjitlrGG
GLI2dOgTYa7nVsL1Jiw9JS1zQ1q59vf8A2XBpojqh5mGcCMYLXmws9pon7XxtJn5
zSw2DY1pJVvR71VYab3TuKQvOYtQr35PPebt/E781Cbww8ZI++i8MGult9A3HyU+
awyRKoJ8OQ3h/318ukIqloU+XguQhDgfU6ho0tfU1Ar5VCErgkk1OVItmckFAO9w
DjH3sR/Vn/s3GVf+414ikTxb3ROVEqGmLIBvYhC/zR1Hk3g6gVajwyTNHjlAKbuv
K7xphcSJxN6rHag3gKyHQAbMuyJEEhWAM97tPKrJ/O/M3EJB0VEFw1g4gfxldzqA
qEOSTXoHTw3H1vW+LTsaVMeIJTDtRJVpqs8mIRyTLFwm2kvUYAObxzkAMjxcWfc4
p2b7XDDgr0wwXLkljTRsYI8EMgJANMo8UEW+MIn1F53+4ic3Z81EdmIdCiZCH/kf
TzWBrsNcedL7mc8UU/2LAKA+orTvoIy7TgAbhT77oNgXbalHhlQ0N7MFwG6lMX7k
Ryu7VnlIctE9fx8cbwHDCnjs/QkFRbrM4eo7XfKxPpPX7sVHX8i3mVNGvpirlWVt
TIbZW4QM5pNRVv2RpdpSVXeYyeJY7mTA6uWqOHIQN6LWpueSWweSwx1AUXyHogxN
otdtVvcERYgpfxu9FpSOnSqrQVKt5L/4HE2es7RxFzpJBJriYLh2H/MCKIbL3aqG
In3vfDAPxjZrw04IoKUt5pZF+GVj7UgM4sqQ+7aZ0bM+ZAqi8DaMw6pX4hR1cSgF
rigIF0HNXacc7FguJKtli5zlIN0uzaUv+FgQ7EhQ4GyiQ6LeX1gzLx1l5RpdYkXM
qiEsto1xdaT5jfHNzyC4UY5E9XqW+wrAsGAYMeHrJJThugjfNQZc51s0HRJjvTOm
B8ke1HZE/dNZV9UnN0ODv3DqoZsHcJ6DMDFmYYKqHnlGktMdJzgGqxRNZYZhO0w+
gBpdsNDjwIkGR9ds/FcBRzq8K4LtMdPWvlpY8wGZGn82ZwuK4/VPAxxshBXraBNs
2nhRklAbrtA0soXXRxyrxUXsgLsCxzhU9CA2JErcqYhZgc19mmBOOOgu7ll9AUrj
v85aR2sQ62zHpYrgJtNkbV2ZGUG1jc+kkb4IfOxA0EnBTceLMCvS9CsBDAVW1DOI
kS8ISHS+IXabfGwjqjn1cSPYc26Ucgoq0iQaEubrLoAoCI4MFU5oZ9jB7eym7bQO
05UArEb8Zok1Mas9ykwexGSoDNTv5V9E4ur9Yy/p1eF3oRqnF35j/WtdUuu7mfbJ
lZ3QtJ+JVYKHZxdseYKJM9W0t0hf3LygvlJVPM2FjecAmtFh58o0BGq2dei7XHKe
iDB6KaSyIPDvYEEq7tUUY+vnlogwLun+WBP2z0QXAz2ps2kX3VESQ6UJugC/dfT4
60hUhXzwr20H5Ci4OnSOSdccFeRZcbKMa4Mq69w5DQlQTpNqAi6lU3JT8Y+FHdai
YiXyq2DfSXTgt3CxWdPB+Da87ssxdQdZQKQvwjEhtp8O8HtVyilnCY4osRz8/ewN
HxC1632w1YXAz4wsGlPLITLINWKAJXNrYsft9H/YHZ9K/FpuftoEtcZtkWaqhPe5
n+NfdByvk8/AP28jkwttu+SI7ljOA2Cu4GSFdp7ju73hmvrHAGD+JyG2lpgfavWL
eFsHBnDqKzMMskpZu6+iHVQ5M4zEAS7ccM1ErfYdJEzP9r2J2WMSqpngXreAAzQ7
QmNX8Ya6KlUnlRF6KKhmZTwQq2JxCpNRP3xbs/KmJ4VHO2eTtBTBuZNaErpgt9Ns
Ut3eGCRmcuvqDok2Wz4BUPjpCJNuGDia4+ErCpL+lSKAq2dOMQQkTQvATuZkXZkn
+JWDhNUn/HoIUPN7q7Xngtm2NWniq4V7kYA0a4OiYPgwZy8eJ9MY0iMmpJ5xNNMW
SX4bUNDoeTQXYlwYQ03nIxhFAvkWwtKfUADHD3DtHOjuvNOGniT0GBiZQjraJKH2
PZI0zXQOTCF7iz6xBaqX990hmjWmBChJOx6OD4Ciwx0nOV7pnsHHJnWiAX/qQZAj
GDwyA4LJZ5qRqWl9j1SQi4bb43U9yhc0NiMd2+/Uacw1IwD9moTyd7bdon/3Km60
eNLOrEzBmQM/Wpxz1/10zU9GGNAbmShx/mazzvRH0NYZET0CIqUBd/nihLITl4kU
Qburiy3fyYGAT0Y2EqCBm//EUaLqDGZiRmDVkaw3Kcpze+GVSRbjlXCoqV81y/P8
Z7kOxvixkygBV1I4WEo7o/rxyPyMgYkl0KgfrfG0YxKcr6Lju4k5yRwEE9KgSMc6
ILvA24PSlwu8eu35WjUkVkxeKUReYpDUiWB4VWh5FEpVm4KS3HiO3mFX8Uc8irVd
wpSuLH2g40GRSWmJ0WCHfdJiywXwbqZFHtHtFYv++67yE7t/bHsFWULypwbA0jxO
gpTO4JGIRsCW/2QBzwls4PIa7kUrhzQghiLwU8KfFg9xlIFEdafm95u/LuIplpHh
PmIMsq+WN9k+6SHq9jmoJrMgQGZwgw1Pb1ABu0OqMfbJbHfg8alCOjHGQsdoNK9q
7Y9wHLYAzzDtHDV6NBJYQDWadjkhnGLHwJpUFisxgErlDsI6MOvZDSoTApu6AoCy
N+fTSAjLwJgwzhdOCwhsZDpLMa/DWk8ltII/+vp5L7LjgjgVerzgPlrTXfooAwjR
GFlkFH9dEvHRwgCVx116v0riZq5eAH6hnxIkS1tFXiIgvuP2yYVZnlcrkeu7Ug7t
g90fjWCqoP+d+m6+oubYWpYDMszGwmfsUnAT/Qr+Q47GZ6mdmV+a1NpkBFCKojJ2
4CSybCpOPQCsWhZIGa4CHMyFUmqICexicOApDsYLX0c37XumFnTHD/JWXVMccw0L
r/s6XKVnkjtHIUlU8JaNUF2lpL6F2JXViHfwAaGOQfVmB7XVKUh9mYssaNs7oi3v
nYS76bn7TihdNm5yGB2vVPRMVmgYJX7A6Hd9MWRHKcp2QMynncNVUoy7fZblN4GX
IhbRmdNXPYCdW/AuiYCoGjIW73uHpi1OYExqnlg79EOGS3olecKXZYLCrMYraIGi
jkRgISzLIWU++wbFR/+PqiK4qcDk5qjWq7rtRz3N6TZR/jy3GVlWiyGdIZ8K76W5
43oorf2vzy5+Z2cYTvt0lEsx3oDsg+e4v72LOxBZBtDkh058ZHdPhB2Gw0NifyRU
2fCOx0TRyFHTwR0K9u9sea1hgnwpZmPESQhS2SYtuO+Gq1Zsz1VaUsvI5Py7bXCp
VNgUDbWeXXANIgZWGWTc6GsitLQhI2p5iesThkHz3yGt0ZEcRFU7uJP5L7eyjqUB
yde3lIGdLXcW/YDEJiaxONexyMmmoqTcveCsmdnySJFw2wjjOOJTMdAFJDPkTFAH
8RygYT0U8pVLvYUimS6ZO3URcNyc6yRhyBLMimJK08sCV4IDxVwy1+dEFhaITY49
NFNgZfcigEB54uuaGq+NPRHRRiOY887Nt/jjKy2lCoXqBvWgaORs/aIAGOyG7dNY
212yPu7DmEA0YK1Gvc6ChvRncD7KLSXjl8xj5ZhI+68S+T3qHPGYpcmfFP59WBn4
YjFBxX96lWJPK1Uyya5C2tdLcTSeGN0u7a3aLivTgSckiNOOurJa8amqMBkCZ2Wd
kKCtgoEhK3rT7YRH724tZPeD+TDg2Ge1L6zWd9AZ288le9N0kX55ZQQFSrLwfDYs
bwXq93+8tQhqUvW8as9oFNip3BmeBjzLPl6BbD9tbt76Eco2+sLOZeh9Jqw/X5mI
Ded34Z65r/r08EJ0uQVpiy//HPfn+iv3YkEU92smOvCAFze7E1qT36KR+e12aZ9j
xwrVwijgwZQI0IF9cdcJW2fKP5NW/HevrYcqLL7TseitWuF8QDOR4/yvloeWHqyY
SsBowQHo+toxt5HJV0cvQ5Tr/lbsoH8f0+a26v8CzmzBOTjcrk5CSovaphsvluLZ
x2mraPzGFME3XOubmPziSw0lFGBCX10QKGDP5hZp+9SxJySE9CQxO4+cNuCQqjsT
ftoQQ9WvKsm2nWXqn88fl4CkkKMmdt5lDO2v/sTl8dDT+z5hyuCDqwJMMSiIreC/
9vidn4orQQZ3BzQnrfrpT53P5rG2krguepXcwYqdUTpUJ0gWjB/onK9M1DrqM8xZ
i4S2DDrpd5K/W5jmp5x4ccQv2LU8n6oC6h8sg1RdU6YAG52YmszJUy/tkqkzywoF
9ezLUSW7cAC1Ft0DDHB6rG2l4/WjzfmfYGfYtoHcLMKT9RHfqJ5jQAaM413RXczE
qABCVseDZqIqla/h6SRLjKLcacoJ8sJndvfIfBd1wEWd07mE2b0OXQNuNrZyCXVs
ZLV543SXWK8wvU3Sja8O71THVFl3BpS54VII6HxGaCBKtbS/j5kmqx5hO2fBLkU+
dXyjr3zayHiF3FcRkWDJMqPZ5XfyjiC4IAFPPg4f6KWWIv+pIHvrR9G8tb+S1YPG
KhzO9QGwRQt94gs0s4b4w9oRdFoybWxGCG3j6D29sd8kcCtcJkSxVx8nIuJwc4LA
26aeFhiR62549nVHPGCwoH8l61VnELCAWZAVjezB3qTNwPfP1plqXFmbkPk8xaI/
JeBxwFClbPlwbtTjD2yItx9MPdH8BP2O2VBXOTYkIPfXAfMu0NEUiYMRvXt1vk0K
pTLlNNTH8zX4GpW3tEwaJu8E5wICnKBAR1xEUf4A+oG1aZfjOoZehKPcLRvCQcXM
/5yVU5v4JhNK39koE7zkWSMqXUPEOR3ihztV2TQ4vXQRQLepr9Gaa0MtgT2Hf523
Q1pFyuOusmJApoB4KjWFKUlvyKcxwciz+2yRjl/SAJ4IUg0lMxKc86mLVFFyTSVC
8uPqX166w83M0s63tKosjpzoR1j3m3EJ+LRhFL4iNxDRVOA/zeA2gKI8n8Jm5lD0
/tkGMXD7SQInfFlKfWm+IRc/7cTJw4IV6B6V8DVvNRpxpxBHH9Ra2N15LMupY8ox
9dcNmerIGehsdxF4AEYd1UdujgQDDHAKCsY7tSwn5y1Arz1hc0F2nXoT7ktkCJk7
h5TgHn5xwztlkPjKNT4vZvfwUlzuOftg4QVTjJ3QdH+byL5UHG6FUauNsoJrvWr1
cpsEruZymsewJAGQQc28kAxFEL7jOc86GSJHYJKtkbOTpdc6nqc9KREWIZuXGnN4
91Zc9mNp/E+D7siqixfAHNiclKm3C4Man4lvlIc4QjFUpb00A3lBdP/BJoU4CMdd
fT94wAZgGOWeLIPmi16YyTrLGFEuGRBdviJ7uy6kg47qr/wCxWMWqx5+xZRpJhue
8I/+Gxxrm3OYG5DqLqEpY3QAJxXr5NqwK92oUZ5Jw9Op5/ZU69hzGu6Nlsl01tEt
d0A2C8K1aSlAPGULtP9TbSGbsGniXq6wHt9sBOTIjny71gZYe+SnnJhYgr/LdbsG
hPLFSCR9GgXml1oYNsu4Ie2o/1vzggIKQIrZmAtEvgkCD7dq6044Nj6aQ3Orwnfv
ZI/+DpsuUBtlMcOmg6G2/dsLr/d/oQgAx5TxYYz5Mi8/1XQYAcIigLgtWr8qKHXW
y9JBJCi977gY8aa1MFHLm8k512tNAkykH25C8tPvXLD8P98FxWTHo8fWS/wywORn
5OvoKr6zv/JETwTrDXE/SRn8UJof8W5Q75A/M60558ZpnpTPbg5Lr6mfdlMZpQ+Q
j7IPuq4jfYVFafeLb8Xjc3gJRoADkkozX41WnvjXsWDQohSG5F9O/H6aZJgkyiMj
iRxIPhe//DYAwFL+Ed6XVFM9kev4WhFUyf2e3+zaAVRz7By+nKPBuYlZPUhJI8Vc
pwl/8mQAlkv1KaU9PB+83iLlnkcqMUZK6N/lvKVnldQdzkjNp7afpYoWOcWeZy6a
bykfNpQnfYwqO4tCgEyi15Rs3nCffZVO6Moc4FhnU+mUoXoSRF/GQ+WhCe+l7Lh3
plOCGaDTfwSiimC8RUhX5oWRHKRTiJjhNiUxcYucXealQJvep/wnSOHZoln2FzD7
lpKJ1Hz6OCx+hr+JZoza6MDnCBNwpo9WLpDHRbh4DkVCRUyF/CweOZUcMT7/4Rkj
E9JXSKDiZue8Eqd1ubsjvN3jf2wc9kuD3r2jj5o1m8BDaqdkOKg9W4NmNOalzz3X
8mdJbukd0/GM+LxQ4bVGsXH+fC9+L4RFszmBHUwYHHgWoLqFY1RhvvvlReV+BVla
fOahHftV50eNjjHR+NME14iH5k1VPwEpe9egaIBZ3l2u1pUE0JUlEiOYX8+n1GQU
U0AORjbW4a88E/JOvhvqwP509XDG1dCFjag7Dk7rZLusfeA+tTXnNqxU4TCpHpVf
Dv3HEEqQnqdU5Xb43gnZouIDXuS972mlGL9Faf5sp/nkSl/kvQU3yuBj9ThDFTTr
aisquIkYMGDdjyTHZEliNgwW5mQX38lTcBlJRSY+SmoSzd5eRAsR/EnYXG+MyPXX
OKS8bmYXbA/fcr7UpDNtLgq6zR4tlAkNwT3kttWjuPHWmgvn7u8oJxRSW0LoLn6w
bQY928KWzmY8Ihj3wAIJKqaVG7i5ewum4PDh+jPFaOKoVeP9ocxSq9LJk8RJ/Oe8
NXCwh7ZCnrkk3gT8t8exK8Wurk+Lji29Nymcqv6u0MaLv7WD9pG56MNnhprc/Ud9
0gJWa1rBM2RFTI/jxRLTmoyY9uKeWVv0c/21JogUrIl66YiHrI8PYXWQpcacU878
MzHfpxsKJ+z6fO44WVQGf0gK021R4SDO2NZHnyPzdMQrRwSV9f8psH9eYwAp4SWq
95NGKnmEk0QjYSbSfP0cls+7HFShe8IMkCeCoAjw0uCGUTxfH4Bu0XmvWZ1exNpf
tJYSSce1riqWeKkV1kp0YqenWcNaqDO/cCTqg43n6eSG2bkHuJ94Z+NQPbbhsw30
ACw1E4EGZBXjtLD3N0D+iAkLlMlipNmTb2eD+CAVReB2D82B3AKaMzqvw8N6Xftg
JtNcZyofUTVaAb5EYsc63r1aG6UtEf2iozOj7uX2inE2pM9GiA3wAPkVU5uFs6Pk
TerUWftcSDSLcmyZYXXiYlWOWGVSi4QLZbDjsQBETsCaWkqRpllfKHUgXoN5Eq53
tz74LYEWikBGmG+fTNaQaq2t3cwP50ubBKHj2d+K5SOSZrIka2svzkviuCUzhTy/
rYSMdrRrWcUQ93dTDlgNNVP1utQiAs+vbaQ7kX8hq/qs0W/Rs634LqnmY0OE9+xx
pJjvEH49OarO20cmsTKS1McFDlFiK9EfKKNHj3aMc8Vnpgci7vwzWMCAAhX/QxBI
33rwGAMEv/mz2/Qujpxcpk2RafDZPuunPp9iVVaFjlZnv11w9+YQOrIm5K3V+0O/
Sd1c2ZfBnsxcZZLsIcgi1Byviqmoa5C/sKCW51RoQrbT6BO9tTZd86Ay08jsnok3
EMDyil9jCuXQ2m20P6OiEaIpnsAVOHqT56AWTilaGKrRooNqjQM0qIk/A8qtRLzP
Qd7vGEThTPv9y6kAPCqTz6fs9RP+T6rX6Xmp64Wijl4WseHj8fYclv1DyKN4L3aA
CH4oliOmg7cSFjCuRU1vbEYQTa1k676B6GOuf48hCgllD5u/WVFiwklzAcaQYxpu
xzL6172C4JOPFKCIny51R3SiIbPNTSnsb6Ag25kAMFvrCTrLfBWzcZ8kpiWW/+ec
VoswXPgOp5qk+ytnwDN2hIHEc1xXnhTFTfm6DQ5O+jGVp/CpL4hr3UCvj0WzvSxb
p75Mk3DMLNt7jAWiVp5F8hLk87Jlv4iG+mhX6+AlARN6BhoD8dE9PBNjXPitwCzG
D/WgrrksDVMO7pnwhKmEdWvtzzNp5DWsRBas45XMfEVo8EuUGf2JyzHGdytIucsJ
V7NgMy049Ez5Kyl26Zvenxo/OZHlsacXL05qpsVsTHErpjMsraSkPMU2Ra+qjseF
CeKmZZ3hqxMqiBe2R3Ws55sb8on1yNhRi43TqCu4kC5urfSCxI4ekZVSUIbs9Umc
aT5E6khyef6dPCAVFc9tTepJuQKq5YkzZNnvS0POENw31JhgupB3W7Ycnjnyg6Ha
QXaA+bE/qE4ASd2WZ8IXex/bNbM49TtYwDAoOvPkV7PGVxrap9gg2uvEhT3/VXQ3
FFZzShCDABshnW0qbVu3JUnaEgMWT3uK1EXJXuQT+9bdXK1wrnkSQ4D58f53jB/M
hnm7BsZK9o0/NOmypBXmJH0DgYpO00zkyDIoXpZ5wNCRQ5wmLcotF3Mgla/8XOTJ
IoryOVV6Z466uTZmQP0MygoA78hFWrrZPOVg09fJSfZkCJwmiD2Py1FjVBR/LkNF
rz8FBH6+K1kWebuyUczrhSZTUsQdel8JsCZDRli5uzDcPEG6rVjYM9A6RU46WD7h
pie/0LFcRno4LBldQb2ivNCFoCGiZfaPimzOgazrbHVD0Sj9+oAGz18lj+bBFAj2
eByEZmkiMpKDE68DYw7MKfO9xrXmfj1mX9hLLUBg0GGSk/xQzHg6zfw9UiJCrQZs
5j09DUG4ZRTaordB2JbU5UUeM3cmQkj8+0+B8r4LqTr0zd6wAEWVkWfxUwrjH/Rf
wOT02QRDICX+JviFmTC4hoUDBHNBo+jBxQVF04mTyunpB2Ihp9cV9i2+DUmwoNzC
UXt+f4VkBBF1V23Hr2Cwq1dZxdfNYhI1f8xjLHzfMHklo4Z18HsaC+zdLAdaZ7Dx
eOvzFdA4CZ4aqsnRMKLgfO00/edx7bIfhsv+utEjKzUAGB09YyjBSqoJz+OIuPho
peLMgZrLN7sBuzgdrv42kE4XqvfglHcSF4MeoHfCoGH7Imi5QItu1TB1ExlvRD/C
mE4SOrrWzMQJpcztPZp6gBrIru0I9AjpLysA1m3gzH3E0sq/AkK/YV9/fXFWUvz6
GXhCHRLp0vvmA06gkjvgGm4b5B9nMM12414GyfyR9LDnHb4DJJdx6Mx+wixuWQtV
LocF1B1LneOcvDN67GS+tttk5oiBlxXYPHNQtWp04ZLzU+tV6dWG28OrPe6tHRE6
DprxU/hGQzfKu6L1vL/j/RNrkGswrW7e66nKSy1fDp48zm6QfLrAKTWLidXRcrxr
0Z9fFZILKXFoMeEmzoLX+3LEa9Z0ltNmWbsOQs5dxecgA0PQ+C6u/BDLwIS8vLCE
XGby3Eh8ES4djcO/VBXlp3ltMkt4DgIH5vgoQIyUhQvoTXoruQVae8qLB0LirFuG
XYurV4wazjNm0CvL59zsu2ip5in4cPayf2gfLm/F+BVLpRX7SccyBeNnAfkYPVZy
X6QBWXlrm89p2vvkftS6G+E2TuQR1EpKLkTT/4TxuVQVTv8JK0Z+V9LCO7UxuVH1
7DFP0THA/5FrvD2eq+5Z5mWMyRSv0M8rY8waQYqTKRJKFQ4FcSDAQn8VZ9dCGWCp
JupdAj50WcH7GCdPwK0qNLgKOKWT7p8kH3Y5o7OGPIg21LVSP+srcM/Q7wRjw8GT
2wi6iWG7212MdAleSS/m8jzxjG41iBxHXakm8UjTN1OGFu4jjt8ERw59nI7R8r7C
DomvnCRJcCr2SygLvQ5Cf3zT3oGiyySUYc0Orp3YKCqfnUHFGeot0ngnEyZJbKqn
QuyffMDks1WiRG0y47cIyhL/mYDdgiR3LJiJEs4TCR16hHXO5IqrNsBSBFy/Xy3O
C7JjY+DB6QwrGwmZEZR2Aa1mQV+eawURxidfhxPEGV0CFKR8NOcYpFk8BHKLH7I/
O/Ed9azByGIuSd8Ft/8Z2W7oTMaaqOB1l4sTsfb7BoZ9dVqHILHm1xYmVsdQXRmQ
qxSeKt8ahCaAepmHUZJ+I6hmuoaLk1K/YPAUYHAGJzVnUXHKruFrqJZ/qA1bvV6j
V2NTRWUkjU29UnAO1zNjrgpNmBtAVAP10LnPSW54HPbritMH2B5ugwf3zXYawSaJ
Lw5ZIProtruf6JU8q391GQh8imzIGbKwmWWA1oE+aDzp7j6VYpFOrKv/uEbgMnTl
FXTo5M/MlV3DNuRQQYrMHMMYyrdR3sRqAfZ0iGD3BMAvzEkwu0iCEmQe0jL7KlHZ
HC5m5FdhF+LEVDN+TvE4qxSTp0t2/GG1Tbzt/aaNxYQ5f3lxLG907xKGNis8je41
VKY22ahpN5rseRs39riI/VTbkufEKBoqz0oycgAXqlBXU5b8S3p/5wrAtS1WkFDy
mXoFM9ANJU9C2R/t/2mYbw9l+dDNRwU25CdmLCEy+1G4Tdo23zo5A9Ng2tFZTtZB
EiBmJfhgzw5sakA/S7EHPwyot7yRVmeJ9u/d8jNHXeTOqQur5u7zUa1QrtEOBSdz
KuOoW4xHYs4IjqGhUM4l9jXlKbuxTvnjFyjIENlgGAAsuar+lS0EbF2BiYDQ5YVz
UxGB6oaLMmThkrM8Vdamq9gu7YSqRJJ3QOqygjqFHs5hH9sQ3d2xztKYaH/ymBw5
zZrSivH0UlR7R/1xFbxpQjXzQ/1sblT44cf4IwZjb8rzrUtabF2KCxO9GN9jVOIq
3gJrBn+5sPvCYkClWWGZDJm5vKA97q6ooTfBdK0Tw/UPIRGDIod0ZwGJVqg/DkS2
xb1+Tl87zkoNJwEilKA8zuqglbFCLfom2PImArNnkEhaXcj8bP+ONItxVT7Dj83v
aWMvYYoYvXrFip8DO0bEhcEbSyPHLxPfg+UmLb+Goz3/mQTIcO4B07k/PgaCFcWv
7IInKD9i83H6K/OwnM2sZ1cKkKk1CnQqxN0BabrC3aNPyGpHbr+6sx8HsSKs0yVg
yR7OM20xnUPRp2j9hCJzvxErrlqw8KH4LdqApR3rqGw3ojAbFuFcuUJkkyXwkKyp
v7Aes2BCqt/VdGjgDPtA/1Ovv/ioVuWWXvwGOai3ptYGrGUlJRwUIobxttCaeLRm
4G6zeKA4T4xajRNbpP7yuwzhcGX+yKmLPlZqVoHvQhJauOHVjOyEwbqvsa1xDYer
pPMuAiq5cYKVHqw5xyUp43dbg7QRWq8jW3TYnr4TmdzdZS/K+oFmvN5Oe1T4iYXh
OftyFgPkpUqfsZDUP6/qT8O/03g1TRiLiQNl7XMbyTwq8OP+slXvQkcgN7QSr/oK
nomRf24fNaEYw+zHlW2h7VY/pZZ/vvbIvyDooeWxOSIoUF1bI4/k+R7yAVutBF/K
bSgzZyZnoIPo3akPxeZ5PQVI/OP7fy0p28WnALzLwE5wJrBrrkubjoXx6eFrFtu1
c3+Vws4do/27jKdypPfApHNAsCv4wgIr9Y8Qw5zpeu3WSxefW5rfvGK18FnFY0YY
ukaYnAPY6pjK9aRRMf1QyW5GJvHA13jlkSAg9GBb09gd4wNxlWu2V/xmWD28KGt1
A1jZZznIGguIjUbGO8ZwqSln6aqyrQ+IrHM51B1MOonaVJnLngp/kcPwNd6rS5JJ
rN6M5byx7WloLmkE+B2ouEOnyItex1b1l6+dXTK+ZgPL8U4pliEDlew6i2i9dsVA
bS3kYqHJT1zlgllwHDmr19Pu/Pr9WvmI9B3kG6x0KBc1Kpk2FFkt7HnujCS1RPTk
oZ7IDhcyfCBfGyOryvOOqGqN82+Favdv5ZsSypA5HP/GmGJksvnUwc1TWJbdu9yu
uYXMH/fc1ZWJgznNbD+JMx5NZBHYvHk0xAQJLBY7bXEckF/spDlG6EE/mtNLci76
8FroWbU1cWSnib+nIj3NTAACKnAn7Zp0O3i/YA5+3f3oV5dziS2IKwxmbHIfTRH7
IckFR0WaCEB8jl/3Vg/aIRHAn5C8aYu6Bz0V086N/+9/vhrViYmI7rerESX2+Uyy
4PJLvbtc1PHAixZLc1GlSEfixHYFvR5cr1BI87umoOV+EXW8dKFv75yEl7dnB38A
TGdL1ZEQQhtkkCAqBTdfNtqbJcTm24vCp6QnSIh7nbJ28eKoBpFGWCBTuz0eoL45
Ex+LLJm51IqvClxNHfWaaBsJGFUehbqMYO39OaEsIy42kQxy/ViKw8YcE6/TCD4E
BjLbQTMIDkoJH1zCKCElhnYKKQbAIx9DafudfvOSfESXN/8zasxcslLaSaqR28vk
HxLwBbwXumghV+jB8aZeBfpWmQfLosqpVb8Pcb97/fa8kAr6fMstWWyekES6d8i2
2ayKxxKY0WN4Nu7x36GOMf5JegRtd5Bv7gdPyEAqgomOUk9o3ArtrIvBs1lAC+ZP
RZp8f13D6hD68sM9eW4RKoul1wxUgDOuaUYuWb3Ti4eM/3kI+WrOb6qaiaBKYlah
qlXxh+awsGgy6XpxKv+rNLaa+/TXrcV3oSA+LilZvjLzt6+7ooVyHmc8t5yU4h+M
XPK9WeC7CdwJj/MZ86EbGs+2aqb8wJpiLJwUFyEdpoPfVpgSex4u6K46w+Qo/kv9
mMESi5q2uI5moFXkCZMLdsKwWzQYFBDTHSFA0XP5xeQTYyNPKUIULpWBQp53vSMM
FkBzY+ZKgNwY6Q/ldVIClsc3uXPQcwAyn4XlAzjNArIt0DfUXsJi6oUWXdKaGECI
5QrNT+nK94F/Vslyx/QlFIgkhHJRUFNNVp7DnXmIdtdiMAVhc1ExM9FgGRViXcJm
rRX1AV6iPbWaMsuLf/gfhZasH28JXOZ7xvu/F3JgUc5nyrNp4uWxlPM5YJKkZnqx
AezHpR4j8g++2/Soikbawe6tHRbc4Haqal0mBEDtoZqBIwZaS2CdskniMhSQDmR/
cboJ75yWOvKMc2bCoZx1ypE1mZupoO9ieoKmcf55mrPpRb87Vg15IQq6WPbK/Ndb
oJNsMP086kuGhFkPD4/2It/8uoM6hiP6/typc8cyxvelsqK5JvVAHrNPKqS+lHKy
XEUdUHV6B3WVJh1w6AzxH/STYb+yYPwu77N2nmIWpwZo2e3OhglcNnDqhG2OJtlG
x1OU41wtUdHx4hmjmEsgn7BLegW9q62/JxDJY9ZqCqDCQIPqo9FcQjSANlOPVo8U
kkrU6MBZ1yHtL/aEqFaOBicslNA/zitr0knLxt8ORJDyk0ckcVDeI4YqwLyLzeEp
JA1JfoDr4qbeStcXGLVbAW6dCw/gSoB7P8+WyjKYVeGByQj6V/x4C9RPk49Ksxvy
iItj4Rh9txwqM1yTFiTo5WrY9G78baYjdpwq3/nHh1uB6Kc3MKbd3JBWh13ApvAA
KJpZAcRtrcFkfuk52PT6+88L8yVeuKseOQZfYQDPIRRRPSfStcqWzom1PZP4QyEs
95Ili1t3sbS20iiK1vbnCB1ty8yn/CNl06dwh2b62lpRti97UlFou5uGbcfIKRvl
L1SHroakgDXr0QmclCXdt0xqmxl4UfBaoUlcORSXhPINgLE2YNDETSYlYZ75xMNR
YxOngYWCOxFtmP0i0WXXDMwY0h6YPGhGX9jx2kU6wY9eALH45LG/EcLwFNvV36VM
eK/vmgCyGJ7O9o3NadO4rRDjH5q0tDEssKzD2SXeF4ilmNNnNqFYAI+XGyd6O4W9
CbIuy6ZAB4aKAUx7KFn6MHeNK7Z4uY7yGNfoD104qVMWEAH/IFdCXy/ef3sRUbyB
28g1A3wSu3fv88n3MC0ZpXnDQzm7zPfxpryr94UPG8vAqUUrGMsPw2N2PlIBe440
XDJgAzwxyB0pNZqrJXM90NWXFyGE3RXQ2/fN2izXNirB+2eE9XrNltu0TkTcFMgs
B1FUY0hd1cwu/V7uu2VaS+gVey9a+9b+0RziiZCh4QjfINX9+RJ3zsSqP64yN8mR
33Vq5IgdRKWUwpn5I0E4YxNGwZUYrXwXTW/tLPKz2K5sgSP30EzpewR46Ob1lOhG
2hyBbG++vNIQ5SXJwcuM95jvPRKqSJpht3vbPvJvtzwy43O1zBdGunXFKDxprJb5
Wj6418mJCd0RY29JrKT57r3nE0BflyVZcsevj8cEw8XGgIEfGGrps7cJkIUvH3LG
8DGZBF08W3j6k9d0vKPiSxO4C4GHf2CATJj8g9EjZHSNCqQ0KpgjMgmlmL74ty5G
izZbHBS64XpY7UMmu4qJeSoJ8dodZmM/1XqmyJOtQ/gFt96JDK6fo5DROXdSHhLr
w7B+xGytBg+h6DRRDo5B8YT65EMRyBna8mtgq9kngaw0wUzqVXU+Hz80B5lWxLyZ
ceRGLJgmpinCcjfHHh7eQPhZ+UQui6+sT6H4985TvM3NPWMl9byLo0qYr/RTKVUJ
q0oqfY/Ew5rioJc/EA6Daz5gGBDM0kRGFhjZdfND+3G8PFfspDvAfitFAmwnawAA
eBpefPkRxmqGXlM5O7CZVvHFkjKFmrhQtBXLKjeqV7YoWXXict9J+KQBgcK4IrTw
AEaV0nNzpn3DXDltSzeaU8PGZ4zu3h7NfLu+061CJ9gNKZBDhSTvYEvq2BZCBpvr
xQdLBiRYT6+rKZ7wMZ13ORUctVQNUDHxH9yORS2CPrHmXHOeLg727DL0Hx+2RvMh
nhb5WUHzydHFqpUG2+DvJTwF+uaTDwY6Xp/NmNj6wkOJiTtN923GQqfOtJEhj6g8
q+E19E9NI1w8w/UV9vEMjW2rCQ2vm/XrWEiOzhKVD5sMPkzJziJhpynVdIfJYQWU
Gom4OajcuzqKA9Neu1yf1mrc6XXXHd3OLs38SfJF6WtlmEh/9BAR50Hqphv3i7+a
VuEMd+Uh1Axjv6GUb4qv24nSePdsS4n+9kyVep3KNYLV+FzawoXwenNHmy10/Sx8
qnDSDa1xmyeNG6WHwcezZ39BH8ubVfQexhjkQT268/GxUn6brihk9XzcVKPSGjzo
ApBi086VVizhRdAce6FWCVG4RQ9ecLv67kT2zKCJx5Mjw2I6UGpyoDtDhq1X5/QB
4PJkulP/EF4JBLUQrTL7o9O9dRcxKGMci00NUWHAhwrkEuJAl6DPuWV5+9gM9sbd
NCLoE448dyKgHp+jDiTf9Gnrj/viTNsOj8NlSfofK1+sa7xHNQoF+i8f0TLuNuUw
iMLBGja6Jm8iV7vM61MK/OFKuyhFTIsKvdulL0swwAtU+owfCnWxsGx5Z9rbFTQg
DCg2cyKg5fFPI2XQo4+HtNk0tYSsjLS3mtJ/WvuyB8o69tuO9i4a8uZBCNP+nj8c
6VmhpxSqYfDambdeWi8xvv4UuXM5DL0UetuVTfQE/2w6O1AJoQ5JS4LsBjyB7Fbe
YdMf1g8zdrlNUIUrSDE/zTkj+ZpAJLjAuOCv8fjlm5ikioAfG0DcmnmgXSqa7Zcp
IRx0CD1YQvvwbKQuVeP3cdApSVy1+k9qbknQWYEa4bAVR758Hkd1WKTfEDasEnbg
Pa6T+GEhuXuaRerMMF/WpMMhzYgvlMbjxtWO9Hm+mI+ExLut8ZdhDH2frAPoxnKT
C4z/ndYij3wOqNoEQx5CNWYBjTsjXZ8/+ScNX0i7vPdVSBtX4CmZQG5iLJYhdFEE
d6Ihmhq6fwW4KKasjngxbgwGKxBwaaDeTdqleUJNSDOXBGoK326Im3Zf/75rYbQT
jReLqhBN3sc8jkjPz2qyumS0qjjTohO0jjDIMHMxSlQCdEzzW5dbXHpHt6SIa15g
zZU5HP/dmgnnYrBD0SsxiD5xWTocdKC+b4JZkWPC2SkDHynjUee4G8PeWp0PC1wV
uQziOoJHYbJU73KJPgaFWJvUNLwf61QSbki43dET7HxEG567VJBVb/h99Az20b65
jahI0FENSOPcWw1+pczH/FK3Cn9wZhMrx20fhGR46QOTh+xgwM0geRclSOuD77Xu
2HaxH4Ox2y/k4JnrqesPuhdXbFqKzOrTqlfP05HEmKijl/wm0uW34CIh3R9bVEZh
UWGMXq0yo7kHe5Kl/P85/chy6YeK9wYOXwxhocDbcVa/0GUncvLcaJNsmK7i79By
gTC5qMk12VLHme4NdydGhWxbgIRZv5/As0n+q98H4PEjdFNvgptVXk8dE2XMOmZt
NFS/YOtLFqk0TRHXSOy5BqvsecVykZM28HhtYkheo6kFNKdk72F76akz09S9ajuA
Bpq66bhTbiSMsDseHnFDYQgWL7X7RPXZPPPl//sQ3DWgEPuOPua327AVKJQJynCN
W/j45m89nrikb3O0zHZ9JBc66kuQlv+1F/FlvX9FIhb4mq7jL/xQ5N/2pRBDFrcy
HxNIp56BTtTE+70/pjuiQ28upSJXjTdEZ1REbcVWzQVRv+qQmKr5RHUB09MgHfLl
13iaocpB4Kr25QoTbz2qG3i02uPtS1Wd/yAV86ZRrbG3V7WihDVgSdtg3HJ9l4MR
y8ThcNvPlo5Y2rZsvjvGW4FIAwQadrLSptJgTWNhLT9urCzGB1qEB5LvcFTrXd1J
ZtITsvIDf2PbuoTLrVvj0CIUmJmbts0Acq/NZsJ19420Gnj0Ld+zxlP8xMVCxER/
xOAVRWF3bAYD0721FfdMiOj+ClYDb/Xr3GM2RGGYQ2FRyIBx2E8N/5GSa92OowTf
ipg/MLfuUz9lHX+9Q2YFeQ8JmbGAy+UptRu4BSjoDde4j9tcJtb5Yqc9QXipVvOJ
TpGgKMnWSceEHYskT5DPB/jRUJfEhROZPuCUoCEudjjkHpF0V6T6s+w1fBP7QPIq
gxnm0/8MNnjX2HimudCmTodq7D5Q0p8GStUC0EJ4ppRJvlhz2n3k8vKgR2w2AFvI
Currd0wAdBaDEbLNdCMpCLrO5UwYvLsV4PWc+bhgEilSku44Vfe8DnfXJqzyNjlw
A6kFKpMNzqWLnXFmRMf+BKGfqlQltXNsUwRH+wdzZAta4q0s+0hzj62HW/HLDVtD
S8Uu1bN7anwQ/XKCkZVJkNijozY+Jz6yGOx4l88pl0y9PkiKjeKNrbMWoR15lKUD
2ueCsSTYdz8qdoDuxDuiWECGATEdxBKeesr3ZIe69elVGI82OZtTOi8JurPdO0Pa
oVUQj8ghClhhhbbK4yUpIZh9CdS/+sj5xHI4wiaxwwOpdi/6TKiacLLBVpMR9/nX
64msKNcK9DKlM64C1CUtYDwm7zaGcKWwItBi1897d+M4kz9NME8jIIiLX+0fsZmX
AxumV26v7dO+ug0tArnuUDtP3tAVZCbZVT3mQOCHVv8+mG+Dgb0z5YmETUeUQmCh
vYWPOueYc+LtWGOAkHX3gUH7/eMQPU7hXF1zO4S915aXiWHrRfdyCxAvguAgqiN3
br+MJvNcTn7PURSlzf888MERRbbzdFgkdb/H7buHDi8407jIJBlyVtkId4AAYJ8S
xBJu7ezFrg1D936DSL/BjN/rwVHwiOdy7OR0ZcaKw+pHSgjsHarhrZ7V3IRrlSxl
1HarjTEAN5vEtUYdrY3+HNP4DHUXd9A+r1LYN114QApNaxVeKk3AgNSjocM4QoUE
zakCtEMSSHSho/uE5qD+eHLluy4DYESccRpGFzNIL2ZhWM+yGE8mnZMvZu/2Xodj
ZF1QsejwF3jbkVTT29TH5vCL7tNlcr24GTMEHNPe0cdrs8ZWFW5U6pvXdroG1feO
wuB4LxV/yh/B/5vv/E1p8xcCdcLKTZEZxauvzEuypL6YpjObm9W5HsP8MDoZaM6/
cHtFkqN218y7bypHxK0HKt3rl84uls9knWyltqm4yE/yzQyhhYXz/x8n8yQuE5yA
d68tTlHulIWb2vD6BJLVsiBZCZVC9W8IaE5PbDVFIlzBJSdaATe8SASVbBNcWVc2
FZBp2dDBv+2sTkbC1OHw/vBGtU79L5/FeZr9mGmAZtZZX8QheO3/Ga4MnfLuRDB9
7y5uP8EOfR0p4ndg/OvMc9gIJUmRPVBft8QYuUBePKf3kBVy+JR2232JcqgFr8Ec
AlL2iU8j1GB0H4efYGnwyMJPIT95hRl2VQ5AmKqCtgjTDdHSRtHNMbrc58vNl5Pg
SXjIwHVZpwcv29HsfKmcMh1JaERWBgowfndpIRrV1+y/R+oLPRUPL0J3Ym2Hh17w
gtQIovV5nJV75ze48UPG61pNZJbLphCPdB1xwg6xBQN1/U86vicZbsxVHxzgZeU6
OOevEFvnN3VcLRI3msiTvbV2J8uB6WO9cE+C7isEL8hrxfoSn/qdEHCZ0A/i16GX
Wi2sAE+9AFN7sbJrsggDLK2vnXDT4iIv886XqQ38Zodt+30HJHYTQO7D3PjgAVVk
hP7HsFvhE5myyfXKtsrugkdPoOVdTJhZ1Na7E9C9T3W4A34YvxptreBfHys7g93i
2zTHTodqaLONEgfZQNm6dTUIfNNv9WVt+m9T3LlqFQ5iitlmYuoYJ1I9hkywv8go
FMnPqklpEupk7U39tacef10THnbw6Ppk6UPNA+bcL8rHh4rqzKAIyjzhmpLuqB1q
zEu+xXzKI7clashn+N/69AtCiCTk6sOb7qox/d9ojGrD1pFDYheBRAFbyprfXqK4
PdM3Ie3CF0L8ZAEqWvfx5Q8bgF9CuBNxyaOEu0w0sOyWVxbfVK3L4MtXXXQX35ww
jLUzsGik92UGl4FVMHTi7mdqoNmdoLF647WwvLnQkuQjckmQkBZj5Lh5FxR1D8+3
LVwo00adloj5zh4h6yIwNoWw3x0+Gac7QjMdm27Q9JNsq0rsZ5uuSheBjVr9WaYk
ARD/5V4vhbAJn7VrF105tHbUMFOhYLGRg1Uh1vEJElxUNgCFg06Y8npygmrRu3KU
l7EaszCJV439uBsTNCxeRNSgjnG4jA3QO9ky2XWVBb0bAhl5Za1P2Yv4ktgjFC9c
29RU4QtM1RJPWnyVMugpGAdUnBD+gExHbMNkm0dj6baMW77aZj1Ji2ZGVPpn0pu+
2f+KRFUMS3BgyPONCKizfZovfGo1pwopsdDTmWtNGKixVDkz0BDkq9JwD9/BPVFY
y9TmLN/O0wv50UeU7o5nB+gX8HqqKCZRONEfqWFt5KTSeN7fhAp3kCg1i8WoVquS
kA7JAwDIsHE+o0SmGEmH2RiMP2Kg9CuIbRjdmJFoCSIqqYX5HFwAJyGqVew2i/M+
Jp4wdleDzKnsWLLIt8nl+of/O2fBqZsD3AfO7SXADyeCxoxzbaH7TtRFKsxBAYsS
BhMd6E9ayi+Aixyt6mFS/x7hHJPDCCJAORPuOnEOchUpnK71TeXBv8+vstUofown
sVCpV2VVd3gasfipm8Ra7ohUl0sTVM5d57RFfww16/m4s8SnN6fdrjfJ7SoZacWm
3PzcvcHDYivcp2e9zqwO71m/Q63YQt3lCqeO7k9OoTAhGvy3eywSNEz6y65sv4As
apYZseqirZ1nYGym7KJjkXZECAp4Mv/f2F/woUgrgEdrTm5DdVJdunQ8ajT7fUsZ
bIuUc63Gf+e9kRF0T3rapfCVoJvPSmKkUouffpOWcaekEuYDWiXzG+DKIdVs9kUZ
rddvOKZtw8Ck3XBYE9rU09N84nqAAfzZ6bq5y9TFxmEBDyWDFzxZHrh3gkTS07Vq
SkDTTF8W1R7mR0m0MOPVj/MhiVlVQPoHzSjeGpVZBUIc0Gan320KJKpm9FZEfRZM
liSHuhS8b1fSCIvb104HbpxDVxGhxnNuuXjAVOgx7L1aV/4cMfMkcb0lAUOE5Wq3
+3ZREbz3NNIWnbBd4lU40oUadUUxRpLGXF3na6KNdpvDIf49/afxbVFG8nODuDtk
9GLmPNVdckZBS1oRQmJqatFVgNXX5giarvss3MTjyiM1FRJv5sIDuB0ao/BSW2n1
G91y4DPFqJL6dJ8aO7btJoNaxB/SBX9EmWiF1z9Dy1Q6IOAaAa4tpJzrkycNZ/l2
Ik+T+Df4y4hVgnBpDIsBovyBhniLRey7/fo5Ya5VQv63rQ5mqCcO7gSygYUNsWPX
Dr80ElxO6Ai00Y7dRs/Du7FFdKN1LfdV7Hua4ve1AVnZnsxU9ragNQFRXKIS6kjv
a5ZWPQSKu/0MNfH9Impi8VERruWZJ0RGA/9yUcn+OcFbhAeKdUbIw/Cq/xttXbaV
sglzS68/qRtBK512yCcjLPSW8azXCxfHPgQ1lKdV7/Zi2geov3QkyhY0RVnh5goY
llwazkmwRe1ccQgpLWtPqG1PszDsg60bNmFSTA85JAyV86YVIbbc14tY2PQrvKiX
2Q1EEfF5Rz5aNEVk9C8N00KwafsvRrqe6iNwI8QxhkxqBrlhMWSYSgkoU3GQ/TYT
taNu8xir1w9eB024BMY2mnTTil6N7og7rAWVlLUxtasrJKlP5HnbSMDhHWBV5+Ha
CH2JcwhcNqhPIlfDrdxssA9uKVFyfcCEpOVN5NeBUo2u1ctWaTqZmjc4NiGYB1ht
8KuCiuoiBYUd3RJES+UtxdFcBT1OWDHw7YzJC23QE35nWR98pkG82W35OhIM88E1
uJwUr94QJuRix8xBDhPsQjmtMQV9TP0zYX/fnj+dR0SFvYKh3o3MnM6QyQijyimL
lHSCQKS2yHphj++3raq7bRInJaSdmFrIqIByUUsLvwKPl6NR+uCHdOhd4dzgoAwW
YXrauyC5Gm7M9sZAU1vfo3IV3/tOVxIud4l6Zchg+hcS6spgD0w2emR2YRozkSyY
a5WonLuVfZHWzg6ZiR54G/ykRcyqGwcOYpSKd7H4KMF/vKQ0/KnR8w/OWu6Aj1Ch
u0ZqWhMFSUJu+uvwGRE4ZAyYEJ0L/Qou70I/QWOPnaI5uiX/HvglXdDIpjLppwfF
aMmZT/9a4WUbCZ5/z4JgrvthLOUFELHKhZNthqlcadkaiobYPTegLqBO/kY6ZNPE
iffi4SvnC3pEFhLESiBvu1lLtv5S0sSV45wai4eW+HpAZGaLSgYLzlnnZ5e/rVE8
1ClETS85+LLr1xO3YaAD1tXf+B7qIX7st+FKh3L70LLwOjcSJ1JANxVAR80YV+e/
HtfqiB4j+Y+lzCrlICvGkIK3a2oAcjCiq+G6Is2nt3f+5BD/A6iykzKMDaKcWS7X
z2OdITSoB05q7pvTcaInKiPIiicpZiEGjjlbdHGZML5Q6CwHqwA1JYFwT2Q47C9i
4ayLyxU88B1gBApMSnkPOvd7dO3yw5fCfapzCL8HlUI2niLDttXMZp8yAuQCDufO
UqJGmwN5npLqSxINbwV2JHsyZbUWSbLGoPFMJVc4ByS0ORIwoi2KJ7tZVE5ZwF7g
GmDuZshUvIcQA1POZV6LUsBWW4m+1K3933hlaoSkQJBnrdZBfR9SzgtXnHg9/c0H
qaXI+jfyRcAnK95N43jIYVxI1GCWMy9Pp+haqvTwZ7qZpfAnkIAoIGEMiVyPoekm
Cel4fGQePzeb4L5gJ/+zoTjxJuMdRDdLKy5SnWevsL5qN9LUdJnLlbli/SYAo0xp
xTKxrYFKCOvmHMCLMvk6R3mqV3/Ny5bYy9qMScS1spjEBOjUEG4i59Yu8E6u/HKH
yGKZkiAYGXbN0FgzUcUDkh0Z97RtNSQGtXCfYXUsTeGS1x118XpzM1ABu6scqylL
Xuyf1Yn9Oo0nqg4+pr1zNXWn7I4Mxt2LabTuBr52aB/eD4z3v1X4Oj/CSXHl8uht
q/J7Hk58LLSdDggrkjxhtWYLOgWJelfcrHyL/UGbvWv757oAgLKzNw1oLNuYO5r/
7t4p1t1lQ8k9DjN4Vr7TWTdmPeVFxld8QHSpnOnWDoj4vOmpMIxmDRyudAsjEGPm
ilmpXiL85ICzxNnwFNTcd0xzo+5fFD3DcVfjcYLnwws/sg2hrnzRT47BlMqpziik
nCzJ4/Atnp042u8uw65sBR3Tr8S+xCQrgUSlUEcQmoikDiwEqRrr1Yg7xT7bS3hl
/u2tCLWuewI1hDBFlru0MjI+DyTRm/yVtF1NILmoweZDBh7EcWxKMkNgaxWz9AaJ
3DDvasxzwT+Y+U0BEoHk4miYMkmQPpsQ+BSL0gusNBpkKyCJBFzHV9/CPc0X2tWn
hqGNX014fY0z0otZuB11841YKTm2xNI6xBeSkejm9VOTA79tlq6Xwl5r7gwr3gkO
W9+7PlDhvWNQSU4rzd29s/Mkb10EZtfgGZWHIJFLBq/zw1bwtX2DTMpW4lRyZRX5
cpA3FHAy15ZVqyMUqiEH96iPh77Q9gqx7jBrgbA6x3KCcbrL03slPyHLpq/UBIew
M1cdXWEwUg2cCTeBkAWEs2H32pV7WtwZKk2m7HK15LTK4JG2Mxqap/JYd63Gw8fS
b03oJsvVtRTsUz/vSZ3+E7JM70ylQ0dKQjwClBjFmEE1w6XIzyT2GOdtsO3FUcbA
T9ngCkCu4dCL8nCawysMvbqxJV/7p0qRjiiXiZUvTgh3rvSZV3qm0myPi8g/Y7NI
JCVHAVAUinm3ZJkXSOAylc63cRTdRvB6k577eRG4n3Y41Irjdh1p94Tio14X+DEM
0avL87dwHzaES9ow4IEwFP0IoX7Se4a9rXc6OLCWwUGOi9y+5nVbKLkFsa3JGvy2
D6hriWOFFHfhUVFy4nKCAl+yHGMMHPkaIFnjeRjnIdiSgtRfamMFqgUbRmAiKI1N
ezp48GaNX7W9hKwK5oguuuvO3AtMx3zEsSdb10KrcwhsILVoYwPLqZPBvlRcjLLu
IWkMpzbtSN85aR+QP6LhV/BInVvu2gmp1sH1x2UCJuQKJdbTpCF6opuNxBZ54OFg
ObChwkfXi3CpPC8OJgz/rj90jWpZeNqh289C2D85eXHI0jU2EpRJn1yUuke4ybE6
Vs9UZ3nnpk4yVxRIgtwnM8lrhDXfIRUnYpsiHEwkfIx9OoTRRjJA1zGbyotd/AOK
Sjt2oCuIbu8ERyA3CQ68hYjTZEENSVpHHTtN/W2Ql5WBaZYqbknM84L5muD43FAB
Akifev4tRXQCtMPE0mK06RpOl151zUWGw3liLgne4MmS6+WuD7ZE6PK7xs8ZhoZR
xBlu4+zEXJoJKkCuhCRGp0nQJO8wPKD/0+nrvqbcPZP8zyJVfPTTUCg+VO3jvcFP
SAJjcFGsWGWRiKCj5/3USF23nrJUcQVGIiM2hQOzTWqh8pI0/Xax9FcyzWrMlw78
5jtHm1yj9c5l1K825tYNA38d0j5B9XIodyz4Uurlj41bBYwXssLu0xC0wpwE8rr9
fW35LUZQPkkWpwQ2/gRhC4p1nbeG6yyCzQdoEUxnOAaA+B9ZoZ6Rd/7CTmkyOW6V
e4tyBeSoalFs1vNTZYAqJrNW5+CxITxos0QWvC6GaLY+IP6HljpfahBph4OhyPlh
h2r+Rp3BmZCo6Gbwmi5keyzDMT1EB/58bNDUS3CgRihSIFnMGhfIUPBwrLKkRyhn
2mdgIbn0n0PxBB13AW4/y7LlU5CJcAFszPnFnTO0GL/Cb8mw2L/Zy3ZW7pSwKEVo
n/Iv1kwTwIHnAdyiswSek8b32+PuvoPyYqEb61wyt1OlFPVrmtDbupXwexN5p0HQ
tJODCfV+gvrwTxwPmPjeAEPe/l/Leh8Ac+QK//WKjvVuQxNaUqMVMlqHy45gqVTS
GzkukTrf7Vy7lEg5/vksGhU8PpU9iM+u/EEi5FghHHxw28EuNE14GUwHNQg3FzcF
ZzjXOY3O037ONSA3RtGRnD9+1PqYfAgnzA7EmW9Rx0IKRZktqhFboxtj4SfR8bHm
pIHSWJOVckaqrPy3SIsFLsr9njqkzn/r0vkZvhM5kM+vyPngFjRwetDhr8uWsfpF
SzRaDILvnSgpOzzYUroOiRKwa8CDRrsZHwveJ+740BXprEEuCbiMworQe+ar3q+O
N6bCySE326CR9S1nPIYEy+IWHD0lX6WKSUqIx8vKfVI3xVXhpr2g8TRVlzWAxiSL
WHZ7reN1JA69HKVbutffqrh1qQ5Nrz2jn2u5j44KPsxOStpUvyZU6uag/VYjEbSY
uXorIf0J4txNFXfLW8/v0fQopBKginHfviiwA/7oMe+NUql9ITCFgr+Ev3clc5GL
+t4CQvsjxv69adgEUuGsVu6azS82YmT9lkszpGPyRp5Krjk2MtlHfepqOkwJUik6
8ngwlb40AdwBFiY7SmaQyNwVliO7Gt5h+zTriau5x/RxZzdiUUBk+O+jUEewIyx5
BaNwhU55tOqDv8t2/U2sazsruy38FFCxsImdYDm1UI0dyS1npZZm3Ipt5h7D3h4w
VounWRSf5x19IbJynYxf1dggSmkqEq0LMZf093gp96zCxZpCqfZESFIN/tt9tHZY
yVA5RUQuYPMRsJ0VA6ba4xNUhhGXmFFx9c2ngQo85xorff8+iEAzAzG7u0VHkXYs
Vu9ZPUgDnPYF0O6caq46Bbs4TYObMRkZoxhRFtDJhjgysciB3sESf27n0xbRoUwO
MDDwABUbCE/FqpUrTebh+sNbXtQEC8Xyo0IHx37FOxZYYAZ1gVrt+OZmUu6SYxDK
SkBLwfHDNGzprkNkIzo3zyBttuTK3aIW8+pgIinBkOCjA+DPami7YZneCXScQUIx
dayCflWlbd6yy9/qpN0mpdy8p2bpldB5hxsUDH0UPFbWMDs3/HM2t0GnavTL4kTs
shQSbx63feNBVcTRTgziV4B6O02O4aEyAKf2bg9ITgvCdqnS6sT8fchlsriQQTUK
3Gnt7NhAbWVejp+gmUQDBDZh8mcnX3ZKlQep1sVuBTHlDqfnSoEnkivL5WwXNwTj
pTv67GQgyi5tHiqEfeIU+lxwhcm9o9Kvo2hiYJAkuric/yTFyvp51y1tWREF1b+P
KVebt2BrmxC2CHspWtOwqfD9/Bldt3AxvQYz5TKZZXtQ8eexabK1+HhAMeQSwd9p
Xv2b6hIqMunlSbeG/VhpFPNp0vMlT8bKdNtouFPMF3DTI+LhXdEHfcSiNPwcm5xl
xUBH7JhsJElYiZ1ZuxoHU+MOqo1S1pNyaYwP1OuHqDAYRiNqY8Bu8U3234ooc8jP
/klSwnVaij7+SKFVdHrZxzUNewglGboD/sB6QZwxVgmjn2JGHQaHToV542Mz2/3p
pYefEI6c6+k+omn8BOFaomVzEisajksBb0a19vF5luIwkReFeavq6JovhhsQE/ER
dQTF+bC7dJ0ocN2yw+GXb5OeTtbQqeFh7PueqIvA7vqmXGjzpiRHAhYCSGy6KIpE
OoxcE2CjzUtxIxbThLO3ruuWqzx6KbxbPlS4YXacg3Ha5r20hc9TGRHNS55d7kyR
fcIgV5mzW1S5jv+HLIm0+jsh1oGxUllc2atdVu9tPMfPEIOImWc6Vzvn3zH6Z6AL
fRE6pDeW+tis2X0fbkeJ6w4RkGvee4sNReWPo0cJ+gDs3c0LzlLQ99IeWBxDoTv+
7+9M0Hly7jHOYG7sRBf9V2nBaFJqb2T54DxwKevd8hbPm8XFzGe/x/8fE9CMHqTK
7a1dQFuMxvfiVQbFbERHqsLTlFKjPv+RplzyodNWKy4wrEcp5Znj/75AI0MvMyxE
FI88F5py7z+Kz/ineOymDHQeTNmRMrzgGPq6kKdyDbGtar3w0qWnrab6qg02iRN4
UBUyIHaEkC88jvVBKORFQXSavJ8W9pjgAoDwDsnyGDr3D8bdT2gP+E7q1BiG0woA
8yBAhm7e5kTrC5gDQVQhgxWQrLD6XVmmsy/9HQk1fPIAsmoFOMWSRpmiPoonk36v
aceiYQTbXbecoJdxWIm3BcXFmNwfl6anPPdqINo7hhGURODI0ikxP3hDQl1d5jYg
gaDbi0pvlKmup4dDa5d3PR827m0GgGk3FtdsgWxguY9WBxp7V4eNydjkyOIQQhK7
ebGiMM5XwbNE2hyBrMfHOcKnSW/a9TPD/6gjotLTi9pxPwH4LrFcZ23f4o7L+C59
0gYC9tMkpN6rYT3lyRr11jAcC9w8NI/FrTWzYwZRuqFbOJ7gRNi6Lb/vjPqSguFa
TscbDeYCyXbY4nBAQGaOc0Bd448Y+pw1hvJfQxRpkA3zzPPjt0uS3SAe+toXSZW3
O+H1zfvVhn+4CCY2oK6S7QGLQ4MPZrxK8oRKDA9RE10zElHtrMXawHOqI1Su9xZv
QkKVoGGRmyGDDtoi2BNLPXVmw6i2kMsWIZMbJ8+UgWJuV8afCgO4PqpwY3T5lnDp
+MKjgsWknHtEPIHQ/fcUziqwXRa5Z+V7YfT8ShHTvGNkiZORFQ8QXbDG6eIiIs6D
9FeaS+VBJPYaG5qz/N/qsvYYt1+hv9OeO0pLZ25gpT1cTZ1+67J9Fme+SurF6Tok
HDIeAZT/PqotHlpoTRWmoebrQDLHHDESiRNgU+i9+Innp3DEyzoasHydHKAcmNko
ric8ktfnQzUUN0BMY3c9JUFOGQkl6mDf4hFfwoR1SeCbSL+f+VhxqbD/v4h8iVSS
rNVDrZeoTJQvzcIEO6ryVlUhykd43ztBpH0ntRDrxirOD6bW1S6l4XOu/lf+YEiH
W/ke39ovYxyy8b+VCLa1Lc/W9bH0VO0BXcANzk3KMk/5RfpnJoX2xNTGWy2LAw9k
ZDSo6KS1UIjmSqRJtvvybeR9H6QVix2oJUnQtsQkiVbz5r3BRR+W+UVHyDB5oZKb
c49/YN/vjVygwI8lccaZk/YzR5trC5kImm2Koj1l6geC8gpyc6JsDnMyn2sY/lO3
KF+P9BEndjFNZqHGmJ7wHo40yxYFHDXALiT+EMR5dzGGexh7a/7paztgZid+TIS9
WXPqRejnBM64BBi89pZvG0sJsYK4CZaehE7cBHAiPUIe8VF19fcE4y44KYZC6P8q
2j24ehHaG/SPKzIRS+qYb0aCcXdo6EZ5xB+SUO5ByYJkREBuw6NPyWOBMJ9AW2D7
b9CNxx7XYyTP+3TaYPxn1VesBg5TNNyTdzRJyiFwNr+oHx8GyhitJbm1jlmiVaDu
nG9a9yPAcHleSLauSQY0758exlcIrnqdR0enmEg4T3UOpQWMMrw1cxri5BPaQoXW
sNPM/HChB16TN7Fd/FrXRG/uzzwdF9MHPRmnuj39sC8yoU+362oNJuMj/jsFxCyA
pvqS3BAh2luH5gnDl9WsAVKnCZbRKQLFHLxcXlb0oxLpSB2o7tXW5BUOb+/o6vFD
QZCJHO1gzuBzisKwdMv+H2K6z/C7Pn+pjHGpZw52qIUfBbm8FHueTGYIuqk5X9Bs
trdgF9XUksUjrxpVgM6JxU4faWo14TcECtSKXxZYxLw/7yXauhnPYhbNiURZC49f
wPd48VVOmJz38709tWwuypkz4JxiUXK9nebrVL5bwdwofSMy5UeZHPJ2IjroD25q
VJTHZDrJFU57GYgyoVz676XVKZt47bQ3Hstu2j/JGsUyhPKXRZlhTJYcdMH0t/oB
wByFO+Izrv4L4NwdUvXbPg7wu1JgZcH4Hmfu8SCnpyvG/qKXkn5Cx6uWEPwYNs5o
0LLpDPmW54L+rhl+tGs5M6PfhUhh6kFh5y40+Ao4whRgqrYu09e4acGh26X3R5OZ
lTRMSFrk3y3Ers0L6ZGH9xehOtzlg9cauab1DVYHWOYeEEYmVNLRf3rEim1baZ+W
FJ+7tvYRwLqeHGfVdexL5UvbvhncL0oubqV30+BEOKHY05mUOqLIrGrN8lSlvJG7
kq8tAqSyvQuBXC11XyE5VxOuLv3cKhNfWm3dDbrehbctXW3tDcZULdZFZnJDT0Zl
CG4jv6iVE+n2ONvQ7wKu7/rud8KIT12gIrAKE3u/BiRTBA1ofNDqiK9uEkgCKUcm
UjwvwR3XLULufociS9fIJFTdZwJfW1G+LTO+ayt4iJYZeifptqXUPCjxJaH5KC6n
aVpAPS7K0k57LkM/WFVmDsK5KiLQAHbDDJsYTzoW6B4G6LYgXgb66RHMh/jdo6VR
hgzgSAn2brSQfAKCFFwOy5rwoolOB2olfoHBxHWEr5ZNhutO4XwDadt+HHYy8Tjx
q/YkUYzvUN6A6hjFwvsEBgtrTK4pR4OPsbngyDGDPGSKThUf3u66/dsHkBjh2zOn
u6/TXCXoxsfsZburwJngeXGvEl/Mh4wbDro9L8qbYuMsRBCgw7udYRek50bExL6i
j/en7gSJC5/xM9rZl25eWE0AQlr3LHD4Zb+j1F9Z16dkFP0F+1OGNkp1jw6z1MS0
K52QUyARTjf3JWqDkA6UbJ8UNaq0S/GiQrOqjMgk78fhHkHjV90Bh+hgXlh7TisB
Y9ZOJG2tT7181uh0Iq5ubuz2yxXgZE+3yVsI1WFfre5s+//+IOYUyG3+K3ov2nXt
NPwVyAuGWXXju3pX3rxrf2f1+/Nb5FDUfJZTG8l6ZLIINihf4VADn0PKMinFKatu
R//WTHhy6xbcfOCHQT6wCsA35rjlcoxeaw4Bn5ukiCuJ6WAknrP7Ohc9dnEmff5Z
8uVaMFvGw694c73lfvjsOVMXhtLaEEviVz8JoB2gH+AcCeIKWUjDccXvpP2K1BVJ
HgXQmknZiz78DgtLpoKu/JJRmC03or6jvlAcP/qhdtxh46RSnaO69k6FFAwD0W1Q
w0uySCoqAJRScsq4k1g5wsPJsQDG2sfSKcPuBUPADY80EsJUtMxKsL9i/q84EO/J
wSwqpk6glsnT5LcQ9JuPQmuIci6VpK+cHHlfHqHzOs/gBbLPGDmE9XOd6qY6jBms
ucJJ5Yy1HW7XYVXSz0fKsTgO7Auqnuphzd3kUMrawrCyBh0PrXoqBlsGsXczcshL
qv/VtbURXjMEoiA2+8avCCFOIJ7tC8LhXNaKZzW2AL2CgsMtBpASF60EXlRcBo2Q
vbKdodj/s4kzZdxG07a5QP+LMHsLQeTvqNa799r25y/LUpFlScGz3Ue0WcPT1f4M
UuYXeROBNN+1Aq/5GZ54SiF8b/q9f7qlaoHOMV7i9BcJaGGrLIAItxB5cS4s5/S4
vhTzm7I7wJDZU1E76S7NtIj0v/JP0lJZyAbq0nZjLt2hERmDCBQmApqnG6icW58U
Kn0zU0VghbnuK/jEQgeu2Ig99eclR69DmIVKKNJlYFVhM1HwP2Rt13bHYgq5subn
4Wwwr9bU5d/3oQWMSwTYDbm6DERjcD2dGNQwn1cdpw+9L9fUGlYbaDsA2NkiW17p
uVeEteYrMjkUtqZYx8fo9KZdyIHBhanx6PRq2DLoBWU01VaMa5zwyjjsbV7E89PN
O7TaQqUCwHZaSM5uNcpsCO+H6YD+DMg/j0udbH5wfa/Wbch3EXXrh9sKr/pTmeSU
WrWCtHDxO36r0ernk+7RFRaHEuriXHos5RFBiPbw2oZNgPfL+s1J4cnhwKhC0AuG
yOldVAMh80wAOVbOhK01CQK+tb19veGLrU3j0rgu8hdkrA2xq3+Zhq5YiKZx63QJ
IHYANaNt9T0Ju03SehAe6wHtrfbNLy24ByGdSHD8/Ls6MYeBJ+6YdIDFAJU6zifJ
yCbnnSm1/2Wg0XalK7rDm1SH3W4pxG9vkTVtH/7TLKyMaFzrHFmqt7UfNE2UIH5r
019ofErxu2Krt+W9v7hvc3wnHqI6hYJXvqtPVgbQvYVG0YwLIo93oePoV+ZzUPIL
VcQElTLqmSza7cILM20Wd99GuCZQSBJDZjikgA+cSSonr2o4mNvm7V0bQzmFdBgV
WXb4bnwxwM/aLciXad9EoBy4bMOtpSLBOAsN6SsA0QQmXJmlhJFsU11+Pr9J828q
8tzTn7fCjzZ0Q/zb/OlB/bElX2PSzTXCeKo1jBJ0gKYfA+XSb6zwc5a1dQSgGUxH
tg6tw99o1F5Lt1TcFvwgXJkOMCduqRVN8NV/2yFqBTIGXmXOmeIPnVZ820yvfWgK
bNR9h4JaTWe5EmDuzP9pGZLtwRt2DlvHKJCGbjzG3o45Ze/fGBT7zdfa93BUfNL1
eEz6DaCnehoTijTBxDNslT4xZZoqr8MgTWe0zeykMWcMgbw7EeNEBcXWihSmPxSe
D9UfT1+aHuV7HwWXhVspZQh+P2PXOr5lcvlqYRVJ8pJCBceS34A0EiRT3jkbJG/s
h2rV6e+zWVuhshCWhMaUND0svn70htAIX1flo5Om2dKHE3MFnXNb0IsN5LoUOO7l
5tD3QE/wTlY+BxUOL5RjGitIYquIbRRBEFFnhxh+xskrgSBKiDU+pZvRVQdClZYj
c7SxEYzX7c3UblA6rhS4lys5JjVlCnLQvOPzCWJfTXnWhhunujKPJ3HHQdPAVvUH
byRa9KrCh4VydZwCxmbKe4Q1L/5+0jWksBouW5YF0PjHFwNvOMfYXBlnj0OOqb1W
WdeIS9YcKuG4yONk7CJvrki8XqST2PSj1pvsB2fxH/QotzjPyZMytK6Ntf/9wtUN
EqVqa0fUI6s07o9s2C8t3JwrpIhVstvDUOsRNVWE2oaxWXf19vqr0yiVmew+pl6Q
qglzjT4W3goslJt6YHX0wKrqRQfZlcxVjvI1iuJa14w+Fs5i/g6DIop/m6E0FfCe
hTkDo55J+Zp3sQialeJoshYx0DsZXCFMJGR1dqpRjUxgoLClUbC/6+Ge6sfiRmP/
/t1tgrv13Uy6//w2RQ3+T+oOJP6EEiZvuISDImVsGYGiIjhyOG73+FuQxe1uAluY
5/lMmdZQUzVgUwgrV7RddHl3NklHecPk3g3qcFehqU8dMx/TZGhVdF+Env5GrTLD
LMpkseo8GXRZ11It44H6i2Evl2flCKXkMmNMhY4KUyXHNM2tFy0KyfbMwD6fhUU1
2G+w0b8Yf1QMGSNv8rVBoS6YzHZ6PJHOoa8nhR/Xg57/DIhobRAVxwIXw6Y0jkVs
QZ4xnhYvYK3cW9KHfq1J31HVN+01yUV+V6YlCAm4vlQxtIQ+NWtrtq8TyB8zms6G
C/Hu0A7eMEi3e2KKNlRz3BVQUWv/K07BCP5yBM6wFrBrJ4vwy5RUEU7sEZcYmNoO
Bwf2YV760k2Jlji527/1w5kKyqvtQPxO44nMONoTlX+HFBn9qPwZgskf9nbl1mW9
E6OWdOgVpjyg1vORh2sAfbQdYnx4XZ20gpXQR/0+xGJMYjrKN/n5Nhdqa0ZMGmGr
3WkMbQBQtlyzCCJU95wSIP7w4fJu+UmcU+fS/ahnwON3AhESJDUpburV8814U+bi
9CxTASTE2EfnISMO43znx1Pq57ahVgRml64A6ugRnwl9E8AnqkKOLzyFg7CTS7gu
jmATz7r7L1QUKDp0QHsr/cnGXaUJP2qLwR1ohSonhE1EC2/Bx8y+wSlsw3sQMmdp
YPSCsvcxgCN+YL9APG7PsDSo6FDnvpwveNKb4RC3aPVwhCY7JsU0jmwerhzdR6Kt
pX8FRsSM5pMI3VuNX5C/l4C2APis71Ci8D0MERWnCAZcUqkUQiuApLNV/5uOlaUY
GM2YnWOkK2OCLrJNljhZfXayFV7nRrSUU4P7m7ezCfWwxbxu6ZdECBC3P0YdF8+v
Xfr6TAnXmM4VRTaMXXr+ccSkLFBLGMewW7ogLMbYeaEGrwW5eNkheYQ2L2osECTy
EkC44G2OD9joDzNIRvv/18++VlECzlNad3548UM3LPMhGoAAhpDSpSojNcoaGrNp
tG8iChzXJRCcsUpXt6uuR6kaM/xm25y11jHEQRZbC0SjVIDx6wIwwYtljplVumD4
c+9ZypeHr34HkUut6U3u5Dtgj4z52cpAdDBK8CWPpaG8sQ0laTbS8PKv6gLqscd8
n8Cd38uDTUddoiI+meiBAu9cOFekmkPJxkrSBhvQ5THmf5cVNXE1hIicio0JBnwF
J8BRs+2SJVEiKC3oxkrLnI/ZgQZAxD8JZCKASAlf8fW7PnllC/SZLPGXOchaEOci
jKSWPLF7VIyi+cnBwhhSLD+m9HdctKO4+YGnViITYBruzE0RMAFGtu/rFPJ/jV7p
PmyqL+Jj8NPuOZgeCd1QTf+8sh0Jizbss2RBTIUF9qNNgEOkw9bWPuGDswudzVSI
yPDhtyIhLI9/bAxXymqONm2LrHw/Wu9h+3+GXuOonZLWLKnhXFermUjxv9E8Kr2X
F3v/W9TOXk6eWPkkIFHzaKzku58MDCOsvnQnDSPjOKfcZ1WpdFrqkDFjeNB7a25i
XM+rfLDj7ad0iAvzWNGDVeUDf3VA2txTfysarc7S9hzNPNjqcOzXaLNnY3k4WXUG
C7sWd5JZiORPsYhzBCf9ynJtemysKDMO7Wt3qPZCL7HomJNbyUXeuDHPX1+au0dm
Km5Z52G13sg4ggvNrd2VP+QZSn/7RWtdBznJJbr3VKGuWS39F/AZa5i+E8zHqUDJ
FYTivK15P6UzKGeatWlrQHxKs95achFaEHg3rsS4odlXcgXvcZp1Yzrr8kh4ugmx
EELW3kXy6E1n+7LlExU81NwOHF2N4FZJmhaZbrAzU/Roqt9SB1wvgzVgS48vgGiC
ikvL7XXSVBVeu5oeDNhNrR2bL8uR/vAV2muYeupiX9K9b2ayi+bczRlKs8kKzulg
TbhADIjD6HsiyWWpAixLk1T5e9D0jIgIEK/9gdHQDwzgVyn2Sq5Ez+AN+tuNyJaH
g+h41j9A6R33Zjh7CMgNDehLMHlX6SpHupeDXg5YoKh9f44ln6Pjn9O1/pn6AlRB
gcA7VP6c6WQ2PyUVI9m16SimWcLep8Np0aJ8JrExpTL7klOD6z6qP4KZtTR5TYeS
Bb2+7d4JzR1AlVHBFaenmcQj2ezNqwdo9aoU4y2h+sPY3+cm41sjdGKQHvhESDNt
7+ODt4/3opTpO1mWLlDEKwia6iMAuNFmaggFGA4Db2ohEV3QNbbbkTk2t8esnHZe
XaQV8AlsHcvciPbptCZHeMuKZCVpKGr6FMgWX0nJOHWjk/G9et3Bm1nJWBHv6Q/e
j0gPw2BDZb6Td/NsmBmiip00oVThaZu3QvAT8Xz2T6PA1T87DwmGo3wbQB0K4ekq
rqM76NjFvVKb2P9Dpxu3JnV6cseSA2cXO7EzTRhlxYdnefWr8lBXFRQhiCw0krR+
8wvAC99Ffpyax/ZabJKyEL1BOXJTBtpylaFc3ilpENy3jLjtZcH75AJQneRMLcmE
Z01d3iv9iFz40rruF2rVJ5hFK0cHEjf0RAVfXSWzgKU4pQQLum1kvgPQzlVS1qwz
0ZL/UlMid5CO48hHdg4QwSFpmwZ5of4fpImVKGjAoIb3JQFvBQLceWwih3pU9fAb
RKQqfz/d8Dbr1nWPr/veNrTUC+JXSlbnEfm0PNWXsfE2Ik0NgKRPOKj/DY3d4aGA
T5OWregCya9dIJli4KKTPl7TmL9n3+edqni2XFKHLs2aYg+bQZ3btIcuNTkVEQ2C
kmp20BKHwR4+8+h/BcIptphjSJ3cIlpFmr2nmgMq0kSBcp3Y8+N1xKjp7aQLzVLx
41DciYoEaN6p9k6mnSquvAoj8ubWH4EPhFGJzt39i7TAUehwQRe1JJrQDVutA1Q1
oSeMm+mwp76bvby1h3j6JgsmDcfeDz2uup1es4k0n/Rz70f10rHgbZ/cCHjzbqOX
PMQtVT96jrC06dI/TDCjRRtjMKCT7bH6y6WaX4PcKVh+eHM+1AcRnO25BhHXVCgP
hJMg+U6N4XCVYdAg1w8LD2t5CVt08YrN+XTwg/ciTXBDlXMGS5ftW02usB1Nw8Cd
QX6Dv2WQjiRJAkOug2syl847DBZ6UBASWtcaIGl8xycB1QK86bXEYx1Ub4UUMU95
dC6UDI+dHTLAhpee2MkGSZ308QA0Kk5HYYG7oQonTFXJ0tZCEaFccFxbSAcSsTxy
Ui3Yt549GSJSMeRJr5L+3jKP6jTBOpCUygyrNpwS7ihMk497k/aJUsXOpA5OADbn
69ZwepFikJIBdDG+B1FlWiCuSgegnGh1rkX3BF7cufSRkGywith/hN9NnrBFj8k8
Qmri6xyCUCc1HBBpWkyzvDKpbakFCVyxad4JbdgQPm/ElflF7v2dIrue9ZnHIah8
OXOnOTHHP84aQqoJgomEZlRILxhlJgU7RsU3VFHgJQ2XlQWY6EwbNThgsi2Gi4CW
w1PKcTUfHDLTPoPTc+PkbxUffWjbGZGj2BDAlrI/RUMyjF37jdCEOPyn5QB0KNt7
s9UQCHdxG+95SVjdAUxwtBtM8l08xtMOJtLON4oh6y2ZWb9C+BIY4yVcA1y/rLcg
BEVSv61espQY6Oo8Lqvwx/U2rgL4jd0W4vE2shDddle9s6HFaYrjxkzrNRtmX9rf
B4MkTmAh2JOMkfyULQtXj5Hbrt7rMUD9sk7Rg2rsmhacEWsWiA6k5Lbm1K5/i9xi
PByEXzFZZRFpIBn9ILAqLcAHIOZzzhMCGxKwbp0FSs5o+y2kJ7/SXPyLCsxKmwuN
7wFNEOXZd7xCz3SEaVsEGGYXsZCu01JjZjWLr27ir3ZJjlbyVPwauH0q1Hrsw+Hb
+euzkbqYLanYHQYqDEGB22TSfi+B5qXuRLGza8oijKnKWDPt3CQJsrs4fqpxzTir
9lzItk6YIp1gCLWThcoaBXUm+GWrm+26T6XDapG5bEkgAvuKCVPDEA/Uzk5fFJE3
ftFniyCf+DnPMHuMN93CbP4LHEc/1mUkU8OAzxpdMU/gcCjhWudXL9U1JPY/Q02p
Rs0vGNjpB6L8oqHyLdjjMhnIG0jMPOomahcvS1CvzUNBTt8kG1z0wau1OUrCqmq9
4yzNnXkGNScpbYSVH+34Vs/QkLlQFlUqpznKV70SxbDvJp6PF5JRbCQnDiCFBgqX
s9/o4Goayw8WiyeQBcpsfxWVITZnCTDxDjS71l+amGKPSaXJK7N4VE+Sa0A8DXEE
eQLbdbP1J7wdm7kVBqqn6I/h49YWnJIbkZgutocLcXAaC1TOcsY6CCIbdAhC92kE
pty7Zbf5sVSaFPqNbA2AhwKb7QI+CjFH6Ee/43lY2yvYh9ZGUHUbQizaHwhmURLo
GAdsk3LtJgmoM3taBwJCFR+hJA7wcPdNh2HYbBimbpfCSnf+Y6lbnnE8o+hZt/0H
VMYFX98QMdZd+ipOgddps9ddqbCkZWOxCo4Fc1aYjyQ/rrMqoR/DbX+epoCR+Dsf
2hPNLXB4zvrriEy4wsFAMMjxG+ceu+k4azHRic38WNzD+wbqoIxYgbDKB85yyIWQ
TYI3s4rC5G0Uu4EIG4+a+7B53AG04QaJjMSWxDvq2n2gnRZYGFqL0xWsUkcV883M
hlrU6OmrTG1+4Qff25a9R6o1Jiscb9t7nXriyh3//eyoSC+Ll4BlSh2sTgJmW/kl
qnNJwxwA8nXek86v6YTXWNRYlQkVtpcpO+VJxpUFT1ZrYpHEr5F3i8eq528KHOYA
XBbNZztwY+Kv5xiNaLyWrvnq6XN6K+6BNUeux14BFvgO6Arr0zrxeP65gYY+aUO6
7FH8wt+EYj7CORhjhQkUmHKW9dp5zWnYLksiOgQP1Eo3O10b93stAdhjs1tfZn+m
214tgRtM9X8sQ4diDkCBuAFnynZkGBYgeN69gDxTLMjIICCeRfJAg5Ji3Ms0Xd+h
bVOk2gHardoHh6jc5RaCDYIeiJODJ8aRq8m5qI9Gsvh7yl+Hl3O19gw1znlaSXzZ
fdDLVd8M4Tv6QU/kCm63KZY6jVALbJhO4y63uSZDfMTImu42FE+b/iQ8REGVEHAR
3944oOOwV0HCYVJr5It+D2muRo7a+s2mxQC/c38RkyP3/WJl2WiS8PmWuGnWPiqV
UqD/ucJJhRyeulTYshePPwg/DhOShxPTK3XtKVPcHYdocB6Zz4Ve3cZLRztVqgNa
ov4N5vM0yzjD3Lr17O5EVaeGcl8KHuQQ/dPCX28FL9okaq4BgBIm/p0kkIq0zepH
7RlFzcxXNNYIFwfMprUq1GXxtiQkWyt612inWLJH9oCrDczA37KysLjy7ZTW3GXZ
/OrBF9Hf8xx1Xifg/N04/AioVdwtP5P5SIpvUChB73SXgHt9N8T9vbacfrzCWGSq
7f0AGKH8L10FHNIs5p48IEC/cR48ikzEnP5LJ2sHSZ8xSRZZdS8a2RRtyvK+9g+s
KTkzmvUl4heCiX72yZOulkO9DQ8OKlM7J76bHIY8qVa6o7ZtGvf9mWBcAku+FfKd
2sgRfsw58xx9uH30DsRiDZMSTX4CaoMEZRlwCdt4Hu86o0qXI0x7JkJlb6xPgtNd
oDavo942VeQIfSHp/EYiHvnd1an9cQSJAlefJ5ncMyFonnaXveYUY6A5e+f/xQV5
UaY8oj9gbYu4FAAslT4lnEoKI+Apjx9eptWjXw19tth43T0f6fcAtYu42fNsyFNo
LVHqKKxzlH4M9C8w+1Lh4+sPwKQ0gm9m42ujWofJaK5/IGOitW/mBgIek25dXhmI
RWPechv82oQvmid5R2QhFdJct7rBKaSgHXewTmWhi4lhZJG+0nBHqLSTkgOsacVF
IthZf9Z4SdK+Q3nK4ms7hZFQyM3mjKt2lgEztaJT+Sj5C+byZyhsT0O5sTbDVH3J
NF+nTKCpu5r6dlAkPI41RrMJyoZA2vYIzT44rUMEvxybuRqy12mwJejxi7Gf/V/g
uK2ya8GJwJw/48vEQ3pe4eaQd3yQkR7RFQdtVXyc5Uc4tmXc84FKV/6i76t0XytU
0DJL+IXsJJDqlyW3VGfzNXfLmeu/mEu8ls6vOtSu7APzLWa7mafr4+JklRcRf8iv
Yw4CJ0G1vTDtD7k3vt+/grYMD0JKw9SGuV98mnU84076GdB04uP9kyriinNEvyxk
uqt7ltsYM5vD0nromTJGB3BfYG4hSkqgNhGRr4/b0KBql/mOXDU9ODK9s394rG06
U2PI91c6zAeT2TwP+wLAmyV5GBP0KyBgVQRZNDGo5vQD4vQJjGOp78vGxEetlUrT
FRWKJjdNfSbiIHeNkMxDlnYjywm7ARDA35KhcXTmXq2aAabZe3yzPfJtkrQcmlm/
5bghp2G/s9LJsHBdVfSGDHsvSzl4idYAXEadNM6Xo9KHYKy3ArxlHZsMkAdJafrG
2ne3tKZYDludXA5eMwIgKjWo0tjgU2qEpA1FI3MhAzkfDwW/7bcvuQxxj2XAYqRT
fWbQejm2VCUFLwBACs9HTzINLnu5ppOpr1kiXufjIgr3RuB11MWPHcOTB+nXf6LE
8f5yRlVZO0rev1UfFeImd84jogdoabTlK7LzDs0HUAh4RdanSRL7FpC/jFtfrGgU
zKvccxHfcqgRS4HZQM5carHEaqS7XVgb+yXJCStAakgKMIIsf00t9agtdIIkZpgo
0HmSevDwsDIH6MPd8er0PiiTBdAiUZaxP7AEdHRozYLvVwb9ZhwPfM9o/thyniKV
BmOaf8f75LAx1QbvXNU9B534wK8lMyiZMgn02RqTA6rFMUtV05AvRb2I3oxEhhbh
gBvxtqtDn7s9SPKe46l/gmzhJ6zZ3Qe9PKa/lARLuTQozDRMKhSmHn32qfdLBO8E
X+FEoWWkb1Mqc60q11bQzCQwuDoB2a++wjJNqm+IP7BU0YcmY+WMDmVJNwxcoA/l
CdYqRfiM8U8Vh6LKKcf4PGT65D4/V42uC5U5Gsnrc2WOSw48l9Ktk8XRXUNcz0kY
8WhDyVOTGkBW70mit49cbtMGW7v1FEmlOgIs2W6tuObt8MS49T7s1i8wObeadYLf
r4TaHFxHQgu5nK5b+TseBQStETe/rnHgCkqnpI7IEdtsd1vlvidCieq5hF4brg0M
esxIqqkJMfJ+ibKk5ktRCN6qseUihdq4KRfGy3JWmz9j6XTRHlsnDw68kxN+XMM2
Sg0WVR/yo4G/+uxVYmFXqxXlJvJUtmbRsOcX28eR9Nkj2VXsqP6+Nl5TmXE1oI8I
4WJBZIWs4x6Hv4lrR4AJQFx1LyDwzKQJ4IVOOZo+KmSDFwQKtm8/3ubFBxzdnphs
L3hJBaom+CXxZyoF0JE1Ef3KgxPR0+Vtehx3XcZp/G64yUh4dOc5dfM2SSYfVMei
GtClcPMVpsA161+BrdSiAhQKCfBQ0MjGLw1sbIQCgkCTlbJzCcKAW1RIW0qLQa8g
avLFl/COcVxcUVGUngKeVBw7Shu9EpRQg4hVxo1oPkyjddxrRZxMzG2fXsgwserg
4GS0Y6ieSwqdH6a7vKzcRqZY9P7K+LAClL1zhu6MvUh7H4idBF/HdY2BlFTXnIgh
0wgB5JGo87q3IwgVDxdcWYC16UMJVdsvnzaLKVdahdS+LlD1Ei/OiIqrKd9GXKjy
mySWG+tbxyu6L0ZegUXSX0UHUhhj7e5LNhgIMzVpB4gtn3DGypYPlc+WSTV2kOCq
dX17w0R/A1+8/MVQF2b8WMglaFGHTm8IIzU/GRO3GjzzNrjhqrVSx4YnhOHzkOUc
88ukFayVMv7+P3rd8472sOpmR6ojMPBUP8tyIs+gAgLjUvGN2TQWwOIQZx1yhlPS
yfnbj1xqUntDHdZGx9dGE0etFR3ILnAYXz/LCpqmVNLMLuGh/z1YhXtqwGkglwzH
zEDvczuZ8TkhBlG8ZNJ0HyVP1+oE6iCDn/A6Afka+OJhvTC0FHtbkarX+hxijf7P
3paLcxhdPcgNmE7d6tCVimskkcX3yAag+rio8UR02EeRi2qihm9/Su8VPG7Q+/xV
H4J9/sDXGp4dOqitT+jTQhYVi3QeIGVJhM8HVf4V4TH3w4QSKa9HtNLMfdwKsPdd
LV+DYgcn8DbkLdX8DPReuR+IXbqzu0MC4FpHaRhCg0SlGDg/clsiMXGTayQD0fNT
RVolv6ehv6aerrurLxyhy58DuoxEfm4k2QnNAHw5nOE7xP4VhY4J/+qAouwxjElc
FmQsu6sai8rIPwRwFA/j0LDPnN9WGstp105k3EHGkj7MNmSqD3iq3+OvooU0eQLq
gpBIE/Lc48ndxfRRVAg4jZKO9ZDZ6A8wMutbXYe3n4Q1eTAFbomgSTRU7p676l9s
VQufvqFN4RpcY3v9Hmg8aCDHbHtRbYI7limE832oAWsLrjv470vkwTfV2bu1B1dx
Z+2/K1eJOhNSNsULfZ2k5BlTwaK2Fei1lXE5GZ7rSIqJjaRp1fqCDGpBI1wgOvZT
Sj2fEGCRPBjt6vtzP+JGIpewGbjJvyOSJ1BZxOOtAeMDXoz4mCQ75MRo/CYoandx
KkFdkyaYMu060UDBp1979uuWRBIzpBpP2+OTUgphk/Xe6hXaFT3jhaLT+l2HGeoV
6+yxIIzMq3j7K8Grwn8cIa6+LVFG/TztXlP755notpcRO4KuIPRnkLLbomWNs+Vn
AiMykSM3TSPHFD/h/Yj97qne2kqiE/qjQqQl6KwzKMIgth1zXl6JRKwAqTLGmsn2
zMxxOFBXWm11xhpscvuLJeyS7Kc9orCkVV3O3FpAo87+qus+5b3bPHuUsFkWBha4
jfc9Hs1eXxQ7aBDGFQafaGpWLgAeihGMNh8IBCk2WfOJiODzsZXF+mmhd5tdmhsv
4+hQBlLP+bz70S/s8hivIA7Viruhqv/6chyqJg+oJPsyrHOyC40vJMsjMdmHcxl7
unPcXy2ZhVYTM0wwIXn2HvXAzBbZUwt70aSZNGF0l6pfIx6MlRvBSS/9fYpd/qeM
Xd58GWsEjjDG59l0HxWZU7n/ndruQV3BMwDsLvHsPJqp9SzNYWHo6INNABHGlq2j
BhJJHT1ZN4jhbfnvgiFgPwOPGsUBioyxyr5lEHGC5E4Tmmw8DTvswxxpxSyhNryU
ZwZrT+NPhi0HG/gLGqxaIluD/7gq2J5P65QNWEU8RWtFe7haXO4mQT3F+MqZYgFs
Xd/mUqcpPxeF+AOyYSIxWP6hr/CYwIoTkoUrg99A3923w6Pi5CPQvKylm72kYEri
JagnpSji1NeQ5xGeYiyt3dlpa39Flx8C8L5jCD4rVvMeL9ckgpl5YNsmfyPmfxiD
E1FHk1FmKaqFhoqallhRHmYMBctOGDENcfW4sjJZmQBE/vrWLLqdjLIkSkLbrg1H
Q2PG22wBG+8dMh2Gc9A5V6zI1kDjVw4bWElRCP3xXiqWjCrTRzpOkbq9jVUovBym
LwcsLe5LksZwYYXEzVUmkEM/11eisXD1gYrhBPth5MO4o514zTb31a6WwOO6yHMK
VzsV4EnePwIm2uVUhOBAwvqialXCZAvuaOZuQr4B0Gt5/dIEARuP4DdKHSqldphV
Jz/ktp6tsn63xkpVfA1+39u9DVK5qIf9agd90fnMR6DOAT+/4IFpPxK75L/XiQgt
UNzbWdQzw6pgkLxaP8+tYnQOif1QKo8uimx1WOA0CCOOiOEzak5yNtqgfPFvP21q
M4kJjV5MBwsv0MuTkuc7T0XhWB+FT9UHo74oMt/vQtr/SPPK1kB1nBLLaEBA3kdj
7w7zhTG2iqW3/eDNTbYTnADbZnKzaLBRdy0o7Vg50QOdFi8MSckYGNYrB6a+7LEs
L4DdasVirhGuTWWZhJGXGGPTnfxvGn+d/DS0fPtKunxQcF9Qd6CZ4tx6gQLUywqb
G/uYI7cy4LbDsMiJTOeCzxXvgWgl6HlbqEw1JQ9MBMb8Xyd8YV9CEDL594fB1RvY
CAT6wz2TkIpUnMiZ0jHutSZ2MBC8GDkji/yTke75ohrbUDIDt3CbF9tt6t8kgnNL
knTyVwwbJeeGkNLj2Tt6aHLzzMciqo3jotxn6rsuEcamt58WeT7Vavbu/znvyozF
lkP4Qo7G/8Y4Nys1DJ1K7TPVurvF66WeARIDebAE0aD/K4cJOidD0zlrNOmMAN0V
pWyWumChJdXwbnvL9cC8JgsW5tf0ZYNLlGz0JcVNu/riYCnIFCKD0ghwec5hHu7j
ocdcGNTa3yfXnqzb4jYrW+mlBvk9zu984FGNz1otcqKn9nCRGxKVknQ3wMB7JcgB
wCiAHlCrA4jBU9Z+s7i0ZmZq/Tgeecsuk1WFUF4Uaadkg5n/tiqYK9mhcqyq8cb6
bv0L/KqjKxLpzcXp3cqebQn7q3R3XVSlGKc8evy3wQZv5Bg4q661YR6gkXIMvf/o
biNH/6c+AEJNAoAtM2QDrHU7Zc+4qmqJWNrC8BchhRgg1ZCIGw6dQfEeFLvfltQN
fnSCeIm7LdIfD28QJLILVazTzQXaXHNBg5rsSZjMQwcM6IB+qVc109VSjxivPfkr
faAHEZwzEKkq296kbssp+1lrN7wcz1KFMUuDlcodrxzTK/rdf5HeMO4egYraY8Is
ZTMqH4dKvKVwYKI33Lcfp1IFWW9j21XYnDrGwYH/NdDbYkxR6xP9WMpZ2MJDB399
t0Uz8+yp0ZOmwPaGA+5St+IgAj5mQv+HCPzprNDwDFgzu5FkD6aQx6i8iuyi59+J
2k2lCwkAbZLKMEhBHaSVsDCdU/f6MyVE1BgV/kU+SITPhqniCl4FxUfJMJH2U3ya
lNwh9cqvBJGnvitfa4Dn8rEAKYzj48a9mP0OYubz08dJrwWjPmc3GUgdsVWYP2+7
cAHiYksmhSzMHChudGSTyBTo9R6gC/AK3FXPgCv4RoDG7xjRsznAL3kn9IHNbNwA
uJWN7Mv50VVUnhUBvI/Ql82gXtCEaeYQpsjte0juPhZzg/KY827xhyhbN/Byp2hY
uthWB6b9HZpMBIKNZ2ZLNLeFhaFgnypp29bba+MNEI3AfpkzjAt6IBxKTK7JxQwM
XAsFooJNBYB4MNIhN97HpcuwaVBF80LRydHv9gqkuydSBPAYBrSAGHggWE2sjhNs
HScjicqfZs7Rx+cMzzw5xhrD7I8bnPFJUSvWCBW2K5Ac151MJG64spDqT8o2umOr
eHRoX33m74AMVoHkB+jm4pZ1Ta6GbfVcwd8O5h2ul5MI8CNqW5aJrrE/cxVS2XKN
036h2Y4BRkzexnL/KCV5yjjeTRnX9wgtTnTalJHtS6bTtT0+HCljX6gSv08QuURr
U8ruIJ2+MUtmuCvpyIhVy+1Vb+3OTeJB8BM4FJWT9hAdzYskiRwkS4ZI9a92ufRf
qhNMvAx9bKYOBNzfKI5I2hb9NxwfCLhRAeGTOOMWJNFEtambjTxdFIqJYWrYKeGV
/T1opRyasGWs5oYpio8o1zgQH3Qt9wC3hCuhkmxIoDyV64mZcHUSDzpRAF1F5hnz
AZfUKUe7QZDRUNrh9rZYTdEq93AkjSukNeQ6sczRaHDrPjJpFex5cT/Q4qgLKwMZ
H9uAs4n+GtEMg+g+17TGtg0gXItPMemHIF2HaqZJJQs5s+OIP5gvTvHIn7NXxyyu
Selo7rXFQiHIRUeCoUD8sAayutFFm6Wd3GKIaoe1FJb28y9lp3tM8B73UPmVj2rP
Yh2zqSYMqb34mRLr7w+oV/zHJWdVnwVWnoHgjzMU3yzpIXO/x5rmgTXwqNDphRp6
3T7EQad15POD5TtWX6+8XOun+r1H5w/cRodVgGl72USUHjkVHVzFbAt/gffIS1gr
Un4TZBbgjZm+9MP08aAyoNDCE/iBbnlL+Fog95gSt12d6tuwasLv6QeYSk/Z8Z2r
FsDWn2Ogn1KyBar9ijbnq53xnnPr8OcsFKAUALBH4E1kiH+V+82IlIevVrQfRj0N
fG59SC6FaPWwrO68ImxRG3A6TlEDxURd4ly4GJcR36FMpCRtEymJS3gqz0aIrjlb
fHA5NID0QqAw3Ae3PdT6ltxgajtCSYGZSdeESft5gbUy0RpXlk0ORRxlV95P1Ixj
a9z2UAv01xAtzoDSEcJOzbG9JgJzsoQahdxzVPILDjODYPvUgyo3GGBqCMrpj7+S
d+JYXnnvXkdnmpuAPG5UKIyWJhaGk1erfGG8wpmoJE13Dh0zsJrmlYgzmYVuOpg/
nsw7HJ4WjF4WPNkh7d8BD/dAq5n2mqzDVWAm9eUJ/Tcx+XVofM7vdMNYKAL4qF8W
iuRO2LLIFf/cRsWhf1YbWDA+DCcHImMhNeTREJeiuHA6wrgaJKDh/Lrh03ZmMUkq
KsHIVLQz5PpK135BG+jvf8L609I5O/RW1D8aWFx99/PhzQoz7iClhBgf7qJBlc8W
ibmbLMqWWqSjRhBkSX9uA3/COjfEXSWCoV8hNwi6+3YitLOGy4xP292ESV79DfCY
IbM1scunym85wIVktCtPVu8FHSp8ZPNyx9JK3J8L1Udc2sVWC0u3R8z+ieUv0PCX
7VV2iXB7fsyBndj/nmEBpvv2ebmiw2iMywRniDzYjUJODR9FI10icI+xuemugkjE
AWZr+hbFKUQqLQvxzKhDw73RfQ4yVVsHU7nerxNmF6UVFNoxPVVOx4dnq2usfwFg
mh06HiZ2WngFCT08vqZelE8IfNrYlgsTofYbcv2y48F80IwpMUV3Q8GHsJ8afoyU
FKAR8n/QdibyIF/tzW1px+OJob0p7Ens5NR8lrzh6QiYhI9+yljTRqheLSOMBNCP
ot7tFm5R0fwBzGcuk9wHAs0WL8WPXiw0o8KpgI5sUtD25OlplQsF5rqy46ypTuqw
gkz6fwqSP1+QNNIhxpR7qCMRO6qTNm06UAn2cBQU/3RNcbsNY9q9nKiJbLaeYIhd
lfZ37gN5LHXZzKPpSJJUePfuvQpcv61ZtDXlcr9VG5utobtwFesexBHgRgu5X8lW
SX/+S391aJ7ygl3Y94CJirfD+6jx2aGyZuN83NCpwemr+pzWh09T4/Fgx5AKUGCE
r9aMHDe9TGqe3bzmHnikKZ3x1rEIwPr9Erq/OwLjJiKSo/g03O0FsrYywHDfCG99
QZebiZPywVL2jE2peT1axKtdX5csKQxDdXM61xCh3Dr1fVKAdDBdbZKg/FUjiy6L
zN5mC6YodZToP2bz9+wUr09N433JhnAWT6iSV/dFaGHK9gdB/kNStLDUnYszpQyQ
YyqOi7VUkmmmfMeD5TeL7XSVo9yh6ir6wmz8hLmcRaDcsZwzDliP4C08Jw8fsSt7
jyMpc8G9GftEVxHYFz1DnsnPko6GghIxKghwXO6IvDlxMzHJ9U2uP7BlJJI6nScw
6/Y7XJWfjJsl0gUWRzA6CmfYN8/ZB8f0xkB9R8nhWrtSJK7db6g1kIYsEzHT5QDQ
cDB7eLC8IydL8WYKLAjOumB0FIifObgB6juOJmFpuTgXs999Rvd8EXJcXcH5E8RC
BAJ5ZmYbpJtu2L0Nh6KUfuEAneRmehqsJvaKD+E6VTJb32rwosMwSNZqC4Tc7hkO
sEQxPknGgTuVidwK9WmUq7DWyVWKweip+LIxcTVJDjr68xRfyGvKaQLVyrZj5kyP
5BLeBnrbN12haFjyhkhuWLAZaKPS35hHgV0gPcKxAew6KvY4d1kh8pV14ZyBzA7R
13RolTRjexDKX6VKrAWs9z6kIbMTJMQqkWxq1aLofFEVx1cEwVdpLMBdrBt5b20V
/o2cYJPzg7nyS1nHuSHWQmbCiJGVR7Pr8rwZPRJ+XGu+RmSozvROK7vfeAB6+Wae
NyDmPqC7VVYpdnbmR8IBNyaoSoRcXdmerPUVyS17bN+5o/yg2GLq0zBoNaSVXbPf
nO98N7jf4VjOzYjLEUOxrfAadYbZu0A8kOmmHKtNfkeKNTO00sfenMOOPGhrq1Ci
oaNQRMQ9Uwh7rBwphMZRsxgfw6iLJEUaYLlFGX/I/g8MjBSyQF8holzywhD2Jd3R
bvW3Bt4pKYe/lOCrXtAqei5Zu8Es9BZIrNyVZudakrBSTqBOSMy5ke1DSMeekGnx
qsUN3yJ/J3JwzJXowbVDI76faC8vhgWPqnEsbGRRHaZ9opm53XBDesTiXBjenFRa
rY49/McNAtq+BzqexJJnY/Op75OvBCr2DmzTIcmAYIYBPdnO0DQ9IOE0d6JiNqtE
HhS8FYs7gO2St2eNYjivjUPksimgaiNLbP2RFMhoVQMB+tu/WwimXq+DKp+mRPah
FhTlFb++8xGVMu/bo8NbYQ2EJG95Qc+JXMIVzi0mFQegGi6UxQLyT54jg10W6UnD
Fly/jGcXvBFdiEIrIfmTC0V6SwaTa7J7BQdZK+vySFqiDAMDocWvwu8kU40cM6Jq
HdimkT1ixvkQxdWbckCNeepf7Ayn+BINZv0nYH27Ezt2+TzqP3o9Z9mAuiy8rxqY
0yMzQDh+4UoNCjTfGH7mdyigz5ZG3Vb/SQ9fwaVWW2VQaaXhwyIPA+v1+ywf8/oQ
y7PDtq3HAcfey6Y3UHjL7hwxfkgDXQRqbodKDUEHQqz/sww/VqFqRVNCqmv/q9JR
V41/UK+7UghVWRKCWJQf5iAurGIOCBN9FIb63/G6OqJITe0PK6xabCaZCcDLjK/4
lu4FO0qR07IdkXvQdIHYInjgays680QxwJxxM3AEF55m8YBrzk5PauueZ1dmbiqh
PdfyJsTXFrLv20bD40v1HG2L910mFzsaxYmfy7p+LuCZypledmUmcvDkK8EOMiO1
QVsTviCpk4XldW5EQKzSsP5Ih6TDBYPPavyOebc2OmDOkG8Mb4uXhOKsQFlSjO8t
xj35HXbAPdMnd0KNOKi19z7fRnLyoj9TZbeRrFLmmb/qlVhZFewQGjJrddeZ9HWB
R475b/hywxXzUdUyRTt1uY90mmdqhJ/bzBxdzQYbFW4MW9I16bVmyeJjzJYQERpf
3Mo6OJpNTuB3MZLHvoFVQuMON8rZNRscLiGKB+eV/COlsoP8t2hZIJJbEc/rcCpz
WrskyR3PHLzrTrhuY0ZU6D4tYFMxskmtkdQdhdaozK4PN18IcgaLWr+F41ZzfiJP
IndKn6F0SfnKBghRjgU1sJu0pIbC+kakRSOnP2Y6u3N5RaFijQbGA185ZR4OT6gc
Nia7dNwck9qwWxm76hTll7GlI50b3QAHx+KCR4gEHdG+Tps2zC0F8HkSAhNDttnp
2WvyY4PSfHRt7f0ctvLGHeXFQYoT881iBuzT9UydpR5v0oecYBstFQSKi3xFfgrC
MjSuyaH6FSt2mSMR3fRcBgMqeQCa+bkhACzi9VxDbCmmvJo+Tg/AZgTtWfooD+zB
bQCHTsHH3fxpQOVnQ8ASNa5F5jVGDWgGBR6R18wrxwu/Z4YmH4p0UK28gVPJ3y85
HPJ1q4y8FUehV41A8jEJ43wCc1HMW0HeoqfAXdKHxCVKb2JesImF2ir+vRe9gO3H
aiKh/oc40aDDg4mRtH3U4p4JTfByWCIJYoU5GgZBPSVUEUH+a2e6OgFjOuo3KnSv
7gMAqKtkuU8nM/xMB8clXboPf8dH22G2Jz0SZy44HuDUTg1CVgFt4cxttDDe6n8g
o3PT6/cJnAQqQI7RHQDR64iRtNJVeiJUZOADUcKc54Lq7PuQFNdIAt6o8XsGqmEw
HPS489xXWHoGdAtI80uqdH9FCqftYC/kFjB/15sFi6WsENUMU1Nx408/unEcUaTb
s2J/fCRmYmzFA9glf064zivxW5E6bq79ouvoZfJAE4yW0ETxfQPR2Tm/kDYHF+sK
GoGInAkeXraQLqfbFdM+EtD27ySbxs0ZZoINPbkx1YZYG8t5a/cwHpE695uAX8rT
mBtlKQ+rYADFLkAfbHlUMQx3ySdPDrh/M/LyzgafP5SQVHVRIMRmkMfzhS874SuH
pVr8PxGqitHZ6UG31Ev1kZIx9jHxBia5xABElq0D795X/4rcPSWf3PoQTZ203WKV
nZpqRnqoTmuEBtV3jTT1LlXztIYuA6O+wsP65a5+bwQciq6WuiHKszryG/0DNYHB
jXSJDp2F4j64v2w4rF7hZm77SnxzfU9wCOU9qsNKb3q7wsjEDA3qrikwt7WpuJfA
ISrd+2xuy9dJzhAj25n9wUlV95Cr0HSvS0s+x3dIcocwBu44GKOFG6644Z/RckTL
e/nbHpQI31JhUberYg3v8+R7KNiYZ1SVlRGo3YYmbeUCB1juLXd/bCGfMpGofiTk
0vpeZvTM4xuAU57ChkZvOHjAuJ164EqyNBmTzmsQt/YjvYzBZKDnRMLUDkF7uocJ
qjjPO1RfZ9GeVFk31GkezMH7jR5eceM9o2PDhHxPwLt18WwOz0PeurrE5XMMCWtT
nr/RGzQ8TjegllKVPsELqQUVwQO7Vpsh+miNgLGS+ryZXNFipVbR3KDLCLmwvpBN
TSj4UxQnjy5CiBnc2yvhZV2SbCL1bn0BmNalZjp926EH3/4tULeheNDr+zJelXWO
UzjL5uQMgkiOLzhdvi9H3gC054ZzaRb4tdpFZdW/aGA2RPmJs5e/CV6Jmx2huugu
j7bCX1fqfAaTPhEGHVIywrIsBgNhoL96CNaQFe1wGN1mIEz0a+aRlMhKBXl7EFOo
x75UrFalMiGFDv6H8iHvY6DIK1T2UW4gazxJcxEUPD3bhT6igrHf1l4Qa+j6AlWd
JQh2mly/kywcW4JSJUq3OLwW0EYxxkRXAQFv0bLW/QL0H2XUt03M/8CiRnzdv2IZ
vfBCQwiUAUFVrTaMgO2GEF76JcoMZc5v/kgM5EBcwpzH8ehXASXHIxYiep/e8Ubw
bQeZd75OnYXPZGXbvRWY3Me97Ti9zTmxz/pjCOqJtC8Hn/MOtjx0XICZ+e0B4AxJ
3blOISCrOz8O9hVbbvprvUyEveNT8yyvS+qwGEA2NSHCU8tJtx+1/fpoOcvjTO6m
b9kO42zwC8MDNlWQ16HfqqMrU0NvukYn+2NmnjhEPPRgGDNHUh6kLBH3Ms7o13tX
F9FC6PPk/poRY1phHQmoFhRKrRYalwp5uYdD8WVsxuXo/iz8cUPm9IdZ5Pp/FyVt
FlY/J/SR4aHXrPa3SB0jegDPSmQlX03k5nUm2iOaaUMd8NOefqyFP6VgBKDQKeY/
NUiN78SOhFmpImNQQ2iC2sTTThgkw1oXrQgc5fx29mJKM3bY+ak3sODtfviNxDnu
NeWfpcuaTMPFJgjiE3lKt/QscHDXp5VIuyHYPyz1QpRWuDOpBzY7I1oyaFKJDSm+
6gwYpMw0zTlOPZxQPq42IvYc/k7nXd5IXjoTWBoOUopWWR+ZwyXvF+qBzBp/md4h
1/FlrnE7Akd8Zv5hBPsxD5Fp4yeY60dnseElyWo81PAYokVqLzJYUzbjfIxlaFpt
tdTmGVP6IJd+gLfK43FqNRQxGveNtjcA1rtPnNLWNKQgO5x9SkrvSiE1Qccr59fZ
/uNNtxi+fXpUzxnHARhTacXeAkK8qz4+ZN1gJCu/O1sDi1Xyb74PlgXQxIP526g5
ET275+/nyb946LpZKohGO/Xwnbax1x9oT2FO4EcPlnkU2bXwOJfBgbh35ITGA3e/
Cj+Ko/gBZqZqIWmQUIN8gRz9yso/vL6WHtuPCnZCTOYdhfKaHTQm3BZryU7zoGqt
vHTDlGnVYiEIxiZkHHEMTXrjRfVqI40e07s3yJbC9YbD/bqqUIp9Zpu1RqtABNNA
nngWaWdHdOoo7sX8rrVMiLIxeSLHz/l5913n41+QkYC6tcNZ39iCOQwF0FtImMdb
i4WCPUIa39h/yxqc30jYgYbLeqpY6CzhXYnd5uIFh2S/OdAT2+G/99aOVG/SAHF5
+f/BHsVj+xf8acoQdI5bto9Au56pwcHoFrtCX3HamlUk4OyyW6pcdKRxP7RitGNg
DDO4IrCrR+M1Mg5FMDJ4uiuS9gjIdFtJsvlKjKJv9S5ObsXbuX89sanQVmXMzQfv
0emO9Tp5fFQ8hoY3Ue4lUse/lTw8hdHKnGd48AnSpClUBbREbAP0vmD/Uo6ewiUn
xT0EdoOswogFwfO1KdG4YeToR8rvO3/cmqdUdGoLiAVy404j73pOtknXmrqQ0fDh
H5DDburJRE/o3kUk80kYzbTORn/zCRIVkHkCphvWgnQH0nyvCqNOaTQ1068NMiaX
TAI3QuSrqn+z50QCffStd/42uXCIjQlquh+MSdm6Cg23tLR/xsfGw1sHZddm+Pna
lPKM13cJh/PfCXJFB8pgQqtTblPzw6f1/t+wveJRanJFV5O7suSvImKCD4GFOXHu
DVpOCuRG+/UDGBtqemwr+PDRaNmDSjbV9OPPNbb7EZPx4Q/fmNREsL5y3ay867pU
JofZX9S48RdqrukQOkbdKlbpDU8GrMryTTx/0rlKUoiW+8++VQLjMpw7Sy0Dp5Xo
DFite6vWBKfFjwRr7sO6NR+R2qowFFdnkBlWSwH5G++Xsg4rk7+6xxu3IN63+NHq
KgswNXLauiJwLouZFG4dCXGr9764d+1OqjTOKfJc85qxlK2aCnqNIFA3xkMNXWe+
ZXoUtYgStxCs1oTmuHT0S5fZu/ISsLebaPyKptbUox0KYf1LhQLNToT1RUwLVQtr
iEpK3qw3ljGZnXHcu+nbfWC/aPccM7VnGKYl9BrwpR6Ngk1ggdkNi0tnjYQMX7b8
yP7qyF30dm7Jj6mkhc7r1inSDqpKhWphybED5cUea2vlMcfO/a/di7bBvKGzwPOE
F4q7f3chch7YvxETc0aJ93pmykVjsigFB3GVLik6gNTSPrTRIy03/jllnXvNFTlo
Er4eMiBpeD16KSJOTtpqgOinXZeGD+DqsNzVSVbDHoHjvFaXef3ka6ewHmcyg/Qu
SIPHMTysLCuvUu7vRUcT63oMZ2t6+Kt4q5IC1aG6FUg/M/jVKi0aqb2orxQ1gLit
oxzTh6/84oOV0SCn9D6N17IIxtD7H8sDrjz8hIklEUy0uxlbluyiunXPNg9Yg3Sg
P/lL5scmXg6BtpsOk/zzvfZfu++aKKD3zII4/F5K6ZmiXlg7ZeF0y4LM9XqkBBH+
rT3Qtcm1slkjkTW/B+CxibecC8uV0TyvCTA5kZkkP5JOdy/uaEEn8JLLyo6JE745
Vkd+TnNZ4MV2pJ0OsMfJMfjXPIPFrVsCrtZQ4Vm/WkziEKE7+ov0aR9HFFTIfNoR
R45PE0IS2Jr6B07gVX6xmgQPh9E0vCj7iJg9yuskdVdqqEgYfhpGYdApMBrbaIQy
eQ+JULUSgLLWE92YmQs0IaoPzH0KYmrBmis0Xas8I36Ly1f0SiWptC+2F0O/7bL0
g65/P8LMJDzCA/2XcYEsvLz2ydadG/n5e5r5dg6TX3rPVLvlf3iHMYpu3xCOz2lz
zrGL9ub7g39QUbOuz0UGNeGzfCBGV50tuYU5BKKlmTPaLCvAQzYinXQX4xWTEYsW
EwAzYI3yuZqOtzGqjqBza6Aih6K2iD374NJBsXEuix2fl8U98pmdFDYF+sXFxJ+D
H6ViQTBQ6l8vugUR33j2Yt2Fgo5zSnmc3uT/IFBY+kA9VYYxEE4NN7gTiKhGDAQU
/GeWpLAI+RgELD+EDcqqEOxSEkCNDL01ROC2AJbalzQ+BGsGho6uSQgORyYwaYcG
1GMDYImjN0fHSCQP0poTu9W8GBPJRsEI05VerU4LkhApRvm1R7QVHKV/GLccjBxJ
/89wdfnfWM+GwAdA45COnTDrlr1m+59sVHGYMcM+eKByGpV8KW8/bLQ0cQeDIx0T
WvAXmmPiTjaDD1qh4+3ZdcgStimawPLUzSnZp3bOHdU44GomY7mLJoaHfYVApTH3
3fx4U8EGx741FIQTCZ4Wrf7gXpu9dQmynNyYkcKo3m4kMRaZyOZwXM4pkTNRg1UF
v8wVkIfjvQ5kNYA6WU2kqmARwOsO+Ci1tBv1aNJSwckMRTa28Tofe0oT8x/qgr9M
Zlep48gUFzl/PI/ZNl92y7nwlavCmd/MB1B22nmyX5Mj5fVt6L9nYTRl93Wdq5LQ
5YJgIOBXonIxE9QiWeR/WsZgTxdyLilPPztXyKM9p/Yt2nGXdu/lCa9EYgPz0s4J
0fTfcb+sMTDSh0C8y9kBQvGuz2BAMlDs1kZ+kdTjM/X5j2M+PfbSiEo3vR5NvB8Y
MqmIy4Zl1826J36UirHgM6w+PFlT8nwk7wSKh3KKtuSrdcMcySiV4dx51i1xtGbE
333Ecojdo/EYwIidCi8AavlAk+T4XwyxPSDEtZPHywEgMpO0pA2fn9tNnCyamLND
8EeeHnuMN/lRHu8vZcblLZ+cStdVWvaR5uTsEj2+oLOJpG40f/Y80H3MbnI/kfGo
G8ABUQzcWo7g04aXRuO5B7oYoBNduDm8qlFZYhhF3MOAN/CbTBf5JToQBLOXfV8d
ND62eQAwUMNHtOYUqJi9qk/4py/JENtlQXzcPhZBD6TEr/mz0vTFdyo6JUBTzjRU
mCQXnfv2Wki0z/Nf2DK474Vi9unmDCqF5Ok556wCHBtPZ9TnBSO/qgRDUkOXntd/
puw9X0FpSMi7fP5ckMU6g3RWvGQ1ulsLNHI8L4Rg6U9Nx+2JDUVQwP4tFeacV8Ct
j0MbtCmWH+W81Aoj1DCQ70reyTGwHGM7Qb+Xo19F1ZRzvVR6u1HN1p+eIYcj2Pz3
0ovxXh9okupE/SWntKq0uEoDvfES74Gut3jP3CZVM006RgzHvkDoQuaJXv52TXZO
m4PDCy42MNeuIQSmsYRGr0VckmMtnsuJAJ9h1jrbYe+dcYx2SHX9RSaBGOSYHJq0
krYYYMLtgfqTOne/NjCL/onsdnNhf319a4l8p8+n+8vb86ZgmD9b5boXJsT1T/1t
oZYxfDtQgI/99dLLmxgZjx657C1GP9qEbq2dV3wS6IybBQK2zhmgcSblkLygWOlR
JLeCwBtoG7rNgG6Hqggt27vxIUt3O75+DulgB8zfACYQ8kF9lZ8PlJc26wFM/62X
2odhTrhIWjPESGZD4Q5829VYCd13ENPCyPgsAXtyNpkr8quU0MfCT1t5/VieLdfh
xaLyOHhOJPBFoGLtiDG3pB41UuoFgwvs3c9zMvz2AjnyFIVVY1paAYWfC9wKACQ8
a+3OqPDFUkiIBIheoGt3efLGbpRUPDeOxIAiaseh7jbQqcmfFR3T2xZyrA6nXUHW
Qtk46EJ8SH3KHz76A2cNuY38AzlCCm6tRO2+q1M8FsmXJG47p9U5JW3fml1/UL9F
68OOvaZpgazB5gRJ9pO8voemOOdLrNiZmnd/RfQUFWAQq1mEEkId88iwAj+Um3P5
ykECgUGN+sKvVBNNIJXjR6Xt2DPp/QE8sRKpyd4LS1KG5Jdq//6gf0GtstubVhGk
6eWn4fK7ziSlFZx+ptnC0L5Vr98VxJEwtHJlm4R8RvOZGHW+7BM4ZqIN4Zpc//TU
QduykOE/74umP/TSc4rzSwoSqlWGqsoiIZzQcIvq//OiQkQq0kZZMqelVr8Qst5e
naO3gUh4mZzqgzujkQlw0R/q2OtvrMhHmMowr52BX/yvPq2SgiWhY3/ZIo8edjNO
FMrpPgOeFoi15lErbNNoVxFeJmSN8XT6G7r9UPcVY+sAEWTJXZ9PnNjC+W3Hgjeu
IxiO4CN8SM+CjS23Na6RK7AayGwRji4Sdv96w/KNJvqz7KR4gHtWXsMnY3niAvlC
JcJJ3rSkDIApUiDBivTIpnwH96Ix1CFdkdn3ydlQTRtfYYK3NjDnGFFZelbgegFC
KA1Jz22QPZ0NUitzJqcqXX9ML4pR7h2bk0I0rYnt4Sp1nuNfdKFLmVs5zZrD6f3u
S2nZN9Jircs0eSH+uMrIALcaE11RvvovDVMG6iovh0g+aUK9Fzs9afazakCZJkiB
RGQMS3TnwtLNod0f5cVlVJ4ZPRg56UM5bCeF8mJzp6ivkaPjkdR/tTc2EWvIWFJj
uFtk2EeuNiM2z+jHik5K2A+0qjO46iiKmpMm7kl29r2psphewpQsQ7aUbfffsYCi
3nrnVweCdw878spTrYCH2fNYx81zDpeyGX2km3rzRZWer7utyp+g2i4NdsdVOY3e
Ti7ikm1ut6F4+0f+jdyl/mOa/L5u/di9j0U981zljpvn6DCvyzuDTlyBhjFkhR6I
3ZR06C2kfiKHSunX9nmL5c1CEyNqxAbifGb0QYRSJamSFaJxap7gSszFR6Cx8hjq
cLNOoK0iecK7YEVU2brC+WevB9CRTv3Dc1f9rQ/rDJvOFkXLjXDa3AWrF+uDLQ2v
tQBzi1WBxCIIINUGAPz5v1UWlrohxEVwH485n86cGg2tRyXlMQkU3gu9+hUhJEk1
s6oIV79/8Wy84dReP4qclugRmDh2G//84uJ2uycg3ydNJPzBQRJiBBxslrpE5J7n
WRqOr4c9k+U05uHJJYpgdrLPul7RSBHY9Tyt5maJAkzanXQBCJ1kqfz8oiIE7+FD
4jl8Mf6ngVebknEPbTtqw/fLzYarhC9+Jfvyd1SP9K/D816fe0LZApW34NIWs5Y7
oNf6AjjVeawEqtz6KARBTURyMXcc3e4Y3AWIlclSmcfTnx0NI8rZLLO8b2uweYNc
0IE0ESWj6y+jcGK9lEsI/sOU1VrJ0VRy/4xD/H8gYnYYJwNtoZBBiBdzSRqSiE83
MKWGxeBFAh4Udf6ZhBrXnueiNzcfBP4Yh7ZJCAHzfP8pVmWT8nW8YwOgATiGQ1Zk
/XUeLyRWDYtAajLdFT/gn1E8cmbBW2zKxlR/J/SPr6tZYflLCzXGUoPdTVIONNrA
QVjzSZXcq/iwkEiHr1teJbWy3aok1NcQtoxEQ7EnDcDM5MmosqFRapeI8HhMATAy
vIf5XJWEGSZ9E8wohGyYeB++8H6XUB50lzSckn+2PUJx8T11DhM3Qd2PRBwZ7uS5
SdmIwZoS1hFs9dfvfWA+EswY0I2U3+iOMJjuxTrGEveD1XZe8wSotPgd5zpvbu7o
687gr/E1Eve2Gc8vKFkrBze3Zv0mofywJrybGwC8Wrzn3H9YDqmNaYP0c+NCXaaV
9IAYObT8Y0odpEexogGPJEkzYyqSG46OV8HqhgSiVxVUelVEdPhCZS7AxxD21MJU
S9i5GrufVigAjFh+JDc3ua3b7CVuD3Kf2jSmGNxTn2C6AwtJgaeEViRp4flLll6K
8nG1rrXzT5BvKVt03UfaRUgA8VKxJjSUfftc/gjxoPJsXCB961UVH1kkWP+larDy
bqc3LJXyVD8OP29RXarxmW3ephkOOP0lrM9y/j0tJBgALGSMZdJ+FydX8nXo9dlO
ersX1ynuYjndvI8bjsd1QNCi5ABn87kUL73iEqbGxrymB2cQv7NxbOxXLWMCkBdI
FSNdJFlmnQ9Bhd+KOuXUcYIQ1+VynEPabBh052ZTiR7tNeq75xMhJ4MZtuy1ofkm
oh7mkJyJjIiKRHIwyCcxTQp+BeZFh3rS0jHnEWsieOfBNXOunri14nb79tuKn0K7
1jU4ltEyAbO77VKL9krofG+Vr4li/WqHnXoB2J0lMi5qgZb5xxmc3ITjGuNt7V/j
o41B6OwkehX8yxBBaWdMLBFTlReVr9VZAGnnf0w7MOD5nh3z0ST4aHMr5YltmKu3
STd5xwjT26um0zMguVwyNsGn7hxFeDvx5cYRjM38kOz0/oJVpyobfpdMjXUTIrbV
6XU4+am0Fdwg8P+1a4OERpygg4p25Gmj4cPkkCpVvtgKUKedjm8d3WKTbr75bAr8
90edm15E7o3WObbcF66iVFAsF8LNbFTn2kriTKooRGBPLHxVjx4EfeO5z3wlltae
/rxKMM+qiLu4M4NAgwfsORd9XdKJr+ozGVRYfUfOoYQL+8MKQ6I6y7npKJnYYQiG
VpZoYiP2cdoAw2VvNG8BA4jPlzc5aWpLNyvihN4Dy4PqDYhtb3OeITF+0PFznVKL
5ApSa8z9zpLe+qQwGjKhA3V2apmmf5nQQnheofKGy500Aosp00FlnbsSieJ3dyuM
XMAX767QzOA7MgyOObhvpUTKwbSiCV1Bqu44gsYyOp2eh9cB22/MdLF41bJe2YU8
WcNPgl8JXJbXKS4W/HlSp0K4ERm+UsVsN4AgvLOECDft4Fwfeb7WL1Fxg/h+NodW
pRG/gr5crYWBQfmGaN3mjRHhVWwCkYkRYnyn83sAMkN6ZtFZCUI/gObZIS06hgh3
WHaAx+8eCUtm3djEyQhIi2ivBWjmdjRpJDHwChOtyTO6+w7pCzdQ9FADUYPiavgP
KE2JUgjkCjifDO/cTn/N4fG76sL963qLOkflcv5o5zl1cuyF+QtkLxGWzSZkJZIm
gIPR90atNHgFYEuv1pEKbRwgrHwjNSMYy+EQLXdv9tV1IghYhiSBCyfVGs/vu6QQ
QN9wiXkbARxeJF7kzhiprGiduFBHmjmEN50gXUE3iPEue0CM1h3aMNP/SxXeQhTV
OLnDN2CEsBBUqoQSbsO+pQBQUx/yPpTcSCub0NNpJJEe5KqZjZDo2ejn8/BsfrLD
skwsQdGrHSHpVB3jqmZ1QHZgZJ2SAqdDTrRhdE2Ws1NHm4yTEBsoO4TxN1r4D0Y/
I+le1sNcGIGQrSm0qlKsjvYtb+e6kge6Ex8WsueWcdSskP6oA14E8AI/SPkmKeF0
mB2yIfBWikPsUtrFpzEMOSTmrWfKUQ6wigpntsd/2Hlw+AKOvHXNZSr1s0e9XRAk
XZ3eGZZsgyggmE7xmPk7KCR7usPY/r0cSFPW1bh6LDd+UEDRXiwnR3NO5oxY6xHh
J3h4xlhZXd08eVbStbnrXWAJUMdVIUbtPI6pgTucZzydVW+W5mdrTu8chXoVTwne
BANCQU1W/EYPRk8W2QU6pYTCFem7MVWzdxqHSCbRJzTvzjG86p/gZRROEoy/MTQ5
GAxOLOq12wVt6+GfWv//6SxPtkO75b8+vRb3OabDQLY7kena4vbQ6Hm4WFmg4vFy
hM/5OpY6dRJmWXxpAAG6P7JijBzSlSC5np9dwGqCxzR6eF9UFizVXdqlCX5t/Ck4
gLtIVXrXF2dX0gwuuz6jaDl4oGMWerA3VSAKOdvLa2scAuwhAofVo4EdC3sxHcFp
MU7w0tMqeXqi9pT0tZ6l7jDVjfEE4rt4jrDwiLngaB00kefqBG0Nq4dUcbaeFoC5
GPqu5G/zK7fHPQrm3fOoASzXCZRmEe32joDucNO1JBxR75ZVbo+UHsQ+TaHcnXOY
/uXows+At25yf8R4LsvsfTbeKISuDEmveG+y7iK2+9BwLSyfmPAieZN8z0Bn8BQs
B/l4JjEV7eH9hz+qcs+fo3y/EWZXnWiqSFswMOoj87n1JRDUmcvGUcBcWHCFS+Ig
wXYi5H7kXQFj5tGKXdlXZiyc61yxNqog3/Te3Qxvoe1ZK+74nyqj+kfxcpTzProt
KY8ytkJ5DkZDSRHsLy//FGWcNtvQarV+bXyiTTUqJmGNLAJBbT1olnGXGSGWW9IG
DG6HFOBQuBavAKirbuFIRZ7iVL3uXzUCxWm8YKmU3CtPQe2917346bJTBfXvVlmG
uPCgMBCoJTkf8p0sMO9dzIxGhIHgCiofNLkVzVs06VaUCddR0SunX5EANuHYcsfJ
zM3p1HThz1Fmsf78q5XRfmJL7fE72BAL7Cw4xAPfospR4SYe1gB6dsOiYorj1eTD
7j+SF/8tiV1YSfxxR2g6bWZwxQ7r9JR3ZQqOIDPtRFlo9T9hJvjgXiSnTZykhbLo
cTwuQvRHDc6EW7THP0mOPmVbIYtiFnr6hZjcpF4Ff3+EdxwBdLCLsn9a/48/J0Ep
aemh2Y7AJjRRc57sX5ynJaqwVG1999Sq/yTzM2IWsDWFJuuWgt0de4UQPRxCINS+
gqjlvcQjVoiiDWqV13doneIfopSkmUVU98RoHo9xbnJbnckwKQ53oyucUHVGXc/2
NR6wd4hzWKlRzvhRV3fe98XWCWuvaeOzbxQI6yot7UtknmmB/i99RGgYTDeHJNn4
LIv5ZrrXT/r2uFLWt3Vyshjhyo694K91xZWgsj82IkwD6zjQy32/ySQLLRtRQS9U
pMWdoHRkNeRksKgLhxbekeVBMqFh2Jpcu9Z4++8hzGDL0sgWmSi0F25wPMHBlVCn
Oz9N/YcsrJ+LCO3Wykz7nvLB+1YAP3TGk9EglBI1Gt0L8etRfvH4/I/vh/GmzoGg
6FkqIRRM4poEp81VrPOqX633umZOrhmLCfVCuMFXxixw1WEI5hGst2PvVOb7egWb
5SvmPlUtP+FCXDCMaIsCqjQ3TGSUFEd5R9/os/ukk1h3TWPbTu4KwzyIx/qaL1Gv
DwlY7+e6eJLcfAWKvw2j/vkrsOAtRJqTx0LbHfzFIaoOuAsquJR8jNXCeSEA3aVR
J38lBWxJV5Gdav3s/I0s2RsGl8VQyC0jXKobQggUp9RVtx+CFgXwHe/HQ96esCGa
5y9LeIUketXy+8/fh2uuld+69zZ7s4YMVf9pgo50Hcpd68maGbpWHDXP5/g/wetx
HcYfS/E+i2WCuDViLH9f063BT8XlDGIrf8sgf1FYFRiIsHIVxPt6Spz7+pjHutj4
Q/piM2RdyDL2504bmsjhBFWHjCdEC3XbqCaPT7n+bcZEQT266mArCO12+OaQwvjG
hWvHa5iJrbGG2dRNCZLMTnMCIrhnI3oa998xiGlJCPhI6FwZdXRaCvGM3LtPqtS8
oKhZu00ktnIe5nWsmEX3pPLpznk8p7tMJydaN6OXsmeGzRvv5J+OLbGPdbJTf1b0
PbgEDvKBYIb8bYBziYRLoaK6RNPspxfLVZ/fBNITsBfq68CbjSHX1Kj4OddA9xqc
yanRQYr4OXtsEKVAF40qOO3dRF3iSlq6bo1m/RdkdKacPli6MxGlY1uiosHcADUp
+hdEfcdMgO2MN4E3gewDCvHxomVpLRPeHZWcLKBUrfAbVvWla60rXI8faZTEEtY3
1HIX3u0vC7jKXAlwatL/bFIdCE3GRGW6ElHx126HTXuV6bmPNrlvGO0hLMYwt8j3
HURskdiYtNMupzjO2V1IondgUzpAd+XaQXlDynaFMQ2gpclxJPGyruGV2dSefXdX
Xi6UOpnqXi750WpEugmhbgALOha6UV+SS1k5oV63z2gN4BsoG4GoSN8SaAsvzO6W
9bId1wQYeOEXEm9whPGLUGCH6kZHMT2BwBSPoxmVB7q8CtZkUq57vFs3TyrADsgj
6yGYhcZC+V7KYFeAdH1q8EW/HRwMBPETzruHwsoY3qZQSgXf0+I7pLGvCPfHYkxT
km4PWdKkV6qjJaP1Gundopqs8R5IJpWgDpRw6DQdxA+M8vAwUzVUoAu7VMqGpmIV
lpYY7g9OiFQPRzpbGuz4ms+hoe+KgOUPfC+sUHalq413zHWUkrONtJCBxN4L98Ml
S+CWZBAki4vNzPIXbk/h7bvHOx58pN0FjX200Y/o1yf+d2LQrH3oNiD4NEVJH6bL
/FJ0hz4vOD6tHlQd+wtFPMj5mx61SdmCfOUt0+Oi2JiXkSWvzcVnFRkqIfT4qp9I
tlgw24EuVSNkxxA3OY/nTb/u7zGHLZPblgkMQSPPf6PzolxHXZPhgbUNxxYX8/aR
GPJeFzTJJhx+Y0IJZBV/yqCW4ZHncPfE91R3eNUdg05HRuPhfEtOFvWVUdtEP/Tb
dBxrCvR90uH9udqdZGUuokkMp7gcDK1qOEOjhVuwdFuXSHuqiVTl5qD1ERj1e2w9
ZyXcBXGRmoYGom5tRZh0ct6pILLy4fyvKjYUtCBEHzGVJzeouwecFrMW8BDWM062
CqgcGQS7MaXm+mq1XayNLAKpwVFpiIfVkvWzAM49yF3H0macSMRQ4FPM8X3UqENN
nOn1XmztTyzX18Jg4ZE3VlZglgDOqYT9VREYa1Ro5DJc++98NEj/nqsJ+nzEbL0P
eQ2xw6X7q/0QPlaM+OXs95y2o8TdTdDw0ZySsB8qWiKOhbwPCb1M/jKv4vl/fyJH
XnnAf8xq+fddc9HCy8MzywCijHhPGrIIf6DwAT9SrtidtlUyUQhLQdHVk3E31DT8
+TgfW7p2W1tAwQ77C8wmZ9u63/j8Bd0j7X9Zvsnltw+ZXgWDk7EiQNLtwSWNJRLE
eBPR40a4EbHPiDnjeQ59uK27wC45GJdZnG7NFd0qC256/jbdB6J/brgyaoVFajkJ
fZMEL6eB6yVeswM4uXKdCIXyEWZw6NS9fR8PE8kibU1QZEMY72wx0czgJbQxyUEy
en2YAcLBhkEVp7D2WJKqsASxw1KATJsVBoAyaBfEdYQzMeHO+VJmYgEQef7rK4/E
A4XbkhS5dYiAup/JoUJDyk5xwsgEO1f0VlxnW4jx1n04FarvqwoW3q2nYvKE/nZ8
YtKStFWHSIPEFC5mH/6L8MxK3/m5hupZOfYUNFAopIg5zxx8grVVN5iLJ88dHoPb
R8u0ap5Ax3OfEN/gneGAp30/XKeqo7d0Dep8EkPKMfvueKLFJpdgC4hrKT0/he8E
t9kzpKXMcOFLbxlt5lHKqDFp1ZGLC2++hziRb96G7a1bAL5r8Y/5qJaGp/AXxXzg
fMbAu06U9q3zosIqrOKBamVvVkkCF7EHXzVlbWnBUiynISDEzrenNl4fLg5u8fPI
pv5ooB969jlk6ThkRGoz+dHbu/QvRvTsF0WMLBpW1uBb8gzjsBwW339MZEgx6mQM
ZH0anpLu2EoVGxJpEvJJUnI4J6bQKAY9gVbOpeVqXrrqlaYMair1oRLtxVE9lZpT
hwsDtsBwaUKWQPabq5v2+nrymTCWZURmbWuqaSxvroj4GsTBWIwYEo5aCA963l3N
/HIBaJNLKjJj+dVmkjfIDTZSxSgoyeD7ivXSmtxxIgyJ4UFfU0SgWwcA6K5IaYJp
+spKRFSppNKCtcTGPs24tHKWHHtjcVfysqTegzUld8muswOZeSFGR4xh+JAoseoi
ylUsgK/Bjs2AgiA5J1JqEhU9V5ojE6z/YQR2F5EKblX4XSCahNrCJS2xAplBotnj
TgeNtDR6PG/rmmmjbOnOQg/BQBuIO2ScqLmctGCNfCl9fbgZfVs59XJbHX81Lk+2
y52tmFxVSAGU5DciW/gzReUZ4l4rhyZRDckiIssX6UGQAzd9nJNL1Ea2eFTKnR2v
9mPMb6+mMzBzFeObO5ai4uj8pe3JcZwLGNfZcLFJX6HSeNCyfq4t7dPy2I9fUgBB
yvvYYKsk+NwJFi2ptohh1mv7Jl5DIg/sCZcyaQwPWWxuM9KTXL/fX12oeNzxRAyF
T9kM2Bkt/GwPwXrmP/enLVZXBsZkrn7VG/3nY1rHhIrDfjdGxOLKRdjTvdgs4C7M
cGNdeppdsN/AaDdd2CBDIZU1oZ0xV1sQD5bJ1W024OapLmyPjpADRCjASRS6vpNK
kLXF+8Sl0DsHY5bO5yUSxsikFB2rpXOFhVU4K3t41/LNWT+R8WbblNdcdtqxBg6r
6bvQ7lWGCmS+qKKzuyiENsj7Zox04ymXkXoLC/HJVJhxVhP4m1sG5Q59atGCesxS
xHvES7fh3UPvVUjZl9cI33gqg9gX1wAy73WPf6TCOdyFeQMx7evCUqhy4vfXrolc
O/U8aW/L46EYn9SZ+sATb7dZThVHCkx7b+qhG/Z6Eij81AMUpaaJYoyMYbWTrf5p
HEXjQ+d78wpvYYkRChjkn/Ex+iOffm8E/sSDulYW+ZTd65R/1NiZ3ZHFEWf5vqZG
tp4HH0Xv1YuB5tG4Z4DjQHL2Bqg5XJXZ8o3Bh4CcHBg1gVO8jIybKmdogqGOfQV0
vxy1DhLc8Os2edS3OM+Otm93uh9syCbbPsEJU3CMbSY0kMbj/hgwWJqVJc1W9Nka
zVhZv03Fy85aAG7Zu0InxzWv0KX9Zp5Iq+QdKhS47x2RmEXDqwhyM2HKdPZWg1WE
hHoBlHiWaM7eFwW0xoby7ZiJW0fIJtqwanRQaz4oCwMPBVOjaeMfXXFsLS82T7og
Ni2Wd/NH7vygrR01bb2KgWns61FHqa6IhuAuekdSr7oQztRltza0UMkYeoNpaMvm
9AkkLgFHqlncv4eZLMwEeqL4npRJX8zaqSxhvSlf32qMbvHxXl16SvvNy2C2Ze8V
B67cSrT+jJH2giNk2p2nPnYQqBXa2RHED5CvsNWeBV22Nv/5OsqQvWnpbbVQ+u6q
SLe8E1JMbqeU4pL4ub96Sh8JWL0bQC5IvT5qNXRz2cpX9VpfrsR97u/ybGH9wBnT
tZK+xExfrcqqLdULHAaRUbGh0DeoGICLqc30Q7jVKtR82FAhewukXLO/WHDmxaib
2eZ2JCvHCX7NmHblFd5DOEPAYN3fS4qIrekHNptF8QmDO+zmFpopfACnVC+XVn25
7BtlmtJpigykxBV1KD8RyGoRc4XfT84ES/i/mZmQB5wxD3vqXnVqePQNyGdo9sGF
+N8JPSLWaxH2kQe0mjvAYsE0c+8gISxVxrqN3DsyE8RgC6xA56FvGDE+MukNTWXo
gODFvHqEhy8BBTPkPF8cc976fE9x0lLa8ESSK/eGQQR3PSkx4VjKwSpxQF/H+xo0
1lW+rOOqFlyI2bTdcXh5zt2eICSaLn2UtDcFauZpq7StrUsghnPyW8uOKI+olKE0
kLLPaGDLOkGkmOE4ZYtfLNnahSPkUTfa4sdcta7tyWKxlLVty44U71zBVs3LDCyD
6GUVxBIIJ87Fc9IgsPxFW70RJSaUns0LfFtt9GsNqA2pgQrzhSH5ECTbNrZA5hRf
bVC81xZp8f4BY4YGWASatagYyzpBiIvW4QIHufaPudjZeNeduqCKw9O1f/Az43v2
4sB5lRNymxL9J03JSOQ19zS2OOTToCKPcCpNTLgCJhcQ/5vR8bRPgwjHSwGybVMG
LCpx1XUXyJU4Sfmb0vdL/0uI2atuIccSi5QU+ibaNi7oYl08ZLVqZ8Yho2g8ohdH
Rl30Mb4HKJGdMOflSwZDp6YXIJJQrd/17Y/RTFituBGfT+4T4mF4H5jZj5/fof2k
ffMOKrHy3g4fkby4W2Yw65E9Cre3OMnqBDn39Hv3Cd3FvxRjNkMmAv1MhITBoB3B
sddJ/WOqyYhAVV5A+mWx7xylh/1mx+12PJgkuGkXe/5x5kEvdImvPIg850Lx0hKS
vbgN5Xeqk6djhuv9V4ipsmM2hsGQDpxmpa/wGi6CSr1plf3GZ5y+BxW32vQZRqOQ
aSDQ8IRNrHZq1bmBb5FJi/H2RL1uHOAvn7Q8CNJZ4iZKcVAarcGHqRKQSqBaUfA5
BeWdcD3JaQOEafEizcoYW5ebQKiI71gRb4ZDRarvvUhzE3QOSNvLc3OFdSEDaJRU
Trat05uo+iGPjkHaokCerROI+3tEfUC7FwhnqHI/G1zVd27NYYsf+J6ybztMRxjE
ae/lfmKtFR+t9EjSuBJNuNX/tvbanLq1tg24kcLSTlnpG+ckr4CHN+O8fJUHgDW0
h7NiTu5TW7N+XTMhgxMpgUzmsvslFreVvcqxmZWDYUcDP0o8/rSis70kwx1ITnkm
TXyF8JHAVw6kzuD5DWyudk0RBn5C/0DC+R8hER7qaJ76ixTfl4mAXsMMBxqfrj+W
piRkH0CbFNkIhX5BJj0pbGgriZOpGAerD/K1hyHvn7TP1nGx8tRSp/m6FlkWzn0H
l/k7SsAsBCknWSLPizWQDaofzsi3/yTyraDN/DNM0aYP68nhw0fulqkv6U9nwxj9
gmrbOROZL8K5il5odNC47mjh4Go7p7FTmdjQdHVRLjdyRavFuBhhu9ZuaJmXgBWC
mDnv2XsAOXfqx+WGLcCfzoKA654TLdLtS97AKFPenQHZ2ex9ZwrPZgiWp03U4nXx
2Ny+wlwrcU+Z0wgUkJjCeLG2zj7vyTscfjSK1TVcDIAQzC2CVvklLaTuMK8wT5ZO
WI9hKMUGpz/ByxS9pFojGue8u1J78xU4vFn3uDv0K96VY86d1UqPx17Av5ktkogR
iUUvlcqeS0HJ+bCkB69GT3oAMPSIZptHysqQaZXuPWGOlsygpc+G/PHy2r4AOkh4
bk+6g+VtuUs72xhhv0FXal+OYBzEqGnSD6BalJoFBsAw0jy9JyGCukhnNDBDeiBC
Dg9VlvMuXcUUGYF5DByTycVwYQ7sZIy/c6KzbsUSrTvxvS4Hb9U9zCQTYd2i708+
s2FJKgdx0kHNVAda3licNZGqGWR38FyOzRppzFqXKzFmAoyldjcviUvTuJD17l7g
pgSFV4puZ4J9kduz6dyuNLfghBeOJSYGfbTFjkEQkR4oi7xOjLISgZxqILrRaVr+
VHV8bIm45ohYNau2J+ovtSqwTSPqNA1Z5x+lf6kxi9GUk3wCXOe9C7isqYfySH53
eHV+fEGLgh9uPhC3ovBVEGeloWvL3yr3RiiDY82DXQe2rCJyGddcdvR9WGSxN5Is
wTcMrk/+52CBrf//aKwAgHsaLkWQ4NnR0tATaY/sOFPeaLNJIX17EQSZin+H33UX
ZZuvyG3nkKdaLRVIWq/Lf30c0JCZcylHYHoBGCgjArT3uO9AWD7J6fQQfCKOPZW4
ISRzXtuTnxIgVelCyjutIDeadOqWhGn8YBOabOrv4jhTVbOHQvrDdCq6Wf6LP/8j
DdkNITyrOqNGvD0+b5rrt98lXm8gbHwNacQuRUVtGEtYH6/sOmrrQuKdvTLnxeMA
yti8c+dxbnJz0wet0rr5iZQAs5bB5he7lhT2rfbp3+YclVuFftZXi4rgTgS5j10e
jVKeAA9z5SvO5JRGbk6gQshnvQyyoYQVGfMKwTwGU+7fjqWaGSjjcQJhC1jSHtJI
+wgyQxRtEerW5OJxkhfEvma8YzzbdVII2bvIDOTHUG3ChIWFR/2NcP3vvU6S6b/5
I7YwOGua0Gqp665pU1kYG8b1eaJyGU8nKEWUbz8whYebFhTErV7CNzrN7tEIVKbP
FOfdzGunQ8YsF6d5sVcNKQrMmlDdto4GmP0HQ2kEKi1IeqoSbeOAhBWtzFq9uvbs
PufGylJcTYEd+gBlVd1fOaEK8oRB30Zc6WL2Fht+6952Il3co7dP3j3qWs7EyrL5
NKGmwrI8vCq+4iKI5pHBKL1qrNhC0h/yUINgwccPe6/CaNpXPkN8xKxxduKaiA6F
yCcAxJhg+tQJ90Rp+nOypfC+hN7tyaZsYVilXL/+Tk5KVS2TgUakzSmuk3l6+6t5
/k7bl12cKfD5UQQiQy/aiWffW/i+XD4L77kNMNEXi9fPRs17dbpOhrSzbhQybNPK
6J6C7NRlPcTQOzqbIBjJ90M7XPRPhEFPV1sfkHfnFyxkfA+BsqE1uQCP/DjzsnOb
bFbj9Z3YqZ03ePwbP8/aUlXlwvkM/2IZhpBmGfJBWXmeIMjI+Rv0n31gtNpbi35R
kdqo48bUaLY3w9vChtsycy3IaaN8FBDrQBgOJgPOqWhtfUu6cGMAPquZLGS9s6HJ
UyciTEh7CMJFjp1I8Lifb/I61loEq2rZXDvX85Dxi9+TX1fL7VPfJBSrFlQ24lEa
1kxIP73AucrfrvKT0d71eG4yDan7uuo/Uh5QudfPo6cI5IjVtWNaqwTzBG+T9bd7
FJ+xJrYbKoa8DSknDvG2qTlGbo3zT958OgAmPNnHpBGCCLOkO6ECk/Mq9WoiZxAz
im5fiwyUOlMAShMhWW37WkFYKVT1ENr6ZxWhJzeVYYHghPn2WKvNGsYY5M1uIb3w
da2IfkJersr4BPpInLBttLD6sZuBRRSTdn9r3dFB0ZHzb36FhcHDGLy3FP/fSVuz
NMBXHeh6QBKKKkmFd7ZQCcgumiXhCtaM3bbhb/lqTeiyJU95kKnqJ1wq+fFIuLN6
mrEtjeaxkuC4iCrrc7VFbQiyUBjsORcPDxU96+P4jhGN1kefkhSHI6f6h30cEEhW
vxuwgc+hp/XFoWxt4s5IkKuf1PLz7Ii83PQTZcMbeJC1TEOspYlL0Hcr09DRDVla
mZf5KrtA23O2ZuC43RhuKrZ50VP9Vwx8TitVs32lhfFdeJ5Nq/8K+Gz088JPyQXe
ra2SlW+FGxKxwfxZy9yLETRlz6QSL2aNlYiCTae3VZJVHhBM8psxk8ry4D3Zdrv2
wuz/bqgMTwDFb+KzD6SPbFIoSYRCkSoTCmq6OZLfP3DKN5YTbuFZ6d14yQY++cV3
yJSR2wAC5r77O3o55i02UJSW45nRU/N1gUWtAZwrUjip9WVoWEsL8Sp1Zvaf5GuO
/qV9/gnkm471Cx5jWgKHJ1tUpTvNeiqENpBD1r4bgOLqeQ7Ty79GtTQBg+yHTWBN
gnFPJ8VVrcDgYNLd8y1LybUa2hWJJP0PR9IJXRrfF5yXL6ZUmZtDdgKf9GGHAdTy
M9PaVzFsGTOFPW7KfFjBfv7FHwc9JZhJicd5S77bvK/83QoKGvvaEhLYVML2cE+F
CsQhr6rbdY+SucpI0RpOp8gHt4yH7wSh4ON6VrYNkavr2hF9xqrBlggoUHTN1T1y
844PWh+ZrhMlc2jmm0X2kXu1feZXykWfYFBlqU5KYpW7Lx0PBUogUGlnvO93mXqr
B5C5ToczefZtnVfy20omd1p16HDr6dXxtiBfyR5SHskm6bO46lFW3TpHqmVyFVoK
vkAYn2r11mollbKuldiGlXcpvtLnmT/V2Tl+ma8V3Q6uhtO2y/HmVbKFgewWuosQ
UN2exOA3AhXgBMXk+nDsQM3evID3ynSNgaO41OGp7btcoF2LKvWcY7aNxFGwXg63
3SCpRqNwI+7+xw+jVxIdpLmdkzoUPmEF7GwMzPKB4uZs4l5ouS/QLXuAthoXPhbX
dQ3Zkdl6p7jAxroKp8D7uT1inRcqW6GLNBuDy7ZXJgRsLaP0bj2TcbI1ElQfboCg
CMfb1sWNQ2dvMKLFArTvQB5av/w21vjTlvKApGVMdLfqimCESCGl6MUfe0I0eG2a
V8zZpywqoJwMFHRb6+L27aF1rgTPL7I7EKoPBi0rzQbtosmN7e4dSEue/ZBr1ALh
xb90fIWZCmtxo/46qxade86kdQbKl1mwl/1UuZh6i2L8UVcim1XgRpxu/N5a76gC
1uFVipSELHTjBHxPuWRbKMA8ZxxV9zVu9wYbR2SaqFuyot6rQ7sawNObaZMRgC4K
cTOxV4kVS6dWAydfW1DP//RywIo8ui1SnKJmI+ss/mVQZdRhrC0emcRZo2//h+a8
wLNihvOULCGqsYuGIuGO6zYs5065e11vZI1r+McTktIMtIdTPkTS3hTZ/1y/3S5t
RmQ9na5AhiCG37V6U7JtHdSPFxMHo/S5Vt6nwoELkFdiotxsvtlQap1I8eNrdV/A
hddSUSuZzAaWrCNzeUdVaxQocf5iTrK5Tcj78nhw1BuJij2BGBJNwsDLzkfVLR7G
vX5ORrimKBorFwM5Q95LG5SPLEeLtatrdS6mgRPSFWPCgaA7xNw2rcy9Lj7H6XJz
OZXv6OhceQHKTXBivJKUe7N101tAslKFTM1gi/FJ7tweWw1vpxpVAMbC+3ASEyjd
UVowb/ZMuUqhE036uVsqs6OgbMyLK6AbBhi5lwSCobUzY5sui5Dc3K53FWOiHfAb
NnlAgPm1Q4b317Nvg04uAXXFwTg9oL6mjAMu/Lv8qPkeXr4EoEXYTTyPlJ3xy1ex
5bb9JDB3oXLkUASQ2sgdTYkDsoqJYj8niOL5anZGenUjE4m15w9nDsZEz6MmQ63B
Xom40ZZhc7h9KtPY3gviD9hTMrMp2oK3iZfsZPlxGVoepiaRbeWfXWjE8O1K6kEC
XeWIr5AhXBkjckLHyjYnOSBPTBPdeMGR1b9YICPKvdeytB+z7mWCC0cCz44WD97H
kbp7v9pwjQhVuq8ODg9Q5lop1C7gnqvihqswx1pUufkePF98h3FaJj58nPhTNbrm
eGQ7TfzPEtcRcD0kwWoLwe+GQ8WOOvISmEnkyOVkO7Prm8fkKMxQbQDVu0PRqytQ
3VgeRfI8RYzvakEKujxj3VUmbDNf76I4sAWDzR5f6egveEcRobM3CGe8VUkIahVK
ltW9jx8LXf27NT4//+JVmhsITtM+62S3SiHnH8Uf6VF3h7ocXF8XxG36/F2A1vo8
h8T23lBhZfdt0RMOg9axjuRR4Kv4IkfcdEFq2KmHokuYNtqxj04RV4Ya8hUz8GR4
LJ8EIh/XtIC5yzj/0hKR2NymljD7rbBdEyDCt4M1Oj5Z5Bg0RSwJrmNBGsL1+Rsx
SLTVy/KKrgHSexfqCpeeykkQcgfSlw32qG6l4NiQHA9KPE1+G/Zgb7aUCQC+1Doj
6+aUqfli5YmDz2IJoJePPubgXb/735SI/uGsNxywWMxA7OjwtLjbq2juwZ+auLQR
OfK8vVybgRidkJ3c8SUBzA5YimHWmYvzMavXo1fmF3pjjhzWPrcqidtOFiQNtaqM
+rgYtducP4maTlxUL/bu7/5fXcIR+FvdZr2xxyekTZA3ARCT2BxXLSkmYIXGcsMr
2UPEPjTQBUwFC4TIs+qNcGRdZbBLKDPkVc/I3huR83SHIpAF5wyGANog7Dez9g11
Hp+DTa3zF8Rrezv8D+ytLGZdfAFwoY13KhJ7FCo6aEXAoKtdKjwRhlQ9Ydk3+Oej
kvKd2K8eToWt4USyIwh9Mnc6Zg6nbxTFK+P/1uZwvd1EAV9j19vQQPDsmadkfMYH
KWi3rUwQvdroIYhIwPH4+U/MNpYwewbSQ+YhhwBglmMbdjKzAuYprchXP8neOr9v
ZCeB2ovWSD4oNr8+yQJkjqEEvtPUvcmPQDAWrd0qHwgjP19AwKXyEeNJLPsfb3HB
EqzmiJMqucvhegyU1lHKGgega1BxGoPSYVhsPeQmzQlyaKUYuxhSy8VLThr7UfDI
edxhhZDp3iL065TDsfKi0xHGcbpT0MCyvFLHxJSs2HgP4pcd997+TIQuvwWRlJIK
c7GI2D8+zxXC9wB7skwKwD0y//Rot3eOHQLVg+I1rEcyhs7F4rVAVbpzI3EcOZ5p
tCaDqjnpkDQm8KElP5ozb7tPRwgdhi0di/hNWgEG2cm1NnuQla55iJb6zQLspkow
Vnl2u1EWwDsEfZnPXSaCX054/xxWGjh6YQ2wfzwbRQH0XN8J5CwzUcCFT1Pj7DEu
1B2DMr/N22CXXr9jrfF3gMyUIb8aqkhbGXJSfd/Sdk+tR55/O+S2jgIdy7igmE1y
tZM6qhxU1DfK4GgewmmERVOjpNaG3TkN2FvVCrjjckn2mW3IzfELJ/IlxrZ3Dynk
Vs3xM4qEBoNCCwwBTXEFrPRAEGKpOAmz5c9HlW3abXi1UsuL3N69gUV1J5+0QfqB
sLoRhsefHyUw00IZNtqOYhpmqrr4YXkshTPuFuwghr29r/0t5jai9yrqp47S07hb
VrhgWbdbLDEqh1A+pA01Uij55U8u8uCv/l2thDBssCbCO5/pCPIPfbgkhs+6p9Wa
k6L47UZLQGcEZYm19tusTl4db0HjnPausPD4FA5RfkgjTtBI+gEjL3L0E6KwgZ0n
NFpjQP4XiJZnHpL6AgM6gD1ZLzQAp1NpAtcPQiXldZjxiSdIIM+xSk3yX66ZPozM
4qObMP0M3o8mja+ljUGE2uTQpfXHffHNTGd4Szu3T9taed/uvxR8R1TG5AwlGQQ9
fxFYDKNOLZFDPXqvEbZ9HkqmKHP0RM9XHJ7GmDMsYozXk3miP4CdfoUxdew5IeMI
I/FXzasRS53kJK+IX5gsPgY+1Xb+XlD5VVOn6M+G67WQ5qvXxlnGsHN/VZekyt7e
JPAuC9yKVt7sZoxLwwdOVgoAi5+pqavvv4I0xktvRBO5LXKoAwioGaf7BN68K6Xu
OtmistnS8tcwJEt4O3hy2hVROpa79Tt2H54ANJTjvXmopY82hhzCQVqbJ6l/j9rg
PhqPTl3TKTG55vWXjMEpBam6gNJ39xPaXWLVrkMEw/Sp3uQZ6sV0n+5RgALCO5kM
udv6AExBuHQYfP2+ntqJ+n7G+MOIM5xTRHJIr9CXR8U/UImsCLdqaeknvJKneJJ8
XaeCoxLDD+1a/WgNFmgT4FkBR16U/lw0SEDI6kL7eK0JpyfU4qMoWtxG9TJjJ75q
yMdC0dxcxFJ9sm+cB+eWLmNPTHnpFceGzWAn5pweQJyZR3t0bOmqgoTtS/egRun6
XkP4F5XXSPKZXbaJ8WPrXm9bUYPfCmWM79/vLjfBVu7t22eH2SRlQNHHXJz5SAXx
yldO5fuNym8UBhJeAXjdlaG6/EXeHsmD9Ykjq2hFllBiuVPIWLidOaw5ROQSpVqk
vx3rp8939SJonNLle8hztffAFqULs4/TOgSlGZIWJPBeVc1SicWMzRSFFIOD+DiX
klumM2XdmNELKYDIcIhPZfsF+N0HRELnhnWW7yFw72qClKlS7xP3vOnfX1owi3cN
FoYS0FwySdc4z+vOAc3EV3FTnzD+bVLfSszxRUXiis8ULAhRs9HLbN4J6aIbOFNC
ZLgDNFUK37KmU0W4IXfwh9nFpNhoYUz38Zn5YgcsC98Lj/haurHZrNPfdmphbKXb
6qmIhrztYw64nq0XW7qxq7mVsFKeyIYu+yNgIdzomZXNDCqn6DJHNvF2WjRDggjo
1KHenoO7YgB5W4DreG4gcLFx7bifs3lnDe5PEe1x0dUP9lFu4lkBAr4C48+SLKNp
sSWpugeNq4Eam5UJW7n0r+lwwmpdb1w3YCL6YGkan3rqoQtN6AqGl4/gYlZ295TQ
rnd1nBZg8SrT8CRYv8uTaztpL8nFh/85non2TeXk1sJ9wIs6XaEfzq2GXnR69P6c
E6JSRZzBKi1NKKz4EvmYc+1tzsvRDChjULHfVBGoP3dKf6wOje30lIg8p14Zod5T
i463Z38X0BXx+6frHnq8NmA+dwXb4gVFDfZqqHK4nU3bFMlVVkghm2jpaP4UuuED
XE6HnoQtIhKuVIlPwy24mbANzBs5rWwZjh7Cb+PRjZf00Ggz39FosXwfhn3sd+2D
zMveRpD2oBYhP92YVeqzSOt3noJxHVs5o0wZBjqxHxapXSGkwp2V6+W1vzw/y7X5
TUmuYFbiEmQQpTDuXKW+vnrVnX20YKakl4Z1UsZXoEhXggv+ZGyoGR4tnT9MaAWf
dlWXSzSp00qSSSzlXpHiVni9irz4DNot8A3W9QwY350YOZ69wGSc/Kd5pGJFNRQn
HySbbJBL8b2vg032PFqFEhmyAi6/BdOtxcH4NHYcKHe3/9Aif5vTscIFAh58yWjy
mokrvjEmm0HEsisc9ZkKQK8k9DMlWFB5p2DU6ceTTUmrRsEqgNeIGH+9HUjOqwP1
KdgFQ445gj+p4AWR5C/E16EAD7v9sgfiMyGAmsRFknoOvGQMcrfhMOnaiAm491Nq
PRO0nwLxUhDtarsvQg5KzhTheQM4KB2iCCVEWME+DvEcI83biPmrkZl5soYCJe2y
rVFuk3toqlM7rG9MH/pRu9INCBxrVWXSJy2xNwD4SJFwNi7Mq8aguHfBRGjMuaPF
okKxJhJGj0XCPaTQwm0Ne8I0vGqtN8zJDvsr5Drkt4UNM+ZqUBxyuQetIWS+vIUc
P5F/4FkOGd2LeBu6u7hvhxsy5ELxsM+U1Zkuu7apirMbdbN9o+8KH5rHM9cTC8y2
kf/d2698nhLeCGKK3KXrzwjYGFL7cb94svjW+6YYy9gXkpmjY1rk4hnfszPrJlaU
4ZOcPY6EqMhgaIAXFj8Q0YXeP+Txi75yZBqrPZNGrPnPKIOEHzNzDy4dpBhOcKkh
Ep9l8H73dA4OjMR5Ih3ERA+dqTF0goBygEkeszCxdrCD/D1HO/gMY38s+bI0gqpE
7Pkja5MxXERphniDSLZzi2aGEruoBpwl449Q+JvlABr8W4+U/m161helRnCrHQDK
9ZPsxds79srF7RKlgrkIVnEW3pz6b1gfOMpprUiWaJfBxLjKUWWCI9Km2nUEvYWL
Z5ynWzXui9/ma/r+pSqmLIxod7EP/SkfkTUE06yh56eUeBWdNM0rt6075j3T6NRE
O93+tWRWLvIFTGnQARzA3abeRbHNh6j/pJ0OK8l/NL0T/P2Xj2pyMN9kxIVXwJqr
oTyI0zOfP+It3T0gSZ7iV4LR0rDEhFms3W2Rw2IHG5n/nhTSn84WzCh/VwKPpnrX
+rDYlbxukD9aLC2rsFhXe0ZhYIHICeSwAs/zMLutz1U6MfwxRnXo0H3U/g7jyii5
eE5IkdI0IJ6y/6vYqhI7Z6ZIfjpbsI6tcKW6E4TaAkZ3QTiXJsVfKrOHSqXf3nLd
bwzhp5mKpPKsWueKzeI/JIDQb06LhU5NYW/vljonOeAQ3Z7XBNubolFwVLFFcbtB
LlVJYpfCE+gB6e6SiwELT8niRo/SJxUnVZXp/WHCrcSnEhjol55Axh3b0g30KMyG
lv8pUNyd0Qz5duN04EbcrNsqBgcSIOwI5tgK3NVPrRgz2EtLE6TAHLK4Zd4kIY5c
43pD43/yhSt2t6NkTTdMz7oltwcPKT7vbFYO3S8uOIbUosmetfOpFqMB+rk3uXg/
bqncaXT7kaUlRssf8xkf3oibjWq/vFpLuat9/uRMRBYo1SoBTsw0mZFh+mx0H1sJ
hyxbp+58nx6sKCAzPxJ8I/NkW5XExLn+fBSBkMxtDkCCieamQK6wLYgUD8lC0MOK
kARiiMyxakSTZtw8vr+5sziVlFlXsyfX/p0/Rlf+WMNBi9QFXvdAT54L80+qkWKh
j4Vrdud1s57GjAAToDhSjALsOtyIiZJFBxEGhZOX5ZN02ypqC+9bZSX7rIN96rvX
y9+L4Se54O9kS+H6B0nEZXqdXTn4cPO7gDBAYKcEtwyNeULnDDShjToDJxWH3mJ0
rN0cxmLI10sXhwACMVGh00t3cvdEBKNZ+J7EIta4a9TvTSkPyRqztAm0FrSCqBNw
Jm9rD+PffALDzLOVMtIMES9iNWYvsVjCxkN3bgDJoYs6VkcWbbCqTwszBZfaGiDW
sUMI3U6a5ZOIHGxvwQP6QKJYeX3gC4rIho2D9+LBz1iVb+WXmTFR1o9OM0AeISXO
Gd9XbC9d9dVwlXOZm9PjKWm5JI/Bzam7lQPMbj8kikKyp8R/76hlBroGyhE5FVfi
B93zdXB04qKF6pAVSJkVrQNBLxyZ9oIj1k3t9p13tQKkJcP8HSFVQv8X9pqeygnr
wvqDz6yEXhXG6KKCRsUNKiKVtqfhAAk9GGEBp1krXLIJA1q3KiccGXwuyVKTD8Xf
zMg9vR/HENip/vy/RYhDUQCi1/tqQt4zLajgLFnSfMLR+bUumVmUaaSt9/D+fcQs
FgNgWMa/bad6rNcASNzaP0K2OGbnKzJLSDufYezMZYnIa+JVCg61wK+x53asHFSb
DK03jWUyXkxWeeWo6auY+NgpnaXkPie7HuIolwbSlv+T3R9T4iWQ7123wStaDclx
n4DalHiNnN8tSMK7AB8kSb2icRvBfrdTufIdOeuBsgrzmhFfteXDAykcrO6xzBLE
lDhO0mkvwK7I0oOcNEFNCEaW858i5tQmwLpgRtxSAJnpuGY/Pu+FPDhj0+eOJFL+
hwD9dDqhVde5LZZE0qOx9ra53rpXUrmne/Fw0R8PElo8YLDoRouTmL8NwE/TH+kY
tLFOKOxTRGn8s5O6PapqUDzjPIOEOq0zi5cavdhpuPDn3/aurSZxUlczrPM0rgl0
/gbMhVF7WcqRB7Ds6X+gs8lu+L1iOgj9+mT5IR7MtKPIRbQ1vhAb622fhFhIkU70
lzL//pbctz2GOoS7EvAHvCEz84hTm0fZAQuQNnj46ABLq2rhGukGKvgjUyVVuvfF
L5UEkL4DFgMKzdbZoZ3lQ+fVaqkOStIvht/JlQiZN5YUa+tq0HJLCFrpm1HgVR+J
IHr0G/6Q7EwJqcJ3n4s2MvXANhnYBoR/H6Si2NzObnhnNIMDkaDQI8fnaIowUF4q
0XnVfj8eHk3WZzUN0bZHlCnVI3jBvhb15t3kVJNuHp8l593+rGn5X+RTWhpjpZZ+
wOUxojFfoMv6YdvxN6xLrv+ax2JiEP1+Y++C5vHzqqQo9wJrNuDLlbtxkobElW84
IvIRGiiMpXz/4jB4EiuITeFS9cS9oN+68H35AVtFN2RPRz237U58n4Vz5IsEXYER
/WQPzQ7vMSuczp0oPEi+Q82hzTmL2pzmDtX6JZGTTBoIS/Lmv1O67zfpdYNFozxn
TWShgW/suA3bEK2zsklqTmXQUmN6EHPGkKBtowepcGF4SUrd0veTzzMbeBijjeU6
jD3kJC7qWDCOdjW4VXwauJYgHZQsluKs+qXiC9UvD7x+UuK4cL5cXB5bcaPnzK7S
Gjk9vZLX0MUhFtoOhhb6r8eFoV8VBcwvGWGkVW39bpka1Qic/lbaN9EYTKBjHDMW
JdIiAqXsDWAI1eoRzHfP0RTlnrxECga/70ORpJstQU16DkZkHcr/e+AtQDh8yjsg
b90+HpxdJy6WIFzJnPaM/JSO9WSElo1FEmxpojYevgTqRJCtu3PjMil7ElvBpHdw
8z1EQOTryREVLL7yyR6eK627ebhN9sEirtEl4rNqCZjpyMc0GAMFSp8dGxwLu//9
BlBZCUeAVLjQ3VO5y3UCBlyFmhnkI8AL6EZtzqjYBLBwUyxPAhIVgSns3+r4kfRc
PHIkBAsiTIDLgkHBsheFCDwqGxPMzHSFL25afYwFmkptjDlcXogqy+e4cU1e4nMf
iT55N8WC+IAavK32ezwDiBDchrJTK1yblzvmqcGeogHkbX5s0MsRh444Ue8v+m4v
ucVWx12eqr5pHNO4TBhQa2MOyRa06VRhdZKVS9G9+raIn5JgLVQrU/15o8I7JeDp
Q8jcwOPyxyCYF9YkwNWQBJNcHEbL7NAzNkMbsw5/Y5hFZP9DRym6sPnCSUH6mUYF
QSaZSTN3zLC2XpBp45djaKjasaa1XL+bH4YzlN03tcdj0PfxneLisxGFL++ryH6l
Vyar7gE7HbEM8OKqRZnHSqrxWDYn6LdMXsEXNoFTSVbQ9F2THFdWZa3yl1m94StY
DHjLdlbrHBSuOiyNKTnphgYhrbWhxnpNWpN5D0OYzSBe726ILjnb4z8Zcxib3XJo
c8F+tYwvXcYPm6GnFSAu1wbw7GHavH03715iUDnjTkxnBe6sRFSDBeVHc1KsYqMA
eeYaNrHjBLkSJ46x4G++6X7bqg7vEPcZd6l1Qi4HwtsvypdAfqQcNgvqI99cxmxB
rzN4mQ7oM3RrEE3yxkEwfV+0/hfo77UhVVUA10ygJcy6uLRU0C5nOcW0QujycmUU
NwB2fzgY4dMDp2uDv+/b+YQUuIXbG60faY9msMRylvOArrGdzh28OO/F7fP7k1V0
zeGNEMq14235Lx5Zh7/7dbElSu7BRiStuxkmPmNch2WCDthMaYv2Cm4hV1X9GCYK
z0SNZgID1DlPsp20+qz7B6fo5RLP1lkVTkgklqXm4XlJPpDDrrGlter1jqheVAad
CNnkDG6Bn2iI/zeJTq3aoGgwDOEDMM0TVooJKd/deuGvt2uT15I+oL+KW9GI7mWu
H3NwQvYOpmnVeV/2+jhjVNrlV380znx4UlXofPl5EeNY45PkIE2r50cqFCA6YkEM
wy8K8qMWCjTY2r6Ab6XsX2SSdTFRBHLBRJUGPfvL3S/CODMLMSUaaBQVMfc9b/H2
h8Jqalei5tb1i2xjTm+VPCL+3mp32+ISOE9vPmOU9QqVuPpltP8fFJYc81a6sYPZ
2wg8nfgD+ROKBhOo2o3TLyvFG6vssJiU1Rf9F/91ZoXPykyuheiBnWSVAKNWx9bd
yiZNNksz9S/XWH7JXsUHmkfpq0VujgKtMOlikixfQNereo//Q2oAIxOAoUeH69x9
MJp4LEaFWMGQHZfrUFy2HAod7t9/dQEIxVdhlZfd3GUXkYKnJkVi6PSP4mVjBLEg
PugjRi+2IMrx03YhGybxYs9v4nXc/sQDZ9/gljDfEviG8LHim9jRr96BX5e6kvHG
gDNxdVYKE2P9eIQ5+9JjRXyBqkMXL9BB63h7qbqcH0oNt/JJFuid3jaUydEl+qhB
Pu7vdk2s1ywyV5uYBnp+fDAZlmoAAHjMClnkBi+tmT6EYWGaNISKpE7aVgIMph/8
tfanO1R3uLVhnIsoSu8e4MaqO7bZ2GErwjozZnieMX4kL0ThkKw1sQOdavukZVWV
qf4MB5bw7IEPzhYFfktZhsY1PnolvRn9j5hzqooOaLQfB0LBXpyIMBDrVM5EY9Lk
SPzVWkK65qhzKPF5vKnO4qWkAykW9qJMvK+YIOFPuX7Xih3SKdYeq+dCew7f/P1M
jhl/hh33vXXBFvwMJ+jNpLDPz/3vbBZr+JuAjPQXON1+CHrlXV9hXSkUz/bryDPE
kbaFEEaHgCfUCvnOWDG70YQSsjyAWnmCGo3yaWbTnQB2d+3TaB1LfxpW3ugoq+SJ
Y9EU/INiJ31UCVekYp3qvCN0sdeq80oYy8Q5dqWaGtE3rcZ/Xsw9clWYYMdumW7k
uQdv2/oyu4fa33srerMLH3K9O0HMI4lszkrmbXrk6em5rfBqMZmVwtI5IPInuiv9
OpcsRZYCN3Q62kNYUpkXeRryod2Pg2KkJJ322T9cclwf3IBhKYcAgyzXRsREJUfW
SdtTKLzM5bpALObO+gDLQcj7M6MyVUlakE8NON5jN9rX9LgXP4JV01VVMs2EP0Js
zQxNhNtNtYPKI9j6zwaFs8Uv1948CD0dpaiHMUGGZyeR+3ahjZFfC7DaU2VY9XEx
9ok3uyqrcRAC4U0Fq4rwLPZKNF0A/0yYvFV5HJgKmjWx9JO7Ept3Dph71smhqUtv
bKlaQzFhfBt4l7ZECMs5bDdRQdCY1Y8JRrmUDqvfEnUz92kAO4JS8Wsd+VtvnGME
J0V0bY2uK6YuNqGzfl1Y67APjVJl1CXuZcJm9dbL8e+/QK01Wg+UEQOs0x8FxASI
KocaO4g7nqPnMrrbKo4jMtfYvKvxs7olgUgri2aE2UlG4QwwrMKY9PEX2iwF12AL
eoxIXX0r7CC4pydIsf8f3XUBTnGMbBfnNDwLxbzZF+sD/0PCMIn8Rrjx5vnavGPO
D55axOzALwAO38FPadbIWJdPge//q6tphpMSb/GBBvVEtiSSmnQJSgJss4YbdGZ5
K0fk8S/55UAmqrDH7UDwJJUDW5Mb3iH2VHEhfScwN7FLUTOV8hsvfuPM8lITxrM7
p6NNKKUvk4ZPXmXjT5cLOZsjosDhCLhR+sGhYnusfyaBcyScSrP72uPCh8aU8d45
ezmndeDFrwS5eb/oqXolWzoqQwSj6Hf+IVIf+pqRFLCmi5fZ9Tv8O1M8AYMJSCTm
M56Ay0hp0+wMc6rCaOakKvM49wpiGqmwUG1yOaVoJLAc8apw9PwEeQcxo+BxdBt4
L2dqqK6Yvn8gZFkfIEYl3Zrjr1iJwxkJ0xbSUXGt6JX0+o56FXtv5Pa+m/uQAITl
R5nDOpf+ow9ffZiWJf7XMefZzI/HKbbYhLy1yVAdvaA8AWF7WV21HanrzfVVi+mX
/CvAtIWMcC/uB2XR0rAxWgqsCXOAKp20gE+GyWd2T/8kTIWyV22IHvTlYVsM7Anb
kZBzOQ4Vy8u24nEaNiY3hORdiL1ccmmjcFSA8oCynheuxUPby2+0MT0IyjvKkKOK
TpNjyuQEDLFacEso6Q/cIgbyZ6spAbZKeFRHofEXzmpiNOzIflOL2n6ca2Acs4pg
pll7uWA+SE1K3PQTD0OHwt7YTJo8tlID2cHyZCOF8Gb8Ax7S+oRC9//N8xKVSGJX
9c4sGxtlNgV/zq1+opN2Nn2bV3i+Ppkh3hJIUYu572n5zQYVQ862s9wY2NuJORxu
e0l2wzFHZJgcDJ6nBKUgSOv26yfXdIpXY8aBB/Wjhj4ax8GJYx7p8JKFhDbnr38+
5XnkXRbtz/zQWJW5Z1ufmHjaWPQ/hREtc4f6SR95IHn7Ii23HL84TOafI2NWAfaz
xvwlK32PGdasPkVVu05rWWixJFWT/jbtKY4DvB+8lOterr3nxvh+4LN8MddJuVsA
yint4Rv3hRTTMTr2b+JCayxKrKisCMbqwoZS/stXiUJ8XEMXRakefiQId+MBs0QD
jVZxxKoBu3qXcpJ2irlZrjAp4XoEVFdVHdFDjjCC16qP8iaMeKihU2LRtrPz7zAF
X5nUwo3jQvIfBaVQZcmtYfOr4wq40lYrvS94SC9DRfKXt/oHUPb+N2gn3YO71veu
1XDm8u2hCmki7DqvmeNCfhh/w+CrAGCsfCIkTrDIt+Fu0UQpkZnJDo+HPPraM5fj
06MWMjH1Yxlt87bvIUJEmP8wKQBSNwBLX7FDZNTvzrq1+Z8VuB2u4Ar9x839Yv7u
oRtBbsbeXLxMfkqZjkZJBRmn/nRHicNL1hlxZAhzq86wuL73iQD/aoatvD/Jv+hQ
qClveU709iAgg8Oz7gtTY9f26wT0FUk0wcYkrl/ZZOs25j3PBNKM4oLjASIb7MnG
rieRwFtWgcBcDJov7gdql4l/I80PhOE/7nKScvDl7u30Piye1PKWfqAn22XW5FqK
puyKUf5NJQ9yyLxuz3GIAwQHhfqhCwhVH+/AcVBeJD3QJtg8ypAK2q+vqAMuYc/K
B0QUakywl3t98rhfny0nTgIPtiQqnAnH4ifgLGQtY+eGHXzjOeArxU9TLde1jLWR
Rom7B+rP3Lmab7miHYQIrq0UggGJ8pQMg4/Eey3wbg9Ksi0AOWSiVY1X8Gl4TNgz
gaAGfcx1ZoZYtiy8HPYdcqm+ghA7uxWtIgsqU+QID8o3j5oOLqfp754BNlLskeTg
wsyVUgJ//QgROub3+uQYNYgr9LsaQf6TrRF+Akc2xu3dKSUbx4s8RhX6g5T5MWzz
NyLXTpGL2Qwgkk+Epf9am4QPFe7v3bJhDsNXFfvnebmj5NVsvu2fVoPB0jl9uEBT
d1tEs/ENTLqatpuDCUz0HSqB6QseuX3VxoOBseWcXBAvbskxqHGSZThbQoe5s0v8
BJzvzTZBCkTLj+JhuCGY9bu2frTM292W9/ONZvkbE4mocXzxCcr4ae/DU9INyJZo
gCtixPXSZQ+E6G2yB3HcWoNGa5i/XpKbXoZo2kay/Fj9fgk0b+VETAwJ9BA7cSYV
jN6W4fsWfg+WxtWGEsh1T1HJeNtDe5dW2XEDBPJtPqhUbVm2w0qZEr2hprLMeJkl
R04+rKIZW9OqovitSHwxUKQsU/fh6Z5I7MsFDV9EUeRFl2obR6AGFZ/nSImOgg2E
3llfL38T7QAk/lqPpOYZajh3KJTjk1Vc33BeCV8cO178iCqERg/2x2PFtqap6usr
r/R/pdu8YB9oTH2pqgIs49XJOzThHKtIqT/WM3x4vD39ZEbQ+ra60IHwa1lKwFjT
SQjlYFI8Ul5MgONSJy6v435RN2XsPGLeMBV0ocYI5Ys0Rxl8EMMcDrVaIfKSWMZ1
D13HPKISDdFjUyfHHSVr0J6L8QImXa7B6tG9w5oh1zFgrsCz3iAbp5lvTO2sEn5c
GfPN1c/wOOOXaC3hiBDRlE7dY0mIuiLFjrBg8rPlh7/lY7ebCV8fCq6yKDVVX+Ir
cDLTimi8QYNKhMzETa0fTtAY7vRCnT+KS2tvzAdTmDpCQevZmbd1E5U3Uz+8KBnP
Xt+Ymc0mjNwag5wFXb5AlbyejoSY8ipmrsqwmQQyncXl5XTnlFFrXuLpjm8Lgd5x
9/qvXzF6R639dCo2BhJtjlviwcNCFTZVe8WNB4sxIuiBQZqaTAc4vFtA416VoE1o
FOHPXLVxWpVEVhqpk8Ohx+B6yyiLUXSBa/QJuQof+QAkk8fm9cwscUGG5btXEz0i
ruto9cXCtjGl7XjJxVIB2ONbfnBJdrcQVXV6Pa7fepCdEKbg6tUo7ZEkk2s3WRQ9
dSRi6NmL+5tkAJQREMfktNM3H+rGEv1Jm8jTowxHiY0KNiRFFiQJ/ux8yiPWfyk2
bxV0Q1ZRAFVqxUFzqjk2upBvrtKZtp3MbXV+nrN8nme8Ke5Claro93nuHmo1aF98
BM0pM2i+RYHT3Wq9QnsfdspTJhIIhxqd0qDGeXxeuBWTM3XiYH/VuMPFIgM8NIlA
79lnV0PC2o/VLqU8fmqLtHZRXtW8cOg4t+xxG0b+NOoSMT/kcOWO8g3MxZjZrgUR
Fj3JXOKxwdbXKFRg9XBLUNKKjU45FgQTjMDLpgektjrcgUFRc9rleKsPeGNdzquc
qayeQtIxEQPfOuSlrFzcims5DbSv6H/qjXkGyPMjbwvjvhRl1UQzvYdhrMJjvpP7
wip+RDYYOINpNwEH3gvTVNlbNhjFg9M7/XHsRChzJ7CnDTLI6+AvIwZr9vwA1JL4
LnVpJugRlcA/8AqDv8djDM8AzUcxIgsf62XPOv8e8YIGea2lMG56V5gT4VvnlGHH
GqEHxdRYtuXZevjxXLQTq2NPbKuj3NcNEdDbHJ9HU8yIn39PHdG8Vk4RyH1LAIWO
0XukDNrwktUJr8mZOTXmci1jlSZDntd/oQVa291OB/uNK0ZCUZs5RE2F2Cx1eZp2
GrG8+y1v9/8kN61OyzdV3B0NX3ojln759m57xaxamkKhDERcSzZG4guFacqswoGh
BIj4O+YG4gBEQXSL1cr1YatiuLBAL8EVfCN8d+FJr0bI4rgBpWiKZoFLEmD1dkKE
c7yANQ5Iw5lLDnDdMoXnMDUkB5HvwH0INKHSdSQ/rgSiH7hdRisQ1rwJ+sT8NiCj
K1QQvyMhaplbOhB/FSpvK94Ryx7Z/KVe8OVbthw01KpFeAPn7Wu2tJFHCOujR4S3
j+LZHQhvemCoiVbmtwGODrjKfDiQxIQz3vCciTTLZ7qPVbqcJzpXcpkSnFz1MfLC
eZ/MGXtPiPAkMCOUTZExgpl9cHaICvWbgc/w+E8GbwJS2fefL9fhXAxWxsBgK0lw
4S+W3lWQ0tQrUElbekZ1aAv56S5QGvFAEU6cFlXY3HM68BV4gleoiKgRJ31PaLFZ
f3J0e920ApsY3p4INmlzux2gcr0XGHkepGlkGUmKPI4eJly9ZrNwWDh7oximgax1
6T/UbbhdeprB4+7bTNxZOpQTI1D72uVD46J8/EttdorxWsYR0/oZaB6ik9kgm5ZR
nI3nx7ZnVqKd5C5CtMYEgN/vfP5OUKQG8d++HkpM/fRs4IPZuP+ubjfThu6RV/U5
43KGv7hwARV0asHM6kDDHShuccn+/lMywjKFKwmEl3npx5SNgY/Dra8xDEs2N9rn
9jevdz0scW1/bwSZkl8nsUJpBMvI3Tg88GP9meHBIFuQfqHvqEgjySf19Z9JRRnt
FNBX9suDlHGbAyDDHvvthb7mvN2OxKrHNAcN85YaEii+XLmPjDnEk0BCeKAEIZim
rvfmN9yBDIu/gkcjgoewejvWTFh4/exhi9IlH26ZfhOMBte1iXGLgNawY8lSdsi9
Zh/2lOfm28XOh+nOBuBC3DswJwbGQPaS7oa+a993uiq56xAbZ/EDW1ChrEW44yYo
mwqOpPTGG4wK8skB65J+OQolxLmCC+OR3gLyCV6JPFGLSoPVQ+uSqdloSV3HJEhy
VHJgvxingmI9yUU6zFn6mKgJspLxlN/SANZjoTdyRrokwY0zdppEGTc4rtkYpiyg
32X6GTGHO28cZnY4ydBH7q8o39balvcW2XNcIlECOsiBSJGUP7wGW78wE/yT8a4J
2pQiuqNm6ZBKLfLR4iPg9tOkfFY2qMf3w88SlxGUBGRwm5IDGP73vfSZQzpNYW5U
4lUV6Nu1c5m1+UoacJGtrr0JIS9a/iIS5OeICZQEHipPFP/e9GLL3VV3uz2ONKki
T135EV1aNoTm6l7K6a6g8QIu6ZBDUXE0B1vlEbNxaOReueIKn/1XooMaPKVDpVMy
1NhNisyx7c+ZGD8nTTcMb29zgknrSBGSjNu+xd1ocsTpXop6ufurISnDtiPekC94
xZWa2Z8sO5zryQi5A6V4G7Xxw9zjecf6OTQOytPyySLyvIpPQzEFQYwNXIpvREfP
OMlyec2EUA9f9AJmRzNze5+Nu1e5Y/+fy6xfriEMi0r4Y6dcqhqs+ElHBtlnh1Vj
D7TQYwEPBq9idCX6rdjstvq6bVQxJ+EHluH8510ggoIk5lZa1ld2UmO9AB3qy7vt
hcigsdhbNHW0mAaZh77Dp9YYgQtWE+vgX/T4nwKK+yxmUoFUZzxgXNUYffoMljPu
XhLfbU+Fiebpc4Y5Eqe9/Lam854RSXIM1fthUy4+miDir2OS1XYtVsEmgdo+oxCc
bV/UvnjuQRn2dOPgK9GKfzDL4/Smu7b8pzxX6SZlySoZgcGLpUgjJ/1CSkVaIC/U
YHG2todj/0d1F0QZJskrc7EGrrTFflbp2dsgskTi/USNi9ndnsNyVi+H6PXmPWJp
tXRACUcpnFmBCyt+MrzUE71qkeXDEYJ3CO7C8dfs2EmjosGfa/qt073C8j9COphm
Nj7ha5xcjhnX0p4vrHMjtKfkQWAQ0Ysjs/iPXq5AgZYgIfAMnRmZtrlpF6kGBoaW
3CaxWRjfzYFFxH09WEFcLYv3C594Kf2FgxS6/JcAmfAHSZpATJNLNwv5hiNoITbC
lgWyv9CJAMJm2hy9nOjV/IdQsQYRQmDKMe8IeDfqr6i2p1YRvB9zYQkRg5dXM1HC
YmIytJm//r8wqc/5RtbrYZNUYb7KXq9GdZYdN2OZDJTFY7zqu0Vd6aKuV3A9ik5B
NXtKPyeu04JSJEP6DUk/yfe1E6IxWWL6JaVXshw6iE6tX5s9/KxuVsHXAl1/z6bj
8wE3yBlTJLP5ZDiJbYZHgj2xXhZ2W6LXGiXrAEbaOcubEEo8kac1FZ10mS1oBZLZ
3dhX4ZSdFt0fZBofAwdmdd6848NFv456sS9jN2akqJfKHdEOx1zygdAZD7te9EdX
CyXnBsbo0c4s7xsf0K8/Ks7CIlsdo9IsU8nQOQeG8IXZzhWcx9JVDUIwAmiBCzx6
SpApjon41zF6e7DBGksnL3Mc1nYur/SMl6nAQTbNdA7gCrT5FmRJdEwIyUoEJoRM
qh/0zNn7CBrO3+6xECFwFqmqfkeItHxe8Doq25TfMAl9mPLndg5rSJe358ywBuTS
m/s7jBpYFo0M7kQBw01w0WBn/N5cWfcJNhi6I6qWehTsLfSTk/yhUBG6zsUuhJwf
n/D393sYEK4hWywHiOd59LCbrOG0vuc2qtvJk259u1GpHy+ld9e/6ICHTd703a24
7AYlcJHv54fg5ktD42920oT4/MkjMkn/pl5qK8og5nTgwOa/GmljKKAQLHFVX2p5
QMSldGYuXltV29u7KVgfeYAa5zbvj4zCq0egbFHXjOhr+scYAsIYoYPmge3+gt+B
wVLVjC7zM7tlMzzi68hRp099eBNr9nQS3Rz5Ib0PgcceR/pXJux+zv2OD15h6bky
eonyIV+jp++nzYwE5yI6DTj2TLOriPF+rfp3swVLTExsb1JmNytHz/xOw9+HozaG
b1nT+/jI04VFYqbk6t0IWDb9rGBvoQKrfxZO8FpFuGwsdy3/2+Uwy+ii652CLMjf
Y9InaU9YGhAoclsG4uu0YhGufaLRVBBOSEHyIEeehcVKkFC+JoPttw5M4JkOKR9w
DFPXBbUiQkf9SD8H18EwjW4lqdRQ31XJYWOohFB4AEg9HyyMsn3UGVje+gUF1Pmr
QPj3zw+m1z1SVlO/O7HqGR4FCa0RTv1QcHDJgHcTDLvBMx/3wWw7P6d/sk/CjbDt
mN35NtfGo8HBvg/y9VZ76DYK53qRfRzi1uvv33CYRY/aqOz3wkZPCbNPG2PvNeBm
WPdQ5YS/HCA3c+AkCJ48kgpwIymDm758PIbkecqpL+gpiBGiuqkoDigZxnxJRy16
RKhLycSF0SAWircMbGdUpxbrR0VXx6hc28j0URgEFrJvuSyviTDupNAbTU9a/tDK
QulkKBfxFv5w9Q6xC1AGwgEVUEqRZFbIkOQUul0dAjvLaht3vSVHG+VaSIYiuglH
TNbeDGJqAtAmiB4dqs8GcLFbfufBMWc+rxN97UGk+eptB3v2ljxQybA6x1+hOSbm
xqm8wb+BguPM/FjZXcksZBe3AKdpncXP+nHh1iignN0kbhCeJMidX3+cobJ4wagZ
5ve46OobQ5VDHWaNLmmp+bo383JDFSBpTOOj6NuHKAU0TOzieNNG+DxWWc0iHQ7P
6l7aD/lv9uDeBbWH2lCCuuCL+l/p9AHT/DKcuV2vQphuqICVA99n03THIsPvbHB6
wA2pv5iKSNug0I7FRy7A/PfTAkJc0thIfIFzQliTl217lyr7i/zxVCpQdcagdtxo
C25eAIh3N/TqeuhSZ9q+dO0zo1DQKQ7WzGIKZQtqvdp2S6RoKAl0LMeh3U2SFGsU
uStWa3HYhluvmSS4+XU4zEAZ4btfuWVdybPRuy0RDji6+ygn9UREVr2NyWRMhM/5
zJ0+8snDbLj0l3P26ATAHhEFScu0+P7LG/3dMDUqy2IItSJJAgTx9QgP8gfPhpBp
EZEKbB13WbhYK7eJ/PYG4gFOORkZhum/yha6hfziPPO9HmMkA+oZH8OhypYrxK3j
ZT52hWlMoiygMDq3Oulvkj4KWx7ta17zzwGpee1l+dmpppxzSZFREIq7573c+6Kx
VnluH6rsCpVALBtR3rzwcf6WQkm8vY4PQ13KLI+rmja5DK+/5K9B5K+T/Vf/VrU3
6KNmpYqgt7yAelVm9DgVjLoT/LZMofIxYc2v/+IWIcOCaEYfkw6viejqs32CUYlD
ey36RHl/+ZkTx2uqkebTz/Ejbnmm+6E6hawUeac5hZ2at7QVDIVeIqU4LTOcgTCe
KXF3QZz/MhYAkI571YOAlrab79trxO1zkKKD8xDBuNL18oJGguNwFq8/VYTz6wWd
ZNWHPlLNJspKX4HMmz6StinmlpZ8d9T/T6wDkaM/JIT/sVixQHTGrN7Swr97lu56
ie7zxHmbPVB4Z7wf4KKz4dy1RvlvbKZ/tyNnOCfaG/u7hIwBDxvvpOshA8J7xHOE
TaM9EUgrYKXARsQXzjS3y4TA0l3R+GhPkisfEik0XARLKhgfkkPT5HxTx/9Ov9E7
KBf9/g6fUObuVl6ZjVgwkbl9OljjiojJrKjJQAnOoJgoFqu3+fNPf2MWLf0WxjRA
JLYUmCCS+ubjPMP+DlZxQy5/LLMSNFfHr4+hMm7zlSB64a1y1e78VruZb0bbU3DK
i5sOtJErQvgjNWdzh32XACoLnJp+89eFj6FMviSO6HNaQTxck5e6ud8E95srJ85F
gC7cj5T35ml3IBQnGmDFAh/PGa4qIC/M7dEVVueii0XGBKqlGsQsI4CVCIN4xCxk
4Pi2NKl/9BLaxBL3pjA+bNu/DB3zDnpqhURdBGjAd/42B0Gy99ftAgbYeqtNZ1pn
MkTiqw402WHT24STrWtf0hFJAIlW+b1/h46kwfQmd+Zw++Uzd5GngMybWl+wOm43
IY2eKGTDVtsCdsoj0jjT1MbLcFmpPg1LV/ynCwm99S6H7GzoFVjsqf1c4bkFpYbA
FAMs2Lui6+tCoP30zC29Q45Oa6kiSjWB5/OhEBMJqdV5+tEzkClmYLeVhqhOrEsp
3Kdzzu6WTqc8+RyJEnjw1xSj/eI9zg5msMwoINTEs27QkdJV6/+ZgaweCGAh7HoW
Po4LMY+YeXhXCXD97F6h/2HkGsDXgvbGoKz+fyuqZG/gXw79FmodQNn9kOMOxNPV
UvOGXe2Lo7Ji/OzcHUraJFSt87GJ8zgPQD4dqFYirbONwO4NlMoocJYEFpwFCVkC
Lg821KgsCXU2ZtpY6RQvh5HApd7y4CrrY1r8M/7brbkKs011ZYod2YXXnBRX1X1b
fa5FwShxKthCjFe2Lhbb/CPqFG8V77NHvaZjabwqIDgKdBnJYL30Z1BJScprezSz
QReddDYdtM47l2L3/1JZ+gWUUw2pnAddyO97SOcqXQi2ps46VRGFXl5W8bx+oo2D
ePTOI8O9bfP4rjjO8LUo5gnWiafxxAkCZzQPhNlD4AbPLQCekzrdCRPzxiScXq3b
WWblvipOOnFBof2VmORX/yn84XBEvfxLudxKLFQwDtI32KIhZaqBUbkXTwtCen74
UxCNSoKox9V/bXJwRVYn+PeR0PTXYGhPJ/kwzw5LumKNX63JTtduO2BbNytWzE9T
/8wRfk00xugRp2MhupsufzDWp6iYgFtr7Tlm6bLVqYfhx2lv3yhgavwPuM1+w48I
mM8hsEL8CaA29ncS3HIXD0iaUGvxfQGGwvAwtryZU+EDjl1/++vLlKKBwCVUIUp3
AzLXN6+kU0Wys4vfiOQUoYp6HglUJxFL+6zgKc45nRUIkKtLr2tUhYwIm9C+/l49
yiP/dZ6oIGjjxGdSiXdyr60TnbLSxDzB18hvmzJQEUAisF2iwkzRJuBLFq8UDvzc
QfxE7zsC8hUE0L7FMUSiFwnHyIRWclrLEDuEoEC2FV2SnMi3dAywP3UqFi/mQOu5
AU8/mhGSylEcBH4SJ8IvyMaJO0Lpd+W8/zBSQiUg0y0CxxWGLROpCLgfW2mf0Lli
rNb0wHjDB/2FeC/aM3COsbak4+yks9QYgz2uWpEBe9CL2FcGn1Yz5hGVRjFoxzES
ket5yQMJUgLqZVLAsjIPge2B4YeNG+K6j3BjyfDQgceHlW1fP2KvpsPMohBqD0+q
WycqMY/eoXCXeTsJEM8gBvv5NgvbgAd1DwTSVvOi40jofxyJGlMhOdou9f43d+m7
CjyV8qInaOktMSLoyU3zYyvOBNM3HGTSIYW10/wIusYvrLFSDfewGmMMUdanJIDi
uZ5evbNZbONB9V8SNrc0a2BFgvNwe071yPkuYrRCgQobNXjvJh+LpZy0SoJGARjC
Nz99map0iW7GGIR34PB0OxIkhCWMCY/n7YJVHz0s/eEPypRtdsKKX3T/0AZHFq2H
kt2JJoEShBDXpSe/P1pa+aG4WhOHmYHTEsHKUCUj3y0FUHVBMPK0ibqt5hbuNDZw
B+9pWDsJOoifeuzDrabLIRkGXIfPfR8Fcz0ZdU3gpDCWxkLosJ67HuXiSzFf/m7V
W9YWsTifcAScIy5+A6ZroL1KEtQLSEKYRW5vWj3TC1GhAAvv/+IbiNQ2O/4Lo0dN
f1YKO7J/NukyvCfxIEL4Zi0gNgIcQbi08zocp85VNlxfdh52m6qZj4UT+Vu9qaMs
B6P+urspLsNDjb7E7laNQ7DDW8j05mu5kH8TNFR4r9PmSavVQHL1tT7T4J9vM4GZ
5bLVXT9EGA/cks9hJsLDqlZpqo57fB/tVH/kdtXUbWBPqoqOLDzyTwc4OZZ/3Z5g
3jO0sM8NxYQfDY/Ok3upcQOfD/ivt59EyuYW9oiLJ7Qf9TsfisCGRWpvZcsyqHoy
82d8NEl97ZXs7P3ybXR9NrGFsZAKwsC9GAavQcYS3cUNJTxYr5xmJeqlmNa0Qm4Q
c6Gd9GUUQ4858AZocSTJL18WmpYcL9UEom+XGlsppHI/mvKOeLnf/znXMpHg4PyN
HDvSyTwZUsLKtujj6argSbSvTjA1VUUiYvdIApz+66tCNSVEsVlP56+o7poXu5zn
Oz2iHdHvI4hM72K8j2xY34Uj253JGmzsyRCyqJgPifG0WYRGIY50KdcOisspBF7g
BYMUpbzdYqWQo7ZjRZaAahcUGpkW540evULwiTCXxKm2mF/AUQsB4I23fmQ6rwKt
YtUmIXlV7+5GB4Ug0XtyU9rKyfHqHBO4UmBksMytLSaqPUgujBOCwSQATEzjyDdn
PP/gyGnlm5sARS8dn435eLlj/eS0f08taQLejM659CLSq5ovZfNtSXtr2VGOixZo
3km5P4loMO3B6GhWurZl2+ZEWbYpaFInbV4aswWGrj74VZ7Aeg+qtCd5qQltv1UU
Q7nfsj4PaaUz2lUnnkAOHpRCO+aM5qnaD6l1PcjemsD0KCMGUY9C4IAA+h6ryDhj
W6mhcnUeewWeoCdVuAg4C5Ghf97iNMPlX2fmfugLoNZGteBdM67frRRwhtIbFsZ0
NbI4pllQu/OL9TTUxv/lVy259f2kWqkcE931Boiv4VjjtEnLx7BFgYTvmFWGI27a
pSJ/DDE47owpsIBzfKjxyQVOrKdPl6msj44QR3HmH2uTrbenDg2BxbVnRVHNf79x
jcTRAkYCZPIDZjciey9GBYCnA40qLvbJiZt9IIyD2pgn5jFhJFLuIUX6PmrCz9SO
MaCTM8ybhjzIFfrDo7cU4lrIyqHcFjEhXKtScZJ2bAzYPKrs2VuEnbtsQ+t/05RA
Dxjm5nBOpn6HB+Xo9yfVfPIykkgTfn8yBnjSs/G8f4pevp+lxyzteSiEc4b0uGQw
yONYz/GIstqxyy1BL5YQQCh1VOjm/RB3oFvYdLsImMzTIq6/wFy+LGWT8uLId6xw
UQ4N7dorNxeNYuXLILCaMYSOluJBxdgg/cNPFr2TW8mUj4MyT7K8Y8aByg1jK0IW
5aXGYRZOjpHnXeFLInIYolwuhsuXVk+nAGtu8fuqcB4t+agEeeU3Wjky4I0H+0g9
Uu8bBgqCGMffEsQT4kI2SlEaphnswR7FWDBfelJ3AwkW9G7fS04ASRpSlFq5lKiH
xkFsDYswm8OpkGYHDJAZdrRgfQ3ERGGIwEZ1O2hpqVWuvsFbMD63KEetIcwE8FHN
JR2mo0fjVak1bn/lUKDGpY9josSRERgvU8iGFXZJNSD4UgBuMefBz3/4CZJrVKot
qwJGejQP0YUBkVq+rl1ohOBccOMGiViVQDyaCdZVMmyUXoTtEdDBrcXZcsZNDARe
4xIlCu/46U8ZiZkc/ey3Gv5hOHOHOcLFUrroAaz3cukEQEsPsSfuM8Yqov11EZs4
RZb3eSywz7tO+nh6Vo1P3bxZ7wSEsgZhw1VKTd6DUzfVBiVjF1qN2m4t15pz+EwN
pzmyvfTn2UcmuEcVF6m0IEQjgT2b7SHwgICAlhFp9pq9lmjJPxnEGzLCnkkblDWV
6xrYBxslg6wNqHcmVeEmMg2Bj2D7795IThw8oDVjxSK3oJNgs71wmVQqmDsAmcII
xuGKBsdA+0muoXckh0x77GiFDKbwH2rZYEhnAwzOkAlpeVVL94hBDG1obJb5wC2j
74hT/27XZwHikhpDb3zVtzJTuy9/fGyFJzMWjZarCJ7VZAJZ2UhWDNzxWK+U2JdH
DoO9t2l62ENj/tIx46jXIPiiGDUasO8YFsWjMO6S+CoWGtRUJKVi2nunBBtpOKr0
AU5dot739lOx1dSFLdFXcqDnoX2E3T6WDdfm9NizEa4bdeXwuvj9U5rNutdEX9zr
764Cv/rWMO+8DvxLdxJETmj9kjxqYnaZtz7P1lQZwY42T0pctCvIH02R/G5Dm/I1
rRAERNzrzpFioDQGN6573+UbHnFz0bLeKXeu2gtG5Opi84fP8RIViK3umGsdOqr7
vp4j9tcmoTvlRJ3fWxsg1UsxWT0wOXOP28hh3Bn7wvPi1GDrx99TYRPLpWNPw7WW
nRS9oTCDU56L15EbEsfSGu/9IEgwmSrCFQ8XDITU0tE3PgIBPAcWxU3NOIM8uo8c
JEbqNTJ+tu/hQ+jBribJ5HWatd8/6cACwE+HPBZg4ZK/wiGKYZOZnnaf9xJfXko6
nkm8V1w2dLgNDtHphDGcvK37Mgl9q3Lv/PqhNgwGrj/aGpeW6vgAEg+Dt+v5RZkw
h4m+3aq6OXswGywyZVp5dO90mkm7+b8Xf69+/Vv52fKx8ArWkOUKYXIVajGUN6P0
58oKcEGl8ZBJDIE5Yh55uCGAe+hR2u6iv8I8yMhC3i17G/j049N1YtGpd9iv5bdZ
KBdihjQ3rlgq7PEBb9wo4maOGmnTfq0Rvaj6Up2im9jKNX24VAsyDy77oaEkRlvG
GByBUKiDXyugjqIu7n8Xww4F6ey3R2e303nSx22vRsALqpql4Aheh3dDDzMpmabs
jCpJ/JrhlU/l3AYux04macp9xYohky/VehtyW7k/RAMoCiK33B2lQgM7xuOjuo81
oTuXGe0KJcXhWiG1FzFqmB4Z2OESr9xQYuemZkTu6vud+V5k37cQKW6FkYiBOtr7
N6E7YqGwkL4T1HaQz7li/xWY8w5ZNdX/Elww82aTfPxjwiK1ILENVFYDneXK6lRL
cxYsEBDm36Yv/G3EDOBZ9O1Y/nBJLZb6ePJEvJnbqxCFAIrFNR4u5eC5Vv27pkzp
xLfgofj/9lSFB9dDiC9nfcsGHawqKPdoK1Wgj2HTUVIOH9SvSHUvQwHNTthX2AAc
Q3l2j1dvl7R432P4p6cLObDLnu7igInuvTBR5llCGHExQoJzMRh/wmQS3vq2BTy0
s7CAPixvRhmIHUV2o3un53m8IkpEPysovYvqShSwrzxO/9mWllrI/qB9+0clHJUR
KMoWQ4asZETLyb7aI9EC9DwW4OvjD/xwaAH+gRCtsmqdRT8imn1fCAif+/ZjrmFC
CLbVuo7G5xeQbcTIxObrP3Sl0WlAPTjuEElY227HGeu88Cl0q0JtFlKeGTSkaK5K
MGHKTznnLA2YJpyh/0GJznbsLt6rBZqWvCWqn0OYwFzUVbSZxywp55k8WhAH83/k
lapu1SIo/Edh30ouOzxQ4YAmGeGuCsVtZPE8EHzzE6B+n0u4JPDvFiEBK7jotWdM
JerxgicMbLc490DuxBZNdNwXysov4DFUG89HmJ3965Fu7k8OX1ANFXLsgOVZguo4
d+RSjcQRwgJ9+W/Aol2JjujkPZ0L7BstdIp4IWdIFUopZoqsv6MhJOEAbLkpv/2w
/wxi1szPFaJLy1SVcKoqyRDTDDm76K91bwT/3khAXZ+KPHBDcfwm23aN3e+nVL5Y
wj9cfd2dkv9hiyfzgV64igheVEh8C855NjIsW+QIBf2tRCNA8+180VIIdVeZcBcD
zWSe8h2Io9ylZMMYHTcBIJgM9qA5uj1jpshBwaPyxqMcbZZdCQwbsfS9RgWEmWvb
91zsCSKEqcllfa2LRGc9Jf9O2NgYnZcp7+EEJ+ks6ei0I8FQYmE3SjcCdBxx9LB4
FLj9S04pD7fQKrsvDuCpoMMJl7aPewwYdq6/1nshTNwv1LOMPVJwBrEZ/7KLIIqr
tzzAnu9IK6WF/95+6WpgHZjQju0kptoePb/Js+TVavcZXRnLjaep0mCh+Ns4qkVU
QXXI/dOz5fVLo6YQhpxVjwLaM/Z1Bz6XiKGhkMCas6Rxbw/+zkrb9HBu66XHUwFg
Kmhqojs3iKHIJiCNxDKZtbgZm5XOoWITBUg4A78CNhe2CWmckof07G7pTdbMK55L
0JG367LqwfRPvN3GwcA4NELSmP5iZTBQraO/WcES1QnQuHXRfBRCdIn1dYT93l4m
tLP9alrc7zCsB0aMBrLl8rk/F+Ke+zJBahJtMs8Wn611l4zwW36QIQ8+ooxnWinU
eRSayQ6+j+Zs5IPJdfrH0Tcpbqe1IgZ9wiOcRms+FmT9vDexWVfdP3/bNCQwm2rJ
sbfcNQpShe7jihYQSOkLIZFV4lfOKYoVKRi4rO5TuBDGCDnlkWpo+iVIk/2kQYXt
z1Cr1Qmgzpl3TUHeFZ5WMYcFVPS7FJ+sHgH7cQIKyTYwv63JOg3VGRQL5lSCbc9k
WfQ0fAC4uYQRYVcqRJRbHZKyZRDNEE1EHR9fTc3GZ6Dq/HuZdg3xFH9xvJ6Gd3XV
m1CW+S7LIwr+UlzoFHzK4dq+1dsRLVZsW6bvRbKAqLPVRB0++eA3sMEo3wyo83++
c0DZmYNja/gwcE5fSRgFELq0lohmOi6+RyIlH2i1NcUNv7Td9Hz3+Hr7n3PDtcXL
2l7woARV4W+3f8DsIfy7YPVKy7KJPlLtnjlS0WLt0ol47Z2SRo70ImlYOb9BMOCP
0QsqxIf1MjDWfcUFlvRVtvade1CGZR+m4d6sndJB9847X5+KLaDkk6T9XoeD0akB
NmQKz3UgV0onFLI02OLthJWnQgbAlxinU7PF7myvsM8ly6UT3VCkMOLJ/eq9Ilul
flZu1oKO3+MIFgrlizok7x8bQqWyGiK+lrxPwpinZihOg5VlCIsddU9mMukpK5sI
fPhV9vs/yWNgknhs9QdIoTdspLk6ZgsprUbvZVi2C05xASbxHiTx6ZgJGcR7xix3
hwHqztrV2Wx5UL2WkrfaiYKDdDci5Y4mp24tX6onp2pq4qNQR1MVmA+iR3qPUR+T
U3rTX8gZz4wWis5lYBpp/5BBViXjBeZf6zLwPBrVaDV0zBcdq+Z6ND74h/0IuBMt
Z5hzM76ZXXSsziWFPx9d1tVssWYlnItLfRpl8/hqbcg/WvXUL7wbF4cdeOzcUHjV
0/AUfiw4TBlqKwnjUOgs8iJ2VgBidLI6sdn4S/nCI8sxyyk+338zCjMIoEwWU3cC
46uF5iNHlRUiG82qNVqiojKH7oNdF/gwG0iB4GEs2uJS7CsnZ2LJH8d2XKd+RagF
8Wh89CDG1bd1rI9KzIubjWPljBEKgy3Fk4wWf3pxZkxOMfSvVHhMmtxaRE3Dfp47
ahLyfjfozl1DOxjVPkGCVi+JGQ9jNiHqf6HEjyu7Wt8TcQ+nRjq9dUVmx3+eowot
fMR6UCqlypUPuHVjYoN63fFk5jm9XGaqnzed7qGWOVYkjeolsb/LyfKsbxwXv0Pg
KlsRTizpw2HQ6VJC2CjNQprOBvIMUT/dJgHEB2XWeM352a0tZ/uuXK7v1VfAErYY
/rvlQiRkdkv4n/h3ZhYHnCUWKfpkT8Y/EvRaiJiZz4sJDz5UZ4YTlwrNrKCDwp+m
9JNSdtRxgCqtL2CgS31wjcNpc15YE3wglBwTpsXwJoeO7Nirv0ZB/T5Q6CUwxq4C
/c3d+R3xG1t3Rl1DSOKHkJ4ACRtImUrJgCHa8Jf1aP6wFwPNCx/3AVrJvGq/UiXt
w4USsrVo1fIPz23ZOR/918jxtHoKyzPz1EHrIw5I+htLxXgPx9jllegOfXjm3QHq
PDl9DDJSKv20Kge3tYGGbjuwsZU4bcR8g0G4fe7EZb7efeP5ZOQRt1wNK+ZPrccN
ZjCKk2+Fe+IoKLNpQCEkxf/MxFMdKm3cxVZR5aWMLNj3KYdv+/KG8zbdikQh1MVM
mS4dsVyWqKM4jLRzoPGeQWMw0HzbqxJwYR8dcxFzSU6rhfCieUqIcHIYrd+L9AfE
nRNLsGjAjnRWCZVsIdouhxH49WmKupGn/ypHe+wYnBJ78IpP+3Wpu35Jxrx40biZ
S9YA2u5yVP1sa+XroXcAPW5CdvnzfCu1imAzSOuPA25+K5g86zJLVhAp6pdjdKzW
BH590zSu9PVqGABu9RaimHfvO6Z6ARwfiqxgJc3XaYTvr5us5fZFg+bg5Aae6vLi
RpiiVN1cSMJCoxpnp0xB5RMajksLe1DI9o1dQeNIW6L+7QWKDKkf3VlG5ahzcCnP
NXRCUM+0sS7wU/ZXdbxNBhuq3AnqisH7YoZlyfcjU/IFrb8FhDKPFcjoTfXlWTIP
5XsjfOV729DwBG6jk7gr9x5WABWCxhsr7vOj/qr4WzMrdA3ip2AqlsAZX2Rsxycz
/yJzrscC6CgepD5o2z/9YRy5/xi+M2e2v0BF0B6ou5JYXrazsLEbxbjcX3P/XqxO
Be1dx1+yJtigPGkiVfHDlmA75DrEDz73Im0G7NDGL3L15SbDHB4NHCswzzxzXTBW
9nNBFD9cZ2IoSxabRro8bN/clh2OPhEzi1FcE1cXZIuFE99rHLhnLuVO7uDuyqTd
rCoZ3Lr6R/PSXuxibIbOtqydMisw6mkaZ7ZQ4Tf9+gvC7e6/c6iEE7rMFQWYS2cx
XjqcO7w+UR6eLLQ8tWv5bvJuz0x93Sv+wkTr+UV4h4YLZzyaTervAJXJvlqb5vFo
5nHV2U5JQNHFjRs3sBTrBgmoNgYxbbsF8h0x1j3uSGZnvriP4P5TNAzpdulM3+da
T3QVHDBPm2NSzMch/veHKWiTfofWrR0IlFmXyZAuGlUJMQ/I4K29FnLA2FmxJY4W
LO+/D3eiatFA+Jn+SwLk1k2u8Q8JCQd/uP2pnWRXdixQVah27iPdtSOhrIOpJ+ve
ObgWnj4a2Xy8V8klktppM1K05fbX8wZVc+fV7f/1DZNeAbb3U2ULu9JP5mUQKufv
K9F8Dhx+1cULrcdX3ghpJcz2UrgY5+QLFdlRU9cL1PbsjhGj/JNxorIHpK7fxi63
+KsMD7TexSNnwHrb9uqy0iSvnCjY+LO+uJe3KRNbUwGaiQqppuDAxO7ZGl/mfBYj
YHsz3Q508XIXzGbdLVOQMM6kVCrbcBLNV7vqJeM+3NfBUCKjZQLnHq4xFMqvhRtE
MXWy3IFRt/qt8E3V47W5FXivzhFZNKFCp4ndKQwhVGfy9AueJhTRasnz53AP61dg
laIB1lXrH3WaMbRpFHX8ehnlXXBTllqzSfraGC3BoTkzZvxVceuSQxo5fhNp3IRT
L0jCyo3NVXuQOlqYKP2APCZxCwg8HaSgpFrvlqUdaZ8DEbytNEVxV2dDwXgzjMNQ
ul/zXv/1HL1/HvDkhbYdFv3ZK+OnTWd2TS8JyUfPuX/gW0csvLetxVvx1Uaw37xq
wOQ1cOxOs5PAIhMQsj2GZskutzBdc5tuXpIWR2x9/KlH79Yjdg8wxpk9zxX8aHHq
gaGdMDxXfVa4w/+pkv7EDUMXebMCpisb0mrn5FWD04ctBQwRErOYBkKDGLhpvapL
aQPoDgLW3VH4feQ0Z49pyITCW7OIkNRcKGe8qpbXCFfjf36idkrxO1pE6fX1d4T0
9lBTTF7E0cd/6oZcImuaS6gJ0h8SNqVRJb5uFjNHhUdqxT0vfWNEQTqJZEM2JqYL
WFlA0TLV2CCrkVWIw7OZeXXNXB2Sz7RcwxSlEAGHwcUKZkPJ5GPtmYNGSk0xsEpW
VMeHBbzPEqSFnj9ZLQng3J7CUnoHvO+MBV0MXanD/NWDXWYZNahg5mI51vgCnjsH
jvMbeLVMG4R7agiocY6ZRE38w0WV6tA9MV9qhH5hs4aihuX7bZrsOj32WWjFaE6r
G2Qg1R6W+Z3VR3Yrr1sCELJ+uPL5O4aqORo0LgxPssD7cn6M/A5Asp44I4verQ6S
IUPDepJIule6lrQzKrnYT8qwCU6fRyMmbZDrSuCsZtHTjb+BN+ZCLyO2zHBs7Ker
A1lbrIok/wT/N+bH2T3BA1Zxax36Fy8ZjCqVz4go8aPsORYNVD0oIUrpRbR/RtNi
4p9sm/o9aQxr9DO+HXpS/ATLzcvXXRn6lveOFdY9o5DobWFvztnl7eypB6LlyA/3
lTwyG5kuortDss0PfiEe4+/LwJIfR8BCJecTuB5C70O1q4yAFMxLKnxQ+Ba0p+8i
d0OvOLuP9oybLdnmUd+GecGUT+KHuGXGTlqjN/H66Dncj3xZNHxxlt4Mj0SVKV2c
3wJXrk3SuiAkio9Pydfd5vz2NCiBKb8h2zwN4HDlYBzXlejp7nazhPvKyRGZ0T5r
SAEZLmw0/ypYKSOBoG7tjvKzygK5/BoTEyeZJKe+8yvFJnVvpZ60vy1+pyp/S7gq
LQJ4Kjv7lZQvsRl4+ptvvQJ8qx82L5y8BYVjfK5kupkTyUehYJk87qoqmxWZkNi0
neFQBF/BjaUFlLw8rr4KTOsK0zj0WhxioyjDwb6ThW9odLCzR1LgWAg53DLh+dyu
WzchJfCY81s/e2qcKOZv4ooui9SJ+J5yMBOY5BtUBbXqzxohFrIQWjwZPNTbnUFi
23hz4fbFZyJtRZ7ygpZAXSSzbHRKCH8sx58kIlrPbZERLlNIOOLugmaHlhFoWLDb
KarB1jgdMPvD9CHUMmq0jJt/UerEjFEDDHmnfRVx+aCDbKgEeKTBNzStTODt0kKk
SfYZ+5aEldaX8oI6p1iASbrnH0l0Egd9RmaK1wg4M5SJK41Er8CLCrQX5oXyFIMK
zPINgk4W0y6gg6Ck3wZXrN4RthVDY9otEHkC5QcC5KXB4Y8tpVP7aSCIMJ48d2rR
ZuTkLXDBRGGc96HsKvDtJn+hKkOFU80UR/Ft4qZOHL8aszljzS9ykRgGRtVBMGxq
8RIzOZk4/U9mldZvvPVWOCDVBii8GwmHbRRiFX6rAjPeHWyBKtdJQhBfVJ1GhHAQ
p5+F7pZD187SEm2ZzglVcQ+NEtepjzfTAteBvo/uRfGxuVaVDnqGv2sZJ9v/b7Zz
aI+d8X5Lr4YfJvC36Qw1efaK9hHTz8tvPxAX52zjLFdkYpRMKVOSHE9w5Ha9rcTo
24lnjKWlGc2Ze+ZDBVd7vo5k2JKfJUH1lI++d7nsH5On00PS0cLdAo2QobIUD6k+
RFEIV3Ymo8z4GsGykvlgXIW09ctiox3nvSucuFEYvVUX6uwBm8iEA5MtmqhDnTHC
mVOwb0+O9zNBKvYq68kM4pxdWNG3kiG2dXS4UPYyXiNW4qiHw/1QuFTfieqN8urb
pEgj5bQBryHNZPN0kGzCcZju6ug0w5TG8OexWCuA5o0Tq7TOizTrPPjY7jmxrPGk
kYYCF9BLKSNPzA3iSTK49uF8w7xRf3MwejaRVE0wUpI67pj9nELJxBdNgr5VCw1l
R3J2ygX6hM7jLdrb00VhM8c3IKyzI7B7GkAAWOdraXaB5hOeu2hDPw/ZwrbQEVaJ
zkdReJTBUDucarWhmosiR/b4fv757IVfljEfPvSPCiA0kUNY/MWGOM2YEQUKmFp2
MXNv1xX0kM8BU1h4bWsKB2LYrMlt9L4q6HlNy5wQO/a/Jaiu1pVPCuadnNkHDKqv
UE8J1fBazYGE30kFauV6lYewOQVEVxO0tXwH5VoZecYIKfPyIm3lXnOmMVhE8ez4
Cu/6lwC+JTJqdVICoztk6Lg89cTYjxR8Dltn7C8Y8Six1ZzdXC/MWtOckkSKDBhj
gxSwuL9WfwgMU8JxfziN3WRZO4WcL60ejMu6xOm7aypsFFKtEErpMbsDiTiDuTRR
ZgTge3oiTwAgjTVhtMBItQS+MtxcMDVmXxb0Cs6quDL13qBV4rzmZZyIEzmqp7LE
n7gfQE0X+7q3sDrk+DQgFTitwpomL4KLag3okjE7xWcJZ9J1TTdUmyy/Np2IjQN+
3bNwmkT2GHkSqHidz4MJkGVVFs+LtjdRHaH2lldQUdTem7Op6AjA2KkoFj24r2JV
gR9fsYYWfvXL7gs/StPAsm2NxguUINmK+7/BkSgVs+wlIcVdN1/0QCwqnEJyfk3n
lEc6Ua7ob+/sk4h3bSumQfnp4Cb++68imkvl+oKP9imJasAxRiqVWALp7eof+u6n
DR43mfNuqLvlnA9xaXczpJbesTZDjZVQ3KywcHpfggvsyQtP1DOhkgkRRqxPdn4e
UxBvv5/hPzvL2Ncorm4zIn/YOR6QcXSorgZduhja0vQ5Iribgk+F37MwzDg7GcCn
xmUdWt4XyPSdyMDGwIxBD8YZA6VwabowfwVMLK7mpx0TFTaYj3xzOLatKclN+bqS
FB+9+6B9R7E4+LuH0uf27kyB+qG0gSr/2OgGczSdWBSqI+ZoHxT0x+kun8VPCLdc
xJjyEhZ0qDnOdC1pSpPHHUdVNN7BzSDwtTjNcfNRprIe9I3R8FSbOPq+9EKVkqnO
qpIr4mCGw4cP4Wd1x4j3trsScMcZAuK5KEEasZHIYKzW6EI2KE3gAzFkWrpmIiio
WhK9jskRV9d5BmWstmBtA9DHNUGb+DFoym6CiQYxIhZWReuRIg1Diqo/i/AJFtBE
2WOumJU2sY0UX4Onm79UizKh1htkbh8VQpcepotUTp6C5C8oCOCQ8VDsrQNpb0a8
HRy2nnpyiUuPjnK3vfqEx55VduK/pAzj7tRKjXz2CFyp/MNIDij3hHHszmWSL45U
E2QShM5r5U99XnKXmpK2mbUEGcgke6cAYwkVx4SmVJe5Ig1LAZoBIoszlB8ICWyp
gWggHURmjSfniOWcjUDCV1n6Gm6YEy3hJPHwM+VpmyYzgdcIa4RuVZxU7ut0ZZCN
jBd5Ynb/BLp+f/ww7PO83f/BT9othCTnRnpU+gH9dbuftaVxCC0gWeEb06H85SG7
bz4pVcwGRiSJAX0O7dHmN6heWUtYC7y7go0vAATNAZXfmwsbZdo27H4wgMg7/OLh
QYiAYSXVOUDtcFcm7KGFQ1mcCkpl/4nEBhOlBsWEyIeisWGSkxSKiIMF6goTsO4I
ZSsqi89VLwaYUkYfVVOgKBZuIDG5RvJOJtaa0VGKkvStddYRw4L7Wwb/AmwyAuSH
U5bdAXK+CIwAe+3Mc1ZzgX5oH7rfvuC+TFqyVCBuBGe69hfZ28hSBAqpQxAPECXY
KbCiJq0qVoX/MUs4y7wForShpaZIiYX2P7gyqZeItvo/brfxHqCrzfbTWaGOPlT0
0Hx+b+I5MPUNL1RmHe8QWC0foUdwkMutuxGgpn/KVHT0HJXuj1ZmRDwJtFcWmT9h
KzhynJqbK5ylfrDt/krNecebg++2zCgenJT5zWqi4GkfDQWDrlaeGs1o6JyBPC/m
laD4fOW3m6xg8/PswpzaHRDX08vwrel7wNn4e35jyCuoi32tYvwboac43pcixw6I
Bak9mqg92oWLaBWgy2bdudICxbyR6fSZfHpI32RrXrLmP7dSPYH5rpVLWOfWiUs1
hPvpuFHJgrVzFsJO+50TgL2HYjNBxM20rshytKVCXr6EOA84lOQ4ii69xLD7CoC5
L9PZsY+Nvg6XoVGbvmk04Y2iCUOPrzjzxCIIPIn/nwj7uucW4aVlHL8tRzjuAb8E
E4OHVyCqLs0joEjlR6p06n0+HlRtsSsZ9ktM8Ng/37cNjlW+jmlt534NoNlcZlkr
E+zN42tBvXesUILZCTx5+jtjEWH/EqKBAnd3bku5EnInObfw5MsO4BO5FUNx2C9g
omCU4SmD9wsQOhIAN+YmgLvlgO5Tc7dailDCOZTrUQZT0jglGbZzE9UqrKxNlq7m
vKOqNuo9ns7cisE1bG/oMq756vwtKWd5VjVwoMv1vNL1dTXU1s2yGNnK372NW483
FOjm4m2LZK9cBgRbVDhgFMwr/3XljdYH/jFmpGX8A3iFh0mAI5wMrahb8g/dRBJx
JGMLaDjxMZnRmZ8dw9/BpUJqW8WpbDW23a2wDahaaNNcXLuj5X4DVggnobd3lKyY
DiIA02J7QJckUMeFLNulLslA7UlZXa4ZTL+ZQLJ/7UlxtNjdbIHgNJRfN80VeLB2
O5B0/hMS3uNiS0IMCHHDho/vroBeay263h8AumwdGDqxuqLvgt3aRDcO1NVeR/5h
aZe0IOEPPM2zbu4eI2pg9zTWdLMLUlYpe/CuE9pbW7I/rjABwKAvcsS3uSAaQat0
ssGPFR6uy8DE0JFG4AGCs8v684CnPmcWjf4gE6jEzoJ48A5jivnylQ2rkCtjE9Iq
AyeqFDL4mkRBywXPPjqM4PF/Y3mSwUi+WgnMXV1/gbeid/fKwR5zkKZjtuJqhqp4
Gt+yOG0pLUDhHZTAdXbo5Q6AoMOIma5faRdF2O4VckDeAzBx6CQCY/p6rRwj3L3a
WmSYs9Acs8nLKuXVxuTUvH1saWxLvSRa+ZNQJJTxiBRfU+WZJYXCY6UFqfigwy26
Yi0b1TfV7hpnNxUGGe1XBDkRiOeG9BVMvaOJs1B5aYhpyx2K/jirdQdCcsyXaQ0u
hIO5B4ktux/p8bJx8PfzKHU+kjaOhmNaB/Q2q00V2RvwXkYPl2XJat4IQEouTrzr
/Rr0+0WXF47vTIJJi8nihDc5jb7Fygu/h6DYTynm5H7py8mLZFdCPIcvUT21gPiG
e6VemBxM3j7F6t8hdU7dq98ORljw/I3TMmrxZtBP8lVR1oCgt8yZumKBzPBRSpDo
qpARbWSwSj1Asdii3cTQCbE6gAaZoMlppXYiZlcPdf/sIgkMJ05QoAQHO9e4w4kl
D89SBkL+43uxKX/rSgn/YMYXBY3UmWZEPaAWw174Yt9RICMMo89mWxqoXeTAPj+F
oUr37KO6UZMwiAV8kf/ftLrkkBpldQ7AIaSGvvIC0bHssMjUsBw/aRBy9KeID3NI
Qo8/+r2Pc4QrplsTgm4fJhZEB1g3hg7c4qDcQrDh3X9H9SIVnoMTzz1JAOTvLAf0
YmdHk7g9zohzaHrxUzW6PZLdAkNC3x3rrWB/SZEOlKSdJ6MJLjPjA0Mpe4eFjP0D
hrx2MOmqkQFvcJdxSy5oc8vqw1NM54JP1PS1sghJZT+o35HZIi5HaLZ3K+jiPfYZ
xAsdeSq9Tq/VRNdnIMZPiRRTxfVi51M0Vp6Md9B4RUIGwI2XjEpCY52tzsFUL/t1
dBmDQ1C+/QvYxcaQt7PAmRVNiCc2kG5FcMKtI3X/ojg9f08sudUAG6tgqHHwZq6o
/WnByn3QVSZaKdXXV8omdJA9n+6fGZSr5yEWmo6d8wPo2npdymcwpEwWRZkjr3WA
Lzc1uIDmKhgvL4UKdCumFFFj4af1EvAZ6wxGhXTksuv5KwsnSra7tlB0oFNMorRz
gLK7QbcyUGYgRffYFq3RECDJveKRBeEKNHsTttFcffnEyZnOX3M9MCBowBACNJGP
2w9x5EZqz6017gli2z1BIbsObAnPZ6xDYPAaqq5fNXPEya5VLxLFlBQyUPGl/P9q
mN1D+G3HllZzbjw9KVfHYP7BNLUc//CcanNfJ/tltmeXbKt/+7loKvsM990HWZmw
U/rk35cNImsqu68EUzUD5d9tBzC9cjjI1UqppxylB48+wlmM9wD8JAyHWTmy0FHc
oNIzMkpIGkyRIKTJ/HG7bIffwOAtkUCB9NO1CkDR6Q0hDv3trAqUEo5uMnm2XYqH
T36cTDYYAo1O9HHb65yHPZCntk5P/mCC5iAsW4tSTEmeGGuovZJRuRnCDBFFfVtU
kmJfK8LWwjfHANpOFcEcn6h7OuEYHrFQIgm+ub21mG0UE2/ACM6XTChZNY14Eyji
BD/krZt1LfOjZu0k29Fh0RmSRPev478lNizzT9CVIQH6k857C57xTjUxcUGNimlF
t0b9yd0h0YW3o1mtBbRbv8InXZvG4shiEIUdX9rBlLek2PSsjsXM2kwNyv73k5j0
qoOOICe34T5KO6TcoyZQKAM8TJUSCoAvgJV09msvTEeKxqyPy66lccrRrKPFgL8p
6aIFBGJJIxyWARjareA5VIvefiA+ex5uahLoEmkWqbbNjR/lQaXIKdRKQY1Y8Q1u
Z954PfXMZwUengTjzclAIduwb2nIUbxNfn5sXRmvPELkJBfCwcUfYmei3weCXTgH
SO7OjdLj3LVn4urUkk0kXitwIl82fyy9Cufn5nnfOiBK1SnfTw1/uhe6a7NW7nWT
TUNQUMdN7IRjyjIgGpRdQDCh1lknNnrjg9H9OYtWv4Txi6idmqzIDyqPEhpHgJiv
9kEAs83nt8i/WdxHn1geAQji8fMz1PmIEKuucC4F/ijF0yqHV+R3PqeUt2bOAus1
6feQWsgSYcO3MEX0MD/aleU3j+Nah/LLEezXYNk/OP5NIdmm7u6cn/9yP7ohQS17
glgwvPx9ailP3z0kGQd2hA+JZvgPzbuwTBmdiDrU3ew33m1w1F6NrxFgaqJZqG3H
AX2cm3X/hG9vARk7UmbHPvEd5ITs9lv6FQ1vaNpe6rG+qqS4+P+5+NXma95akpSI
JB2oKksoQz0NttXZKaHIOZY8VRfuQAuwI0CPWMx8K9wrFJTzJ588NMDBdZADiyGC
SbklMOdUGDsGA6WBiiRmRHVuqazDE+Wpz9Cvs/gG/m+W7AF4JiyXQpG21LbiyS3C
ZEaKWxMiGezVyJWd5dhuQEtx4rJselF/NpMOxVEuV2G3zz8LmRbl5RTyH7WkWjKV
d30QsMN7znOUVgLtEYSykRGw8RceZBwQgaDe2vXrFdUunuDs4yUjbEaX+Drwodmi
UP4qCcOvRsPhFpV10QFHypwZIWg5/w58/fYjqxKC7MyulJJn5uPmY7LCyo6LL4ZK
BFO7jojSMpHp72sHrCd4lcgqUBTr0boLQ53qJ51UpUvXg1qJvYBUd6owIvEJbyrt
DAoaQGk0OlBIeUXdY/tAZRN8ULEOFLnyDXCT08S1VY1P8SIx4HyQykMULHLSlCXX
kr+lBl/YG1o51tDn0aWpDDpeJBHCLY4VMqQsPF8xe7q2DM9LiQtgw6Q6Evdy/l5v
8XLppfYSZrOh8OD5YJyIVjNKXrcr6xYF5wmDMzD2zgukc3dxkJiuKH0zXUss9m0r
ayjhgC3Sdaiw0NTqx2CWFJRNim7H9f8MwPE6CCu4PG6BWxA/J4uHVMR9lwwJmkH0
wMAtETBQsxunT0ZhrqfeDvrB6bVX0PB0ihZ+A7esY44PfkiBAqQxn3Ix95bwcEc8
/oemsVuOPT/v8eBsYrt/ohAMORlWLrzPvgPBglNEGet/0gg+O1l8fHF2viu/xFte
omeQVmmvPpMq9sM/mLrhjfRSwzX3VeENZDvImQX3qrJIJZlJADXJtRhhsYc+0O9a
XUx0QFuqe8vQqu5rEIN5Eg3cTsoFf2s6wWUzZToX+XFXSHAy6dBbh0ysUqkd/14n
1DXlCHG27GP4Aqqa1QDzibnOvNsglr1qiahnjTkusImYSdq5sNh/qW1ed0Z7/6RX
mg8ms88TJ/ENJHNz/Q97AyxvrSQ+9Mv0S/GGR8csCOwqGS7805RGM5pVTerIHJ7q
APVDR84uEQ4s+ZFbosYMHItVrKD3jBNhbfyDpOiXeW1HCDhKdcHrm/z5mA9HoLVC
fqu73K22FjxY6dnEfaGFEXS9F1mrFHic2C/9nPy0NXmrxqNSNeIVx3YeuQCHSwSM
aNXE3vNHUZpAA90OqFusXD2kE3MWsYAoy6g047Tf6wGS9AnIUph6idolvXKVnkGk
aaIDTOlnrk98+RxQtNPpDWxpKs1CXU6JoEQR7MJUjX4+5kUwkTrUDIv9IHDJ5mMU
nfixA108ykhQxoCw5HtvO+/m8LcXZKfJVkBpUuT+Hp+CUAF6JSzB+ptGu7eUtHNM
zbFo16+Md1KlK5vxIdX6ByF/sx+3NTHURBgQuCDKAChn5SYogXsriznsGpUH7hJm
m5IMqQOvsGzibmW7N+jRv/Vnx5DQVfoQVVPwVpFACoGuDVcTbaSdXT69CM1adJ2s
SHztOpfiQ3qs2JMp9iBo49h1Q49NDltCj3JEg6QenHddey2W3evmFBZUr6UtJQqQ
+XbNP9ZMKB+eY4q02SjVkG67J3C+714iGhjs0fyIQL8S3jMOQ7/RMLAQAHKfHeGM
EOGV0akiCla+108W40wSmrSTF8yT+OpnDPQ4Fy043mRC/wlCW11MhBwqM9mgFl2+
r24fVl915scfep0AnHz2Gz1ssq1+AeXmJclYV2LdyQAnJ8IOLhsjF1218g04vp39
1y0BK36U3tXoGTL5NpFopyPvmkSY3s9NktqP4Uu79KmqajoJ9tfVFtXGtXyQLCqu
awz9hkfj5fba4120g1ZkfV3vOHl9zzgwpQaYXo2gsfQwk3k/YBh4vULffzSoqSLA
FSKUTY450iGhp1dEa1vCIfPpnmhoyxgXQnmLsT0Mj2HqIlafn0JYgS+aw50JgbwT
IySnZLy/XluFJ7AqXCmu6WhEqYznuBa87a0/WFyF2rSOQlVL9LI4aAIwfaXIdp3t
bnt/AYYoiNW89MySW+WXjRXj2fCMhGVXmALd+MgWkm1B7XQcFMWe6R+1jdXaIOQu
dFlfwon6wp9wX3gisjZB5kQyqONn2CcLjXULEuXUbcxHL3aa5tSi5TunLFnrDio+
leKGk3qwAEJxQoAZO2/DXSQgGQO6nFgvFNCkPM91OUZucqNHiVqTL5kM1JDtjWUx
2a14DIKuNEY7wFoPDMKQcppxp/EQePlM18gYr7Vu2GVeXCs8+PrQFLsWVyAli5S7
voSM6VZFlW1f/mOw9RC5GvsGVt51c+hf2tSHD/VXG3ivwDsi0AFwohos81OfWfKI
koiEPppNJx4hMXlSLtjxQmOyzGOBuC9bOMsEJd7Da4U5QLm7AnatAIMcBDWC9yLZ
zirRuaLF/QC85XNd4GsG/ivVUF5D3dD+/6aQZ8LW1ehMivVCxn7cFYo0RvoEnvrR
NCwP2mULhZcymNQFZvBpcf+Zf9Crr3jKiOLdPv9DFlpUPIZPCLafFBITq5rkQ1wP
le4vOzLWjvZPCt48iaL4LnX5wsNRk0c7uAPn9vjl5X3LecwFHHPBJBFMfkUb1wiY
aVnfYFuqtZNMxtCngaZIG4ypJ5mg3dBfv9exhd+YXHOGLtSBy7dM5h9a0fUdJN01
MREcEBnCbEmWs0Tht4govQRyD+krWzOd68+S+Me6B+KYmrlYCcKZ7LocIevxK0U7
Qk9+WOdsfOiYJDU0NLWL82VAjKR9Pp65Vn/pOy76+EFn44/x0juB0XHs6681cJoH
2unMDKtiiTDq320vh2pkAPkyV7YKNGuUTJC/kHXiL8ZB57dg47OdNzS8VuepYU66
ufD9ix8wr9obIOywett3W0rgSx7toh0SmbyKWp0tUl7A7oDFTL64YbHiCxoYcVu/
RaeAgYgJg0qPscSuB5ElJrGjKc4guDSCHLIatFhy3x1qWvAQ4w/DapOKja4/jnw5
ZcS454rUbOPi1ZuofOb0mTbqYeHspgQhSkOvphi9sSEwdfTZeU7Ioritw6pm0bd6
ZbfJ6Z3jPae4A851AiY+bOAXyZj62xnF95kqnx5gKJHxHp+JpR5ppzAN+AxaVP5F
Kh7VCTJda2a+tSOJ9+/np/UptkxatT9iLFH2FFtcWI6lxogpd8BxTu/Lzjt2n+Pw
brmle9lz9ngvitMvZcDQzUItplY1UFBstaTFcwC5fYohRrPX7TZJ9bJaRi0VTPxk
bglB5D9hQWm7t9pScqk/aIm2R5bZtN4WKLluEnLMdHrpISAX3WzllW/vYYrZlxbM
lycor+dKO0grtaDX16zSNrZk15IrTKSTjRL9rPDTTN5DfOywUJGQ/33tE/l4BOp/
qrfl0qcN3evkSbClxFx30NqFUYL1sGTUaA0kB7B7mrD88yJhZkYVOXAA9r2Wwl/B
eD5HNgo3WZTxhr2Bt9Y6lT/cD4pigjdT4r1xe8CwkTUgfzQfRFU7GMBGCOB5fWNf
9rDbdQWU/JeiDLQ+LiVESsc/RZjSXLIH27OKj4d2X7YFpiZUSeXGmmCIH9c+Q6Ud
Lk/IgZFo4kiWScMbTgc7cmSzPXVESM3wuuL3N01z32ZbbG0uWUnBSPYbB5kEOtyv
8riUeXhb+0PMtV9m8sD12yBlSfZH3Qf4wOLoRxNdCkiul1k65DYmXkK8AL1nVKxJ
X+rniWtDv79vj47cTYV5f86sj+aHpmH7RLfJpNJG7kdEep6NRAIOagh4jOUXcJXf
0F7H8Zd6OFdWkGR+fiKDIAdc8KSaWAixv/ksb0skeWyoO+YSgr6naaCnke4biZwN
5p0od4pE4qEPeqK85HB/oPjPnO2xbTxvg5zY2emLpgHYUb2uNrfcj3yxSgjujsJQ
hrYXgy5Vrpk0JvUhG2rrMio1IyYn0Li2PDXDUnHo6iwpBdpUmAeksGl6wyesP+fX
aSXUiZKFy715sjmmzU+x0BD+6KcfZvn1EhklsJi8ralevI2hsRoMfhNlYcxql224
M8FIeqRYRwr0Op4vLOGM4knQetqgdjcsPAlUJMKtsVagKy9mxagp5g7DXMesPrpT
2e8SEklPFJXvZxIJ3+g5O1WlKKxVEEt9DCqwy+og9wbQN6Oh1Vcgw/eGJ+Frz4xt
byJLCmg3rQ2xRn2kFdDuJAbyaH1ZbwPJQXeHm1M1BPdk/iNVsirpqWHVsOATA/om
jJQBVmR93VAf6+Qa6g5RouamDwwvegfN9AV8PUtVQS27Pgu05UOiQvZleCP0VtT/
ImFNl5l3n1NdI+JXV/zbRz5S2zvvMf2shd+tjcID2lnStPbJaS5D898XJDUN+zFF
bhmcHBaHTJDsQ8W7eVW+3mZz93/c3nn6lLcyIjiOzfAOJwkxdfH7FqWlWeprxQIP
izVi6h21Ieuw4gIA1211lIHB9FdrVxg6QUkl2uFkZWKNrgDjp+OyequZ9ZQ9kWfA
fzzRhfrGmluX1Pah5ToWug/NROTytHD/t+wUDLSpZUPGIfucnZVe8zjcD2chj6Ub
FUMsgyAL2APU8flc/0q3admOrNeXRLHLGyqbOoS9SIE91wa0/55dza4MU3DMNgno
pMASJ0Qhhzxb3I3SSQEofu69Ph86DzaEiasicxhnTb6A9PNcT9YN++KGwRimrtDz
YjpRN9cCPqLEHcHZ1nBOoNG20sjI+39tFGEIBc0SCMuU3QdFu9/W23ilcKHOCN6T
ezq85lz+MTjwUdhznAu6f1ijL0iQfsbvgm28C4QTHs57nalWUstMYmdGXgt9q8vA
ikozp7HWloOhcq7nvd1cGjeBIJSi5K3s0rTJu9OEjkx82oJSaudv80R2hVpHBlEA
1j39UP5PNT4JwJj8+ONDthNzSSsKZzPOljyUqt025KTD330zzVvkH7dIIOa3Gfnb
ySBV3x3NGGB9+8T45SqFqLz+uRrD+TCJHaJvN87NE9Iox+VwVTeOgCzg+ADzJU4q
pSiAAQIKCnEQ0I4wObXvwtZfz8RMSHkzYabBwUvoo+w8dNLn2OCZbaN0o8t7WtEM
qBEjhoVz13mwS7DAc6qVqPCW+vt3jAwh5q7aF+RnoWEmAxBn415nD8inyM9f5Cx1
2s8fSESVaxciyn74zIXqnp+SpG0J7zQzUJlf7Rn/FS6Fbr6J+bi8BV7iEXBKKUtr
4GrVoUKMUJItdrDd9fQy0N9C/tJdSUqc7a6tcMArJU2JIQ4jxEKdgCeBlGw+xZF8
nkgqNAqfr2edkAaWeITG5Nu6Hr6VuNeXnGagL+bZk1QVE6of2UW/CJdk/WgEYq//
HhnWi64C/TYVcODY6oJ+mqEyu2IRkeAEz4K9tFZjPjITTyxVnGAWS3RKCUkAQJqV
Ovi62iKBwVibF/1DcLQzGVqbDDhMl2z526BPh4tBzT4vlbcHGCaXIa4DtAeJw4lM
dHyTrhh/ADS/Ld2CHXRErmNMz0p8w4uZ8QUR4mqhrJmAy0Q0pA6PZUrn1DFCmGft
89EADKJn5YAYyEKuonqMyyl84qw3YQ8hqeGCruT3wVDv2eUdWyRRr6mh56JLICqK
F/UPwjaef4xBlKI9qySBAdbAsIYsvA2sroIuWJKAIJUdisDL9j4BQCYhj44qcLGS
Bsdc/L7ElYed1MuTKrmXxys0FJ9c7fe6z5Tv1FomifRvIt38ozAWYsZRezICYldC
+6Ed71AV+N8643XbFGoWZknQwF1+d21quZLsygFcjvaGGl0KC3KnzETv2h1yL/GV
rQcM5TC/+MXdR3ESgTK/JzoUxOy1QwnqTbXongSOsQq4odqmpfb3jTeUvv3+WPcE
r2OrpZ5W1fLXWB9fMLgtk3USemiGV3DqGp36BFPKiLrLbGb02gjLQo2wYIVZNhJJ
u+xalQrxx5sODerPZqTcE3cjLxuaJNzJlCNShmefMMS7ZfWEf0wuqW2u1qQXSKnD
UIcrLkyrbxAJbwmeHmXAqdPXm8EDQlybHP9kV1TGswfNuzbDHMknYJL6JVBOfQJo
QZFpaxnnhQiX/Cs1CQMKjApCeCPG45TpLTAd4ldM9pl56dE1hMysKq3dD3398MO9
eUG0M+5OdeD9/o/kmb3kGHXLxr7DYsc7TzN0YUB6twyl2TH8v3+hg91q95uUavhB
dKL1Cye7vpK30wIHdQyffpmzjZsG6Bvf8PlEa3p3NYrkVNFhXit2s2lNnGgVBU8x
DQ4cyokGtuuZyAX/EzI8WjbsZlhhShAhWuPv/sdMvtqXn/QslJld+qP2D3AzRoF3
RLt+Pl5j38XuwD+0C88AT0LdfRDAvS3AqWUQorkG33jqI0Seat/eg5TwWR4R+r87
6YQZiMqT6XMk72yMrF1Qsw+eZxRsPxMqwBdDTsT7SEsUiFthmUsBiCxZD47vbFVG
4I9eDavF8i580EkB7SA++JTnEVUhgMxlAv+UdhPgdQgPm6APXojV8XmoBdRaJ1y/
5sWb9hMqCc9j3pqZ8FzrHGj1R4Yx8EoPOzRb/mLB8EB1Uskhs8N1qA9GYF9vk6dt
outGWPI5gjq5+fdmKca/ztUqzcWQAMcQp+bqk9fP7Gt8qb20tO7caEguCddbVUgf
Ul7SHX6YSTO2h3Dp0jmHwuAU9s+wal40fRdse+XpeEZ7lEULdnmPQze+2LlKYe2D
Y47C4jVOlbhi/tfA9Sk8Hzbay5tIPzAV81BC5/hYm07okOgpVu+c7EMio5ZFdue3
O50+hIOpG1ZEx3bSc5rRzZx3xBGPxLe8TFdDqP79KlQ9umR7/rSLQezSmRwVRqTv
EOC/0r9p0//JdqvaqLNwcMmQ/1c/Q53Cxv73QP021oQMplTvMqzRcRiIwfnmEWkR
Ch8ZkydUqY1of+UIg8tUkMjoSgsbNmQne3lvuTY4gpp74cF+A1tdixNK34k8w8u1
ZpKmnmon1QVPcTdftDNr48TBEW/Wt9Az1ADnMj4nGQkOCBhdvwzPp0n0z0rEoGSu
2HqWY/adiXpH6vaBJEqiCzEyNAcRP4MDrFNZQ0F4utEzFhO3FR/djIJAb/jU8cbP
JnPEH77N2dlWiqdMq3Uqh2HZV21y9s5z5XpH4hBXhCP+wlF4n4OCPOF2VU/haNca
QWGc3dt1KQKLqicwQ1+m+goP0xf4NoICjlgbTx+gotTCteBlujS8Q3LiniN9U8bu
QJhbz7ujBu1wyQO2RGjtgN0qo4hBFY5EyXfqBSx5SgfXfkN6JdbAOSPif0DGQ4xz
uDyKgo3H9m3mx2VKk6WI34/2xzNGuf7VOd87M6d71QJtxSY9eZoAQ5bU13fbrgG0
WZkuTsPwck2hY/5JeTAZZ9njYjZ1JFCpjnu9MbzZ19Y5isP5XJhqGtxDkdGAYHjf
+/d3D0pa6cf2QNxkwTpDUvrl6U2jd0MdIN88pJU6FPdSbU99SWx9dZgqQbNAkOzE
9TMEF8BxdA68r7GPIkofUyTHZNMUHUx/LVMX+zs5UKeUS7VZGMkcMztIhcPj3X6t
ODkZVCHZBM71V61HwZyxwTkd4rNGoA8sRu56/wZ4LCMmY8JQxK+AfZz5gupKV3Jn
UF3ZHKgAOetgJXBG1t0led9DCWkoc2MBaBl0KGC16/jUMAEOkBLLnglgfFYDdU7K
583jhKZO2nguNK9tcEppswwwpRmd7OunMm4J5XlmqARD//g+/37zYKGGZzS/M4ds
iBN5H+NQgcOHM92mYYw0PWThBQ4/w2lK7JMxIcYOnVZAXUS/JGwq9LL47X34j+5G
zCukjSrgAmmyM/yq7LU8GBXTPlJZXGwm+52qRqJhziFMS68iFh6izzXSFoGE5fUM
ofvJ72Pq/MPW8rh9w1NjLp8LZ2UkL05X0Ke7g3D7DtGOhrZQ8OOqRWuTi8OpniEr
3YiXBwYSPGQ09GdpeO6ZgSuloqncICUTDAMxC/ha9/X6otpPvpQzjzZffRiyFGR7
svSwXu08/7EUyga9gcYtGkblNv3E8kgSgQIMYLLQ/BFZUsFKBRBRz64r+rm6BNQZ
0s/6h4i7OXZRRXNSCibG3ERTcoIaK62BCPj4BYTAhM2Xqhw5qmLMoT2xzVgkNJ1E
fdlCAdbTFtrrz76o44rbZreHish7ncKkjAGsbf8bNAZgM3GFP1X1JWOcyQw0X3+k
9sc/yA968GWvovxmoKNYhu3dQKZ5jlV/Lw1BHpFF+mIQQCUvWtE8rEy6t4Qk+lvd
6J9roq7opJEVe6e9SUiTTKv0ZZc4B6cQlqbGQWMLuAfjNqryELFgO+2hv2MvaoRZ
wnmCnq3pUlKQm9B1aHmq0fWqkO0u2FjG+EhJbPPoVSpyx1BzSRQhfh8iTaTJvF6v
Xs/qfUW+y/JIQFZs7OOULM/xWljoBeC3UMQgDbfnJvFnoWcwq/4xRe2S/LcYdsa4
x3PPH3qaSh891lFO/Py/hCE8m2CemnQ0VfKm8YNpsf9tDrdA4XDRj6wTOBZcGp4P
/R/g/QA77V3smCdOKQGZJxVbe7zOCtsIEZXdvSoxOYBtOdaS8PbceEtbK51UTtfk
iFAv/DmNykhhU4HeQYsE2Ct8tzn7QGXnFdqkQgL+h8ExJtFWo/vtQgsOuue+jIqX
NZcRIomC/Tz7FFVKGI8xeT/bdiqrI7Uxrjpcr/B5BypK9fI4CCXlqK8Oh0W5RatC
F9VVi5EfbaACPPi5KrHimUiwD5ApLL4H4XMse3FhjToyHzvMXw1X5jbKTZ7Cq0RG
o2s4+di8v5m/AQiRWuSPYzFg5gA95SQQUS1kVDaDefnvJVRVz0gwn76qFwNmBbJB
mgR1kHpTD3I3dHG70s8cuYcpi34co6P3JR8qkN1Zqz6DkhIW++1hGFUZiIbUgHtK
cRkovOMrTGVzm0GtTkBwVdBbppbp9wuj+88NG4AMEnvTDfT7KZuECD2fz7Dq81oO
KdAiPC7GqxS+R8IQ7GVmdCkPoVHHPvNHBCFiIvby6MkSGB6PNDEDEGnp+2lPVxsL
Tu52w4gprmadsm4tae5OBOeFienk9D53aHiVTAc34Bu9yO+E7fn9gqUWXWv2ADji
1oJu5LG/eVYpdGGoktIsJFFy1ZDEQlwkJieldQG5uNl+GSzZG7b/gQsB5g3WqVEF
EgmLHPu/FTY/zAXwSr3k+Zh2HKN+Z0l9VzRd9ABk6r+WaNARERGPmVetZy7EESGI
SJAyQek7j5FuS9ne28ZA0o7ZOFADNU30CjImX7xzDJIj9gR+fjZE9d2yPx0KmuFk
Y5nU10Awxnj4o3vwoq4Mlmt904SIm4YypW7MGP2BSNcLn2XtwkPnmngWLtwcNmpl
ZrUdSUfQCwyxRNwqJpIWHW8mOzBP8bQU4UkDodqNGAa9mDy+R5Uq7XF1Wr4sKNtP
Lojr/R/TM3S3nu6+TIyGYMNBlUPH+UPqzllGJa0ZgCPjZq4kckxDjZ3xd65eb5PL
NLC7nI7JOs9lKPascFffc5wNU3KszhSO+U4WOHCFe0+cMHenjIjEenvNok9yRb3k
8xQj6v5C8AQ5DNAJb8VUxUYEC/nhK3WP++Y6kensqe3DjNfYmxVsf02xZJhwE2FQ
gzWSzB+VHZvkfUzsdt8Wy+w8dBLGuvF9C6o1EYkuzEripE82q4TdOVFcHwUapwzp
Uo/44D3zAeE48PGyIsIVBESjtPQWTdP+1gDcoxo4ihZcwkFQ4mS5MmjnpX+8qvvI
QuFgdX80pNXgXUHa8imJ4ZncCZi0zKSKyDAnHugF3s+TOaEpSv2cKGxdzEY18skH
d+XWWlGmnxI0DUG+YlUAWENbwrgXMCKfxDOb0zTNae3KH2ENRbZuvTl6fAoLp8pk
CS1/NQdsOS+n1peQaQGonvqSBnFroJ383kjXwVVZ4tWTat+p9z4Hpdq3RIDinvug
/r6/XsJ1mOMfmpZZyeVfbHAOUEwFf1NDpxOpV0IeR7Xob1jl2pQvucn9Xs63U5Mw
dwkJnkMa1uygbt57TfqKinAIva1hpKWR0SQ3Y73c/6XfrEkGUZcH38Ktu6g347uk
BYWfrefbkM/IjeTDfB/LbvGAVeR0Gl+l21tgqEPU0yXnJIdTj99QGKUtHEHzJV6X
dGjdzOSIa8x9VKyhbif8nNsCeneOj7MxM+9lgk2MVdXn2DhNQMNdmis/iycvf5Ob
pnWGAiOmIqkLEcM63BQmLk3/2mvcNKPhw6ewcyFoW164dok7jxzAzY15OAkW1czB
0/Bl9hlNHkA739Q+sONr3i8ubFm4X+q2pIcn++NFn+EgQghiwkwB0o/EC3IlZJE5
FW0a4aMA5umRNxNqA9x+kLu88tmWn7oMx3yzvPTbBhbmVGPD7LUCkWA4TdMWr2mD
NnBHQKhNLqqBYCssFWPmpPZRf0L0X4fXqaeKJp/lqCMvSq+08GNW/xzcnpOcu0Zt
/NzF/84tcgTW0p2OQ3gQUZScfYOfph4ywFVbQKcu5KP2FDyX8i2mEt/HEB1XG0Vz
e6/5ekqwlmRcKsG55XV44YySTECWQ1IjcQvtCqHwDHaaWRaP12kh17LHXesPL6J3
6nu/qAnF8wojyKSW9c1oTnfInDJlAvesVsOiSMOWvmdB7H2+7W5hKVAhcXXOPxOU
MnnNcBuzX+LFs0RgtzOuFDsPD6HlN2bLYScJTndBef1FwG/ggWm/+GvpAnaM6bR7
vtUPf28wVrgWY/VWpTphKmz06tam5j9mKuhj/4m45vDzxASUiWOOBLisaofB136Y
TURtAXz+6YCxSAqbmJEDJ4r82QsN0m8F+VV9n2Ar4yK9BqBH3HyjY6g7lUMBmzEw
41Hb2Y7i41miK8zb9znDVKv9JbnjUprgM3G+OU0RpH6hI8X4dS13C5Z1iZThb25R
yeWUpll9c2H9U5uJjRoVPDN3hH8juJw2zDeTH7+Jx8Khd0e4Fc0wvvhQy5h1G9Ky
7qxAYn+YA5xzAGiTKh28st57iRWOlaQuXHCzD4YEH89q91U2Kdy/RXQIceuYsDT2
mmJ298+fK+vBsT3sokjKXtHQuNVdlgLowpkho+TKxb7I2SpjTaWe86MgpPP180h8
KYbZppODA0W2YO58VutEmsMrlyHsxfd6hIgNo7LF/Xwddpa1A6dDHB0I0hpf0nvV
JP5t4+YsnDVzlD9DaRQJBCH7K3fwgehWulSOLyb3tCxdcVY+cAcD0Eyoks/dkrn6
qQDy2guGbqsrsuE/XdTTM6WSbcReW+PLttIvr+/egmIGIy+xNzhz73Gtng9V3XuI
g/hrH38zWjG+UNoKUVBXupLRO63RKXMpgUq4L6nexZVVv2XeINVq6s+owNPocAnF
Cn2bvoQdkydIEnQ8vTI+gbjfSZEmG0RUQnYIgaUd1i6M8nKcLqd4DLHtqpEwpiHj
Ekr0qFzshv83olvVoF4c4W9hLwyVzG/kALDOz2fXsae+MDI6b3ylrwh5WpW4GH4k
RiWZ+h+sx/WagMjOHaFKhV2b2zOJk54nS1bKmMGy4BoFlxRkY57fltIGDqMs7Tvq
9SylHFyrg85l3oEVrP5LvXVd+AP09HVk3SyZiQ42RPSs8EHeC3UWiN8ZFcNBcA1B
s9cCRLVbSG+hY3fvoMwuB3MzyLRYpcgLbOCsEUZw1viA9PTViDbn/nccBN3WfhFm
PrVP9DYWt7Kw5ZwQcZzobn6uBDP7AS2m+drep7TfccgtvFQUOua/+88VCR31ncc0
Gx3cl4YsaMUX3gPyfpnjyAG2rv4amsEMfN7wDp+rvH4V7Y9gR4is19KoKuicOOqU
poN/wojl8fKOCn9NhRgBHd3t6uC1xfMCIyVntDbbQaRQ9oemNUpYZE4mRy1qWpOS
OZdJF0zAsKZMvMwXQs7Csxf7T+0tbg+C5n5yI6zZ9sCEMu2d1nQvneflXx1mw0RF
gnDTyaq9Ho2aDRKW/jxKXy1BVERyOsSEun9N2o42hB6Ub5FoJ562a60XkHaMD4sg
6Hde1XJFXaJAegoR9JCYyr/jhxb6I78J/ocemwHsyaVqLlqLa4eCx9z+gS0Kmccq
A/3VS/h0uHe2diDsEGiYVGIlpRNTRy2uGgErH9ihlAiD1HVwJduc8Rl2UfSh1zu4
Ia6H4a3NdAoCHaLh0qqyRMl/sY9pvyCBpktRBri2M/VyQHzw2R38a1qk4RF47B4I
tjmliVCZgwz695C0N/QfiZGZv0rKaSk7n/zWAEiGLaAL2Fo3isDOhWtcZB96fPx3
+ENOGcY7IaK5+6OPP/ky/jm2j0Pj2o4zz4Db3+/+imGpzJhZ9A4dJIj8OEEvJFz/
PODd564KRd9mbLdotqzUMZvbkWXQwx4pqITGSpfan3k+3vaZCvrphRGlAgmUbjwF
/JXz9/72Fc85fyXnAtPnGT/J2Wzxd6b1a7FbsrOmCnuBlwL829vX/7W5vC6EYHBZ
boyb75xK2Ms/piuBHV6AAyh2t3Sob1uoEQQU76XkPFowuq9lBZRkahXuBWpHX6To
VlUaHEsMUyrfAvGV10SxblDreg3+eWyzrHptQi5tIEAIn/lXh5ZB7Qm3A84/PnlG
OdcWQly59OOJMj+VUK666zCB2JzE7CWZa0HhcVqI/99Y5E+IVxIhxIuMsb6zEmx8
MSeoYMpEE7RRrw3D4JjWYR/SQW5CXjJfW1+pH/rQir+c+8pQqHOV2OHVJxqEHBi7
lEHkLOwf1QNMZRsiMeVFuT+ANAr3oGP9CsQfcPLZ2C8okBn09J68LgPpRVGslKvt
PzKIgHAR+m1HV0YLWUm/RY740M3BhG9CPNVzAuIqp3NcOYPmNZAJssERQouqwHdC
/8zqgys7TWiVxcP7z8/ilK7QFDrjGu0BIn3X/iiPw/nGtJzM7QItzqc72ruyAMa6
RHGxCQ/1JRJHJUOOTAmn0ezKhbFTWRnOvSr2YOD30X4ImdAup9mOsj61lZ4JQwX1
2c0FKUmkK9g4jygQh76CWs94MWHiglSzu8Z29rDKYMEsL3KYdvMMOxriLkWm10Bz
0ktlJ6kVFk9WhFosLau9H5jjBhBrgNsYBnv9+Jukk5ilpzAqZ/moOsJq/RuLAd22
vaUSbWsNCEZzLyqhspnTFsO0qiV74xRdcLqvDfB1+49DiSdsTwIiMyZE30Eq1ppA
rYEq/WMmrjqLZEvIK2RE27RoRZc36/bHEf59f1HHaouKXXwUGMYqYGrRfOJrgaGo
2E8Trbb6r+cxT/Ys7VBHYfEPoKntcFF/dHlcmwBdG7Bi8VuG0BveyPZRNTs860zR
OBT3bRhfUVhYKNGc3IvP5/3yYCIdMwROVWiU3TalIQB7jDnWl3ObuO4GcqXmEeKm
8wiOYR45WFehvcEYD64vCp6GL+R7bOgBctAuay7BYdCsv9rNNy8WcxPdDhv5BlGc
mmlL44Amzubq6pXuRghSmPtz5oj2aF7Kw6Mj2Uu6NnP6wjLQ05D0M7Wjqhkg0+j7
G9rglHMeiIqrNaqZuXWJePTptDIpF7zT6nipS7OmItKKMCLli6JnqSCh5BypQWIf
19jspVgrl3T+48cmSOZwjmAfBo7ydCGPO+g1Xj1XGWIGcCxJsMYyVX7A/urWlZuW
WLkONwI5xL67kziT+7b6KN4qNFPLnkRM0mbQC63Nv3P1NQligg1w6rYwhw68AWc5
lYQCPDbSe0uJf2Vhp33E9S30C29RDKOYkkGAh+yl/dnQoCTAmXtppIADVA5p11cm
fSOj/JGtdOVsR+sn6MZvlKULOdMJoNWcl0IdjvxEPw7Akr0cA2y0qPqj0ZEtKLOl
bth4x/NXvtIJuRXTq2OIq+ERltpcbuwBTBNdros10dHibbePRbprzgT4SldX5hn6
j1BXkKH8SpC4aqAH3IKGxYT7ITqdUPM+z40L+2ub0oTKVoOrl6k2g7EZhtQr7OMo
nq1O0jQg1gp0WFhXB8CdOsHJ3an3QGP8eApkO2qLXJUfGkhqGX4YCSTgAjXIDITM
P4VxMohCgWTK2YTpkF+h1VDvkfJcA8s+gBWCTOxpnEW4BCMqrPdf5denpgw1369d
ldSdhPKKWfftyxM6xE5lOCPCW/g6BIYB8mp3wUFWT7EygtfBFXwLVL5YdNmMirBT
qvJxTkSwO++gV3AZU0yTNpQhvDl9b7GCYSqXu2gCZS8mZ9L7a/2Q4d9EGOgDfAWA
7iUHioIJPY937hbr1P3px9cOThfcIkCDY88KH1EWQcYjJTX19/D8sUDB7Nb62c4f
caX2OJkmFRSqI118Wp8sDvOHwaCchg3MK7knBgvHTRbLxJ3/rQfWIq+4bwYmt1xq
NvwKaN/b3vGUWjZlLwlWVNE18ZDvfBBHpovQ2u4ZoX0n+lP5m85MWn8FNokbWxBa
u4KGLA/iJLF0E7AoilMESDZQCzS7bLpxVQWzERNETWaPL3gr6hipOi+UoAKJx8hp
upLjNt6RwiTumQFrShMuQp7InQ7PRTof9p7oQUbEvWko5wdnZQLYVZcX9iFnCkEa
V3Vjadp6oxjJPbXRdrjCkRAnBWIltLVsBNaR16PrmqHnIB/X0W4DaqZcCHxIlwL8
TjE7PxLaW1F5ueFl2uDb53bI0HZlUxqhnYBwFKxXimIKmY6OGoTkIBQHEvL9rgR/
XP/t9ImlWVL7syy3JIGWEUxb56EegKaKVSgMI/sN4DM6g6FVIlvo8wry8QWUj1Or
D3ru300fcI0p85XWbmhjN3J13AjpP11udGuClYljurd06eHkS+VGg76MxLTQSyZb
Z1h2QWlpqp/+H0HO4dFJgxzPVOXvky6p6WJSqSpV8r7HugTZf6saqUuR5Vq5E78Y
0WhFojkM58mJEPGKWdTHxyJ8Jg5yAhC4AUzst1YKxL6AA1b8yZXRHU5j9qOkxcjh
keBsSMEyiAOx47+1NjQBRDJQcwjwZK3xzucj71rBdpQQG2i9HZg0WNZcOd7CT/tJ
/vYHZ3ftHZ1+GN75g6qD0BxSwXxDj3X0n5XnNJZtQQoX5KAfrRnM16S2Gl6sacfu
odDyl67JFVqBR/I1pCGCWZcC1omOko+cRUOh3UlLFPQ/zi89XOIU2wolzfeN7AGn
2uoSnAhXWndZm148eGWVHwoSwIPwSBLNpCFVG2+BUIzKe+xxb1eiFjvJak2jRtGS
RPJq1slQV5XPGHXpfSKnw+WQY6tMwrvc1ikd1C8xndSuxaxOunKI+EHlJT1W/Et+
FOoAA1pPY8pQMfa79yh9vWM0pfTLCcO1VO3fVbITpSD3dEzQ4Llih1IFV0ouL2Ug
j1K0ejV8Fn0AVhytGAcamFqk9igxRlVC4mjUBuaYZ4UyfDxbNcpt3srQUoVNGGk3
SdwNIEcQUAHSrN59NwXTLpCFakYxZ3GUPWsyLKx87IgyPyNXFSAQHydB2p23gePu
klLB8EP/iaLwufaOMRQxYvDzgZE778RCpWHwycxn76Qle8OPbcHPuglP1R/jsvzW
K3CG6l0lSS45AO7hYDEf2NNXy/A6GDILOTphOU54qCng+E54a/AdqYblEh6+1c2g
opGNC0WR108aUaA29n8inDlTF4PMUS1nD2+Wvssu6Aqaqz25E7TsYHEQq8o5EYYl
2U6xLxJW4i2xDApQ+KD5lH9eJlU43JKRN29y+yjh0ko+L5v/aNAJ3io4iMqEkqIg
ccCZCCHkpNMHwN3UGktQUYLAEqrfhtCzDn3dItrV3j4gYG0LWSR6qziLOzQKmTF9
7a+x8HVK57FnUIwwVLjHOv6yq4vH3ZknQpiFrZaHV3nUV44dz2d3rhqTkSjamwVG
F0gTY+liqn20vdMyct/t0y0XnkjNwK6e6fXXJxpL4E2BFlq5C4l6JDWBH2KBCpWT
s/PvT09EPPax38YkOJYJMnZ/EwaWBCzQsKsnTBx1d3YWW1G6WN+6sYWEzSzrlq3f
yuk5/O19IWbAOaweQOl+cXso4Z3lLSjA5gX0kFmEz1qLc1ZUH9FcTpxUfQAnh0h8
EPzjMrhk3HOgmWsQXI3Zeqx9slWIDN4Mf3uX1FU/VuVtnSdO6MAyq84P5j4jKukq
NzC9nzSY617tFCaIuJIN8jj1/XWEwcjK0t4o+YaOhvORr6ZePy3YNwL1vva1HQPZ
l9m50JoXU8rxSG16qDfJCO3hSEQDMtoF+aoKEEo6p+zSIdZdXLZZIY90Nei2Ykiz
n6kHO3rmC6R1F1yEjLp1mTiS/MBi3Ce5+MPvk2DRvpi6508sxcGYbUe8nt/i9HIe
HEhKp9kCWI0L+7xYwjqrAJZazesVKyfHTGJ42pcod3WUtVHFuyBES1V9ZRxcLQmr
iLucthu4RKUXiF/v7lMegGYUJrUYw7Th+yph2bcurya/ZhinLO281Vh59SWJdyL+
u1nw3OYpCnOXxY3hn5Zs9cuku4JWeXvGn98vhqy8CRhTkc5O4wmGptYswMSk+nVS
Q5fOrZWyqmneCSTXh1SgzdppS1tCCKGdMyceOLLML6oqCi/gR0QryKDBwLmXuEPC
njsvcd60MkIhdmi+Uq470uJr5TJ0V00dky81CZJVO6Ww/vD3AohCe0A7t9kOhql6
waqdZ502dlWFqvlnBI1mNP0P3o33VjSYgsn8qbOK5adSLV39zzVi0r3tZGG7Ak6i
33fRudOqRwB/4DIbCeScNat5922e33dkpFdXX9RxgseGC/CK0PtGlwEstmgU5HjO
M9grnm+W951XQZWt85UBGhwADdPDX8mf1muCis3NlPUgqDrLJ5RzxuZJPYFbPqii
2L5UOSGMTpLDGmeXD47TQsE96jKTPhCjBtGhp00qxjoZjPbdDpV/JzvOrGtMh4YR
qOtLc/ewtDgj3cR/EVLqA40sv1vCC2lT40Cse0sWyuPOdxi3qSs1sL+1jQ+NJdPD
2Iz1AKnD/y+Hno+kEvsdIJz5c85Cxnl5YdBTySyUyi8EHy6oyxPav/Rv/uceJ/it
Qs2hV0QTyrIkWvq8/VBADCZ6U8Gv4sC4YHDTfPrlM3RYasSa2JdyjjIR/EnOk26b
PvW4w4SSK6XVX5WKcgKU4/MZ18nisL8TZqg8JWa4RbaDayW2qf3uq8p6EgZysrM4
hZmlLInIu4famVu3/2/zvOMT+Ab8PRSI2f+fTCBzVdx5skUucU7mNpxTMelYOeqK
dXhiNjAZXcdlfT8tz7qeKRIQ4NBuqj9PLaBBHhW25CX1APRBhKJWBbh9MmB+fvmR
lluSwg6cpA4b1Pz9RQAIdIE8f3kCvmadpwxjC6vG5JrCvYHh8yK9oYg9pbqsO6o3
S44xXJvxFFNIEiuDbNRkaLCPvqMKfqxgBXDplzQbSaZjCKH6LvTN+yfPvOXQQSfF
Os6FY25rbVOpDi5komki0m8jCRht4M59N1pHm2LnhKGp4486ahJyFXwK8obPwPfg
z9W1FHQLVpPBeyhzMYTpE8/wGiBQyWnUcVl7hi/Gy2QBYMpmR76d16obQoryWeAH
C10+KUy1VSENYDkXPvbNJ2/C3GqfDPkn7KT5T5A3yJ3WopyNAf04Dnlj2XSGIO0l
B0rWdhDqm7lXzhUd3lroueINVscScqJW6SAZhePnWj91i0fNqS8GhB3kmqL2sv90
yOKuonsrG92dZQekhXDISpPntlWmvYeA4B4Gq3IUUfr58CcD0TqhEnaYOQ4Cadg7
M15VLgkC1HLwMqyg6gVVKiNeAQ5OjtvnBwKmL5KcZ+sR20WE8G4AgBRSOgj/8loe
I4GeMTvEznjT0rC617VLTZOIT5ULaMgVHb1x5JhwIdk+SsfkZTDFX2ULwDlUMyNY
jCnv8xywC/2SYDrS4NKRMiGXdwaeMwd7HuK3gnSbdBxnTtGV8iwc31IfmqgcWpgs
fqoXrAcMwanjJT77uXTuAFSE4r/ap4caiAiNs9T39dt5YSTS/qodezsWQRusuoWr
uzxQBroTssfUcR7XzqJpJ+aAvtKpMxSUqJk/sg0GBbIu+huJBJPsYm0upefPagQ6
5BFoeC3WrWJT0c09ukfijiqHT04DdZF03zHstyIJV/vLlCs0dQ6lrT2K3fm6k8Wy
CyMN5eOHVpXi0nZdaee/BC195SuuOINsFj/O+7/0HL/8IhiHgudFCKMhP+mDbItT
gaOXbO0RYUyg0utWts82Oz+1lvVsTu+MQN514PdE0g3osqjpYiwqw4ejDwXfPi+a
hs7W+5eCj7TDmQlU/4E5x/I8miuHzSO3eddopeVLUODQ4Z2jFlJbzLtn2i8uViW5
BsZvjQsnJzfdLVkzxwKpg540ifopBUj8A+u0qvwaXtXjqev7Nxyn9NEqd7np6JJz
1lGbq3vJuDVfRGXopvTglnThbGIIzKo8MFftjq6/naEwrG9ZDmVjRsZHvz1fclsH
mQoOhR9kUV/TQUQdNvbgRqhj14fW5/a9JUsGOfTcxzRW319bcvrEpcrVP/Rzxkxb
B8XsBua+rOe4RK/G4ZaTbMXyB3viI3RnbiFxnfRk+yR3Rk3ZIOk7JPvSmzFWLKG3
MPOsTAzB5uIE2OCj1cBvmrZORU2VGfLSEMNiJ6zjg/JwrbN0eZ7ikJNfjor4LDgU
2FYYScIPjatxX2hL13/WFAd776biLkONZAd0ExXQ5iOcMUKXv9S+8ZL+wLXuz8j1
ZG2mR7doJElNQnso0DzZDYPedwXelYF6C+va7k3OafBt+9+qN0H9EEtaC5tAMV4W
FRS5ix4FVcQx+XCY+wo2TAsiFOLBz579G/n+9ti0R9Pkg0Rh9rds9IShOkRiVdzP
ZPKlBuiLkg43p3+lLvEDh0+t3qPysMvqK0nzZjiKWQO/88fZWYbvRIp9yKUg2xXH
iIucw8/3V2SXOe8zyLlgWu+9emFbKMFF4It0+nCboN+qj4VDBzhtv3WvIyHPhc65
NMbqLwNJSL5NYDtagskAPWrF8D/2s8kFmG+iFzOQm+UFoDH9TdmpMABVEFfB+5EN
wlk4quSzfjDTIv2Lss/Ot4LcQFWI1jd+pk4p+9vnt6wCUC0th4XihEA4qMd2ShCD
N6wlAWBxkQo7VFRsw4qHAZbuba589gndSYYjk5LZMZ+BXUvW5XXeaePqDl+163+l
uiaSqhjJEhS+QQidhZf0MT1IhId4IZ306cAhksDsIGscNt8lK7UTTBFOiyz+pxmM
PKOiLPjZ/mFLA+suEbVldr8gwpssd2yB2/nCa3sfLIWxMNYl8BsQ0ok+4t0n7wZ5
KRXTjkhjdXZUDPRiPuIMJ766R0V27QCDdrGqEqWy1dzvuQObNUK4ffiI4alnOC1h
ABHKbOrT9GGghbmdRMAIRMxtnCNa8w1uvN6pKZdswE9u9wJX3z0o/Cy1xiK/EBQG
uQSKE1dQNRyo9xfbtSwum/8Ab0cAFHwyswuq5GLUPGxtjnQzs+n5g7QiZUpRtuAO
wWbAwSO5clS8W2RQ12k7FhtVTZMT9WBz8Zsfx4Hjw9zfLpMasJqis5toZqa8D11B
mMnUQUo4IFHZXy7smxCunMJOhT5r+5uTTXUQtKNAl8DnLWVuKznwPP9YRA7xiBs9
1iCHkEisz/uT4sw88tOf/aGHcjKfl5cuhChQlrbVlFTsbnfoMY2b6fxtjctQlN8c
8pvQaV3uTMVh+5H0A1k9LBiTBdKDeqXitiSCsJOU2K4AGolixoq1ZQyXvNertk+D
qED0OgQG1Mw8af5gHc47O/WCubfSOZBShRD9c2iM7IE5pWrMnb/6EaimZtZIyMxC
SQf18/2eEEl4JVyZ0nHfQfprBsZv2MGq9zWym9RNivBxiNX0beyYn38ax7Qm8jtE
Fj9GOfREx3xdGQgYEHSN9epyCXfBUhIrll1mnvqI4Rmj6zTDUSnapAmQ2UxkB7Ly
TdbSlFSkvdptkIZy6L6CLtL5TFJXMfpA3szu6Rk468i+Y6iuNFmcp/1/VBwQXbqx
JKoKzMZnWMCwAQF3s3t/sMskjz4o/KjFciTTGJ68xC2IwsVpQEwoi17scw2qkZ7c
IrrHPLxuKZHZi3V2GQUcn1EAw4sPRwNq0+gFLqaD3o5D8eQgEsbJ2F7ZtYJRBLZM
EdDO8rjRk1am3vX/Z8XZTBaQFoXYV0L4XwiU8lEPd0za8qIZ2DALS1oj4Z5Mtr0V
70sLdbJAD+lMp1iHgHjrC0TH3dsJ9ME3veNkSXpWfnYzohGuS31DxxHA3+pCClVE
QOQxNER1D99Hzlg67jSnFqFMRD86jnLzOA8oyzmJRXqyIBbtntSJlNhVmOLPFrai
RGBGNQJ2QVmBaeX/EMa5vHtCkHST1lLUMX9ZSzlMtTWVJJ1XhNgNf4U125rSmWUp
IPXq8NOWw0UKiPdpJQyrL4lamoNg3EmDAt26Tmxrm7BiGDDL1NdQOROf/cpXvr+Z
wLXFhp9KGlb5QBvedtjcuenJP0Ox3N2UKS6Xj4HxCbezueayozj7Jfhz6fbro7HV
+9wLvRQXwXYepsJtuzK26IPFBVK9aKwWmlnvq0EKIYl8cvdGsvFJB58X47TArbVQ
Pp7BDscDNPvgRK8wNDiulPIb0/X1JWeIZYwoC5OGA39sSBvhzkHm5n+PA/uXh411
ZGEkHuYl8h8RWktKw/iC7mbd/2M7cGhVUFNHXAZ3kZPwup3r1dF3ynogkMQRnbYB
lYxnwEDvgrFq36X6Qoz7OKACJojXtwlFICDIeoQ2/Xlt4ZCZtE0JCcGp8jZd4kf/
ugYQtHrnaKHQBKqYiWmM2bwT1VDaXgJkOVvSSQaWZL+oGUMNm/S/bNKXuxNj+pKW
ZoiclMwgsgVtACYBER2mHTLmLGEe6VJ5VHNFL5fNt2vk/ByR2y2ePNsVNzXAv360
2rk1B4mAh4lGQJREs6YaOsRl8KfnxKvkuGXGWcZ0Y2RbCJnIXR+Y2/73IR5D5aBB
PM0X7dS5Bj/RMqnmi3kO5G2Y7hdV6i2K+CKsMS0c6qz6HlO4WY3zTDlfxowIKxFo
Gbuvv89Mrsq+acwVPo3uNvr12vSS/poJJhv3AfYRuAWOwmDkb3AStT45lqLpwiDV
vXboMNBl0bfHV0IfUfWfHn0egHCS4BLmduJGtWdc0luOu/AVyC31PaD0/vfnrZz8
PXL2Dd5V1cwL19zet0WQo9Z26yhXGt97A4OTsxpCQ+WzYQD7gXYuH2UBGI1SWWkF
iUJjrz6OxqKtqh2C3RNtY1xMG5sBl00kG8ufNmKdG4y+TVsLfRpDBU6Q0gRaTNuT
rFaKgirDnAnYeqJyBpja4L/Q0asCB0rKrXrrYb0vaHxKVH4fEDMNRAS/UFyIqsHs
f7yIylC9PAIxJELF+BZIpsDT5YiRNpYiZxOJlSm7GZlZegK7fbnwvxIHmkx7pbx+
j73bKpfwRQAZff0sP0/38RdcWleG19G1yypdWXuBHjgtnXC+mhUu41NlN4W6VY2q
snzvlFAxE2VNzmKbZmy9SyL7+I82iT8b3P3zoVr4HsVEgWPgUsL9LfWeVGfsxG4r
xGsHmcgPFLKkPvucsbKEReRL8OOw12vmT8rr+ZJe7bG81JAsKdkVvGNFcka4qEMA
ernGcRgI9i/01XD9UoUVG6joXx8XRZ0VPgDGedElYkdlHvdZnBThEzXWI7US0jj6
w4+O6mQzn4jdjMEiEWlq6ZUcVAGpTY/fhBZUpX073xvr/RxvoqQmf8q6yApkvveh
YDdRVeeveCej1yoDBF4nRGdx8g2Rbbi3pnsT4OvZEhD0hWl+cSeUtX64g4RKz8V4
iSC78oXt6HTEoVq1Bbzwb6dLmBN8dQhq4juA3+q1tu4kAKE7wRtLgsa0PNkTD/+A
03WyCTR9JDKKDQmyVLvpnGfAMDQ4q8IO1rrI2AbRqrGGYhjX0mHa6lCKPOhygFPQ
ldtSKincyyk8B10rFR5CbDNc45QL+sQSMX3O5aYBQBlhg6k1/2etV6g2w6CTNDjB
URoebgdh5yydV43MX/qaR4xgoFuuFtlCTHCfVbb+DRHkFGO1a9k2V1xHUK++d3nJ
8Lai0FWHUtMuqnioxBoPqRs7Wz4TET4AAw2m2HbWc4vaZ5xQitURq24KhHqU3Kdg
HMxHZzS6oulcZS1k6HV3eKXeqmS2qtMSt5dUA47KU+d+KOs5oPo9LEt7ZSasGzY+
r/gRBRWP/datJ5K/o6UDA2+rnRV0MRFPh0gxJJb97eDPoCWyzKOQ6f6gP8nZ/PEC
66Qy7+0YL9wj2ZPxQX18eciOMPEe0O+EE6Md13VpFfVAxFAaEjXVW1fsWTGtU+KC
Bob3Q+rAqn7zEze/Cqx+8ORhigX6b8uW/jr0DCoIHkxFdFwuaccSXNYEuh8kfOuj
RQDfFd2wroblRMI+ephYQxCcSYwpE5U1qfmN8F4A9UPsZ0ljNRXiufXeF1qc8LBS
TojCQ8EcjFRcgSK3Xtoha0+QsFxJyd+pag5UihgqjggpYMgArEVtQwyCD7/r7rEf
oavhUJj30LzInwHULbt6g5gF343r67MmZuW7pNGAyA20EVDXmq/TADQkMrWqU/k+
Dt71RCoY72Fdmh5f1p1c2qLfFZ0X/R00PAfEzqBAz5ldMcYtTkCSkxaXu3/EQYjV
Mrd9ygmQYcCjlxEAausToWio0+8TTecLM2VV8P11ZkKXYFBYuhuI9p2cm/4q+oBc
qpyoGg1wfyNEumMEhLHw905SwZ6UAhrV0vLMzCLf0oRt+wy4yL2EL+kgW3bEY0/G
B7eWjkJwDpzlTXAtQMVio2qsXZNAEazXsdljSZtphgS+6KdRDapInZGxIg7vHHOV
AwUlc/eP9FP5krPr6+iZlCrb0HxcjXIoZPqM0PJM1SJq6Hf7cvQpOb+j6ZeKT8d+
3vTm3I0B73qgJ+BnU1cWn2V5scaJYWToAwRWeIGvREkFd8auMcQVhqBZTBBW5sIy
fVfvvkTJ/iJca7E6icrjbOH40rZyZPfnArUSn/vAEOanX7hbN1Wi8MpYd0l6jIwK
YMG7kNayhnyhtRsYmFpkHgZ/O4DTfZHbrmFVbXhzGeSVIyvgz1+32VVmYxO6Vdd8
G5IoTYZovkb1CXoTqMtookppBwFH5JwR/fxP1oTxlK7c+C7XOaGyIb2qAmT4Hl/L
ZewNM7juEv2LoKkidcuIdTIqslXGFBQxYQQ0J8zwZuIBHEPpfFYbnrxodOTy4Y6k
q/rMBGlN6M6YZjU34X9S6qwEYGn5JoES2PWwzMvufPqPIO72PmdvmkkwjzUC5So2
hMlKRL5cCJ3QAQet0Yc9fjxroL4GgA1stW5tRvq405BMLJc7ieZ9pHFcBP0lIl4T
v6IqRei6SUsA553i3v5XYF0hE4nJQHgv/5r/lgcGm1oHuNIqMdmOe8+JNTADezbl
PFMzX0HCGUIyc+UhcOOjJ+O5648hxD7VbK+eZ+8DbpncBF//NdcR/WtmxRiKfB1G
N16UcUPMCrgEYnSY5pmD2YXlw/dQzeZZFMcceI7TlqPQjPT+BhVUPE+IBE7pX3iW
ORIPw5etxfC0C+OOCMZs+xnfu/T2OW9v/btbf3sgsbIR6fQVReMIle4G8Z0HyJf8
Hk0xmwD+RvGKCUQDApxGu11UvUYPL3rJl8ySurNbsL9V5iQ72OKEURRjUcMc1jf0
GYGDd0bs9R2B60YzjFdZUfTenZ/ABNx2WyXiwyaZjqf7ytLi6cJxNco93YcN69QB
cuxPm1vTPT7zv4ReN3DEXIyAZWAqgUpfrTV7om+oy2cOZyfzoMPr0Cha4UnL6cHu
aNfy0qzeNDKjfsHboCGrQhqlKCVeA5tFtSRYPF4DZGVH5/wWA3iR/APSRz/MRVJq
+9zaBrpjAHuPJHftprcEHYjXpjJdtKSNmTf7QYHsUAelFRa6fa7m1pnyyZxsaCAI
sYshIFzJ9iJJ59ORHGvE/ep3OPQCoODjKRDql2Ue1p9bABEmnenZfwemL1aXvqNh
4qUrzPhZBrAzinvBOH/E6elbexR9YUVG9v5f2kPgaILw9lljnbaukLkvWDQ7Ah78
uohvLPTUHc4IRQAHdXxZI2RBLZmVBnTPR40fylTkv0R2RlTLeXmuMrD9mGIKw0/j
aD/xSzPxWESlKRyTVX8O+CvhLGT8FfGfxePjchzdc1+hPcjOiAmQtzs7uoPUA/Yk
ED/Y7YWVfDtD8/UVG0woNEj3gyEC2mNlj3Fg3W9mz70Eg/2BITUL9Oqvo46lzASN
Ko3sMQn896QE7U7mEVbWP4ZnlAze5ncFgomvXeSHEcyG8S0OSxnBC5rYPM20O/PP
PpeV0EL7YZ31rT4GXa1Jo/tqn8pvyXmKNO5WaRnS3QDfGHE7y/gdfdMYD1KDEDeO
My3HN8WBO+Czl6sVfE9WU4pNj5RGE0UkG3m2Im9Ss01wQPvtTHGhSy8HQFhVi18K
6CCayzoJVanIuohpyJzGIFNv19NLsXu1ZAv9v+jqNTHdOqKq1VJ0hFgdE3DFemYE
gy880aziiJTNfxJmNsD7aToAecUoZE5T1fVUTN2wW6K22W6pTTw5QYDvKI3IiVcG
Eh+98pnaS89rsEEZ22pdGDJjEWV9yjSh+wVhCt4GS4xoe1NL3KIEFtzSe4n/RsbM
htbwkg+i3MdSWwZGHCBXa7Fzt3VbSrGvo88V608o/UamdC49fXVGUaL6SnAgAKRX
CsQJKRUm+fCtjQQPafO3FA8Nf8ve5dMN8IkeoXJRBEzwLPAH+hlx+F2ZEG2SiRup
1HZ0Xi0ymPuxc3xXvkfDvQaY0xxfm0Ydl3VS5MeIaaldpZxDCUo/c21sBxwPnCEi
NeuFy6bhwyOu4iDS+djt+TPmiS9tU/0SSmW76nL8F2lQHbavhhFydLN5sPjbc8GK
pGy+HxG3nHSrlmJBGbVO8rtsgfZsmZN84f/lWgZjt8iwIHxp3HYxdFBn+zLqS7Mw
oiBfaTAwhTex/Ac3IrblKTjJ9Fjh3j1k+xqhk3n5eIfjKffXt0tlA887YSKsoR0g
QiOyRsnkGxsrNgCT2puFDek/+WkoAMXjThxf5V03xxIaNZFMwtIEz8NrHVD5ot51
9z5nh0WsjkVH+KJ+EF86iVXsvnhCV4iKi7XyKzh1Lg4Gok+Gz7KqXW15K6nX3/jg
aLVGv9diodIPOFMJXNKgJ7LSjJ3zkiqYG3flhAyyGiNyhqZ7E5IL8p7lbg39Pt7D
GcY1x/oyusDflmO6jDfUBPKZgvcPe0mOZIG67xiTWnfYpY8T/gCzdRVeHfbaACUp
8rQ/Xzp05l1OhNenkBrcQSne4Qn2YTP3ap/GpQnrNxH3MQoo4u4d7I3jrwqgROJd
xPMNKaLsFkxNpcU1QU5BXoIwyk5gSJ0fo5mxxPpDA6Rymk6S1JrhEYJnIaLi+oXX
pCmNmnh9vw3OZWNtlKjlYjW+J93qxkG8cxJN0VU1+0F1lufskxLKedDVp/0HIJFE
qHiN0UfXkBgejMcfWVd1a/HKsHf4ii1Uls91FIMQFsl2dgo6ZlOJIVSUoWtXS07F
MI3NKaWY0B136un8v3laWnckgqTj2OJ36eU7r6YgaXxyl//Ds5EhCWwovGCTtvX9
x41jJFVgYRgKO9JQWiqfwiwevAktjQla16KSm5E1lrPXIxGz2hxbTLOsWgyRToS0
FtRKcCKlK4zxch5HKW5PD4HxA3+YyaqCXqGZidLp01zDkkl3Cptn/iR7OxJRQg/t
NP1nADkMrMeT4udmN4YLmt79JJ1T14ftJCyyQ3c8DKVR6PbTig6FrvzKla6DQUWU
dJFAevH2l3++0YVT+wXT+SjIeP61pQp8fcrb/Dmv0nPWE4roYB0cM+qTgIjFniae
amoGIMAzK9KE/Ul3rW2ULxiN8CVNRP0DXjtaGaXLJCAFEoNJ6k4MIXB4zsI+JAmW
kHBCugoU6P82w20eOJcPuMfwk1qEE5QH6jZyjUgaCC7DTnIal/7bAwKOdCE3J72o
PTieRkR0qbUkeil8ZOiSXo1gdBWoXod5zoaTVnD5M3vJwmZmQ6XSM8J8sTTf00Tg
ybEXG33j2bkkDP0W1vgu5L8Df/AJQ2k+DgakAue6+w7AuddhmSYeTbrb8OK4UR3A
Zr/NHF8DrjJxN/4uJzTNoKvcWfnm+BvDs3sWarN5IOgiuByqo5XP0XP7QB+ydW5f
YmwROX3JhahfNxhpt3xD28esd7cqQMT7DgibH92+niA0hKGBz/jFLChWh7qnEIe9
r/86W1JhsDMSOKpp6Uk0yZMPSBC5xKwcTf6oFgumb/3ckiiwh/GWK1mMo25gNQu5
unWTWGN3sWnY6OVhyzzDIOaMf+k+xIzxTpGMs7QEjQxLSLPATU8YV84XeS+4T3QC
u8YL1yRbxB28BkfRyNn9RayjGiLJPkLo8vcjaKIuJX7pBKT91LL7NzFEZd22GiA1
tY6XSgQ4HgXuT26b/2AWPd07ECDWBemzxobAWY+R9jlJlDAzy32R+715y/7pXDiC
4htYoO69f6YNxDhsP1tnnJ+L7NHXsVs5SFXDW0JUtW99NsLODE2IYUbJYqhK7NrC
ui0Z8lqD6Gq23qx/778ObqTrwaDNxbkiPiY+P0CN4d5ABbU0n8Kt3RCaPd8n3ICC
YBuksEHqI1QcDbzc32yJ9Qtth2IKmKXnzOVPWBDQRbfp0A198QBN4BzyPNF5CZVW
G/MgBKkw8B6Z6FnF3Gk65juT393DJhlQiKfBrL/FUj2LUKmZ2DsfC5NGn44wOXPe
a4SoSvjp052GmR/evNaFsOvBssECyNegkppAAtX9EmLsvCimL8IuvJOUVUkWvRdd
pNjadfOUCw9watXl7wax9PkmiEvvtJ2Read0wcsDrQ2Q/JOuDN2rTD7MeJ8rDcG6
1R4JDwnqPuyy0C6j7TV8AParBdGwbp8QDe/h3iJ5G5oAf4cwoF2u0C2o7x+3wQS3
HgxsPlHaSIZ9Crab1mARCrZVyrpYP+GMRBLWF4GRXML3vUevORgNJnbnXo0V1MNc
FoP/6GTpsh+gPRLo7N364qwCuhJqP2CgnfNLo6xNO7TQhLdKi8phFghTmLteSquf
TTehQr8w8PxZOJp2BCKK5wDwulGZtjm5L9lvwJWZJUJJhzUrT0kZM4xHdyBYhK4X
O90iK3TuoUrKgaBJeraHYy1vN4SnGmnyz4wTQGsl72F7q9uSe9t9S3aTxlAdyBuR
GZD7Rig+xxC48lv7vLFIIVnCWz790ckYCOBTI4+/MCaLcq1UcVZkk/Q2OdsdQEE9
CdPJtgDh6zHZzjv787PLORV7vUrdNVL7E9saPqNJ9vHVghJmvz1+auR/9WxH7GDP
E9LFRV4RWfX3AeLfR6Y1zYy2o7THx+N0VMaxog9M4LYuO/Zx7THIjvFrvRr8Uip9
x9CQCtlrKImGuk1Pj+E7b/W5xzMWlFNuB1PjSbiauV1sAsE13ifPAJzVx4+P23cW
eoTRSiv5mlntwHW20TmptkDj4j/4q3OdtblURYNk2TkbY4xj8O3uH1IRRlpAReEv
RIOp3M3WO//RVc+CSMfX+g0q7d8n10iBNF0YKxVZbOG8g2cnxfqgeHgd3kl88q+Y
V88jWzyh5yokuiv8Y4xMRv8s5EZtUCpPJGKiqUkUW7eksXR7jzpJrY5RRUSTLVzO
hcBiFmoYpUZicg7B9OF9YFhWrm1u+4uw5e32H39F9+KSLLefVeZimpEyUZI73pJK
GTtppTiO3us6RtuD3o0BbM199PGLWgU+BVP8Q1nuYbQjr3VeRFvrOstMqe4WVBkL
/kG1Lk2z2cIzW2Wlyobr9mMLEf44F5uB6er3SAbuHxvZnmvUgqvtMutbs8rWNiTs
c0mGZDpUiX4/n18nCwn7f5dy4M3D6L3OwZqAdgHEWzGX40SvHYbP3MRPlzzTd+IR
76Udv9aLBj0I5+so8Xzs8JT5u7JrlmM2HTDaazwYxm8D2lHOCeO5V3auRzZXUd2Y
QwFGqUl6O3G4MWkwbqK4u93TH+mmXcldLkqsRakoqVr8jLEzlYj9KcVB9TScRhQL
DiXwsiyhvI+0OnGWiV46FpXXLG919Vo97oHpOE7SjtPZuyIyCW2aedtk57RFqkm/
1YJIt+DpTGzb0kk4CWKfS14PoiI24pdDKaUT15AX15PG7BWGTHjN1ptlZJPSKfx1
2zRA1Rnpo87+gd9mGBHGiBarXcv2dI67uR+SZ6seeOZDKH8R/hDQ/xurI/envwy4
imbUv5K0Ahii5/CmRxs5bxcY9BS4oIvIi56vhJ8A65j1U9bKsxRNymaA3f9h+ydR
r2iHBlqPWqWTqflC5J6QpJWFkAXQW8Prf8Re+5h5iG5NGwjLWcojcALsQ0JpEQGX
NjdmF2PtTXefcTDiloXyPjQMnTKnQsNX5/x5MCsxNxTXaZVkwy5X0Y3qWH49tdcz
gV9lvEM28Flb8pDd/YiPQqD1Cz25V6Fdtlc9hoaCGbw9W0bwnlB+oCIt5M63eVLo
tBZbhAoXJuknFifMzB4JCjKqi13tBOgRPWUasmKaAcYE3dXWtXCCP/vDC+6wYLWa
NCcnTBfFoukoGQsJH+M3kpJ4r3kdpI7t9wlzAU0t0NuUMtqrCPhWpAMw8dmT2z4o
ktlgfTxBtFCxBJ+8XLMrSUMMBJTSMRjzulW7/CwA+QDjvSK6rt5ai9aNc0eubuA5
bNUbE1pD1Pag9Mw3FKGLtSP5kEsWE5f/NHNIRio6DysDz5swtUOjVETAOtICjC1S
EWCVhpqcG0f8Fk4wtCcY9Sq05qQkBSg5UUN1TJI87cujcN+2fa2KC4BVTIGN6oIi
ZDgWPMFkRj3XdGu5dMPVztv8DWlsaku1ZgSwc2C0j0tkdV8D8YJrWWStZoCtR+4y
F1hN5iQTWOxj5zpGP/Yv8LPKh3aN2lbH4fYXPfA4OgN8RsVAKr/Aa7O6poj2KBx7
CRTJYFS9NkCVdcoWawppsass5z4VmG+6m/1QcIr+poat34XP4MfYoNWzH/b9WI6x
yDzBb9B/u+lqc8+nRMmnFN8w+4b/4GgW4f8iIJRFcz7whOOP/m1wif0n56o82vHH
f7mt4pPiErkcVNZaGj4tabn6t2pALMsqkQNzfhhe4RFDlsE2rVjkDP7yyz6s2mRm
4w7ZfZnQyRWxJO+ETHD3cAxLOddKEbGDV4FOEsfQXqwJaVsGmdOeB/TN+KlR0e+W
OeSeIvuq0I5hf5VZRJykg9ruoQMLCClrVFv7x802iOxPCRGWISsplit/61ICborJ
ZuU4fY+OoEcLBOBMzNpERGW0xRXdjHpAShWjm6/jepDJC7R7kaq/elyvw3wWAp5O
HUt/kyONN9OSDDnqKQ0W8GA7rKOwLkglvQ/0GglwOsL79eBX0fsZNxR0IpnhlJUD
czWa92gFJhqs5CQYFg+xCzIvtJAjBmFe3Oi9a9Zauc1weiRfj2jHovXU10PEs9Hs
nro7kau7/3UpVQOtsX5J7zYBfaOgjDJj0f34nRkOFjhFs8F4rl8Gdo8Dn6ndA05B
5ixbdsp0y1varp7Z6Os32Y1jjkV+jZyLH5PaYLQVnqUtFNLO2dfh4tY1NwyLri7v
xzFzmQbDrozZH7ikppq09tHMsR4gsWIfBdOsLtqv73vw/89FmOd2aQxYYv7dyQF7
Ex0Hp81tweRnJcdhyF1B3PHNh/eL/agNNx83O7HV5e8fNm1sOJgMfdiUmRr+VXhb
7RiR/JVjNUg6ZlDH+dvYnMckDamhRlnI/AtDkKhPsRf5DcQLEK4r3tpao+r1kKo9
OEBl9krYI123a+s/V44X6L2RSURhMzeYvWQBD+QrCo8sKSZq4DCM6dx/9OKxTigY
36ErubSf46g15yRZih+Y7EuwV8gCWHWlynRPW0ZKqxRW2CozUrC9x6qhmphFNlP+
mMaR+70U98HZVoqdyJMkTJJX2VGHjel05z68PxbxQdKKKxOG8o69ey71N/tAmftO
MdZPUJhl6nXO3BIEnTXKMWZHeeUflkhXmry0Xrfvv9HfJbD9eR3MDW2trNTHB0Jz
DrLUyTddew7wt1/xsLPUnIEXS3wXI8tMgo0cYiHipcxebm7voODFHg4P67CDtsWI
WGWEOrMFlPrYBXiWmwtf46B5hoJJanxIe4L5wm/uOZHrJv9aS+1GBDEQ1U2yRb5I
hZi0FHsrndQ+BeY8pngBJZr4ApwkRTCvwDPR1ff4fpXlXQkZIeijfVxYT1YsecYS
sKhzsiT4m20nF/OWSlqE9VOm/vBE1T9PnxO8K5ZkcKuzUsSPTnXcvSBHQL0ND292
HZ5aL9L1RLyI07riYPi8I36V5t99YZCUN9BD+J70dsVXqpoqLnBWD2ZNsNIEwacF
nQOZc99Y/nDDZIc1U922wSxcFLzorwEa2N6r1hRRNt8bQ/NivN5/V0Ei/IxamU3q
1qVH7L4jm2qp5FUNcbf11XnC8WWzAaa3W4PE8nUR+52sdBs2KUsULULJDsppRAh+
BCubnxG8J2hGv1a/RtV+DDL2EqfasxpN66xex5ddlOUA36CfqT/14CvIy3WzVwV7
yBcVvfj1XHLwmZOYxR8S+o4iDdeScvjNsJLwjILwkz6trSe1ADgJ2kI0VveN+3sx
3Un3XwfRM9iWfGLHk88083+P9eOYy1z/A5MZI3e/1G+K325B86+hNio6/sctCW/Z
Ocg2Z8JSPFmmxqpsFHxvbJTYRlzHnv4oxw8goFXqPaMUSL6ezrv2lowQCnKi9/o2
cg23JFBUGEU19HhIYBsOLblEQNNaZvlNU5YikSojRvX4V5ktHwGFGIHgTEbIgV9J
t4tmDF2V/kGRbF4FSOXNNHwKN0YUywEbNFPa6XoR9XqPecg93a1vdn2vfTD/rT+P
DFcYq62UIZff1jCJG2fsFrgASiVhy/wZgCJTapnJ5ezns1HTOc++fx93OEPXg+BO
2SlOnlP2OFyxmptcUhMej/9ACrnVd2jfKbI2JNfhCftp8FIKSxDdohEnCiPAFMGY
CXTxcYv+0glVi0ZTx4UkE+EYNbomuwK9+qVCdpEdEayA+zqv2Seczs63p0GJNg+k
lv99yqrS38/CMi52zdUDdlqaGe3dIkuWjEwWu+sYt4gzQ8iy3ioC/g/t011fKFil
jW2sVLGXF1tV7xEJMmYlVinz4IW7iDnzeh9d1MYahWmVvrbjpyR55f1WN+iwEXxy
LzI7BzA84DEbaTJOecp3io+xgPe/o44cneWRrEWS6Y++vmLsVrxnaYhlWMuDDsAU
nmoyI2dMu0zXXRg8jyfnOCDYRAHwe0nVOXiMFS2qYucygvw2R14UPHqwhF37/8Bv
MpAj+dsDXM5Eh/tQ+iSgBrWSYZufbcpggE+QH/KLFNMUPj1CNXdP6R0T2odWd7J8
vCTY/0A3bJKjnSMmXF4IOG7JCAlJ5Km4rvvC5PeXxlS/lVmYGYfARjh/a9zM/U0s
qsH6yDJFMSg1NkA3Nv23fUz86W2s/3FzZJjHG8I+ThOPKYVuT4tRAG76BqCQDAf+
26sPV5dC67UDi4m8WLz5V8Q4T/kdyzWrQzErXl0sN4gXqELIE/cXJUSfDkaiNXGY
PU1zSsPpBPlAXrJVxi57KgYXHpdPrOMQxi/O3cLv44UPd2qSDib9oNrM0hXRq6Jf
GbRFaQBLqr32Ghz8CPH7J1/oJH9Prst+NVe17WNHvr7bmP3KN8jaCDNeE/WeSE1C
npNy+RwUj4Z9IoaY1dGJw9qoOBCSsN1i22AswW4KPxSBn96qZcv5MEzVQCLKdLQQ
1JwsNfttX9GtSlx4+aUR+OvJfpB6s4ZjnQ58+dqmjEM/2TX2rrW/DEwX6XFF+Afv
m3t4NWWuNwTfsX0i+7gRKAxI4vOWIFly2cQ94STVMPHy4NYT2c8P7vjhl59432QV
JKAUBSjSleYR7eBbvX8YdapS66bGvtRwZ+oIVbVzjRREeO8jitlOF1ndnWP6rnw1
4ZaXJKUGIxkqfmusJTWcvw6ZDZgc+UfYt5R7D4OD1ObNBkoH7c5pakXR7FQYeKZL
ffVIA7Tl4ALF4gejj9Teu1277dAI62mOLgo335vzaOy+z8vNZchYYbUD6DAAFkh2
sSjhMZXjP7DxHD4zYCPZ8zLkp6/uR0pMGFBFBh1IV/Aht/1uZWRJRHeiIzCfkOng
JoAvVmuWbSz4GVYRgWTpRS8z3dKwva+GHzo0en/68tgHYOOX3RZQAgLDBEG0nnmT
ObZZuYPOU847nClTuZrEysnpasmGC2UxdlLghEbkOvSeAhwDOccOb2p5vRuiLWYn
SWZZgvsz1WaDNywcZaYPExO3OscomsapZ8uT/guNx3dFAU46HnSdYlX76PMh/ZcI
5U/3PVHBeVrjmBBJzXN4kiCiidFRpAEgbvAYWZLBcNKZCXLmlAIFfLGvkTMHXDMv
ZtM9qvQcz7Q9g9t9FRcpbaDXiVDeCsQCeaCMobwTGZYWuM1CsaMpQ6kKcrD8h+vl
odAgDdTCNh8PRKeDv8EUSeK4zmDscLK1toAtqzzHI1ylO1MQkFlTq/yBP1o2uUP4
/woWZ4CKRjBpG08hTPv5QzFCV0stsUABSo3BFxC4KguMmmqD94n8T0zz4MceZ++G
IprwWtnQuwFA2DJvdjsIBhXKdcTD02QNtBpLZDQHzofCDXkaHVkPvOqGQ4//wMc2
W/CddsI8kuIpuLi2Q3N7YA/+TOwaMr41QLQX6BsIxNtNcXrLplPVQ+1aBzz3Q0PP
MAR6PCMwQnpuUjhp9snCO/jsMoXhm3rp/JYZ/kNjh/Ne9EJa0tVto/RNVN57D7Vs
nrsQcTsJvwHP0RoCRf7JyandiumgSg9eCmH2yimC8kbl6/0lluhodvgU6Eut6Xvr
zp2AQmucC/cFoReUkY99wGF1biEeUBWXB8FtG6G60n/I43Ig1DOe5Icqj6RDrdx/
GpVpn2NUwymipHUrHLcSXivmGEQwsSOxd9+m3KjSFUDoQokN54bPe8JwaNEznRV0
Jh8l5TJctLCWuSRsPCqma927ZtOkqfnmcIyld2qxBq9o5doUJH+yw2uI7EqaRTNZ
mzL41CVbWeP/NvI5k0aXO+smex6Nue07oq/1VGtih0ldV5BnCC69do3Jd0nCRNCd
+ZAg8ahHQ7L7ECleCoqZdzXSk+1X1IToBhtD+jrGtptKvZR/CC0vMmQQXCLxKXai
Ts6PyY9MsjTDy7Wql/Px7oRWnqq+kwuGvwioQRm4/flFZPTQKivVtP5bgVnCoe8K
nRN7saNduc5e9LpJVNnIBNppOm1fLZBEswwj6NYVw/kTWNqZ2YDwvCVjxTFG2kh1
r3fFj9XJJ6uXusoxYe6nc6q3EUxvghIxFpUVFAfmnI71i3RBwt13wKhzWkG+wi98
E+JHM9HRll3BOE80vGixWHgfxme6Whhcys9L11QCP3zspVJd4qhtjXh+8Q2mARqN
aeaYmIYFVwZj8Z0pbVSQJXPvTRkly304jjdah9WgvHmmZwLb+jCsTli/MyKCiTXd
qN7tdNmu1GDh4Sj0yKs4fP9d+fhU/Sc7PeB8eMDZduSzRwjNeWI2s3pZ+FzMVFiF
kUG7IQMptPqSR3Cd7JehacSuil5P2jcpOeGYpRKxRkuGalEJH1/hfD4yMGbNJgt+
wmUTJ2dXCLj/5/iF55wX62NQ1/cBipbPzh+vYWZgDqFL1tTBMUjpU/U9OsE1/9jP
1zRUNHU6rsBQdfR8UtSKUZPYCXuXn1d6NNgzy+lD3AT26Ify1tsXSKGapJnhkKyI
cdoldrmr5l4UV9m6Nsk7DpLbnalWMwvZZ5EyiMyBtG4F1h8vUwXjAfb+Wv5nGgfW
HbSmXg8wZLj8e+BmQkTdYBUrnMV91h4AglDA3KAZqG45sYrkioBOFlCCJRA4IDAI
+4Q34epbYRM0Q816+qyPdl/dFvmCWSLUNEvD20ZcNiLIkahJqSLbW9FiLoF7qJ3q
6yqyzo8gOqqz4DrgLwV1X+W6A/jmRe8VSkl4E7QcVNSMydB8qs+vAKB3TTmUo7Rb
Qn44LOqyaxCC72zQEdCKMjVgkEFfv4hNQNR37/gy/oMnf18WWwu8KO5e/jfIdfQx
57A025TqxQ7SQzMUIReEpjBvP2XI/VdcLmWz1/XjD7i1ZDgj84HPcxROaKdbv3W+
Cvv32YDUHocmIzf1zlq5tM07lvkvk9e0Op3/nTcVyBEksrl3ViBeoIkwxjWVL2Q0
+ztQ3YkvPX1M4ByhDEx4C6BpWYjANO5EB44sXoGL9NVfCfMlXyC8h4NlU47ejdx8
DOrSNOl7PKis8wdNP969PXhsKFv67t661MXgSDuKiZzFqOSDxlzO/Yx9Ii1Z9gey
Ax/I/Tz26Wxim+/fXBCH8HzXHlJsakCd8aiyjOW3Z2c7nYmGFHTKO7BwiEZyPzoD
M0wnFqyZpkWGVthAUoQGj92ntDz+jn+1sp34EmjJX2ValRyN6Bxj3ODK7M/CL9iy
dMJGI70yG51n2gzG23cs8DTTIVHGlO/Jt+W41P6x7wxtNZRh+ltaKHCV5MjmoEhC
G6OUR2/Fk8dJqZYllzlQujjAOdYWdp15X+3IO0WFYyfMq7TknnS3pZZa5swMM8Q2
oEseI3u544V8pmM1wjar4SOQpfnGYVxGq6hPsg/vB2bqFoyv/9vcnjzyg4UA4uCT
jo+HJgIwzxI3PckjF3QOA4Zk4DPNJRm3pqzNRGe32FPvUp5hOiML5YMW2XUeS1qi
9MwN6NarTVJScmJP2R95gNRXuYcRpTIqAm6JZXmkLIjCqJf1wr9eaz1THy70JQ3x
yZD7AnBfF7GVABcxV20LgNzD2SaNACCi2dIfA7NR2RbftdCj76PZUf9dn5XkCPc9
s5CQjPtlK6RPKp2O5PmDl4jbIfWC+MaJ1NX5VjJR0PYnrl1Wf/wj7zCOJ/5rVBm6
KIveY0jsWxTO5xVWjWZqleabPmf3FHSQ+tZSX19NH47ba94uae0NpXrtBoSfZaYX
EfMoJDRcGZFyoSbQi3LrK1WLfVz2pLWRR/FXYfS15FE4Sn5Dzt1R3AvWhO0rpxC4
T+En2Xv9+kKltc4XqUaoFp15LJ+YUzLLU0AGI0OKkylMf2NlJPk8/N+dr40for8W
ubyMUQlVGOPVDYBVgIjk3/Z2dD4dmchaIFPtX66GoosAbenNcz6cvzSqZ3BHjQFt
slxzuS74UpyAov+onfjK/xB8DnAc7nIKSQVxCMBJ8fOAJ1kgunBeA64dTzWEDDzQ
+g2DmxCrkYSCB0KcDwqtPgT/kFD3d1+UdC/+ITlotyraRkF+6Y2M2cbNmOfrQ1FC
fib7OevLoLB2X7rBVe8H403E7FWS9zpirF5j2Sxq3LhOgd2KJJQ1bNZ9na5VeRNS
SZQ7JBWMywwn5RN2FxRHzcSnJ+Ve5ZoP97QNO6XLI+RIqwJxtUvPy9axWhxKkwTq
EfdlWJYSjWrN4dWHDAIPW8UtvE5MNL0RsL2H+bfjGbdv9xx2BoeqXKfq2CZoTbDc
VtaOBGgnhBbR1jfbLmykQC6HLAJtlb8rH5VOBs/MlAfBklTnW6xkSkC0G67biwPB
i/kCN34iILUfAijsRzq+1L+s6ljGa1MZJPYr1stv7zw1meJoGnwAV/lsZ6qdumPG
qHfvYSN7xc7G5oenxAEStj/mf2eA8RImE2y5r2nvzjUmWfFZ1JxXgUNBYOHSE6WX
KQPu87ytrvGmkxyo4Qzcq2jOY1C018D3a6As5W+Ci1Rd2eLvTtGBjZKZhZRkIbqZ
SKo2Zwaj7fxV0T3W+FiZgzFpI9Pg/tyso3grmUamWyCASkWBgZts2aqZidhiyqYJ
M4a49excXpU4vQo0LY70rOBlVMWpofs3YQRnVIoGpoi0HZlZ3Hz+4AE4tIjurF6T
AVp2RQgWysQE+SZT8/7XIpYjF22RUTAWQ0O0Zydobbn7A1vf9InV9XDmSUY+C2Ia
AQI/Xo6PisYhAMHTwelFLi37i3pPmjW+vcJHJu6Csqc4hSD/f5NCyl4EUcDkJyHL
DK+WZdwBbCoBdjNAxBwIozo+vF2P9qDCzxNKKThmwDxhqIPuHw+/buqZkhc2lFGO
vALWbRFh03lAZtLqEcNmlwjwrGlqzPWHuyZX3qWK88OB+qZjGtgNZp6l0BXrStJb
rNj3xXhJLjafX5X31wTxGuwTRX1U9F/ctMcC6bYG5waztDQumXzWkumVHpDelNL0
sEmrU1NRv/MdOkjHwYExNr+vCrznOJb2fGzsYWPFSNqXlp/oyp1HNj11Jj4GVObm
n0KEpPUFzR57VErF24GW1soQmWEvAG6AkbWZd2VsH3yOHyw4xWQX8Z6J2NqESgdA
ftycJZFgQO6rOCon3wUIQ3aHXK2b2+edStB6+kRVNb6WZz2TuYsuBwevIrBaGyKw
cPUbaJPQvoUH3+ISlG5w/DQFE3dnGAIzjlpPXjpvJuAVnlvLwne2R4RuQ8Ku+LVW
5g5yPG8i2aeW2f13EuiPCz0pDvblF08PQ93gIUaP8WHTucZ073DX7ZXPtmuc5Z90
ruEp2kWSDlPYBOde7pelneGb+bD2ZjLKLZkoLLpvd6DAy5D5y7+D1m6GBP8gHkt9
fj3gCkFbNeLmgoZOxMTZGgNFpxWNcO1CmDu7w4eACs5QoCC2KK/a5QHJlpToTs0M
0fNsIgZFxWdKekqbUBbM/RgQKpNhPUR5yOQ0vDY9s9z1uzJs4OmfFakp+Gk+UA/V
Vi2imyKOwZVLV15NhDgYnzQdDKKAWF5gkqw9UiMDIGXXs1Caou/bUgxEA8BbMbYG
R9sdbDmwDZGRaVNX85YtCIb5Vnm1owQ+7qMzP7b++gOJKMrc8q2IeGIaqKVrrhqO
2H9Gr6woyZN2yQZ1Qpxbj5BEW+1BpzgVAMOvQYy5d7nw3tSBq5Ozd/PLK/kPzAYa
ckuQx7t2OvImPSRBu2aojtCJMROJ+EU/EKqT9PhlaAKmufUghMuweR5MvhH+jGcI
P7POrCnznJ+iU0rHQJYdNS+b54jUFSEOOVC6jf9XltaWDsckJ1v3bvOgx6OvBVDN
d3FF5d8CKjub+mvGtuJLE4JkLAAScPj+FcFqh4a//d8k9tkGrsWpVZxwi5WgCWs1
LUeHAiEJHx1K/fJyrMLjypX2Y2U+9rzLaNfia8k9zeFGAhM+nlV/I+lpwDcnb9/A
1C9264mX4CxbqcU70Dont6oI7Opy21wrGc8LKLYYbaqtnTjHMPdv9K4ZWowwAqMX
0s6RaBWha8LLJu1/r9vd8j64kLo6yY+ses9HZH788g+Zdfn23EA0Lum6DPnG9TgX
ot0BTbKhWdobT8Op6oQNyLWsql6pn8L6gUC3ell0a3ZKdsuc1zrWyQ4b4lvKAT+t
BijiHUEXuC6hNUC7zMTlpNEZaXfPm3xetD7GYpOGJqyRZex94RGdYcepdYHHa4DA
44snLhhguBLJ+gPyIC/+sDtaXXrkcP2VQPXJFU2jGr5iUm7a73ocU28GaBlr2frd
EXR9FRy7DRIb/eWE/xk8x20khinloYbZkxEeWm+XwjkXFnCENoipVmofZMWVYqBw
qYgU/SKuz3wjuoG1G0mDbJTXBULh8c780oxhNdMR6p56xzrhWjw0TOd8ZKS5jqXl
pSH4P3QJ+YWef9h1bTxey3cN/tEYKKB5Ih3WDkMN5wOk0o7Hcv+mLVS7HCmXdIwh
Gw3fOwWbonZ0YCYulSi5uMtJGy9oEkvYBj28wsqmYmVEtQPFskxS05nujWn1R9QM
MrdesjIMulMxxPERsz04JXF5lrMxhTg6DZy5r1uY7hIyoV9nJX7ZNVvble5s3ytR
OAlaRdlHjeD1mdr792o1vxbHallC/06wK7mE+SToGco+uUMQS/VkAlq8+O3cNfh3
CpRIogowq31eYZ3InL64wihGMzc8K/SnAh74EFjwRx8EbvsQQkF1ZxEAuu2I/yu+
dgdxVdFc92L6tSQzaZH5XIo3/kVo8iDuJ+MhsXCcBSVH3cAiodD0Xumugz7LJnI1
1mGtDXwMW99gXE4hxRKSw9n/T7BthPTqsz17+OjubyLRoHWhSUeYP8m/Zh1i8GM1
1ETx8Q4JsZlxNRLMZcghTWmoj5ZJrWgKuyHhAjXznbEFRcDQ4O9uC6YI5C9OoFAK
xYTMkd7al3jZr+XPG8FSvHwyUofs7oLi1InhdEXm9WxbFcQ5P8TnRMe3poFNC8AL
sEabY6n6I+gs5uMoDc7JOrVQmQwUeJkmegbXKNXslx2/w1Od3pniNu/F+mJ7pm4r
SHiON44cZZJUyiBCXnERq7M/dq30WoN8WGEc9rya0bZz0CuwnKKbR+fsxHpq0zg7
rDNU4aTbFjpihNfEBo2Kx2mn06Mj47BpTEZ9AlB9KJsBThcyNrSH0trXwwXpIPsn
yYEAFC/31awjFL0LS4bfAGed40ENhUMzcW9g6qI2gNH8OPV1MMdl/Gd+evwzR9Gu
Qe/lzou0AqSK5/BvMzYZBZ9kW1ztHttCvvyRZml1GmCl5do/tCmbR4CfB9m/zwVk
Lq73x6rS7zQBiChlVMEfl6vRrcLJP6PAKld9Uq43VKqqoqzcjhdP7ZRWCXbJquC6
0UKu9CZvTijPPqEjGm8EZDJNge8llaGgmNwyXFrNlA4aaHc9kKbnWaP63Irk060H
27j7pVVRMADW6wjlB2zLpr00ffYa2tl5+5ZzErMPfeAxvm2Cs1A/IRc89CMQg7/F
v2hBiz8aJdMbiL1HPzQBr6sn+GRXGHBAoulUsa+pukIHvyri7CGZU3gjVxS5b09r
6spXG+PSA0jORnLqA8/8YnoG1Xu0EMr+D9lTzMPwaUuWqglw5m2ZsdZ2WrzEy21B
sQHvrBn+XpNW1Ux7jApPnP4HPbszDshsDpBBy1GXXHcRx+mkUBzsWQl8F3/LkGc7
8JyYMEYyYVruK6aSOy/Q/ksFieprJVZw+PV+Xi0VEdZwZg3BE6o6AV5uu8h4+sZH
XbOhDXGTp2aubQUN+Qr3gKeGMb/ZR1JADiZxSxvq2MGYBdUx52I1aOVuFSqyP7Ln
OjuWXKc4ABK+zSplsv79/LQkRYFntuXYBegnXBb/WwC3lFupkcm+gBF8nL1fW/18
8lf8dn2NLUpOlzECftnVzICCKAA0BMSBFxbJq37N3/QoH9Nz3pw2MAOYF+ngkG9G
NrRl9FxIZllJCPK8JgbvcrccCz7uV2WxfimTZO3Xztu10Uk0D0O7aKJYESbG4OEh
1PhDVtCOlDTawDLe7lkHicARhHzTNINJl+yoG5GuWpMThv1yhussJb0uwS46dnhK
14R8RggOUTh9kzFnhLo8hpnRY7LHQ9a5XcLh73pDT3v9ENA65nqgd2qQ6iay70+p
Xg55QMZzfQoYhV9g+BRH0S6WEXChyUzAy7oaWnAep+jMiAlHPbSzWseALXEd0XfR
GDu+kneSbLxh+90Q3pmLVctxek1K7W/RwX22Vl2GlopyE0sAOy48dHsZSCc01Dqv
eG01ooIGpRjJMA7b1yObRVlgJFMimwbISEFbtFiEgLgpyOsMchv2vMVLY/UR+wpZ
d+jL8WzSu4reOvjdAkiT2uNmEVwOWk49iIZSqvPsfPSVVRoWZ1hDLq8cv1dAKTMD
+YrIkpYJLaie0ogeidz7MpoSTppeKiKDxG1+X76ZPYRB72fbivEDWQze5IvkdoKA
Dud91Bkt0dMY6RIEf0KCkb4R38KAHHyteCir7kCnakvEaplZYObM2RbAjfakpqMK
TGvgDyYgqGevidgDkS0pA9C9ggxmBA6YiDZXGR4U2qgufoyXHF4JCWhQgIf7NmOR
MaieUKdrGnAg4M3c9QNSG4DtLkwh5C8fmX3NHSIq78KjGK/xnri8yhwbwLzUtKWB
0h3nvVUZzS9nag78Ks2d1V61SkGDqF84fNdb+iXdXKQXUHLA1A459PotYdlXf7oh
5BTopdsX8rMOLN6iE8ml/YFLdaTSWfo+3S7hAJkN+19MlflJSi+ErtZ20joA8rkM
cEo9ElZDHOrIImOTR/ntf2SoGiMr1+NFv71evXd/at1aa87zbE5nIeqiE7MXrIov
1mXt+Z4R74F7JkHmMuGQXwEzRptDWB5SpXe+fzOuWO9DS/PTt9nMWdOCfO2uKs/f
LahgQ4xuLkX8JUJP2tF4MSKC/QgxS403U4Q6E+B4ktDHCmr5DiBkpFTATix8Xo0h
JOc3tz33Xoo/cVeDHreBOsDkf8fGOr0g3lTgbZi+BfF1twcKwoAq2ua7H/HnUIsm
PKLkQa3fW+FiAT0PVhdWC0+yBZgO20pgHowX+bSjmVmu6xTiaCf6D0EFwR2QToE9
JGm7XM/y+Rz0ow5FfdI7CRSe56qmvKwAWHVc4JSW/GPMRSxdcCz5kjX7bm/kkfnw
iv1GbG1HI20SQ7ZzvSc6n8oxc0dZvc2XIPLTL4VLbWROZcgXno3vzunbJ8pPxsMU
eQtXrqrEYV3C1oanj7eqgjtixoG8SNpgiz9jbq3DkLsr9p4TtyzJ2qZgqF78AQOj
UPfiBfDZBm1yHsfnCt5xKWg/HyQWa3TUaJpzRjH8qicWrWGNSdHoVwhVM5FtR8AN
Zc4fE9bpLRV8RfgDsWUcMmTqcV52AN2A4gMHAjTedopUqM/B4V6wDIwJI16Q5m67
/fNV0RFvNoaBvaPloY/fpaykgnKSG22TFhla02TTl+Xu0WaOfnJ9YIRrKBXi2iwC
TA+mgRyQH9yrVwDdSpnwLqrfPBq8az2XBvlupF16087fBefsk6xm62Zw1VGZsoZV
LlBU0wGkIiBrGIn639vSj0V8M2m5hikbJ+As8QK3TYfOwICCEMN5+xF++yODpYHx
pMLbds16XrYRnM18SLWENyuRUCkwBfXv3ZqNw5/Gkif63exwXGu5qjXaxhoMaLqy
crX2o3DxjRXJXz4U1a0OC6onhxCmYxbstmYud+yyq3YR4bwvFzeQrNy5JmFZqjUD
QMi66Ko9YrrjxFHlK19ejCFcaP1kX05gyjMdMLfX1byO4c+OmByufG4RZqj/gwJL
8+kL2v6swzKASZAEIpitsUhI78+WdZT/vCFaV/V25V2PF+b27PvTY3bVvV7jBAox
NHntkyrMq5PkP+T0BpMwkJ8v0k+03ygrZ13i7KLvMn3QrVvwdXba6O25HjoCNVj8
9D1L57bSaoIsL58Jqv67hsBOk9yhDHqd8KyiGKXIYh3GbbdWfKGn7KEtp78ozl2Z
nK9dTO/Kgxnj6IaUMGFsOnLPa7uuDF5DwaAh5p60c5HCY92xA6zvxkukR9xKFpuM
6vEMZgE+MNELHrgV+0JQhs02R2y7KL4Fa8b5uewACpQcR9HvSELF+4MUGXgcg1kz
F5OAoZUQs7sl5DBKSdlF1UiF4697LAIzRXvi+WzSPJOrJIoVHePmripALEH9VP4r
22QhUzhJTlBj1VJHRSBW5rffFn7aTIvYvmw78rNNK+Gg+yz3gAGL9ycC5ibHU/QH
e6DdaJmqPpx0jfHqrU2iNZ4gbLzrSo4XU9PAyqSen4tL5BKEVo5pteD9/JzXD9ZM
q+1RzXDh5+3VGa3zdG4KGuVOJoVPZ50NMCRL1+kymghYbqRWB1hAfahtguzdE2yC
D2lwqyULbdGqCKcqJ328n8J1dHKLi+/7T9oaVme3ouuSq1OcKOyYihPGZjBw67dn
flLLSnoKX7S8djm7r5fnUUJxd/WPBTpyM+C6okSh2tN4iRUn2veiWsRoGSYfKSd4
STKx95vWrzYqY56l3MAe4WVP6XGGLOkWmuBungDzj9qs1rSeJw3SXI1gb+w+uBm2
WGP9i0MriMNiWdYs4oz22qhooQhtBShtQr3M8xymBVYFJuB4dxt/DF2cx64OYtFp
kv6ouWqz0B571dnC/XoZbAaGjqTaRO2KXCTOU/Ig9X7+bfaa4hkRVnVqRsiZRFNi
hhPOQeCOjHPAU87e/MEXuG3x0Jq34ouC9TYiI5xdKq7Bwyzz8PBfht2wjaCSM4IH
4BPTokJw9soJffRjY6epeLf2NYpIXotgkEowi7jiMJ8+2nuxUW1RdSXhdObv/JRC
kt74f0FKCCw+6xrsDry7wMtQ1kd87mP9uHZeqJMnA7zDDjxKwElOn2G+d1MRGIC9
AY5+x5RNqDMcmNGhXeY1OKClZZ0NYVgu8SxYjenbX9d+tCFL6VI8XYVn91GFxbWk
+r7SFC0+dXyAO5HTr7ZwUd2jx0X6uMYI+AoviNlqtE6/k8Y0PmoPvP0ELPiFbvrO
QiByosJZZzg+OtWYe+ROMM91NfSV3qCezb37oaR1HpDDEa4peyc9UYvrvbAxV/C0
es9v6zZt8WH2K6Yt2kYGPlTWhfg0B1uTsENiBBLSRcmaAliwg/ATb3g0qn3AyQP6
hPHtY1OVvmqWhnLaaHFu5n9owCP17+c+QnDeZHmHjkRA0ELO3q8ZesTQOvX33qim
DpPCt3nOh/yXb/u9x5pYsmC/KnubG1Dmd9Cb2AJvxD0WC+hg6zwrTeV8KTo33lbk
pue2XuV9FATdebMiEkw/QqiJN0+4t4qlXHbf8i9GfP0b6Qz6XlumB02Sb6eaNhx8
oWzB54EUh4mcr712uXceFQb/gtpUzzKm5M9Mzf7nJdDZwUUZjMfJqX4/F0F5iugt
tx/nNSZWk4C18xmo3i088xpyJenEji6pin5w2BRigI+EsHx/lAAGaDcHBYQhg+He
vE/m3ok7jqoDv12n8q//J8FyGVi1d3RjVQYPAqLGHO4r1SKsCbsyTVWVWtzHeI3+
Fh4Vx6HL2OIoRxCle2N9umx/oUymeyyqe6IZc9bJn/AnClMkvANzc5azdMT/DDSJ
nSP9lw8dPoVeBxAQuzQI5NT+mMYSlNr2QXjl05RB3qqt2CQIHEqo9s7QfK+JONSn
w6B8HP3ePr59rwQDJWTAyGynOcKsxtZ73T+zmz//ylAPKC8IX8e3aWW9Y6Xh+/F1
z2Fvmm4AQbXXN2a6nTzsH5OwOZ4G8b6QpN3nHl1kRZgWPFb2nKXtuT6SAfzDeWYN
LeODDnu5CA5PlZZr4ReqabaCDCPigN5pi6yj/T8kA2XDxmHb4ZfufgUia6QVBRUx
rUxkZ7W5hne2bF6MGj4ttjc5fsmBEahDok4z/uIL+oIbsO4art/IiWOCtAHbrZfw
+zYtk726XXn4C37maAhurmDforB9xLB/8KUhs1aj8gFML6KVce8efXkmMv8WWKhJ
/M8yycwW1WU/uIoRKeSvFwWWGKN5HJ5n4vwY6xMo24dSamVcJsPtWqfXoq5d3e7u
pFrWVC+6J28/cjf6dxGOJ33Y9rc/F5DRE1O2p7VDmtdusWWknNjN8wqyzOHYrMAQ
5hbLfG7BitMzJCq+7e1OF3CY71vUbDf9oF+dxbg9WppFGHELd+F1KDYIyBFx5TdC
GQd5zdD92R5FvjZdOdXwDmwKINkQLqnyUZANZFfw6UhdQ9XGfgWzfmNRYBo6S3jV
AqLW6A7IUsfcSbWs4H+ZTk+/uqHv3wVL3hUFXCnRXQOaI8tU7vlMenMmtZOyO4Is
IsgyGYh+WrWeF3j+MNClY3iR/YlYpVKVld3nvheA2ODcGULMyUHGzxKqpFYc5Ltw
7rCzrWsu9zOmMsN86km08mAkTZn3MGhgOewvhUtr6VMUoxMIlgk8ESMWMmqjZLRC
18mCFdJnSmOamw9FH6Oo1UwH7NvnVLKP0eZejfUVlIroXlJLKFBEgHadjYaCqA56
qwoC1Z2/0z5ucqnPDgAVXZTBv26bJzPNSZ4wRnwA8Im3zBYGk3F6Wbz9ryO+CfKk
MSSnPYUuVIE83Ury19zWdsx+mETuI7wpFDS1W7OaFU/1kloUhug5yUCWT62QYik1
pHa+NC1kQ4q4w2PzcJDfyDszhpRinm0GW17VMxdxHKdYxu0LaZP/IePME98x0G5J
ntkTGuFaTVmqeWJy+UAFuSIGAM5wT5avS6y5U4cRm4xnCBHxf79sAcIKYGpd31m3
92trcq1GOugpqu898+I1aXJTK+FxEuwGDCFKdrFoNYzcoz/JBSwURxTxwWRxDzVj
nfE0jDNgry2IsoU9Xvdq18KNrEHTyGqdgcgVVevD83bynrkxrtaSU4XIlIHX8f9B
CKJnxLGfJFKhBVdkSnAFduXYqgyEQIOPsn8+LXRRSi9DX52WGcZnqpJQYOizgMrG
INVtKEIhSUZ/828mTuJDc6USsL+wvyaJzeasTEWiSKN514Hxu7oJ0yJKveT/L2Uh
W5Z2IgEc7JL4hqyoVZjqdW76k8q1mO2BvexeVg1DVcbMOohdaopBw96k8yVUVzit
x/LSVxsbsEc9wqSI9L3/6Bg+XdTNEg/xLi3s9hV5rCO54f84UjTXra3xC43hUBGY
ei57bI9Mfr+LrP80pneIPaIDxMirG8mgVG0hzwOHGXlwCv93DiffHQ+V16YTqiXH
Ay4DOIbOVkkIo8Tf+/MciRxKdPkgadvKH5z1OQIYcYAEF8pw4RlbXrkoGXB4W1L7
EY/xekoG8eQAEPUzccLzdz3RcHLpM4m9/Kd8Nci9mIMHc7h1pw29pDO9fAI5/pVN
BWmeCO33CRpNqkrgdCpjTuWaHLnk1c8GG8PW64VTdev0WVZ+AyN7GHQp8NKqzXWg
yYpbfzDqqSop19EhJ6MXzu9mp/Ik2Ap+T6FY5YdXcRHDKDi1H92/asyO69zzWRx7
nJ0JG+r40CWzCXfB2szDho7qzArGwDZNlLV6FYbzmUZhoRzcIBB4BYEHWaldG9P7
sT2VB7yphMZqgzcDNyb+ANBGbtYFjoBDBikk+aTqc2cK1rgE2nQGDAx5VZfV4yMu
kgL3SELVj8Tiuypts5ovT7/FURxlf/cy5d54uYCV8jRaJ/gXFiacB/JWMquM/FnH
5h5Vqp1Lrji/8odj5scYBTepQNfmhKLcEIlul21TYObAsz/qlpfCxJG9K13cme3t
NuJXGm4oFPtiuPA86CZoGPdYS/xz1jH/KJVrohjmEka9bDbcac9Dfv3FDrhP5/w8
lABOfVvgz84q3so7xjnFuLhb5pX8/YY/FKVbtXtXtVBbDvDpLPn894KG6E2XYsLt
QRgYJBqxAM7m/Xp4P+IAtqtAvJdkQDYhAFGLRfiIlQ8/2FA+bPzF/iiYEHG38FJ9
08ve1SDF5Pw9zUqlanB4MWL+qY4w8C87fTPu5XKUgNhZ65SVnIVECMQ75/+JLO3Q
WTYaksfoFY8mqzT/aEZ5csMynOQB2g0EaI+GJIiQU7aY5wSvXOyAl9q0FM6zWFYh
2kB2feyF02DjA+4K9mtRXVo1YRPq0mT1c2y9YN4hjIAYzyJIRa1OIwf0ZOwKanLP
IIaGw4csViIZzVoTgHa7lnP2dva8XVyumw+J7PPtgwzdpLf0HoCMjhlll/LadoK5
50saS59hgVrcPODz4D7mPXwvglBXRnfyhlIXqftfXiBHv3PTCxKukOtgWQUWDbDe
aS6VQAqOw+QxJ/XT1+6ZUjmS3uOtTmH5GJQIL+8kd0DI/xkSXqFWmO/d2AMOrvj+
ces4Dz835frtS/0/AWJtLnQLMli1zFVjuMn2Hkvd4HbLXciISqn50VqTnOXinZ6l
sjVpd5UmVi0Bt9v5LfsDKvQkikKaxsGbWGYWn7gsZxcdijloJXvbPKbwfdSHE4ag
vXmAEsbmUdS9U4QAnMPMEmk2wvTudb0XV2C4sY6v3MUKcLhMwR9Eyju1J+wXfYVj
C37zqhmW/zB7I3QQ2wv4EWHE98HBf3kpkJkwynRypkgNFpKSC3+InoKC9n07B3Pc
6q48cpu3BerKQh1jCLnofXfJEb5QmCT52R1F/W0Cm1+Lhx5lIJlNpHn43R53llw9
j4UmIFQkv+a0LISgz/BlWvbGxLS8f6s+UMPItB20T4JDhw44RPvhyhHLpk4BCmHt
Z54p0HBl/7EoQPzht9nSM6Z/h0tG63o4jNgNx3TsTamNMOhQRv21NU9AH20SGvx6
aT16tGEJf41iCCGjX8SGyFbWoUrYDCWC5VD1MGMJvjM1s//9mX3OZ8PlhcRAnU+r
eccGtxRp1CRzxAiiQxDfYbLxb33PmIKMO8JLy9A7GQv4EsPEXy2sC7DSP0wu3Sbw
Ue7lvFxEnQyZtzE7rRKHkBp+hOIyPa/DrNvcFFAkUGtLVZovSlZSup+XsyGNmHZF
HfhhEC88PlD9ok011hxFRchFVc08EyLANzsNRWrV5EAC7wuQ1a5GWlprrtUAnu2V
AwfEjo2jPdLNKM6CfvqW6S3B0yOoGvWNL6gwqjmEIaO5wuJCZNr1U5Eb4q5b8eXZ
vmYh/q4pKPcKuwOqq+rBAo9Ypv7nf++lhhTAe6DKg16iMpepDKZQaoSYNAXI7/Fx
IMie/rFjinuPQL7kBSFznwstB25QVCak8Nua8N2LROMlVfBf33jG//o2ti2iJSx4
OgHJCc64rkAoo/kpmeFK9+qFeodNVU4yxfKnPTozWUvHSoBss2hBusi6gfT4F1Jq
z4hkpzS1ytL1/ktSldiZ+SV5/vhoGePtq80TKkI8nexp3BWEvqw/Nrl9qjqy5SP1
qsus2afpuxA0pMFxnBl8ysOPdr/rTHz9KhYrpMeI4PAv+NvU7rQV8dPYcx+3vB4R
DOHU5jswm7D37eik6uVL4X+R1YMTBQfGHnmIqKx8gyw5wI8L+tLQGx3DFRVic6I3
JD7W30t7nlE7ML3lhfWYsS56n/+9sCzmgqeHa9JMptXSm28bqeV/+oVoiOsab/df
wX7uSiTisfWlsXOS5FTOezidJ4+b69KS91vyVs5noJiQHYu/1ojw+5Ze3Liur6as
Y6CVCE/ZbRbzxypmfRDE+pCSlc74mmTXC5pd38ZLSRIo5Uhd1uhc/0+RViJ8pJ2z
BEHZfg11VPKQjJCJcYEEtUvx/xQRqXBnI4r/iR7AgtYG8PyCOvZFTpMzbNrCUuwB
JadUlmJFUqZXUTmz2iq+UjqEMpp9NpZbhxPYdPGzjHhP5JxqApCBKr1z6BmS3Ynk
/e1glNQ2m2p1VDcv8IMDA0p95RijGf9Kr5VhYcE7A37Q8DmFp5sE02QJiMveYn4u
dwHoW1kF9rR0OcEX4fs4doHKCfdb9jGdsJB2yPUlNM7vMeaU+tzC7h6Rxg/YtgKm
3a7fXESyjX9Kz+RuNaYlh9emnbOawZE4cCjqPPrRsSSU2zLu8pAn4CjzKqS7K8rH
eENwxPtKJYX0RNC0yEliLmWpnOUEDyB80W8gftbeRwXqz6jO0Aui6o0X4Q0tg739
TQ4LiguPbB8pkqX5m3cF1cw3npwBkH/7yneRXPGQzncl0pUywWcXUV3h4lEPli1S
NActMX75uDb0FJxDdrsszsdp7LBONI5uBM2z9XKraz6SgWpEN3kPLD8k0qUElZRb
I3L/8XHGqZhRa7CtyYoSbF7de8nAn2lcgmTcSjYHoXHJGgBC0wxJ0bexloHQrgxL
EaLXqS65NJwQUfLQ6UAEDmheBxQpxbNOdZ8bOzC/Hh5FA4Ba3UQmeJSTJ09u3QhL
a4GD0D8fdjmv1WRF5d6Lv/zhE2TMS3/aaPTVDB7Kbfl+GLEonAPJLEJdW8WkCBRD
2YCJRE2piddLsvqzu9SVegy7yxYqpXXTWxzoVjsmFtxcV5NcL8T8SvO0TL8ut67p
wz2HBOuKJm3mZfKVbiEye175uenfdX8WXbuJg8XyWUvdRBaVoYr/pqloaERXImgZ
+w+09nBorofixVXI2CdWe2glLI6YUm0I5+N41jdBcQqkRIgd7lzGDxoqR+A4g0fK
dVhaqNIx8gwndHVinoCHECMhHdr34rDkQUBDQfsO9p3cJXUEQ682uEkvBnwgI8U3
UhpYCbCyACx1SQ05tdIrzgLG+rPtthqoIofD+LuV6YmN4lNe0W1LZyvxAuKCP+wA
GSDtQLKQPJLLLhjCWC4kq0cX96AT1jahMhzcoIYdvOANeuFpKJZjRsvqsCTUzrpN
7zpv9KfnQ5Ma96iJSvZcjSPQgCr4oxxWT/72/kVw8gaoawVoic0N7tyznRq4+nHr
g1ahtptk9ywBG4SZgcmt+AylPN4pF6f7eF2JeJF6WjIzuvUGXctybB72l0nd8auj
H/j7vct1aUHVHzva4ABfXQ8G4FD+P+5d9Qo0U07PbpUxOARv7JluMdF1UbciKRzR
vwm6EP7Fnfe41USY+5NvxC76SrzZBq07RYnQDC9r1CqnxizDwQgFQXI8gylFEdi+
hIeRQ2qMKaeh1nhHynRCZGs0V2QaBF3vJGR905l/+oevXkHNbGjnsdh2wTgJM/fS
gTbUGHDcwDNF0VM9xwp3vWV9vEcxhp0DPd+HUZom8Fb4VbkCkZxGg5kVRY2b9Ijl
F7E/hRAuNC7Fxc7Jyc0uGZuNSCtZEAq3/ekMDMhCtHhDWAc1TH4Q7CPYRSzvk6qd
j/H0oVLRpLLBVIy7c+KGSC+XRdfwXEMOpW8MYTdtqlAZh+fuQKZ7rUG2JyL0TTMA
uxlEUzAweZs3QDRZ4XJK+9Pub4+rK74myQg0O8XVJM/5GJSjj+KN84VJkhvAzEln
rVpmz8ers1y3XQynAYuDy+z5Xf/AeyxeiSEqnmQV1eT6EVYZt11bh0T9zUC8pWo3
MQ6MM7IpG7zECPBMRTS0Ywcp02a+O58WPTzmN6Ysf0eb1OWmgUX1uylMN3Uz8QBW
XzpPzv9F5rKrym3cxP3gQms+4yO6qcytyigCJMzUXVu/KXlTNBUAI7oPg6ETwbgn
qN3dOBpjh5T6TLVQS3rETCUl/KOC0G3Z9DeNFZPbGjmWXqvW6dKw2AYbTq7TwRkk
rBtOcI1V61Xn1jfjLEL22Wehkl62qGWLUWJDwfBTSQcjM5MVHQkJ+zcUetQGBSTQ
Srebpwrv/ngCtSyQiA0sLPzLnczhDl+QbAWKSH+ChIVA4I3wPDqvX5fqQg/+irlG
42st8UJE5qWe47dKklP1bbra5XdN0aGaQB3cjcq/rEIpvmNoLDlJyCvOpJK22OWK
r3Ld4LMH3nUTIWTjh+oYxsR0d96XF4ZkB7fw9u9c5iInFDx9lwGwVLMRMWE1ytcG
7aaEhiWVtYHvQjW3Owf8KbRnwF7DJtwwgLCUBWW0w3IA204sPEYbMAjSVQc2KFoP
lYWQtjXWGEbXggSvsDImnvMD7d1/J900ZVzc4LUrNJXNXxIGz6MTNAajy0lhpOU2
IhKZzvHqWRWxTeluY2sq4jXhCkrXmF734UutIjNBrP59QeBGe+o0Rgsp3M2yleUW
mGiARju7lot1ojHM3aRuLeIsWXnWSBo0hNMxey01HcOM1JGl6RRu16/GYSgZBOsk
lHZrS1H1y3Rqh8zCI5AqAYFAMlnljMelpURWWtru9NCInJkxAHkvLCQ8dpON4OKJ
DmRnSNupOhfsCH5o0jaJwkODddC2TSHb9laLRY4wE35y2cmlmcBrUaYXuAsbQsDr
PPWsUzMnDA4E36GTCi5Cl3HKAzDSu37DtHV/+HIOoSy8Pen6o84QdBgj3EUyt2NO
F5Qeu+5x5+iCjwboabaHL+UB0UryC1TWNxCUg1L+7DrzHsIOW5zODs2BeEJd0Tx8
/6qRf7BicSXW+U4nCt5oe/4p7EtgMCovpH6WiER1Koeyg1Io2WD2xqkPLdAA3YH1
X2pn/W0+EymDA97BnaM7BGhG33dMmd2Ghh60l/6YIeeB4xsFZ8GAwFkvM2xB0Zj0
tyhEO6g++QWrls4SXuU4MGaY8vB3cnDyanjTEgIK9v7+KOylTGIul/jG1CrY8KoS
jgQubbHAbUDm95KQAoCo0dnZ/XCCrvzTSGcynnpUVdqLPPS6SsBJ5LbvR7ec+XPP
/e8UUmy2MCrVaCp2woIZLD738xQGjm43FppOijjJn2ELI2CMLL9wmWTE+xjIwy7Q
qNpV8TQoMinbJoOmmuFVvhyUcU66pLhBBoparZL/SS7ousB4OrRj8wKjOv+GodWN
cXB1W+OITS/G9a171BTmfjDDvPUN22pwuiskkpms7yzKoZEEdloRXUPPNvGymmC6
OY2UKHdwr0+gSocPSIw5a5orklYHs/K9tmH8cNbPsZnfnVNwyWNnsUnJluTN/zmR
oWLasPq7dJfpSsBRYbhXByCzMR1VaOYcsjyxztYrTytZdomot7ex2iejVlMvMKte
CTTbHSTnDNBAPzgcDaHfZsZZddQ2UNcKDS8S1IoqfvPU+vZk+T7Q2ew6UvHlS1KG
D5vgOxNEbyfUIxM+IgIlseMvxsMbq5AqHoLdf4TPIcvEWV2dSl5rWvf2LfrreFAB
Ul4HRkjtOj2fkI+RJdnHmGcAM2gpChWaNRyy4Wy2LXEXTirlpt2duQtcyppTAyVU
ueCG4gmkZ+QCW+p5Y/JiuHRA633nvrHOz2t4elgcHqXNBrZlNEIdddsD1v8Dv7n2
0WNLyDjXMceHJSKcjrMj3chLPwlM4T5WRoN4q6bfMIAi3jDjKn8vdXjcbMC+qPSK
spPevugGzUWN9ZExFw82BnUj0Ka2yKzKQGT68NdVMMM47/FQN2SzEKMut/LraC9D
VUjMvsx5upjZeLcua8Dfxq9UvasRLhB5I5C/IAcZZltdsT88iuVCtYXMxYPzzUoL
M8pNYVyIL6c4iGs1SMWUw7JfW5RItm4aDhxteMipf17dBTjG1s+IQI7UTGIpFTK0
v9P9p9vb68Mt3I6AGB17ljknTaJCNHXdV67GAe7pLaC30TuCKGZmHkIvJQjBH/Cs
MhJgPqHdNKDW+aB7guucVm3PiuPEw0Nh5ukhTl0P1vtJ/DuNEwCK2v8v1106+bbx
se/3TYdGKvVucFhWjt1LvP+bY2dz7ET2jdQFapqJkWmMJ+rwYav3s+pfDJcHGZnb
NHaww81O+AttO7HOH6ZWXPvzTC5PLEuwa22ZO+GDJg9QKo0xfdYVwujUsQC6ComA
En+UYFNQI2sWKeRHjf2kUZGernt7OIZjC4Pjs4mOECfAt2UE1ShcDRY6p/USeGNp
vUOU2VOjfjKG2xiGSu8OC3fmh3AW/1iIT/qrVMpTPp0qrIqSHhUOORVo/ZMJbDlM
EEiyZQd3RaJJb7wmManHAdVtGVormsnMEHlVVeQePkRsqR0sZI9ffk1PpdqMTVYH
xgxdeGafiTKy+HYkgjTotuCtbDOkB5fX1RTN1DKDrd0sAEHNQzonxZfwWPqB9A73
ioIt+2r9AB25OiEFp3rNBEFsVXaEy9Cp4Vjv/FYn8RBPtSB9ZwwN69yHor9h6mCy
G3Q1X6M1EUS+NmAtJjUQUF1ZxxxxnDZr/rdL3uZq1flLDFqnClEvEbKwna8uLWzf
3hISUbEw2DOFVJF5+GmPug7wXQd1EclqkGtZNDFuNLiapt5Evb9T5oHNe6NUJsQ9
93Jb1LQj5LF7B4AucBknzHk/btTLwptWTxMJ+fLndQ9CtD9tGC20URfLnJkGlIVi
fEpgvy2+vsXf8c/3+iOU7Ml5OJRDtodhlSdhe3cjbesp9HKfEIhIzHh4emK6dmee
bIr99vnWeCYbXOCCit3ZkJ/CzigeCwDBq9kUz5Fi38auuuBRJfV490zcCEWQszyC
wVcCsC+AltFYeZIH9iotHhJVglX2/HcZsFfiGGTJJO7CVU75VWmC2xw8888HPJeC
icR7plt0X8uRXX5/JLt8RK4fzWuMFmhgfiuSrp2YhK3qHo3BTJs1+PD/hGrqTjD4
9GF52jodc5mwGF7NNIQQQagYDiWxSXGgNr756pEeCZt9a8C8m9zzVmHqGLa6Cmpg
/wKdWBG1m1KSApPlVZOzEcUWaw78+fRl4Tlldjq/LuThGwMaHGq5blwBwjtUIx/3
OJG4ExbZUSMRXjmMXoJ7u9ZId2cGBG98FQRsUF00zHfPJBw4e8hQL8B/2Fu5Kx/z
ylTK6I+GN33eOGA49iheq8nLQIPUix+C+lv/P2ImF8kVitsMavrAbItF4Ktbs204
o8LR3yaC3yYFKzVaIe7iY5g+QYmqM8StfwCkA2piWWvQRZzB/CrL+ER55eCPq8XC
3RtnQSwLUkeqWF56ozL/PZhCNHyk6jihEe+sOqv2Z+Ea64q4AGerkTUhoxO5dtil
RFWBO4cf6PoiEH1ZVl2gjq7e0c9+PgnJorI2Dz7sATvObolED9huzksY1yETJc1u
Px6f9+SOIAeg8aV7g6ODRwO+wGsBcU6hEcrpv3/iCjzPV7xMrBViTQadMYVS21pW
2qXrB7q9Ck2cdUPc6zyEptIjgOkqIYBJn1rbfUFeHpNEY0SIu2vY9KXD8qn68rxM
Guy9UxgIIO1DrrvsQeLbwyV/+GqSln3VnkmdViS4y1QXSrK/8CiaiZMSZeGeLQU6
/cMMxLa4nTKsJdFz23Cw8XLdtyvNNXiz2bygQKAIpM+XCDUm66QeREpG1svNADtw
5KgKsY60ptyJZqzUkggKegC1X+vuafKlO+aTfqmh6k1LSr0wkhTXVks4ZifqJkns
ak9D0lFkQrq4LZWNJHDpHlQj1S7nNJWz444qNdjIoyyRY7QLayl2xTuwmeqiiFc9
5gZoXtvNbpZO96LvvUNOL+W2boOu9+HR41hmJ+NEYvIFYpYXbBERDr761dt8OgKL
deQVwjQ3i9gTFPbiZMuX/uOYFaCCFvnaN/gEIMo9g4yH+zOKpzVKt4KmYwIqN3If
BuGvJ+4lYrMi5xQbuoXtfJRdlYuzh/IJPVSp4NTdEJKN+rFLmkdMw0Ri02tFRafQ
A9mThFxGiFQLz6VnXwmrOVyZt2op9IJDrgRnEl294nruK+De3Lzd/eRKvYUkExvW
4IGq9HD/Be9uxZJUT3HuLjlrdxGAJoiql9c2kBzmSeh0l5ObUw0NW7HKGamyB2aB
ASuIA8llk1C5bg27GvWvboOjWUX6Jt7+P+fPlqi/jJw2TedecAOF7IU9bYw3zoMg
85t9acePxdzwi8Ini2FQEURXmBnUvvqgcj03ASWyijZmjcOD3Eve+JHy9B8g5M0D
zuMjk//x4W1e4eLPmJBf2WCE0ifpUIR3TdivdmPMtSUskVZKYtXqn6XAPiDCLuMM
XzvjpOtru6zmZ9KqN5JAd9eG5mU/Q/A0+iaR+TGHNGTtWk6tmOELNcQrcrIE/zrC
OvmuQ/JWNEza/FwIUEah8oNvf6ebukarkcjoh/VWfjRm1udjVjOKfK6qzAPV5Wd5
wRSdaTmGK7b1ZMNRTh0GSZWT+ZGe+ZEe0X+7f9W9LKH5s8RneXNT5kT/uh7bnlmH
UDOD/m5NTgfoudFCxdVkWfnYD4ow8HXMQx//cVQQS2TUOQvsaxfHQM4vnK5tdjeC
1zRRxEJhEHErNIPPZltQ1w0nZUe36wjswiQJHR5qqQJsraLD0QVWisa4SNxkIOLA
mz21wUUH/KbPJ8Av0xSBK4scS2GvbCEkclXSivxiDMsUbckSZKvd9EtWTAwNCX1P
Q1n4I2xmdRi3gT8J0tHKLqV3ZODjPiK0IgFEVfkex7RRut2PTG3k8y/Oq9l1lO5k
8SwY4lIYoG7k4FNYIsMNjUu8jpMuZUxk2Qfka/oqNoBMvMO2wF2bMxh57SKMYz1+
DW6lQqsEwc7uEWd08vY4x2nnjtSbijkLOLGVETLKosspSu4UVLxkC4F37qUJ5DT9
pque4sgP24lbIr96LjKE3jKXR4wYbuMRvu+6NyJt87P4jcwfWt/eL9PPFMxXk0ip
fjW2/eYZQuAh0chuVzfFeyU4kEpzXjs1r2Sj+gTl6i4QdIx+jza2bZHTc02qUGGy
Ed2NBD2h3w9LGQcm1SBpmwj/U93r/nTY41B26r6Hlb4o3P319R/0HLN2wUyJYn+2
k3KsjKYEKHNWV82XfyEqvBQIIV9IQ+whINe6lV+pP0uToq3DqQJZrMA1Pfdkl6xi
oQSSdxEoTGoMJ2mdWeK563TJU1cUFfg3P/rvKJ7Kgs2VbP/+Fe/6TRbVLJVplSdI
PXCyxK/VvySvl1V5hdSMsaFb5uwpYXzmVRc6Rab95SgjgGkW4nMIoJcQTxrh6oUZ
oTlrM12SGHPI7K/3srKUc17jWy/ORbf3sUfkiTKy2MZ/EzwQK9nrvGW6t2fqEN54
/Hk2Z9zGgHY9sB7ZXHkWbm71sQxrBc80tXskEX0Ai/JWf35Km1e63EDDyT8LisRk
O/CToCtACYsVaF3h2RdZJq6HJfj06+4+Vi//ZZeF75KlWWD3jG8r6wyrDeI4n11W
qfgQwSvGtqIkAiEekeqfd1NTG7SJNRGmQYDycXmIspJ01gVWwHGi26VehYxTBpqk
TDsw6bcg92uOH7DBxwlsAy7uzbf7ixK4S1AQjSwskYto1GwaitRV5yVHnUBoLc8P
ATweqrGTsmn/KAnU1nbULyJ5uHZ9NtfGrKl6zsjKzenIQrn5zbyLHQQNi9jqRfE+
app/MqcCBCAaLhL62ZfdLwcUr7xwfD1F3WoO9Xw4Ixxer+fJqnZckDGo960revYz
ir5SWplKCuYZqqiqe0xAuUoguHbI2sreoINglBbNFdlCjy7DHXVbRdbHGpcH9oXU
4IUW558nBNElsNVZpatt8GftzpzlqiXdKtr0ZcEwTj3WQ5eTXYgy8ONekNaCL7Tm
TlEHWFUVLN9ER6+I64jfnuvGJCJSTaIa51fFrE+tJXHeiZFJSCUpKRmhQsubsF2U
diORq2A2BPsw2B+fr/B/axR4T8u3xLwzcHL5eUlVoYytM3d3b7y5sc5NDNZBWhJM
46qkw3mgTJOFbrn/yZZ8b5cdYAJXn4omlAs9N4X0s9DSI7o3C2/ZeYsPl1CMlkwz
TN0KhI+ePxZwxqxdU0qcahxeXtuoohJROXwHORQXtqXOsCf9WXSU5c5G4+CYUudJ
bbSGxu1MsY3Ti6PQTb1wg1XxMamFsCcPLe9D+GF/pjw6nxSIK+0KcfDY135d0cad
gBDGqgQwXg3tHC0tJTOTFbP+/M2dpi4ErsXRgn8U9p3UBAGm+992vB2tzwiBIy6W
cLK6N9sh1s0dyyCRrlQciro7I+2YH0xr2WFxdhiztbCkSoK/5OzZYLg9JWX6L53k
cfzrB8tQW2euo2rJ8Y28NQBqwy0UC/BM3QBXQX7wObzl+70ROofviw4VtsQX/jMg
/9MRbm6o+kZQfGYIMOEBtdCUbaxIC3C40FkGeLlY+OiAV5Kzbhc1dDtq7s5rXQcF
+Kdqiqaof3M18ODLp6Q9q2PW8ti2MzNZl0rTMHbF0z4Ixv9sJDXC2KWUmIICN+H4
+TGkoCM718XnxZexKc2yvj2H1uYX5xW2umt/rLkSeY7R4O4LgoV1ZPVgsMaEtzjm
40703X2CAlc9ky5LIkVVHB5NPqTJ6eMiDpv21csExeugP3wxRHhR2bj8o3Ev06QG
EvXHt90YEyy4fAti1zACtLpEj2zCVgB3JZvcsqJjJl3T0WslTaIU193KMIH0sgq8
9h9EI6sWyioI1icAiE1lmwaFMZyGNhfSMr74khb71M4TvhBJTkGhlZcAP7EQJ1Hb
qhE85kA+vJibsYr+mj9Fdr4+FhPMJTLwarqh19Muo7tIQgkZKPKewySQzhFJfCxo
cnRS6qfgcz4xihqfBZMsb8lx1ZV/HBiSid2v5u8QzTQITeni21c+ZBrKCQ8tbMIG
yxQPqtTexyGpmcANyyqy+4kDDGHTWwKgvle8/OZmALgyWtQvRJy3qYiMm/zrI05/
0YSIPYFGisoOS1GjLq67zvzAep30bwcbN4+wzg7nry6ZxUV0BD95DDlJZidwoK5p
UqoH8ipY/U8D0wvz1OpBUE5l/LguCtZM+ZBE23vED35ilADwmr5cAII3iTYEyEka
tXyTGY9LCcWTCdx+a3lUv1ZMmr70KolaUxr3xvW5kTeWVuPI2KDulxnoBf2ILubS
6+ApuiZUAIgFcVCWx2GvCV3fpb2eLL/C57Ab+zPXy00yeB58v9m00K1GBmfRL4Xf
jk2RK3SS7bCnlWFifDqWf0lIRNpArNWGGKzjT45byI56GYxjTYSmt2tmnGEbtWzn
8dXhqxDeG9A59Ky5ZGpOhIORBU7d+Ua5KFxZyQmFxFLlDudeLqx3wFhGg0pBNtKR
FJU6MdOgNuP/xPrO5bJ4sfcDFTApbCDmvWq3NH+gB/fdvOm66mLMZJ+ARucJ4bY6
kT9puMNpCf/y23zn8AQi/XDgKRs2fc5im48HQq53CUY8RIEozZN6o2+mPwYd+fIB
EVRIe+5uJQ85i0Q5k25md099fMk11UvxViGvB3LJB1tIXQGvxsRv2djBYusIlNl+
0mHlZvXzFBu04qSsU3Z1lazLABqZrCWj4m9J1BvIppN+LtbmJA5JBiovDEVulxkK
K50upPhK1lS+ROCK+cRz69vBMFcLRSX7iM7YvtBuu4DipxJx7+7dhMZn5mVYhp5k
NMKb1AgcwUo3uk8HjMmb6BbC3KFc0Fy1S2e7wtiUPf1v0MiCaJSEChSqJCGW1lbE
FJ9rEWusL6apDJmVfwmUUjcEaapFH2j8+O48Z6iDQcmFU5pSrB3QulJZJl+lN4AI
vH/3IBGbfs2CMjAhMJwzJa31K+nxdKAbttP+pll4wBiQpc2PlUodnDyLY/emQh6T
CCWjIvkUyDpLo8EgXNdgViqO1TPLlsrmpBtkR9hy3st0N74ODCuvrjRTdLa1kvFe
YWWSWpuuNIyl12o86MuEKBCPn3YtEPLtIoalREXLKKDDTC8Do/n3buCv2iBC9/xL
S5rtiaUV7tbL3fDaLT8Hqvmy0UqqKfARcoTrEE5n71zZEHRmKKoURbHRsugMPe5S
anny1MmhJk9llFP6+MM+M/BpZRfiuC7iE3dHwhK1NrgFjGc0k+gBfn8Nw5hmJXZ9
ikmvd6MfHNvwCTj9/J3N3ZcU1m57rM7D9mkWgOSVyijejKZzKdRw7r+s7yP5F9ia
w4SDnkhZrLpurvRh80wbCxrNhJwQMTaYeg1sl9EOQq5DGauH3u9/tOLPPrTsnbhr
lyA9ds3SztcaOhtyDgFNgLn0orB6nJBf29vjV5wN+75Q2aqGPac9aUwB3/5XCbWa
QDuGaJBwp+zo74E17ElrgjaJ59T7xJupms+lOR8LWbEp5EIcSH3z6pniC68189uY
6bzioqaU6eh9+Fry4Ndg8CKnegAUUHmhOtvubfxq8/g/oRsxg2WRB9P+KNXT4SC6
ymIK1SvDd2/E1CYEbvdBoXzVdsUYCDH5xX3UoLAUgiV63efSfy4Qz7HbwsJwDQMj
HvAMU8ga3ZImY24bAwAUb+xNcr0C8hktsL650C9jPsiem9bZ5Rfz1nUUagO9k5fp
5yKfTbw+bl4DJ0B60n0lxIibd2D6I1kiUWEXJsTLae8zNYNpiTJ/UTpgbxQ/Eo/t
1ZdoDzHutNQDl872PYZuog9S/DdSdhD9LVlueh9BHFLv1rig9NskHyNd1Jq6EV/w
enC+Aet/X4dsBLlFHro50MFfvkJgO7YNOF5QfJVlji67U1s/eiONOf2bJ4PpzU1C
z7i6ZVKSj5GZQq6h8iu5qKaB1MbYFEoDEPW51gTA31xAfWMdhu1Xz844OXvjRt3f
hgd1ZF3jRU1z3QIfQIzehp/aG3TmSaLJzNJJpeBl9aofa6mxvkFtIDp4RukE5ArI
wdj2CsCH9sqkaozMqnmVg7oAlf8w+eGwkhc1XIRygUyQ0P7KT4xUq4xtr7p2R5oW
0hkl9MybXdVfnzgppNLuTdLIUI86TRGXrKlU/+kmwvXLYrsG6crLE9hOCMPjnaxt
156JVD5A8NkSQ6WC1430yOV9eq4FNIS6wpXUniU3jyLs5z6NxnJXYqIUqzcv+1ZO
5fRpSpnNhViyL5FN9t/7OfuMSiQXWdAE+rikWeSmef+v7IETn3N49/3FsPPzKLpE
S2akBBHwlVxABwRh/IJy8JjXYOTIRgD3+vaxAO9T6ggm7ySTfTz4WdOwMkeS/pMN
hnkD0bSJsm1tCZXAsf407X9bVjCGOi2BcYPgvJMQYuEL72mlCFFazbOpMvPJpiIl
5IaYLhmNp6BgYGSEms0uPpYg0ighIOmrmJcth90Bu/jh4soLMEFA5PKt5CAtFkDI
C+wSD2flX3U6qsN9EJxAXoT43WMe0NcfF9IiTtAeSgPjaJHcp818sfNCnjCb7CL7
ySMEMUfH8fwQIZNIvYOtpVwJIMInr1utEzQ3ownxojZtC5I2Zlb0TuPgbj9ZaCV9
T0q15mGCd8bK0OUiLTnC8P7gnEozf1XiZAHLuR/pvfgo977RfWdRNXNByhqh5axW
a/UbvFqNjIU27vQ86XJFSV3blJ3cY7YFS0IgEEF+poVMuuaXKMYSC7U7KOMpLsC0
S89opT6zFfmJggdqq3O22KhUFBYvdbm2qH4InEAIcmIvCDkWkLw/077Ox6VGo9MV
zLTpxOGP4vfGdcX40FRzsTg8v0ij4CAJCkslLzQp923s7UXPCEFAZYikfhoh86tO
Yq3WtNPLOPERNo2Qi95zsiAoQ9eIX03MiBzI9IRahwc0cWS2vBxXGtsH++mTvk7G
JRiax5XC6uHzmuBnsRup38L1ST+ErU8kfu6vI+1CLqYgRA1xo3h1KSp8Jzp/39pa
rzJ6YN2ZOVdt4JNgx2uZRi+JWgxaDWdlT348KqyoJP+zWa9Uri8d1fGxHuMPnQeG
q2wrE3M58hvyWC41LXc02Q60OiuXYQLJf2XFe2sG1x5NNJYfiyVmlfwhyhP+7Zqf
r+fGRvz1mgFTReH5iNqoID47m31Tk+/p5gJ/Asp9V8dNcWjvHLu+KS81YcGrfG2U
zOMhJgZC3PamY+gH8sWDFPnPTQ92WCi2Z6N0L/u3Kd9sbjpEHrYS2jU2Pfwyg0rZ
1Jlp0PCqRdflTBtWHZW1Ai3+amzhGvtlGJxd52c1HizoA2khWx/29pWuplvYBu4c
baSp+gjViqBIONVWSJ5QDltndKkUIDIVt0x2wjNgJ3DmiGF/GSR4VODf+WSbty1l
QAWZmb91S7BCZbIfVBunLtnc0m2RJ6+VMXFZckjB7/rl2FwY5kvSxq06IJoZOeFE
XNI+Zy/YGodyKG09Gb51ICd9DXt2GvZy2gRb01jDwuauNL/NwHQGgRSQcl3jJ3P+
LdfkHkSta6riTEtpJ3MSpYBi0wAUBvTBoFtPkp+LcIyKWRIY1zd+O8KwIvpL6C4v
tfZH4AwUspj0tiglApug0RpWcbe4u2b0SggNuhHdXANdCP5WefEyzFsbvZwN6TKQ
NVqRkXzS2EqzFEL5YoMakmjKEC9YwSivba2O7TjoooP8NBI/7eTksge3Y0GVMpTu
7rs1U9/se+FvlXo1Jcy5SwqCmGpxEwcXJ4trRJ98fM8XyiXLchbf85xSJ1+H6U7+
NGxDLox+9wAf7uRQgyQjeb4vbLRUT3Bu5SmXHeMJv5x5fBypE4x4CFfBTzDLk7Ag
12NelPUXMsDV9vTWZlJYiWVEmTjig1tM+CJD5rk1HO+prc13xsk+Knhp5kmX2WkH
bUY9I+RRdLKXGO8ZkH2syRvfryE806m9OI6WFTWtcIu211Zr0VwIylhf7YbJSHJv
C/v0BKfqpmugmKFUKl4dkrEIXGy+ZgnUAwkP2c3dUsfq5NR2uHYolm5Fn2QnNfbf
M7j4DgANwEChseX7kyyo1pv+kzYLuZpBYiHq2xe3gEByA9Roi4hSl36b4D6EEBia
hI3BAax4TXwBnchouPxzIJqNQeU0DDQNK9G0e4wa4DOJpMhQBFy2Y/hABEHlIPrk
dHuOL8n5jrglZ2eQkm9RZ+2n468zQ0AC5KtKhlQQN7llUhL6OjQM4yonJKoVJ0Wq
OfTKouHV9ZpYVeqQJ3G0Lua/0RgQfbUynqlqSBWDbMW0dp6Wed8HUJAqNSPhH9IB
Wo6qRn7Z0cdn/QotCW15aWOXk0wo2YFNsRDZ9MOaqIhPhHb6xq6/o73oyU9zr8He
S9227pqcrE2+tAIy4MoBagGcWteS9pvs4xTgi9NErlxjYLkj6kbCNRq2HEPoECI4
cJ9NBSML9jOjEkaOdtxJrk1MRmSarhO2NFNo+j38asTTbmhczibz78RA34epoVR2
U/PTvZfMkCfYDz4qUgqI9bB9f4fNvE6/y9/pyPqHb0DJD8SJ4JUK1ID0+mugsPqP
qTL2MR0Y3yw8EdaQQmE8OQ48kxKeXMZZG3pi9ysGZtDcU7vPRjgbTfXd1ZcOVKUT
rQPhDL59NGnaH3geJPAc3p0tWiZgetbcoSvSrsnABMIs+ndbMoCadujgPBTm3knp
zMZF2p5tLGbycKZBxUaYsecJtNtk+pDTEY6cJydF6K3e2K59z0tkUOXNKXv+RZwc
CE8NwhWjsrg9yo0lhP78b6q5oKXr4Cb1W6yij07szRv2ovYzZWfjRt60RhAs/y2g
1/t90RBTIc6lfgCZR8LmRLZxYrlWOadJsZ+AOygJbhNxMq9tuaiPfKTm8BPnZAc7
1+le+cbwyqTQuOaGO/c8bu+H8jk/hez97d9sexjd5MAkoU9eTbtDuW/w/xQuY9NG
4Cj4qRkudeX/H7/igow+xLrc3QhmB4d83UvdA+MIJg9ynYXkMzqdJC+ZGFeAwiO1
LEBDOh5KPgNd42BW6/dAvDRMSGDuDnFI/T/ZxShdaV6/FLdQRho7+vwEw5Cp2Hj4
lKS5+hjyw885mJnlOCCZuyrM5L0fSYP0bKa6hm/sSZucXkV8gqNiP3g4hbnS7VuC
4UhjES0ESIuEKz0WwX1kllEKzL5GMwD50++6S/nARXD1aIj2iS0/a4lozjxBIbqU
j5+9PK0613FPug1tr/x+xl1ucCqE2gw3+0gCmb/RUjLyDjIPp9VzW/h0E+gTV56Z
J+Wa3Cm+LvqHll6MoePnXq9SCNsDQTwVlKCFppq3K4lwLs9rgZssIoxSxONtV9yJ
qD4xx5uAXM7kGJSpVmmjT9X1SdWoT89KDRXbHOJykWp0H8slZUVcCvZMRjzkz5D+
hkDrllwRdjCy3kDNp4G20MV6n8mMrbtc9ALpZxA83+9DBUllZMQM6ml+TaB+2P5o
kf7lkWdvaN1hjcz8uW70MovdMIR+TZtVufFn/5JgZdsJcO1EJ5Is3BFbZxFusNg/
8+ONOJVKv19LWwvU7iJ3v7QaTe6n1aJX3PTnAvGJ2NXiN+9n3UuM0/wkbUQbxmrw
2V/WUsBkr8hR54Crqv15DHMiJTwmD9eIvdRofUryk4Bht+vhE9yUJ99Z+bl+IsmQ
Bx0GbIHYCsFXWgsu8zUqjvZodplAR0Inv7zmPXf7dKHg2kS7Swrt3VBg2e8As9cO
AyFFTYBnWEzChbCvFrLf5HpIW0y4/buQSRiUaCSzKHHwzlKfOySsbDtzEsln27Rf
dSKnOibF6+SAia08A49BuTwdidMPFrkMi28GGuQBZ2bStAilX9dHNDWvR4k6u7eZ
jYH4NCT498RdW6A4O7weaqWJkTM6aSu5voy1vwNLDa9BqySO3IUCCcVMpaam6JTO
DwfkRNTU0JvM3dHL5hQ4Q90XxlsIPhq1OOM18EnTKb2596TevZj6a0kR+YPC1YeU
7iCwlaCadi6xyfNillpRWzAs63w/kY1XfU+xCbvehM2QnJpjf9vMm+qm67mx9gTC
yakgMnMYKGUNkunLdOvDqmkWhwepYOiUO/fTorHGe3RNDZnMPm7pIZVlC+g+gRUA
8Jr+wDlvTvryDgGd2/+HSlX24FYlEFSrEzw7wZmMEU1E5HoTCskygEJvL3ucF25r
f/PRCb167bJMqnQZrYWqFY6ViinJZqCEKkGdOCGFYc0dxCw8LCgrXBKRmk0aI86/
1lC1R1eogK8BjaPNBmUokHcvgtGvWXBgeCVw9DR3JbRGWSSngp5rPWylJZUoBp1H
KoVkI7rrJy16alXFnYHJOLtoO3iumIXYsGePc2iZNhsMC33pdTl7wcrT86/T3G1O
J6er9Tr8nHu5KQKRvgaTqwPQS/hevNvfuXr/MPXWv5/QIpBOfQbAoaBSj3LOON/N
9TZ73I7xTGvNwSMOtSUee5bkfVD8aahlL6ybheKy7FlM7C7uFOZq93cIQw9vJ7ir
E5IOotf7Qw0M6M41TjB36JIABom3mkZiUpfGKGpNhZZLCJ/ybToYFBkj9FYNNB/0
MWgawhuhr5szZQDRuv2Recl/BZhYEtwwot3sNv0t7MS2ZrJ8n5ZLVnSD52jzWzrh
hiVL3TCiqz7PPtZlJFM/M6YIRCphuqrX9h4CYMRRzPir//R+PdnQEdVJHuYdPnJN
cvk41OV8BXXrzGAkeCj1O50RTs8NF/u0yLXe7BhtDg/SVRDCc+kSdUwRVJMXwHei
lRw6VojJeTIvGhfgzdQS4EO+ecoxf06NYa0za6lGqpzonQ77Ql2mzikdHAp+DeMh
lcwit8dJ/24f+gijjjkRtpIZWlTsTRwVPOQXkTQYTO+/GyniOoGMFnmnKtBKTbFG
/rd4L8aW9sVWpQGxxggNImmU45SMtvYaL70Xw9iEAn3wBig7BES882YpPPd9kN4O
D26Q1qvuBsUjsWkv9glHAKwTCJUFnIHZlx7mswXUf5GRbTA4AgXk4yncv2ha8R72
7qAY0n83GGb11MM5a+h7kNXhSBigforpDmkGIwJqHvLAsHL5t7yHJzRZ/Yr0BlQN
rn2HxgI2Sablb+KzOPwJ2kisORi7dV9I7AZLz+8BvrevDOfx/4Uwm0rpcPMQPV44
apkAEuaUfAf/Usa/n/cGojuu1FO+a1GWTAekhNAyVzZjzfnl1HPemSIqYgASgrV3
M5uAjizp0Zm5g04gJHkfsD3ZWql8jUQkfp9sSHDhOcOJ52zRzwJIxIFRobGdd8Tp
UxCU2fY97KWxf0cVWzS/WVWJ8++wS2r3ZG5ioT2zc+1I0bdcmD0mAEfLTBDrDr/z
Dn2FogXodlarRnNOOlZ0aIKXvDMtj+eKYOS8RT+PWMEwZdO8TpfIu/4CXK23z1to
MnqreZkUGRHDkz3leN0zH1Ltx1/yfkEF1rVNWu/gpB68LxSW+55X4Z2QaNZWqsk8
3yEzqn5GLQO1ffIvZdO8IZyAg/Ir4AxcFe4k2UOKkSwVXphYY7E0ixhjfaYJ2+Jp
Ns7W7820XWHUx4nnqFlGEoP+mlj9erZAac1I92VCGvdULsY/zaktqOk72g0e74Pm
ZUYyDx0eWkf8QaOJ6FdtbyJodh8AvhRVQScyhnsOHvGtMusnPp6dW/h1B8KJMLlK
JfyuOkP9GV+xF72uPxquVDDpdm3+NkfwomlD2z1NlyNM4KGCUAA+jnoVrDynDMCL
D/jzqzEslb8F3wcDWhd9mQpmsqGQcxJJ+V3dLBVPMNK4w0bNLUbYmwyitbQ+FUR3
ORI0XIR48Zb/vwzn3NIsQSfJ+h1msdqbPa51xBOjRABPfMwj6T+Yfl3zBXjd4WNr
JZhw4fG+sVuILted46FN1F3yg0Hylqzr1fAZdo6Ylv8iFzf9pmtikModGHkb9Nyf
dJV7PxGg7qG8z7Fe0RL/56CTYzxaX0Jn8VLqahA22IeVLkCwZaA/7DrVCKsRSx5I
4xcbEJCpJU6IhIAgtuj4IQ3LdE+0JLezUcHSq53OIEB/ZEQZ0aJpg2OzTM4Qx5J3
VLR41EfZO7Q3s4C2tZxv2pSoZqKZCNUPgDj8MpYtoCmxzwBBly18lbBhHgqiynAM
43xkctZnSjNkJJNPiJ085DW/V1/1C8byJ3r6fo2POt3wxddF7J6Dl4Hbi8BHVX0u
U+9/eqb8qvJf+o2Ry4Y8GbUprLiJBApdfVnoWxbZyMVNIT+9IdxJM/Zj+Q0EsOD3
BOwIKxtJ05Posb4oltq2Siy4A9h+aPXTQMSy1CkFDmUjya0V3qZhSUT/AYWHnnga
7sxOIOzyWTp/sSoenz+4PH6knDBUrdR/bh8f18uP6RcxncZcU6/OBTjCoGfJEM75
KuEtvaoCtR3G0aCP9aEuhvMJ9YGeRwCx9PO8DhkK+MyiXfCXyryX0hzxYg+DqwMS
1pq/Kp0/w5Pf8y5nrJNk5SaVCgHr/YPSNGYqNh3GqdzsgEq3c1rBDlkrhbN6K0W0
j2rbHvTA7/gbBuc4opdd9omRChXLCd84m3can4xqcgmLRur5avBErvUN5zH6zqPe
C8BUtGpWbWaaJ9tT9kxJKsoHvm6fkr43JVSxF8qkZJwdHbnckunCmbY4/DZyx4px
OukemVOO/5koBsV1ggL+wa2ZXjTAGmIVT+tT6f6YBGWx8sH1bfihMVT8KZvxNJH2
lgWYBytCu/QVdVqoG1LF/Sb8Bjs276agdwSMkpac21z3hOADgb6NSfS2BdhqmIjr
L/P5pT/B9WWWprrQSru29A/8R1DpiT8sW0oFglY74VvsdXXn7Cegj07uyGQA08vi
daKk5v0DYgZ/Fb0TVCdTIBrhqurSrlW5CW4rB+8hAIMNOkUfsaSzZGnS5lQ3dpZu
FcTn4kGsjysCp4nROYaB8c1heORb26qTLd83Xn7b+2XVmkYVjtvt+szE+jXMLKbo
s3/ae7svtWdrIO9uj3cliSN1UUL8FilbI6VQniGbNvgR9SZl2jeomSG8Uq7sO4NY
LwwQ0DGGlrcT8U+jSJY0oucOdN3LUHDnd8S/10tqK3aG3HqxPW6zmCmCHRGf6jXU
DtPlBmw+X/hEDOhhLd3VVB+IRFhPowboK9NHdt5OyulRR/BVNKrb6D3H4rt/CxBS
e8ZwPUbgkeTFkvS8vYZkvfqngd4Al3Ec9kA2eeFDkx99jP+ZKuZAFc5ApXsLwmnd
Ov5Wz2LMrvgncgN/86ykbfgeF0Hc4SSDg3xXwxbXApD79saKLGEeYUsXQbRCyJ8u
mzmxfxQr6a/0egmeujbfvOuLcC0a1/o+2rnXOi9dvAuOyNkBIzmRtx6s3EpMj7RA
qsqVKnSOj8xb+JVAEMqOp/E5G1sQQ//A1tTnLWq8tTW3XJsEqPBCac254x/DI1bc
qp2t5n5jzz7jtrFvKNggsg1EtW3/jbpR8Vew8rM/rVz7GnSxZmWY7P5fmd76jyQM
xYauYqGXCMCw9iouPx4KURlta3x6H0ARsyhfTMStBcIRlu2xcopHgyp53p4xgv8q
6bwAPDV8y2iAXg3XGZ/uFiprjutSm1MXeiWGzN93GnYUKi/Y32FwBSzm6Shl84YN
EP9TVyHvef4gS807tiHB+b2ntJWI9+VeOxUP9pzl/GlO/zyaedwMSK2luxkH5M1w
z6l5IPUKLJiqx36qfVm8qT30ciBe5yzf1G5qMkljYXSEpxYFRwCehEOeJlUWLbMr
Gd+2xterqwZ/AfBpHAfLUQr/O9revVv6+HzifR8Kq41+hkh9ZEg7GZhl1JU/I4On
V1nSPDh3BxPvfkoKv+wiUWlRuRntFJsmPeJsgtEI/KKu4yeL5hUfExYfTT9hLDHj
LiIp4gWOLUOtkz2deDsae5DRXfb+p5fzdIbzRxiPqbJtVG3/zzy62OxJsZwOGg6q
DbUxMo/o2iYGiQ5GHme3FJrlYer4A2WIZcsS1ByGIbV3sLStqbFBsmfNOw3LwYL/
1vGSGhQuIEPgutlcrF9JJqJwbYypdOKgohcVHC1YR/KK7mvJWTZ2FpQhwVqDVvrR
Ws8ea/+u81ky5VsRU5wwEEmbqAM0u6LWBQ/14xucaziD9qDC/9ipWFbqtYSbh9Dm
q4npX6bzrhv0wnI8fE+1+cvj+H+wLwJAYoPRTYuOig41gIR+RXiSkvB+sitkLcZ+
xLkqApO/cW4M/3+LHgJHocEOfJIlJQHZQpmRiX7WteKdn1L3vmisVwa7wVTv5jtu
FpZOP+Y7iTc7Gd5YmmEOStzCa1SAwqVACpmZWeFhJdE+h6s+8ynhq4aZyxLnKLqA
l14xomHMSyBAgehKoc99AWd9A06MBUTp0P711jjyRikPycl+pw3PchQkfamaIURT
ON0kGLoP18wyMmyrjJcDKQsZyfTKXugcpGygkK7sVwxRTJUN1RGbLerCJ1MQkNZe
HyOOa1Hz7J2eprG6GdXk/P4pe49IO2A+uLvBjl/MIRHC4jbr4DtMIUjvne/APBa4
r2NE2nrz13o/Qf97IbYBvtHIOcnUH1krsIVKdDyCXlDUAiUgZI00WMnQkEANCdIJ
kzV9rEbUV+L5mFOa5iU3kPcM0INGGPeSERnyPxSZ/b5nCWozpvQS+40Dsq/dF7yp
pcU78gGZqxCMTobb4+7yB27XPrVAUXSUA4MxKm9aR6avBLigTGFl30/S3yd65hlS
DcOVo+GMyAqI7jDAmRjmank9OP+KTqzzolpbf03synjEaLMuStbIc0X5W/jAmOFb
ge1Setps6Z6E9RCgoPNsbuwCYZ93U3dyvuwAcK82v6yUmYUYZ/PITXyBUDHeeKNf
DmdMTnSVgpxGUvhzsmuDisq2E7JhJ8IOQNV0q7NDONwAZhIgpIN+ZtoeWEy+UUWt
T3boBuiQRizmDCCTLOc32Qwx0en4XeLqrbsUKT5gtwLhPRmUbNWLZeD2OZJEfv16
Kz0OnxlKLMX06vgO6iM62X+Pao9ShFuBftlE5wGnxm18EkIRC84RRDBvk6IXdg+B
UId0dOb6w7GE9osXo7Ig9HjbfCTamYzfQM0CgRrK7OizsJTS30L3ExIICimZAFnr
ikfurbKFpHksAMTuhqbYYgoK0sNCy5P8V2qsBUnE92PO+8IlBudPV4WLOW8t/V2B
wDpnzZbINIZx4fwH7ibaibmQeStttunjVaDN6Sry1PZtBOPabftb5vr1ir3C1JwK
QNidfi6eIaCb/StDU9ZN2TUZs38uZvQunM8X9pQMQwAXLYlOgxmG6Pya1tVstnjw
nWOKozCCkK4mWNuX8rxlCeiqjZigOucYqVzGvFp+QqN48sYE5YWz+JY/jB1nAbL6
pzMve+ufFbDfaBeyHPpFgMbygfWZuTxOk4u9eu1V7+OrYJIo/HhoL70lMf9FaVPd
66I54yj2cA2dT/XPIvki+GgFCeEk8523qwzeQ/EZukjqP3bb5CyE5XP6+QOmHLi/
FhMAjNlKSut7wyhJFyaZod7phiKcO4r8pHJAClq9LgTwM5TWq3hC7WQa3kAOddzw
kI0AShmL2aACVHcWK8Re5bEIACtcfabBiE3POHvupqPjBVGn98lpJYmpInKQ7ir7
JzM5jrcBW4FSfF36wGmMXhlLWnnn8msMXTlb5XrA56VYvtZRdNlx/jPcMTcnwgjR
9ciqG3FZFX0q+qGcUQi8UpLvFw1RowYy3YpPr3CF8dBSK+amGbtak350wBq6E6D9
i2GFNJun3ict/NuX4+Y5xR+4TpVDjktWULhq+GI5WWmxVnjYUo04JhqE7TAN+qkg
O6nM6dze9gw5qyBac97l0WYStNFErRWL3Gncsu3ExBOFk0Gch8PdpeEsWjgrXuMh
Q0oBCUlplxUJ5cb8ua1CYJLH28wFOxJ1RvtH6v7xMbMIZM0cHxMi/5joyJjixR6Q
Vh+afZ9XimavoGwCBcM29JQ0novPrddaNcURQPntDHeVkFPrSUr7M2E8fBqZ/9vS
oTw/8fHwM7t9FGynLRgHOsJR56O0axwJ85Nfu5DUb/iq+VnXlVZ/Jt3lrx7q5p7g
LQC074qDjlY7ksM6WLCEhwXgpJ/Sxw8WBcS4IkeVDwEberqnSkeAUrtXK6dR+yOz
44oeZwBRuvbrhk3XApCaUhYPWCAUcce53QzO4UwfNJzmCN6IbcRXxHwPYUYkpuzJ
R7nSt4qgvQKlMQMu4ULDsQ5/cqs4aRRndzsStznNR1qFZXeKIDDmoIbAbgZzys0K
+R7kP6aYUxTXRDhJvzNec6bGCkodZeMG4DrSrLxZhbKFPhJjw8FIBx1HU0iOSa8I
7Jhk1st7jgNVKSq6sx4pZq517bjPOa15jjxQM/AsarleHhIP+DSDaS9zWJ/b5IdS
8QGvkSG+7ud79cIGlwI3vOgYZa/WE8c/BAVtEtvnkdruU+68o01tUspdbZ/s4Zz/
zQsxJyUJKi0iYxRBG+CMNno4k64UlXqHTwOlGX8H7REz8sV4qJiKZqdbaPDiBMTo
Hwq3gjHHJsXg2h3SqiE0HcV8CSN2Wn0nCY8Q7dEpQcvokoPtpRtcptUv64DtCRad
QH/ptUtu3pRTm2RiSvfDgLvfbo2cmPHZ+/PuE+qg+pR5shjSNN5wr3pguYoZI8B2
Dj7HuBcFE29cB3k+M0TPY22HbEhKoiDIQ3l9K3OxB+KPEDHDyYxLG/K6tc/LGfrn
w1s1cFd6+XNLWKQI1Jvar5bdxOBh9VuLRxFuUHgpTqGpcQ6PfmMH4B+nQBNH7G8y
JQ8StD75KPWz5bAXv9hLlXQm7NxK5BwbBTSYSdo/SMvDqObRF7fw9p/8Yp3FMgEN
pYgVMAW6uycO9PyMzrhZP9eaaKSQcruRWNL/hIJ8ff2NUx1HFJ9BOHhP8QHsm8I/
mN1BuHsdZ2ZCGCx2XOEkaF0odImnkhhkomQocLbQKu0QGjkXfQIUFe6IKgqvdKAx
vewZknCgXRaN/SH5xrImsdNHvuzrmi1Ku3nQZrUoT5Lgt1pJTd5s6QAjc1bdJxQ7
EEnMuWloa2elXXHObsTDRLBv8teG+7aSL//ljhWrMBq3P/+BP9j8B8EeIv7hvC3W
zf/XauQIdeuDmJMlltT39EmZ2F3wzS+dyIpUMkUonNiSEY98jnbHkTk+M1RWeRLZ
W4VdM/EjiZ8xoSWqNhb8e6Ms0uv9y3kLfLyrwPsVMIXts4LVVDFuj0V6Ikws/lwB
nqqdm+BB9JZsFTptatPyQygc3UfEDeULml6CTuKWwLkLS8sU8lfg4f0UhKBO1xzb
N8llN57POmwWMJ58tMtPQ3kAFXUR5xE7zOVYw1InTaqtTWggQ3AThEpGF3tumewy
qk1gl7gd5cEMEYBu1zeJtATAlrA5fe+cJOw/kJn3pBPBzHOH31Nsj3MVPBX8+0/K
OKaFzx5vsn5RBh/u3pqTo88GD7SW59rgOrH3jvaHXV64gVF10oo/UOx/FsruaFri
LK2zNLELRpszVLsG3mNr9tjAjTkIsRgQC2sU/ItswJiYN898W24J+DgUz/D2RUh1
WZif3W0zHKS1LRS1lAdOHIIBfRdUHLSyIl6TYrB0Uq68QYDd3b7aHZW0m0vY9Kil
YNUmRdnPDNDDUBn+Ewsbcp9MY6fcZpw0ie4aiQVx8B9286oPY1+Faoo2idbmvkGD
XwavUM3Ww3l+MFUaSbX+Iw8e3PFPAvbN00A/t+CwmhCPOJFN68gEmhh3j9Rm9sWo
nVO0adNHEPFt50JniZ1syOxmFOgD0NKNKzAVpr8/8AzTx08vlMe2oJBu4mr0vq7k
x0pbRffLcUwX1pyaoNfJDMnhjGZf1+LWpGSJS2Dt9J2oSCNAmyFopLGgN7DoPbDn
luhYqy2C761Ki9NsuHgyx34lSqnA18omaQZmpa//GxItcl+Hjod9cNi3J7FZs8q6
OntKOn75aOf/Wi7rBjaIIcbxrEk6dOjYKsUVFyhfzaLIOzEQNq4BVwqmfNMeLqXj
PB4JkG/qN8Pp4I6jAWsA25bg4D1LCgWed7Xc6Kz/d1AtMuhvUWpIf2NtrRyp4KHQ
70rabie+w0tIWYRfvrhGCfdSJV4g3AQzmJSFpLFPD7LjGISDxUdiagHsJlzs3/SP
ADUkT2zFkKvIN+ay+5Id2TBmbnzRoNa/NI7R1ERxcnBBfBICGqrRml0X6Wo+Pfxg
ezhDgphg7RggJcVwLYb5dgtTUS5weehRSaIyx3wY4sz1Z3OHHkOItEZJbNpWKwIe
3wGC2xEOBjyTQJdJpRkfwdVvK59WoYuuuju8PsQIZpV5bwSyIhQap7mdKPXtcl9b
SeleQyyEpDv/HHoPerAIuIxrTMKP6+aHIowNTCZ+/g5v8ud7lLM77NF2FUNRTO4d
TS77WcYJWkrkrJhBy/ZcqIMRBRo+Qgq4hZUmdfhLkXwKEGFBuEFMWUum8W6ygFyc
nbu0DPyrkPL/1carOxlr48M3eWTNSwwOTHRufYtrvnJ/LizNTfB4wTw5yxN91jNS
hE36F4qPjsLMuyfd4VUS1CS3ZpnloG3wzRJ69alCrUcvT4wLQ+GEoclcIb3qibux
YgijyZBw2Vv+tvUdQRMzG2Xuon0gvWz618ZqJIvQSb5CNimCBK+dXuNQEj5I/usi
08aTw9Hfjj1b0VhN5hJmyoY5uiYhMUQt55bGM8rC9+wZf953dZyKNymWCxNgykBW
IBj8Y2WoBGs7YFKY/oq6xL4lFe81gBndaVSAgmkbPDHXOXLIFy/UuijHAnS9Iivp
HKsHnup+Dpn16iuwQzwCbKl93/GWwtgWMEeV5nC1rnqawNwLDZGW7DRM30d8SdKh
siaE2vahu0WqjUg+1GG4/IofkUSIYdqa1/dJhZHE/RlIaA7GXpXjXTkqUT4YdoIa
ItABTXMc5xJNuZ0ToumvSPsCtD3QdVgkMUAE9ng9mw1BuiEES0VVApJ8bTFedx9M
rydXnFe281N0L4cRx5piGoIeL1L0IAKcmvwEcCX5AKBNHFS9GvNST+nD55EfG9wy
SOoJGhkyKTyHg7H1UOxXljm8KigW3Z5TffmFUMoWFDQ5Fm0/XZzgEX/y0GfhPrYa
w4Ujo57EUc/jAEN54jSxEVhcfGTFM1GDmQswCLeohpj0UgbSUxm0jcEHB07kflaj
vOkFGYdgxcd2wgT9LMj70EQQxEwvttAzsTKo9C2TkzOmNnP06EEZvIhNkgEtRP1O
08q894tRbJMrcp2EbzPOuaqEM2BgHKdsgRDJj9kb5V0XtF9vjtRFnCN+Sc2JnSNG
v/kHbOFh85ETov0IdS6IGgwPxVzcKA0z5sl7puJR1DJcxP1uRQWoEch39Bo+UK5Y
qqHXwDjU8RdY8HOn7lHNo1dNqBKaXoD+VD5THwA22dhsJwArHt9MTchF/2KRRNR3
F1wdVPE9Mo8AYxZA6XaBAMSEnfqwMqZZdu4zcqYuJ3G/jnd+rPvN36sZuUUxaZ3M
bDhqdobCVwHEM0x2O2zQri3NA2KRNHgxYGzgMCzwRwXoART7i5QB/+PBitz9MbQS
S5XP/tMrNVUTbaMXsQ1KjA9Es1xcxgDMuhEia0sThfPdZg6nA0dY3e3PY4ZnoW59
45kshM+dND5IrWAkFH2mHzRH+1TrxiPyhzA+NkCRRmnlFUgklfuQR51q6G869ogD
cxvcQHkf/Uoan7oa83k4GcReCmO+4RGsCBhijcCdDO4GbmZtF6qjnhTUY4v8ONsY
U1Aogsj1SJm6H4fvZK8PIhpf6I+S45EesJSjlOBU9m0Q15slaRZ0C26V5D39cWZ4
awfCaLXQpoAp2SVj61ISqrqE0nR2GzH/idR5YuSEQ/QCsbsa1P8y6h+YjvyO8VKl
V3UWEje9DP0rHNcp7GDs6o7YMUGavKln6RUXryxyxodB9EKjfpYpVOlxAUa7rJZE
Ht2TwDkUDOQqt4seK8Wu3oZT7adio+EQcOdJQfelt8wsUV3oCqcVVtw5S8wZsat8
ik9BirEveWqyVeKWydx6hW86FVeFuRrcmE9TnjdBYLyCNRYctD6UkpFmtr/7C/Sr
Th0Le8K1G+jfBCUKfeQrGjqlhHR4wJxBN0pI9ZHaNJ77aBbTFvA9YorrxqOkckFo
L7FMaGUxpUCpYM9A2NJMfOjoVW32rkyVwUXlRHDZu64Ah7kt5bnx2X6NSVvaIwmH
6ujBOolFvtfXOxv6lDm1hgRn5/lkp/S1G3FjqCbNMcl1ZESXQa+PRorGbAT5bRVb
cXjSoGo+bOcRfa1S3CSHsDvR8oYYvCdsld5Jc7iKqfJm/w4EqdPlXUolz3lE66XK
8CQ6ALALqIYk/dKOrK5Gt50uz2tywkkM48OZDJb4OZ2arfnqxhCaUJ44aWFGz9i7
/i/vVyyDwHbCo5IOOx0Wt7GiuOBY16qjW6b7RX7c0ud4vkXdroDUTKunk6zzt/0L
o7lZH9XZ91ic/3DPDwhT8o8GG+lf/2I56q4afGFfWX+kmkc9/WU73NrVfesld+eJ
Nip19YgTGigIKqBPo7gl09Rj2oMkFm4vIk5Wgl40UCXG5BGkc4WiuHbzbNv4rBjO
HN8gNkkTINED8tZ7EF3Aiun1ePkzQ+MzHd9T8vYwPQnUdpG5EnBUVGm8aU0GB2lm
7WXDubmcATYv1olw1+zujI1M1bS/2PuI9WiC3GXkj8gcub82o8979WZ2l6UH51p8
iSZ0sulYxQkiHAJcgHwbfHGObCw5HXfWMzaIc6W5FPTPiXN+PEElL4kIOXA6/gsg
Jc3wG0ul0U2b8muCLdLQZX0IjN9DfIZWNa9Q2yzih/9SnvNvjYXwy/5/uPbuHDBZ
6/WPwFOMpuIPrFZ3fAH0hXTIaP1eDz+SYBV7mCOMyqBc2UAyH9h3rcQJN1pfNVIk
c5W706cstLPPlc4Op1LcKM+MtNg+Ec4e9oi9qEuBvHgGULPIWP+svD96UXqnJ5/C
ThDDlzt1vwjLKRVhkjFwIiLQNCsgD8EeIgXtQKd8OwEcKn0fmbGWTDX8tyWtmK/L
WOQ15IOD3vp9g2ICnvcuzxLqhFmFc576+FSymRof8l054Ok2gs2f2Eec8dwTK5Ah
/J1tYs0VYtwwkGSNoZsEOTWCMmtAWPXRTUIj3Sq4cz3DL/07uwB8ha/iVn6P1Edr
xWCyl8TsFf3wumiDje4U5Y7WwVzIp0W6BD5PF1e33RHwyECcezqcJE13EQkQ+4ij
nkQsTfAgXs89hux0dCYangrBsJKhjsVtUxZ3dCKd4cK0u+KcEO8TFK5QSWSJ7s76
3y8mnWBUZMXAGinFu/XHv5N99bfm0sxeMW/TLS4R0GdNy+hDwi8nyEXrIk4p39yj
gHaWCT/SOWySkibPoE8/S4k+GZdjhUxNpywsGyuJO8YfqZXC0xKmjcdS8nPSs14m
0Pv9zu1WlRTnDyFVQhThGXpEgtalYT1FbKx+xKVcP0MohkbjoVru+wlOYhO3jJ0x
4hIgz1ulXpYD+ye5pC3Gf2JxcqbAsxW5JZqu4RDT2rGc9wGEo42nPe5IJZ9tb3r6
ZZuAiaVb5ezOB+1ml9Eo0Bdr3hqb8afUTNIi3ny55KhMzlSGfmxNE96W3h34LKYh
AQ/i11a8v8Fbkhfx8WQQaDMfpElB53pORKvUtyDqFuZVLxUa2X+Q1709agVcmKZj
FUwS0rgdsTgjLJGq36ZeywmgeYKj+1uIK1XgjY0yk8zaOgmy1K5RG8N5RHCLlRcX
9/L/RfNXHpu3hKJ2wKgLl9aEMdBp0H8gvhyZvy22etHdMoSzGkOVH5R3AOInoirb
fRP/QojQ0BDp78vgiJ9y2V8RCdqXdXKrgksIBlMWUEGkM0m5gmVrqYBu6jJps3ur
YX9I12NDJsDJ4xDtXmrtOJBgSHyhE6sn21LKEmDeXKZ028QjQQjYEbaPdE9XmM5m
ClfKOySrkG7NufkV0Z5L6bzvj/PjVCLhPAmmOwdrf5rP3ssM4QBQaku5YfOmQQzm
5XTpfnPShqQAKkjKYADWUfzf7MmkspPojjVc5n/dlr5FZVv/MswKL7fWweg4M9uX
DhMj9lDj6J5kIEGcEcs12+WG8I0aehxxK9rO81tFBlwFy1goo5QlUGqiYmBrv2vN
VENMVwl4Xv84SEVcfmWZAQlRH3AweQx4tu95R02ykUKypQk/nC1WEC/hc1Td5Yfy
ka/sE+UoIC8eB5R9CcBLZs3Bq9E7I4iSpgqvQf5FC3yPWI7xBCEisNsmlKksmkUh
AQVW/MMzVAB2rzzmRGzu9wPej1OPWw8Oa6M17wllxfRumSSSCLA/rhFwly3TmHlc
aqo3DOL5NyOMk5ljK1ysx9Mis9NY377ToE8CjCLQQ0hIRwSxrSm/gJPHdWiH8Wib
RnXldgbtl5ndLiFLsHzRm3ZLfRh5OT1DX/50qvFMLobCWdHrQso8iOh/Hy4BQYFY
0XkNNs9F2ZXQQbDH4LSPJQcD8/G5dMKQhnaAbUjfJV0dk2/nFqcF6t8ROyTkRvvG
AtywF6wA3M1/q+MdGmiHJD7NMCmRXi5NlUl9aCllmKQIHMmRQvj65X8AVcai51Al
ecTmq5FCilS2gZzh+BHXSE3It6KnHFhn6hBLm7SJJ8kjEt+/Inq+9f/kPyXstj16
1pLNMz2NIO33vPEpvnlvIsNmkb6/U9QaOAGo1NAxiJ1ETm3bRAV+RGTpUQBQiuaN
Ez9m3KDHYmzafjjaXegyB2PtEG/aGpTr5+K7zCf6M4uofgyt9ZrqPpD5YROGSJVu
Qq1oV+DoYjBhKWF3ZD+CjO3Ih23iTLBW/vb9Ib4HQi5hdvEFPE38l71EWgll5vx4
a/pNAk5X2vSYk12QsBFxWZMM6bF2oy4V7dNsapoKScwdQ+ZLWhU+mcF0sJTjEoI4
MznN/Zdk2rWt46s0m+SFay8/UYcDbCKRARqbzt3w+uiI4Xalq9RlU8zfArRDPnJP
30B2+FGiPmxYmss1ayAqWugBPdnBw67f3ELkA1xyeDgbVsk2TenfFs835iMezZSk
ONfB34sNWmlUebxepy51gdJV8eAZodQyvTxC9PKCmMcXBsL9l0JU7hT3XfcSbpUx
jctEI2OMHS7VMYGB8H+mddima2RU0XwIsH7jM6UwOOG/RhGSII0P9ZHiFDDvfj0u
yAVHcibgaQ4WBHlRbxjVB0R74vJq8DSm1rPVfx2iVk1j6Cc6rUQc4gUvyL8OxxWs
ESBiNj134gJ/w8MH8q5lc3USoYMAb05q8RfS4NoGtngsgJv64jQl2bt2D3xYdCEo
dMOpwXotOCJKorlAztFl9mrYBtu7CB9KYI2EVswIJNWNX863Ag7wW3ff/DFaTU34
DiyL+2Ww903e+Qo62EPjRo0MJdoBlFJnjLyM4WEXtK3bypNiNZ/hk8vojmb3KxoB
amiiaqog02sZTcASVls+j+qAAa6jgYW+o7csjLS5QU08k6kFeYB4hVUhqpPUJgTj
nf1gvNzpvLgzle4rehtFolW+to98lIpN4RL+OEKwt+M6zUxnn2QR6GwThjXHYHIp
m9nnWpq4onqJFw5ctUmw/gPphYbwKAApH0yngQXMfN2ecABy4ByfSPRtx7D6hiID
XlQQDdUH2xNsbpbxiAKiJhMy/UR7835VgYjNJ8E0NsNhrv2YdsunRabAomPiRn5o
v3r5WgSa6TQ9plg0Vl7O21KsvqGGOF/ThpUl19o8MvK3Qg9Aq11aWrrWA7nboYWJ
lEVC2gbQqPDBfMta3tscnP0LbSNjXQaxxRFj7LA0A+01bEI5LpkFkY410iZvQaoT
CDULTTmNGsOKewe4HM/N/SU3odirGtPCPxMkThMtqBqh4RbQAo5dpl3Wt+GMNfHu
EyGe4flXRGYaXPm+lvlwjLviNWPinHboKJsuIchT7Kdi3E+qljltInTZTUmeEWRq
quBTCsi4WFdtvjMn2b7QVHd3o+tXOEItmn6BENOdv1YkIFsAQoylN36/M7xdRt1G
OW4zwANgg/Q/L3vzUejOMFJdVMqZbEC0HnTJOHggaUtIyfM1ddVIJcYOco2bOD+G
U3QKs5xC3+MMKWJ8XjaTL0KpjXfX5/LZAWN5udoqJeRmh1QPl3ML2Bh1BUMVJ04E
jyxAZe7QHkrT75if8aezYQwveFxbwbj0lWp3gO35uw1Xr+AWxA69VZOC7Hd0z39C
asjOymwV01XtBYcRKpR19JTQJtlyNuTvvpj0Tgxm9SkLjlAI9LsIBl9zgN/prDnU
bXj31Z1nHezJRMg4UwdLK11is8joGFXi0KcmmzEMqbCUk3zPgYX/C29ujQ2lYp4n
+xyt2x6lINyjkfayvQJJYnI9/sNHDJfwbntcNboK1Tde/S5okX9AqmgJG+fxWV8U
ObnnXDSV9AhDFKUC8i5krKeQRyj4XeZlGfXCj/AHq3V2pkjazUs4izYD/46N/W15
3TvcC0iLTfYntUFlbC3F8naeQOm+wGBY/Sgch8LgptfOkmBwa1R5PeM5HPNgHO/m
bsI/UG9TbHWHm0HQ4KyAUx5HK1VyYMPevZ5aFPsaJXGhrPf1bWFkKXRwmM7cIgNW
576gjdsavpi5Uu/DVLtPFmwiuGiLTiKfuV7O2V8C4tciT08b58Ui4V9qs+M2P426
qEkahFflb1McwD3wCXD02+1YNOlGevHWwJwBMEJZy7NZfz86aLacY/UHX4EuE/Rb
s0c3cTz/qp34iPIfIpqJqTFae/hA1ASsrkxc3E7/dntF3RyWfUkbXkaTa9Orvkot
8He2YtkY0IgiUN/i9iA/kIP6pN2b50skH8W3KlB4DXavynLerQVwXGkpRYps0Q1b
k/t8spOITGFpNFPh46SzC0a8AIXYBbQkF3pLBelW6Lfspl67BcyVWrFhrpA4Im2J
tvp+P0Fv+G3xPQC1PLDHHgTjH7w2q/pa7Df4kXMKTwBRMDwSFdn0F+aCr0lzsAKp
hR7lbGrsbDcFTU5kZ3HukGKJxmQMQBr3TWn6Hbe/KGYt4nV4p6JbFWgVr2b8blcX
9ZxvYEs16EQDNLy17F05vvSkpDMwmwEmGChqIYfIDYHEgMz4zuX/d31X9q2fvxaD
skp9Le9OYFpPMhtea38VCiPNHrFCsakk2037obhA9A9eJ+B9VZSTkH1MGQmCG+mK
beFZ3yKMXXF0ajTdkv/ycHr5MashQWHWQKptPjz2MOHhi/6zL7m3Cq9GNjJkVSbb
H2OTc8vym1+v31VW6vHRXQ4iABw0qaRDPfGLoctujpsy3kxaJDB6+O8LzGVvAM75
00qwNdWXbyts2fJr1bjRiz0E9gSSlgElFaxpVOYw94ioKWyUFSTYRjpgkeJ6m85N
vdajtUg++ZPWm4Mbxr/sy0hDNb9pSdzMHAwjrTqnP3DwypR8oatBupR6UhbHyTZb
DeMBm+0W17L8cKjLviPR+ZncGBV4NtvnpGkhGY0iZDBmbVjYozPYP4f6ZJ8nuLqJ
hhxuOBmldko+IqGxLpqc1+bCzWVwTJegBkRQ7twLlGRoGZlBr4jW2ZZMkiiNlKNP
VEXUamsrHDSdB96ZWKx6rt8/YiDzEx7VkgNIZjOnBVK0ZPxSqNj7ToDzLoseAkyn
e+6GwMguNdV7VSj9TLWmBpWTir5A+Qmr/4nex/+Zy92UH2DHjH0VhKZ46ODBAItQ
8+0MRKASPzOLgWm2WAvP24b74ZHtI1lgwFGNNY/4b2D7LiPlUKroPD0JQdzirQN4
EjbSJIPZsX+l6mLKkMHM0I3IIPcEIFSnSkA/ZR6trm+eQdTlDFIxmmVrRfNmbBSc
U7qr7bVeaaMyvmnLeuMYSiiUCKw+Mip0Xo07y14r3DkpuiNREKX5y1JfgMsokoUC
b00oVlDa5e33mDYmKgXvZfCk/MCO+HLQzonGStDjBwuQCoATLUhZ72/xsfS7wr8j
CQC6J1t17rjGrZB3m2u16VRLGKZdG2o/2Z/2awE01Hj2C6NaOM9l0Yq5pQerUl8+
2W+fcvOiq4XcRJoS049fDCQE/QocHsPmXxC3la31gBIToh97A8od9KXBOAhzsCHD
89T9Q/gMZBPlF1CBFZQkyMk/DoNFyD4vXuFcmKvKjUb9iUoHdSXUBxG6P621BfUa
hKe+v6BRZyXPPBdbTC1aHAHb1wYp2gKxIB0SAXIJXdzxS+j6NsEs9NIc5f6BIpTN
fxE0wePCgMKAqLD4CqT7IcsRs3JhHzS7e6Oy22ULWnuVXAOJVbPogDaMn4mLZ0zi
lhk3uk1xYuTx9+84CsrNVCJnzh338WjJxBr9sy9BRonqXdLnUUhibCcAZXHrHZ6z
kRJHBAa/UmXACuDm51o6roMoJ6nIepA9tsJjl205lPOboT7CLhlwHEQE0LxLkh8r
A7gA+vRKmPUsCH5sM8VZq4OR0Rd59o8pNbnFMb8Bi33VvrSncX3KAz8Mb3mGc4xK
t+fii1dbu6zgSy3JwoRsXgGdhcwGypukFrnZvwNFf8V3a6prqgitkNQ+/LZjroJe
QHOGVFOtIt/j5T/22o2OC3blOP/i90ChfYSIpHnt2DSLbntD+sFgVvLqTCbVGALv
6rc7xP++uk66GhVcUA7Hve4wj8vx0JDvNIb+ZL2Z6jsM/LaDkcNviHClXw5Z99J4
RIjefCwg4ZgDgVZIPmu/5UwAjp1gMCETnhMFO2qJNdF29bFT5ibMJEfm6rwrz9QQ
TBbZ5xyty7E1VRWM0w/kBlICuY+vLire0IL3ZYNHOTrjJqRRz4IjdctUCdT5iCc/
tg+P4pGaV8j3eSjBRNR9l/C4TPqAFIFt/hrw3wa3GKLPQxIZj9tXW+mXdBBRW1px
vmrnFIhrhCyc8xaktGFlwmd6a2TeQKR3/D1n3cJcgiMqPsfX21Ddbiq6/xE9LYnl
gaRIWRRymfrImL/RVNXvu5z06yjhiTXIACETicpxRuKYa62Ye6a26Yb0/KaYpZlf
1IgQVOGzojiTBrpYa+U88C9k64I2TRzaeXQPmCk3Z28DfCYBIJSHLS/V0meT3fyR
QEjnIHk4Df4Fff5Bf+/LKzAlTyBH61dFZHCRs/D45Csc1Xpaf1R8JScISw6J2oHE
RfgjAEumpQs36B3qIzHGPUHJ28kVjXEgmpnh73A3EkpoDLiqaSFeFAnAJIsyBQQ+
Raitv/4k81wYDaN9feLoqifHLH+CNHKG9WmQVkenKmh6kcKcENUjOnpavl/Z3AB8
a8z4bFT0y1hK1DC9VIyPI8fTfdf55IppqVXiy21BLrAT/9zXinzW5+q9H7wVIuOx
ablXxECZcshxwGnmPGBD5jE8qnbjxUzHjasj1YnutRryy5LB2XdNMi2i2vyhSArL
k0dFOdocTu50cf4De7mAnk5vRfq0FY8RrYP3kOm5JQSsoLk+6qNnvzxkxQoGbvOg
G150G5X0wTIzbs7bdMK51Tr5GWpqOugdQRYaITBiA7zyBuokQJ+Sjb/5rQc6s1cO
Xov0LuAvs2xQnRfCRq9olCYAqcetUStyFu2B0HQuTA2IgF6qgbjslnfmfgkshD0j
bx8lYZH+SOJ4C2eJswgE/dQy3w7qhTZF2F7/ulZUmtPLO8tc22gOxsdCH/BtXh46
gceeLFjUc0BIuNf6kVB5tPJny2QU9l2By8o0Wy+PswMTbxB93clnKYGGh14szr5o
sTdRlkkeJW/QhCL47uzv8loMcN+yq2cP1D+O/g2OLv2YPLOeYeLjCv8OFMIE0uDe
TusNLJDpWhebi3kmxkMOPlrqmYtQofYGxChXYKb0nIGrf37dkjgffGrMgaBTcZDR
iHdB0GlJPw3xbXCpXjwbWptdBDUMCFm9Y63PP/ClQr1aUy6s4gk666K8GNDhP3Va
qJsZryi8KWTrzox01BuW9l7+p3fZgoZcA/ocPrYCTPkzX00kaN5G6iYc8fImAUXW
Y3yFUN4PhQ0KMmW1aX4UKkbqm6PMTEDTn5FEZ+5+JE2xXH0rIfUu53VCOoL58V9L
driD7h5FfJNd9oMIsXRSpBfpTYge28AvbQsc6nJCmnOe2OLdGI9db0KLo+TH036K
kn1336Kg0XQZ6RMF1CGS3NITOIr9Nt1cM8IyTxqszfbm5cG1Aqqy9byMvdqZ8GTb
6TOoxKW/sfMQQkuVEmnvVeo/Y/kwyf3c5v8xsUpsx0Z5ula2CLM8NyuDkdQals0Z
8EnfU3PG3nJ6l2l9a4nJiSTtb6mSjMuojIHpeAj9/FxL38yhDGNNF/a4gYhzBn08
ax845iBHgI7xhR5y2tH9lPHj+XFf9Wz45ntB3WD5BFHIxewMAsh3R44BGa6/y3r8
NKjg1toWc7lzZ8JbzHXdctAjHKFpXysUQGNATYEL1+bQ5aOaSm4+vU/NwwfEFE0V
NxhQctCvejt4WpYyaWnXhPGunYKBUbV41HhU1gyi2rb2KNVIUot03aPXkOt6Xa/0
9iu86NPnYDWcy+CB7VDVxFQSOZ7jV32JKuWDw2JDVmvxZyuhHyrXrRQNlIHlqUSG
0XCMdR4alSDpK+zFe9HNXaQAg3g4hzLZCVljVKZ093Ttk2Swg1v9cgPGa14+c00H
/Y1iYm9uzx/u3k/LSKn8x4CIwrDyHiu8ZGcN+qq5Ui7aeExGAh1SmtHXkeUeTFnd
Zbvr50A3bL0T1cMyy7jpOWZ8am6KcnvylkbF3r/ZhIwprBaT8jIqU0V5M1eqepa/
SWcaLMX7r4tURsMPDtRJ0T+o3xSNp/BLQnei68iRv4ymy3FoLLOc3GbNZnWKgoPO
8fX43R8+STzFk1BZL7DOWAdzSvKgRBg+vhfRwcKdPf7OTnpvXzSGzY18+DYdkUgs
0780RDOPwzCfu/hcB7mba32VSSM9KQStaQJX+MZWyaNSJhMa2R6SsRaW+j9Le/f/
xOY2N8Slo9WIrqUUKSR3ITEAtOHcdK2h5FndwNyjKohSJZRl/SBz41NQboZnVDle
hhAvm1uN72NSU+VElbgaq9ZbzG1YK4lGMd8vrx81UXzcSDcVk9bqP7Tf/SYIcCBy
TPHEnDlQah7kkvZBO6ysMBJbJopO8Yx8iFCRpb98yj2A5C39Ta7EztkpjXsv/JaA
fucdZSMVjylDYsc6snm5RiUXds7iNQD3kCYHHtniFv7hC6s9toJ1PI4GYVyIs9WL
ib1b27dkiENOl9jZfoS8goqgHxleL2jPstvpa9KqRHS7+uCs3w5EsIN1HCIbSk2v
kfaXI9rkk8U9Cz9Iv1i+Tx988RpmKQbthHW4gElYAHEm41FzbeeK3ooVNKXaqu84
YuuOPrOh4ZaOvMN0ZDPKNfW2CksdwfUnBW44GWiZx9XeC7OmpQYZByAs2sTR8wYK
k2fiLyURNCieJ409b8jxcL0Tm4NyXtVoH+SmTTHAgJyzyhtWjscMjdW3pSaqvb1V
V48sBv+JJD85D3Xk4uJHEBUuUKG6R0Nvk3o2KuAcYlBGZfOZahVhx4PfePBcEHPa
luUqmLMAoQP9jtmDou72IdKmebpziwxPEHrag1Q0SJXoyfHBDDlGsJQCWG1fllr1
KlXi7mBwjWy1qOmBq7dHg0gwwNJZrfDUvWYqDgT1lCzCbyXdpjlCEJJ4t5CrfG3H
IvlwGEIiY0UdLOv2Muc2b4s3lG0tlsbE1gUHk8ignhuRzg/BwKz6Mv/EuAaTCdtw
xrXqFsk2NxX2XfVP56IG8jZLa82CE1YakhT+PLjoWvif9IRal4do80EjZxEw6SCb
TeJhLtdfFIVxuuDy2WlDNTRYbh5z5vIDgXxvRkOkc/PfGP6rM0uwNxxP9xcLMQZ8
lDshvh4KoJQt0VVAtWphfAn+BKsase7Qie/ON4h9/5OZ2hPzhJ1XPpths4SGSOfb
32BDXwhvppMYuVGrmbuOOpH1dK1+ioURKtV25aDSFBCj11SG+BrgPxv2WYtglqVd
XqIFgoOsNvIfnWCnQJeQxc1cyMCka8GJVaPMAoJXaJQaqNJHtq2KDotl/VcX+KNa
OS4WMIReiKeF7eDLCsTsNHcN8I+LHbMDrA5TCWeR64WoxCVuBj+i8J70wExrREr0
Fn222itjB8sPWU48WMvbUc8Zuy3w5a4W8cJV4zF16Fr5cXUUOfPCn22JpRlXuyn8
1Lxs6Fn1nJsuPJHtIERtsIGF6Vlld+5v4sbxWBoQzaZJ6JuSo0z1QaMzDYqASUYf
hweIDYHtRve0tlzwZTG2FGAOnruJ2n0x6XR6WtEQAKI8oPIlk2fnL5H9frzHPu6L
wjjGqiWZxMT2qKtzrLCtkbcGcwAx4j1s8kMiiFCFOCAiaIDVYQA6rQkvu808BLqq
nFCbR+ez8MpAl3QDR3D2OXpWE7ZigQeSCjKOnghUAQYYPmxsWN82h6/nSvppwHWN
SLXDHPwvbz/SZ/Oiau+sN43IhzYjCBvu/iaXGKnycyDzTAkJqlZX9y15kKnqz7fe
ZeT0mmOvRoO9wYq5bDH3leFvPrmMVvXYI/7GVTXCC9VthQPOzSbgjSrnelAtfGjV
go0n8ztGc7a3WLoTBeg1/T7OXQy+0CQA9viTCtObFV3fJI9NsnXxBuDhluHMv/sk
7Nhny0wPbRpui4HB7UU3h3Hfui8qcN64MnpBsTUSFw9dAZUT6n2c0onMs9+TfU8D
rtJ8CuHCluMB+EuZY7JJTXDaFTQeU33t3WXQ5Vn8NsdEYtrnweE74HJ62XLFE/tY
LLamOgNm/B3ZHPhk+50AzZdK5RXDez2hVSScxwBV5kthi++n/9zzaGHH8p+a0jlL
kSVsZC+a+TfH3HWZSAlaW/sq0BGI4E8kZGxyf4FPkULkG1I9hU38vb/Ne5Hr9Og7
sAUk/2FDzrbygJjOc5iwIZOlfhTIfAqEvUCfaakYsaLR/oKeqguRBhGuSJjcoYWW
udfLpTaCWdUERQI788GMei4zi4rEJZE1m0O1AojZYYXlOI9nKekwgeXz1Z76KeEB
YVjkLtiHCcY3IECQc8b+vBELzT0ynsZhukMtfxJ0ovD6QK+2Hw5QLulDv4IzN3Ji
HmNzLH6uCr5kgAFleeMbHN/9jDtm4np2dhIFglLxgFt7YIlY52AJTPwsMc/NrWfV
5XTrRbU4qpoSc+o2jgpm+499EBB8PJFmLOb4Phfg01xe8AxcHoaF3tfMXZulIJMy
YEFxwWq5QjIZ0iHkOJ33lw3AZKoXLK8Uy6I68h0GnH2vh4F3v45OIBZ2j5mZfN+E
TSdrTJuwXY6Wua72nNMH8KxzJSIC030DDUkSdHK3NOSKkcTMPuc50X4hQhJHprLL
NHlw9QTLcpsrlqiVJ7To/r331PiOk0/rhuep+Ee+t2fyBzNZIDRKQbXUy+HX9VL8
H5YHaDjysNje9zngfZMfSrv+k6SU+R402ip4JVTAyNwTuqsCQCnQ2f8Wrlh2V0Lb
NRIKt4zTIGOP13E7poaKDOfpTYuBl8Xxybw49EdkDlCMaeQr14u9+dkeA1ScsvLA
NQuV8HChOAUv6t7ojlM6QuTzXRbFkf9dJKFwEKThGqs2QG57PD2ojOk54PMsyKYQ
JtCGlA7GlWE39C3urh61KAtEs7pRmvyQawjmce8+vRdNhZfIC3OkCcrCn4ck67o5
oQulgL12s+LwyQp8VdULYjqQwfAg8HoZKke0/9CuQuhU6Q1VCt4f1hyf3sc3HGzs
gu8m2j9iRoPLskr37bRNvO7aPOyLz2KZCtPdrxZ5Slu6FoORZfA/vNirFCiOanJC
GsAxjcdpP626nOporzozeilOdEMve9/XIwRWylE+anrVTay5l22TZ17LeeZV505B
sSc/3Wwm9Tx1NhQhxaLT0qGYn2EHignkGL8Nx8u95zHqi0Dan4/VGlLL37L4xUbm
ele9tKA5iN1fkxrTRfV9MzbuVgeQBFrAjJoTMDGpl1AAJw/qosIV7oNdMXalOJy1
D5xc0Pd/LPmRjohr0R7HdwJ5J0SoDh0hPVT1a+J/yispUoQWQ58ciE4jCu8StLfV
U35UwDAcyo67p/yzMfYvpMnEZQEfTPiK8nUdVeOn+KuyL32K3K891DDYyCD/49eX
vynOjXskfkWkuATTLPi+SZJPSwXuO8t0ZlvZ1gVglU2cfJSFLlgrrc37HjnA9qEG
rqn5yx/W0sIGDDLwQElNBTa9axAqwpa26/0dO8e5lqNNQgpCLVim7xnOvPwxQ6mB
hPMI3GzA3XfRnePwr2JjBYVGwVdYa8yznjvrrYmRK6DSHkJwA4hxz/8y+c3i6My1
uBfa4VMtjutu4luAhvNcDk3zsgDnlgGoBJCXRkpw+1gTVO4hiMZMP0xHfmdWmVd1
T/VQDb092YcUVZi10HGPl38ZVFGNF83txGDDRRU3iweBEBnxAc8d+TCoMaYS42yU
QYuYYPxDVr2eRUG7kYrFnSKZAPN3DHW+tloKyj1Hiv9KhCMl0Y6Ea7iO/303/CSn
CYlJqLa6AJmjzhrOVR2UHn0sF1oCD+JIL8ZvJbixpCfUbxcItr5kYJjYCk2L+USi
qQH72FG8JKNHVWNv+KD3v040N62Be5U5a4r5ZIYvSsEEOc4hHPlSnwWHD1UI8ZuG
PZ8YeklTlcEOtc9WcUvySWnxXhHaBRIqZ4ZKEgyy6YTUWmjOL70mt0WiD68dtP8m
eTYCHMZwNGTvlreOyB7wVfa/nwBTAHS7sM9Q+ErkLLh4SGmedBhCp7kaI7s6AqcP
VYHBIv2ZRttnKkdGPdrsacyXP3No8fC2PXDpxjkq74SIAvLjk0yaC59k7MfrG3nM
at3GXE1GZMISPUWRa+ApVDinjDachRHT6W2SEhaNUrXi3NR84SlEsxWFjgHhJCo+
s1VE1HGkoqif+Dgrpfkly9tdQngPrH+RcMGBAkGvS9VVhNuET6zPMAuApB8w1s0E
e5YMskKItwFUOLpVaaEvD7B/tAQsr/+647eL6cH5AxIbtwJMFaobrZQlcLsxbmLA
SXJEJYItDGL4zGpU7f+pAZuEOVT9+cYaFdOsNtXh3escw+IW6h6gIMeDSJ9N308/
/J2BexsGExhrNgj8ESA6jdhyQ2SG0PMnPwJTtrBX6BPcnFTbv18jg2QPwJ/mhfwo
jSexyo896XCP263eq/MOnLza4YIjqxeQIJau7MZMUrKdHx8J/IYV1f6MLF+NZDQ9
/GUEjY5Hg+NOndu6nW9z+h0/SqqOPaq2Jyu99JHgtfiSSlFCqM0EGFormXosql21
kRzigcoWIYxk4gp8ZQdAv22BQH/3YiUtsjBY5t9pJi1v+wCCTOBxQXwhBMghN1VB
aHuLftU6/JE1jiY0Pihlq49C+cKEgfs5SPsLHoJQgqntOfrOaskoK7OLEUEaYxvn
G2P8zB4KRe6al1nNXfdOKOU6K/XQ3HgM1X0Vw4awnn8ewd6WVevSQ4GOeRbGsen5
tUVSZfs8SW5SJUD0bRGQwPoLj0jHIDpXonkRQvylZrWU6Ta5KTuJWUMVzbINsWdo
tDWTa47oqEnW5r84jMZ5GbNxpOvJml3o+PlqWyVxyTa/neL08UsVaKXjRvPjOa4B
5DdUGOFhwIUSCduF7v0mV1BHGOgGYR5JTdeQFdc8HDKbQWK365X6EwSeVRE6nP5d
a85NvqGaJYuMxhF5Y2er30L56uJZEdrVExKSoy1uxvoMQmJnxZrtrTo2Nj+w6Ynx
M6KbIYjzLwJZ4mjhh/05sA6ij/maZdn/8RgepLoSYgxUcUFRty0QLCAnM8T2iYlt
GVmPjoO3nD5nkaN100hIHG5jFjAkkgDbUhObnWStSdkWt7K7DZ1VsB4bidkNZr7+
cI5f/SEuY1hPhHsyGHEmV1c9lEooRITn9oU4Q5SxblppNxJxPn+LvOVo8dmpS9vT
rj0AE3W4s1aFLFVANMym7YpXBioeRXapCOGSlSVy5t6375RD207mo7s2oXYCawO2
qzWBg/Q/p+jUEnlt971h3xgJz2t9KUDza7cOrQ0wk1vl9I9WbYj+bXH+en/CBQ+v
ZMEDjH0UIL7ki5p1Qz8xeY6Flln+oFxAqgFX123+TAwj3PJW39tuSjL1+taJY4Ta
JH5od/K6NFqMRoOj0cMUeKQ3Dg85BfJpWJi203Stazaw75DCOs3orMaf+A+Tzq5b
+zxqhWNEScsoyGVvy8YbxbW0dFCSbD+w4htz18f7NCX4mWbthO/18we+cPDXRZDI
uaZHbp80Uhe+S+spetv+/v3nuCyuGHGDK2pVZNbqZY6e2VPFQ56j1kmbpiQ1D0YB
mMA4wIHgh9IiZPY3ciGRp6fQ4gw1WM5ap+6q1IBuyi9GgPEr1dxaYyCzw/93TUrZ
UqLAwGcTnrKQD8AVBODisWsnsRVOfJPvt8sdUMd6ykVQxJmngFDJe3RktuogR1zx
dMQ8ppdTEhnNZ/VWipuOdGx9+768yPBSn+W9NqLlufjNbyiSEkABU9d7gMTOOPjl
jRTu6BYHQJY1TcX6zfOEWwXlb+T2QxaefVhgSTwBILeQa2TK4+wt43h/+9cMrnXg
vqOfH/1Nf8p4r76QThZkWH/+UPu9rN/ymHGgfiNfyxTTrJQdQXf8ezDjgoCbpu5i
waQ68S0XxXvY0ik/lbmhfEsqg6m+KnJU20D9iWpUE2JhwHsHtlcAdv9Bj+fA7bzk
1++SOMG5jEziALLZQ2hCBi90EDKN5QAQExMtx4D8IHZCqJDMUXWK4eDOdq1/gXvN
968nr8pbuKdLNuU8JHYfGtoaU/eSkUjOkysbcA0FmHBEaOVU1cKPBg6eeClSVxgK
iZzBVva6CSDpeCPCEFBsybze2ZkQ6Q0IZQLVDGqsPDMSw/54FGlZhZgO3ZGfSOLg
gZygE227X5gckSWrySKP3Kjnwlz9p7Y2cCUmoGYAfAt0wyU739Xjve2BYlNTpASC
NGZjLsSiyowYontCeHeRX8xa09ViJa0UYX2LFV24DRYLe4Ae4PPX5j8VK+nGA7ut
laERyV9WHB64ieKwsT+SsUJQIxrW1J3OyceUGyYyZ0GVCONLNi0x6srzZbhALUHj
Jx4ryxPBey5jLDIpV4xMjbT1PbZpGGeo+fbk6/ar4OdTNnvEbAa5EdJM6CXVTl9x
eoyGW86bZUC8j5STkCPvBvyjbIfeUjg5CkNIPwh/EfAZQCqNSiGjHQz+go4gUhhD
nlA2pHmQrtKDaMjIzl9XcvFslFTHj6UBdJOR2YEbgc7/pm59ZsMQDUwoh8diqNoM
0N/3kXG6vXl2uB7z6EGgk9Ao7YV6N3nu4EQDrPe8MFiyX/buvBj3p1gy7XUDy8Qb
pZQgAJsB0IhtsmlghR3T6i50rVVUuWHKC+/MccQRabQ+cFBD7HGTGejQdk8KXlSr
shbjp+KyUX4uqjQdROonsqtp2N9AVmzGdaTarWvudHQfuzAkaEaUyApGJFasFo3l
ilqJzlhg7+B1OBn3Vx2/w+bmFbpG2BooNjRIhpNS+0ruueGVkvR1nEnXUWV4hxnC
QX1a71qW83nAWV41zQzqp0nbRkTDlBNcsug8WSP4orS+1s3CcS86bmr+OwTnxaZd
/kc0XnYVoxuWjFoNZYlpSb0Dc4ymLk9USCky8W/npnMo4iSiU/VJkZ5iXuDyr4bl
bObCPjTSR932dAu68dlKwu1rrqtrNQcq8nh026cy8dg4x9WIX0SE5m0PRu8QENVg
T84fkcQf1UI38oGoq1biWNRORSGLnWYebPKigAKaiZyJYHko4DOG2KN1U3QHVwyj
WGq161vMTt5uY/sGl4DoBy3S/ho81Yyi0rx4Ao2t0JfJorsd4dax0FVfPOJwm5e/
Bwy/49gAIUgHL9mvyjPfCkL/jObLVEaE2Px5AfuIJSmDD/z8g5aUlAubnvGxUTCo
yJqGoPA2JqKualCFBH3EcZ2CLHObjaS+D4eRry1RHE2ulfy4Io8D29TN7GHcR57Y
Fahvze8o7T6OY7ylfXNXX9XHJH7nookC+XYJ/ds+447L4f0cp2t7IPHbGl2lnTf1
OrxTjD71jhIxeaatCRMJ69V0pPj0GH091daCw4D3LQgyYsXwByJUrE7xUaBZOg51
Eg/SduI95WhmnXyyLlW7iFHk4tibHp8jI16B8scWTNBAnF7Q9E9E/frupibIYPZz
kOW33z0YLg8bkdVXCeNAlNgXgLyGnHXA6D2BrLDs1uy16OQ48+UXT9dxUIdh8uNk
90A6kxqJxUzo6sgHKzPvCga6fx4t5A9Be56IhsZOlcGdMdxe7i1Rp3/cK2gpK/Kl
QboIueW1cKVj0VZubUnLTI8iCwNWXs4C/xSFO75WeXeijeC/nTBuSaeHZ32SquFT
xxK0ZpeUacLnOUvbdze6zi/lt4GXnO5Hm83NugKbdR9ZGf7A3L2nE7+bM5Jil0Z5
qYedM9KsXZg1NRwwHRh+57fUySWjCX1IwxYsL/YIlI9i1R69tVATUmEOt/KQmhWB
ISuGjsgp7XzgnrsOnViSaDCKYTm91hXqtILAjr6SlS57VVPJ5LnNGh5MBNNc87yT
y/YA7HMI2DwxQ3qXvUVo3wNXeEFjGI+FTvlkQLe2HCMDa18fRbUE6DIqpenxw67H
b43sF859LVy6Fh4lMMm8JVbk0HskCvVq0zYaD3ktNrcX6jFbQQfbMEXqHuPy7vE4
pZRTC/i3gF+sv+51wuWDRXz1lSaNfp9IJ7OQ7TKft4zDGBfL7FLSxZ/NqlJIghJ9
33p39EElBVynZkF/nsAbnZkrPzvKYN/PadOrqPYKMe8zQEypHvUPebDhjD3ktjau
PQ7+yXvJ2BejsRXsYV5UlLUxcN1GT2ZWTu9YVuOdhLQTmE/x2lcuAcFhdEcYvcj+
K5V5yq6Hwhg3KS8P5+ZOxKAz/J7++s6gD8vrWiEN2e17Tn/ZqHCh1KzEdIhWOxzV
goKj2v3vt9tDy+7vgwDxS5xJuztWZFNYhosdU2mReyos/2/fYbGOT5CnwVUx3Vsa
oZI36GX0cO1rSuXOi1EjS5hsHrdINFMy8ozsHpwOK4LSK54b0+zptnI+GCETq69m
7AgVsKUWFR7hrXyUIouL1dhW6BumFxvYL3tHZEBaZaN/a2LzFYcwKnMiVjdqLDYI
VjwS16lYh8Fd+GN/MWuRJHIQGDqzwupC8jxbNdtEX0V9DzcGeyEiEgl1vBj0xJfG
GbeMjOXtG++bRYbXtlk6uak22FP9S10IUBL6EVBiHhzFVGriqnJ81QkkBmz7JQ/0
DwQpXgZlcHNb5ixBqO3KRfxLcg9iWqh4DdfeFtFqDvt0oMEYPOV/T8bb/qC8Pdhz
s12VKNuuTHrNt0GAQ8JTxhZkrttAOTmIlCC0krqWv9CY683E3w0Cn/8v3mHW43Jp
/GO5HmpoUov18tEZ46fVNErLsLToaON8AH4JkTHBwhI3uvIbQzDirzIATLH4RwvC
1vig0MQ/nFh8sDRRLd8oFIkeqDU0DJ20x6lXJRYy8xtt6HxhNGRysVFW0iGlFBpj
znp4s64vO1CuB9qWq9pO37d1E5HQoaBq/NVt0z3apEwuwECpys2QT0unW07X0wx8
bUqym7QxzmuXloFNejc5BasvhVAUyXSYxLLyTE4zp4ssTsDdx5FAXFTtqjR3ZLNf
/4rCtanqr6IO8xXosPysiFMZVhinGNvm5KmgF2si26jCujQN4eNimo+FU1dIuKJn
T/HmU/RsAFxZ+oPikARkjCT1151v+5/T6TJbC5k5d3MFtE/5jo8CIpoPAfeY2Gzi
wOu6FTafsrllDWgclR6aVbt6BZjWLx5s6Bk3ZiGp3sTDmhZIq7JG6rrdCgbEJwJ9
+Sz7bTkVVao6K++ACeLKidPAR95ULKWSnDAbJbpMSOCMT/nHoSJx4ZLsrVyMpDyF
FeIizZ00XioE5cDzApJ5SWdZoJqLIxzBWWP7IXyfaT92d60Svtkpr6tRNfdt8r6v
3UAncQ7JS02qJDlzMtNirLlp+vEnNJIW+dtrI/EvUOKyRjvCjl+FQxwFVTN0y8wu
614ldiPI4JmblBbP3ERjaNiCFN9BAG5JSRHcyqg+Fzka8edSOV4WsiAlvSe8Ew/f
2Hm7UWpKifgrgwVYoUWs9TzbrhGUzVDcs305B9Q2XIMEc98fX5RbayGT1bu6+0iS
seYtxQA9htNROZgX1zY6uRrSx1ij3aHY/CVS7Qf4y/GskWY+leBIPNRZC/TAiSqu
5XC/9aY/VsJVsvpgpVtIDbLX23i/aWpr202pZzszmoqIs9E7aO1knrcEcxqgzOvT
v2gRmxJtL+9h1bTSSKkYwguVGqeB2mPAsuXBsXym+/sXqyKKiTxzKoWXzjYk8gJG
kHORMtXyJiHUVbAIe6UtbOj3VY8PrR+Cb3k74eZjl/S3ViU6hYkne7RyWo7KtQAF
hoEqBw7v1gNm3m+uV5rpPcgoDMRmZcvlk9MRzSA8LpTIs5fHH5ITFYkinize7oof
ULuvtt2ssrTDhtc/M3KB4AE0NuyTYJSRm8wfxrffaYiGKuiNeJ7N5o4aP2j7flud
e3euZTY5ClK/hc3J6dm7Lh1R9hDqu0DTBdf/1wZ5KNh8aC2Ymj1ARAxzaip+zvzs
ZcJ7xj0RWM+lvCPutMKLXStboYy62Ka99pQR8KMl43dEYo+5zNLE+0sKSqfp/o/0
XtzasNP2JnOkVCUMhwzEeWgO55xsHMirb0nohK21NHc1tCErAro3A8YH35hsOmC6
FOoTcu0QTnflaFdlPmltadhH+Ac/9QzsLpjsf5EgGbBtdL19QP3k8vyv5O5Gn2Bg
lEHvJQgABExdazmW/OSn0snBAENgEE414vvclYckOYTYLX8GZbrQRPsGJGQGioM7
CBk6XhAwEV8dInKXPROG7VGT+XOfoZgWHD9EQdqRsHn9dOBKyAdp7yPLLl7JFIt/
9UiIiml4vG3euA8q/AWMMvaSjnd1Qarlh2ALcH/hDlqkTVTEhgLHt5X4mnq6ErYn
4Z0WdJMSHf+YBM7jtiAUm1N/WMdubC6BKrZYwsJg8ePcy9Z2DGgbWRhBL9Qx+prT
HALwGyhdMwJuthTQha5O1Kyz2v2rOVu1pjOVllL2W5HO1R7MiB2GkrXJgDlx8Wfl
cko4QO2eDSR36arLjqqAmBjNQp6tiJK0+EtuBRR0te8pq5NDXe/AGDuRdhw0N0yb
S8AoJvK/Oa0HQE1OT/+XTskgjU0nXMg18iTuZVeAuWCgwhdcVtMrE1iOkF+RR21p
ADAxqJ2PM5SwZwObUZvqvA1UVY3yrL5K7V5zC/YB2TjMptCNaFKnPsWe7C3oty+o
ZBUHCOiwC42qZ8hXBpMJNaBgFQTRTojtYXyVVWLBNGJOYJirotkT5QaoZLJLQQQO
DY8J6rMcMjr8fbc3X3vjVxpsfQvKlb+1kQ6BemkC/w8vYRrdEmNTOVVDMA1194vI
VFETCzXTYC0GMde6f8ELi7HduLarLzKYJQKld+msqv6gd1GF2NQNdODYAKjPTjvN
bF7EBNMcR5X9dHWssmXbVrBEH+V34t9lngSCjrQHwQ8iRFeZzNhurZ+7B34wzZcF
XhFGCYslTo9GZbZ7wsrRf96brqzc6lovrSRdRUp+Fm/GKEZF0xK1d9Mxe6QUA96Q
cXzsaYb5iIHVO43PYYGkNEvo9PJ8RNIlEsd9BlcawFCzy253YqWarF/QPPfDLk0R
XE/Abpp6Gw6c+sT9AZgFmPHx9lrLv2iVdC2p6ccJVWqlPZy2FNin2soZJNU/euUf
4AuyA3I/BU86iGChipkSWNmltrRuc3DXilMHge2V7qR5A8pxRY9HwNRFhn7xvzTw
Wv1V51d1DOKkV/l1ibMtrQD31c4m3UBb+InUqdJgr7xonyV4/jGB7hWcU7bgGn+A
Xc5zcudd8Dq214ua5DoJA02tdw6FbUqwVFwP9Vj87jUQRxOLJFOiV93A/Do3VWg6
1Sng7m9q04yLqlkhnE2c4AsIl7+pCP51dahf1MQO5YorUohmUCHhPMBT9Slq7nCn
cdIArhmFvx/E2+t190qZrfdwyKL+Tzt0V9eSZHWnnEY/EUQ5dHHbMwGY1+pzluSq
CnTc7bKKuJ9opfr0KqLmTE9NFCpV/NZGm/55dp0a+1g8OU194vFtBZ9vOb6L+lhd
ywIQdGU4r63iwMFTZp300Xc3/db/gG3p13HhZoggqRLyxvDFp+f3OzXn9BJTLeVN
pl/yN+aZgDE+mQnWqZrZQhOGRGRWyZXvr/MnlD0hbEtzQZ8NdOqJ8NTFWi/7tHfS
g7CRDlsvhZ7rLcRDrIAoRV38EI2YYE3B5TXeDGMyRJ8OyG9/FODux1z9KzjStZRx
+rdBUOagJxkdxz0bnjCBTqjUvfejUHBygc+1fKsShs1QU1Mms6/0iRMJIRMPBJYx
e7pmpngUxVoAYNIXphJNvUYZRS/vXPc5r3oUTRRxLjc91HtI7r1MaZ+4rosRQIr/
xE/pPIWWCU10lbnqUonAa0YepBa7igk/nvGGbk0Ub6l4mwmgH+GPNS8zEHkwPDSm
+67Ky8UozlppvqSftqSDiLHYBOz61yXJP1PbViQG05v57Gl29g7QqEd0aONE31KK
uycKHHW0N9pDmYEnVNPmX21sJXk/iAALKSC1qjL4LJfgkpvz0mzfsve/pBqB9mTQ
1nsE5C4KRclGR7x/PI+iKYXYT3GLv1vinvJI/l5fCI9VPnIDfW5Bh63v1R/qSv7A
Uppr1+wAxInlXez1xZLCvaHGuXXGZainPqv0/VrsE/I5dF/BV3c8PN83/Ng88Wjq
Iw5EFkWn0Yg0zg2mpl6IP2G67sz7RA6cVkNkr7zzow4bBDXlv99Cp5FtVY8M2i46
EXl17L6hUxZMPnzCLP69YX3vrbHibULzS1I4zKdziXTfjtT/qCnMCdDYql9DQG3V
/I+tralEQL/c5wSk61imkbrTcdKLzWR1Xdoh80OqqKvGC7o1kcPCCiOfHcpVWWyP
V0kmkMZ+IrmIt3H7/2x6kqZPuBXIzTiyT4BbjGzDTK72gzOph48F/B5IrrJKFRZF
lto+3ZswjyLNEyA10e6210EMpdrBZq6+Fhul1PiurJJAf5crq7xrmKyTmB3OcXXg
zmwmjuuoIEcSx/aSWFJ/cRsBdIfZXfPuHH6hh1XcjHxvtFk8Z7Mvjw/Y+2T+jYyl
HtomROaZlgnB3bjdEvhtZW01qQsBVNrPj30gyfHj7hVi7NX5h/d4Yjm65S+kC7/f
lzPAfe/CsGyhgndI11PcNzD0siA9RdoCsCH2VD+nbwkyNRG+UzRCFa9WgfGV5vkO
jWqw4i6u8NCsBfFkih7jicqHKVbsypW3jmmzEN4OqBWzNQUeWf/tuHlswWQcr8kj
WLFIMdaxzUYkY1blxevffdDovNrMVECjibBe7FYqL2w3Isvz7P5BhMFnlmheKBBl
KLDUw8TOBM0CcrEvEF82JpAKSEK0J/OeplhYbekTb5/aL8g36ZwO7HDLz1mbEJp3
AYNh4fNaHYUIMqHJtCS1AtPt5TjkGp2hI93NnYPfAEUj5nG4ij7ewUJ9MT6bCCin
8ZK7gx9w10eh8St57nXxDyADQpYzI1KzMsQ3E5OaVjixpSJBb3ZSOBsb+VRdAADh
dK7BhSAChVqZcWOp9J7fWikiLdD4gVKposfQ/Q1LfZawt3z23iY9Gyi2VTWKTUVp
IDldq86sSk3nrk4k0n7ZAAoUfUyKzFU85iUoo08Xdwtq5xhrC7CKynb2QPg9gSDA
Ru/jH09TV2qMQ2DV1/5HZFaSVSko7WvOGb03G1ga/yu+9vwUvc7xSAfAIDEgOhF4
+XfyYVqojg9YngXVQxOsWEIv1uhN6or2wxXZZ3cfuog2EYBTtSbABvc9OgOKGjJH
Nv2QmANkcyg98h44+DZhzXpgBzgKY2ydBt/jwc4UR+d27X/Tvz6Y2aRsUfPE5TOk
xLrGAdLmJI0fODK3cbn0lhESQH1ErgnsJrupcOo9pOdiDSjXfE2OLuVRrPLvR2Mt
c1gQ3VQ7DOHUuAtH0HwlX2dZRjeoBdJ9trSfGgwVvyHuan0dYpR3FViIoONbZoMb
q8Rk6FHUMKmTA0DPl2fU/HSaJ64f8Z1jHQ8Ypz/QjcBwU5xYEv1VzXxw4wgb8I3w
+bLc5uSeYkKtI02wi7Hp8S6FeA5AT9N7gcr3Eq9QLVbOPC0bxcQi6Z+qHh1+XqxC
ND+owun0r9J/7BqA/a8MQ9MXu9gH1USFRTfzqaOacIW6V5wmlPtN1uhH88UAIHx5
8P3yTu1zMvQ3OwJzLv6YnRShGdwt8dKUz+Kak7srImZUhCXTPMhUboWJMAIniaGU
/qQZaLgqEn2d82576ai0MUtAc+IbUb7qL+21+tZSToiN8A5cZA8fjF2q8fq7hALC
dM/lA7YhIDQYrU+FCmFdwXHn4WzMqOWU1H3NugW+tcKem2fRALTZDFbqhr0kdRMD
nlFvWe1Ne4ZBlamHWE5qA3Aae6zAZ2G3A5uRLcbpTIz3O4B5aEba6gh3G6K+QVCe
Cf8q1mU/VgDR2Gurj0uAa+0toYDdgzaSZvFkRct22RYfhA2nBm0suAY9y9zYXc9c
kyEjTYqP7zCpGY1l8pYyx0ZLdkJC1Bc51ovlxHFUEJoH2fTGCCaYtwMgwFPqH4dC
mcLC9KV88LpTVovY19GGnwiFgJ0FGVuAqvSiugXE5RZ3eDiaFPdeeTLj3WKLkRG2
s2dvDi9/Rg5AtoRsKH2TUOLNGFA+iGJ9atQ2iHA7wZLLsasC6+lcH+Igkfa4Rxk/
U7UmKsB4GG/AtSM+kwoT3gIs96dCkCrMllqsbAsUQ15WsZINiuv+GR0WoCOy8xi3
tdbFphofwFJWqmXYbS7Y9S01GPgOJxrWhek9KXgY6/NKHYL65KQq9PO2SHtUe096
/skvVK/AdMkfrHjyRZgiEeVA5eRr7SDEY0T5Cdtz/NwQ7dgJLM7Ro8DuNXZo/25R
d6hiopTJhChGcKiKBr4u/LBYuQoTXiRukdKHHAk5u3ZCJklBee2P0qrP1Lhx/bw7
NRbBD0wDcD0GUtkzxJvWDbZmBKXWgsML/6T6v2WLaS6OfEbs9nLe21Q2nI/9f1Ue
CL18AUcf3Y9qg6SlxZvgajjrzrrn4qKXQaC9GGw5zJ48Jz3fcuIJ9d7SGtfChztY
IejeqAvFCmG+RP7bPdGmu3QO98mWlCAfl5ZzbJvrOki1RctBMPT75naQjc/FbxMc
kE04OAyD7mb23mIBfS+JjjkV6z8ZX4VgKjGF3kolkhUOxrFrU3NVxstZH6jjpECD
saU+SLITgPS2bKsN9JZcQ5MSgAaNS2QKW7oy+XMDAgtGYHzbqb8BNJG/ZRjQfTOS
koHIYx6StYYr7UNvJMs1g0B0Sty26JPUlmHjmrMuv+3jrzy55t3rL64LkPXerxRX
oFLEqUkiqIGUv3yC5gJmzBaaHbOinnlFaVZwv5lYii+awIlx+zqY2zqdKrWhWWyC
Y70zTaxv3FUHwvCjvZJVRSeK9ADRKOFrUx0VWBI29LEYKbxmasGm3IgfXL01Dk9A
vbi0UeiGppWNUrrjDvBiP7E1WrGZsvkQpRaaHBHdL1t1l+qUfXSa7Utuc/F5S2LV
Bk8AOik3LnpxhYVGZ8KwDG/LdID3wzfI5verimgRbV3TXqA+pCOBWVdcCec3UM0Z
DGgA1wtRT8rfvXmJDNWu30WKdAHAT2lZcJK1dVDnM1BNYgM/taxNWQ1PewLkjcUG
Dm2ElypX7PDhj8vq6AldCjrrH+rAegehTZX3tAZJ2i3W/G06Ciswb69P6A6fIaUd
bNALqqzzcZS+I2OoQVaA+WcDnusN+zx/MRRSDmtjH6lvN8/F9zJhjGsXYHJ2BZ83
UAsxihuM4+lIvxIkfhgxiO6Q191uFp6hNGf/IfZs6JobtgEkoI8JjDzJsgwKxMbp
z5blmOZD+oKLM3pzZ1gaHBbjIFmcwhGDTqoeTOhcY+vNfWDyXQtnRLWOn/4Tg3Xr
nVk/gipCPaEccnrnspu+jFPtVY+ygvOejFZ6LGMJep6JbfpMASXXv5XAq8dKy7TJ
Q2LttkS10i0e3EvJk/VZOOIPJz3ZTFIaez1yoO6TcFjUUEGoHVWSrkX/YgdiZwqC
XdeNeR0FeBhEkR6Kv9UHPtwJPHzDq80mFaP/iu7sLSgbQwU7p6SgcrsZqQ8e3/ax
z4KOrfwUZKfVYKV+d0+5k7/LVh8Ff8+lHNxd4TCevbxqOfh/NvLGHHC5h26T3Jhe
6lOa0D65AwqdDXoswUje0QjT17b00Ysixz6/UiF5r9Be+t0Pl6rDHL+D0lfInFvQ
QyJqEKc9dojpMbd2PfPfiu+1tVEOMju9WI4qgm4uujmW+0md3mWhKC0Y9zB1jt7E
kVOaIDnm9YZ7HbLs6CylZDxlr/6NFVFlVC19sW3bEdkNBGAB7ScG4yfUtr9Hy6li
aPdOCW0AgM/+lQWb25lNjA7dOvBnSpp6UX//VQvlU8bdch4v1qUtPn0WjMq8ckEd
XYfXo7iYKct3EWG4/qwftxBldv3ufxPIofOvEPE038GDlZq3JFiXEyk9skYhAu6j
RQs5vEsRnCIFwXGCB4x8pgcuC+ODxADyJRLJkNUxcUxWfaSI0Xxx88cVLkKNwbrS
TAn3DHHWUtq+HPDpAdndjn+P8jRax9sa2WWGG8POboyMOdnkKGUD1K6WjqCoug88
QbP2O8uDC4MJgOwHdZ5imWiJ+faPCGKidXMGJ7ICEswMKfDKe0O+5rWmi/Yuifv2
kS7F2Ro+e8oPTKHd3rw8oLao/7NLMuUn5YGTLz6AAr9t0Cs/LkjFJjpEMpY84B72
w5sU0nLykc5hlihoS8gXrnlgVbziJNclBQiz2wrfGY0p4uWj+/ORq5ccYDy6X6ng
BBJLD7lCXxkE7G9R9WyjQXhP4LZxzfRDa+Co2CTg7sdBXDfqOcq8p0vxHZOTZpTQ
1ohuXKy/ezuWy4ZAFKVlaqQL+kjAqYA0dGhJ8cZqxw5DdqKmMGYl7JXbULI4CTSS
dKinmPMTywJUcuNHV8Sd0o0RD/Ffz+to4Z4FpPvLZ1C3IzdwPDrvRQGKmn6moDNi
J2eWbHGiiFAl35rWaOYuDylrLvoPNskvp8QHu+EB4sTJmer2k5HfPHjIjNYY0256
wzqRlYGQkVMf8s0+2lYuxREPHp662k36E29jVo4T5NUH59fC9/pNPWMcXmyHMJlK
ATVqcoi1Dk4XhwV6P5R1K8P2fESA22duph/C8BNoU7OTfxhdxehAP64dDUqS3M71
Wt20sZgoT47szhujfZT5mMnlRvcRbnRd6SCbj5I1K5sWHOrk2q8HVjI37AivY48R
Ma5wIVgWGt6RDVhLLKwEUIDxO2pZElxa8VxxM9UxwbEintafneEsPkCIGeEktywp
jgri3eOHIjP14C5Eo/ogaSQMyfaSKuuGroJDqvYpI8vfch5teHNpKMelljhcQQPb
F+nbhuHy+uzVQv9bwwAasa+G40v1n7EjfmTrfOa8bUvLHTWQ5yfxaEVogdRdjTC8
/B0tBwN6CHREmi1yCkygfY0AyOVboGtYSerSK+K0FHQCze/RvoDs2CZ55iEPj2S1
6u+6uQR9hl9xb8aqlhNkGJ8Acjfq3wZg6vxMtgj/IUbpy5w5aVTIWaEz2PzfJ6B6
Bj2Zpp08uRuaPg4sJK8Oxs/QXIBwWwSmhvlffjW+jj26z4GFUrbx9ncO+NBxyT8Z
J9WR7/TBATsVZT1WTX1AnOcjwzMzzUG9vB7nYId6i+KnM6GJAQy52QEIAnNxcLfI
1HvRLzTjjwjO3tZ7pGugVEBysykr2LUKjIiaOpaJQ1fD5I27hocrz4lrEg1ALGqr
CYvdi6DF3eMU8vFxZB9YNDnYeJNCB3fgTkQ7NdvOrdKMhy4GHBZkfIOlolUyLFCE
ek3xpzUhSw4AZbA6vJA+s5oSLJ7cPdLrULGBngDjf0jTakEFchGR6PBtyBKHTS20
8SezgCm8bbe6LJrHAGpI8ULORk4v2F8x+GR5DCjeoyom9RzY7y80vUSW0sU0wr3C
KFa4qD77iN9tQNXUPp9Yk9o/rQqN5zKDRHOMPvOuzREjoOIhoH/VpRZYza7x5AG7
HHNpioR8WRgW8qBkc1sHdeikHWvj+tZp35oONLefnMrHFIW/XahuL9fBClPQLXvp
/TRqWfTzS7N+oyblAo4JLQxKPLIxAS5t8MWbw5dO5vzVX1j62Pxp+tKbN5//ymGh
kFPuEsFQfeplTK0b6i90M2b5TT3u/XVZW2lwcKwJ4iwmXhWiGJ3+Lg45a4y+t9Kj
ioh8aK5FjWOfHjYQBBOUryGYdedU0B0serlMB19tX/vcYZFP2FGgLw3Ot3LbvSIV
Oq7SIOcO1/bK+skzX3elc4qM+YW0XZn4U1zRnC+NOLODkEVDLRfw7RkJ46St51aJ
YP3fCLnm+bAFXCeEd7FKq1ENArN0/D4+fAD4jmciXHWf2MmxI0FtHn0tnpTLzbtP
90jTh9fEk8EhxESAWDeEDbl8H8QMfAXVWXzs2dgfGzJdFA7O/CCeyIYs2S9OV7uJ
9TqyuXZ50nQ6F5C4OzQvNFBJvcJ1Zi9gt1d3rBR/tdrCgTIvJfn1+MpTFzENeoEL
mdwrnToUTJniCBB1PO3qEZ2xp2iDm0BR1m90ZRD3WnbZ5j5PTBft/3OBXYxP3fmA
Pe+ugN0WPai6XAdr5dYvLwS/L+QTC+kvH2wPtAUFCSKpXFt6KbMDD6mVuZqWCawb
obAHdeXkWYMRQOSr2aklu3Gm6brXgf5NpCtpDObYNLpWdZr6OuEBPAw/oEE9KUYR
uJGC2uEjpIxnSr68fxFNnqEAA8AWrWfAq7NzjdNqUFuVPnMCI8tmTnS/CaFPepWp
gQ1Tkv1oZWPXDQxFqBoiTlHjhpeycYwcY2yFf4NK2fRfDwMMYYiHRGDcjOtD7Eey
w0kSRiQMOUADYfuyGHPmktWl83IqTSAJ5esFPiBh423a69+AA68tsjDFIPFCzAxY
/NANWMoma7wQdRwkBY/NawV6I1ek+i97mcQPpcYJKRjQzHQVuDvq0rtnyBNwYHWi
eThl4mnkk3c5ZynDuEcAv8ClmETWPLLE/8/rv8dlBCwf7VGcIRs3upstPyw9GmTZ
fd3jtwUwanDoOSr4qtLMRR32xDh01nXSKTVe8ims3FXYdEDWhamqyx9LLz+9QMdK
SOQkxoNHC3NUyn7ed/4ub0Aes+ObTei5d16uJSwBcVZy4sXBJis7+R6ge8aSUo8T
Nv0I/XCWg3kwtIKeEPsxuQu4vdl4ClGJaUXAJcdGrbVj9QWDJKpP+v6jOUKmrBvC
Xc7Az8M+kpKJP7MfS3eDWdAyE4R20VRpL9oDyOXD0YVGOCenvrjwFaRJybID205+
gfaLQUwGGFkcNkwYTMo5Clc8X7Soa+S44DLGsVUsTU0PMdSnHzdr+/WBtlVtcGgk
G5vQi9uw1fp/qySw5LTyoTshrwix/cGOY9W6b7zd2gY58UYyC4NaNJ9seaRTMc8E
Y4yB6qjgO2tnKDOTY7aLsod+J5Liv3b9pkbQ88BrP6WnGPkfIUs7wds+MeBqeNJ7
ICKKPpkKn4FYby61H2yFiaQUNeIyhx0e9DwhzuxRb40cS0IuZrym9qOmzEElZHk7
ELyuywtE6F0mmNnSd1GI7ln+BrN4N+M0a4gDzHFYeUF2Z461LgJOFuguVPvnzx/y
+KauDDO5O8jT5HJrPf8XJi/W82tVAHMQcMqQT46Nm4RAueBny+g9aJ0W2aVuYNEu
U1syVr/V/80N/Jvd1W+4caaMI6CVKwNVuahUqMz4h9tM/hPxiLGFLndrfD8sPy0z
xP7s20UtsLu6nfKRdJNnFx6NWrA34pFN7fOSO1Qg2tyopmFbJAdiC6k3ANb44EC4
x+V2RpNmL8PhpG/yba0InvyTwKdSA9+h0tq5BheANpH2R/75MDVl1x4fwDy5QWw9
/7HnMJbBzCCy1xgAM7RWQ1G0a8j70ypnyAJ81jYHoYLUIPf9+e7K0OPtmNDzhZLQ
ZpkKDmwIn9id9gAYs93m2Ahqi8lJWf3gLb8uqpk1aGfcF82t8VcJbDFjbvM/dpUk
xR6yjr7buwcOt7dUgArOicudIBSfTYmWS+UyXer2z530ubHnGV4Pa/U4HHgfBYVY
ewa3muTMbmufwXw7tRWv/mmZfPba3d9G7VKrIoEAM4My32Sb8pXTUwT8P+2eKU/I
LWeUwM8zWMJZcbbnoo4NygAz3trAMat2wCAWqCfP89uAbqz8hYpMSm7CxZIO+0VI
6lbFgpHeTOGSm77V+qXmqM48kocisa6B/ytJ9FmCPt0jFuv51+/TthJ+Ye4PRYUS
Xj6JENAdZCfiBKKY4dk85I5fX46z7sGZpRyC/Sv4TYQ5H5pTMLjvyJD/2YCk2gk7
GVwpoMo+49wIO/tZnEpbbJjuoJ+esFnwEcTfykoKAhR5+UBwA89V8hEoPPxJFvKi
4/fhegyK91IAYLb5R2uREARHE6l/+sojkErJ0cnVdKqPq9ydfMIZXvwUJKC3/P6n
78RQlWk/PAdL9mbtpNYNEtJgWGJ0JBaIJeMDpUphVgQbAdO1MaPtnnVTXWf88tAI
ioedKvWSvNcjjPdVvvHrNTSXyh8Ti9HDgWE4oWS3fD0TIUPyOyc2ZdHexMPfFxap
vFjm+7jYuLBe782rsevr/ZzGYRfZi5xGn64Bh1OuqjlwNhj86y1QowsQhzM029Fj
8cttDxcDfWvfjwBKoaDzPKzxq5IqAHHPVR0Hr6QT2knI47VXXMed+9SPaoOCQnwJ
6SswTOLKZJtbtwc5b3bPWi+5m6xzI7HUPw4FVW6vqnapOsIaHQ9IJFlCNyy+vsUd
YLx0Jt0pkePJJ5yzJgG/Y54QWFV0e90uUh2HMQAGP8Gq6szpxlJq0HhITj/C8WLk
QFB8qPCS4S/fRJnnAwpWtbRFnMk/G9OzNNLYs1vyBf5gKX4Y62OR0mLKBmNkDvuC
tEEGHGSYXoO7h8ve8Dlv9fvKM1PfRSTDggv0TiAAKqDLlt4/zE/sZb7rAWkTZxdm
27kC2kPVjh70KsXOE90R0JaaD2xyvfqthuV4e92cp/rfPH3aYQZ1BVPELrYwSkr1
X4zvHFLxMzvM40VXCxG4NWvvUX9SwgnNxXdl9dA1zxbEv1+tFxeAXtIodpUtii1i
JdYvZOoQcrwtVGVTfDIV/E3C1yZM6R+4siIlqq1K839a8MBg91HCfkEqjiNaKJT/
5cUzkzZ8GfJBmD9gCYJhtVyevM796hUl/Bf1UXULg4v6pllLwoAkY8wcH0uAkXRf
9+L6bHcXPzxtCkRJtelYkfafo7IdVxNoTecV4+6KMjYK14pxJS6Zc9pyskhlohje
YNpmC8gw4Ohqw7aFAUWqSVrNOEsdQP46dSutBrMFvSlSBG581AtwszhZcdK19Li3
yJCr0fIgLQuGfvepb2Gckyz2E21Rq9ROTa3RcGEj/4ykP31m3LhUON4rK6TkvPO3
bg6skBJedSAVL7ULhNqQczA+CsOjLFWdCV6I1jzC62/KKSWlFhTCR4qcHowkfgsQ
I5lo2RXC0tD8b5WoV1gthuicLWm6k7MrFRYGfqz3/silAcw+p0qK0vaIew9XEBj8
o+yGVOoqVjLnIK01gkJZSyFSAOHgCCvsuV64rzrZSQr2bsGjD1aJj4iWqHBdBrk7
cTKxF0HQs8s0fqvBHzWZbQVeCc5a/R93zSyvXR9jaMtWnnk8SE34OKH3JlDwk7dF
tMyEtIhzqD6KDbYpmGIE1NeU5PfWdKVCoa7ttUd4RgQotrv9H9fiCu+j1tbq2IQp
hMVzfuc/phu1kVaHJqDqWjVpguCk2vxNmJHGAx61CWIldeXm6geqQLq/FzhIONv9
heGgJhwvvAe38ZIryrieIQc0fI5LJn6RG05RLmQOp6P7rtX36QMEZJ1zh8Eamlkm
wu74wQkWNl6dDc6bHOtTg/w0SYEYWUrJuftIZu6BiYsEc1GuGaiOHrHJgG+Quoad
gKSowSienfPNJuej8vRm1qDwO8PGR3hJ5ByU9F/ch99MAVW4NaqbtcNs1uv1F+wI
2ghRfjZqlPHtuUygx/OzZah6IFoiifk8XEIM6NhWwUV6aMvdQFfl8h/ALk9pWbRP
4iFzuHb6mkIdYw9Pgyl/4NqgkiXm/lKa2T9eWY062fjU8RhOXRQpQQ+8xkb1LKHn
b1/+za/wNY9XortT3BOAd8szLXRHN/+84wwh/HHd+4ugfV9S3za+fcwYXqyTSeSd
uWEJN8iUQXDVB3aNboCBIValbBKY/bwQjhvFEHJnHXdOXduHps3JHn2QQ8mB7UEi
60YHrc7Wfyn+juihyOIogDgZuTfkC6Vsz6kqiiPEzPDV1mvPQ4pxZADEnmfHs1Vq
cyZPyFU1y3dmkSUEtY4kFKs5bdcoEt/W2A3nGoXIDcgf+/hLjnUf/k0EAnm6LdZ+
+Vz1CanouK94p6+D11Z+29sqMQL/Tfoe1QRFdrFmyZIgMyktS5Sq8saoGmAgJhgY
GB1y0fvkWnvYd/ZmUxN8N/MnSR6r2GUAkuX3UGIwfh/+LAJQTT4LeDaimXexRI7U
ikSoA7nYKq99DyqrhD31jfJ0cpF9qnNEaTUZ05nk1v5m1pIY6XI4UYmN75640gYh
2SkNI44jnUEyMT0zwb4wi93hBrQDWO61381KEK+oo1iaqvbtrrgGK4llVbpFGn3V
FBtqUfyFbGVj8uz4dhxwbsQ9pQNHRZTKiYnoSM5NLQExAp9sjbWHk/ycOVBdGGQ4
V3vpzN4S79pO2y2TK60rRpH0EvqlmadAHiQaQN81+527gv7Wec9fsTbg1rcdZDfw
QK8GSiPjmG0mwzxM4EHMBhIEBTBuik6+mXho5TjlB3gIuAs5ADvwBCboPw2eu6kb
flvLeVIjUmvxChKXxi4Tth5UWyylwn7BaBaS8AxmRjVwozZP0osdIoVqZim0yLGC
CRKe0msA7MPhKrn2CKZ0aa6UtvQ0Ud5Qmowotk0JpQelfg5LsjL4zn4agRbG/O2s
oYurQcj+i7HLR6IULacZ7Pk43JKcqQUc+JewN17WdmdIHwqEzNDjW+8QwIv8xihN
LXDCTYsJ7LE7uTljdckCNIHxWX5XmJYZaWJLNDSE7EqCRHYbreNNcNXLlo1USamG
bJkESwaZPURps8LtqGLkZkMisWhwIABRA2jNp4fx9zOf2HThwFaNY9QDRNuex6xj
zEo2GLecSR7UBs3qEAqn58KJRVgOmHA6Hq9iKfz+bcRdWraJFI1hKLA9Y1mv1gY0
Y5vWJJuHzzAKuddXLJDheD1ZUiSL+0ULIDQ8SvBfSnI8VJLEAmvbqu9Gjyxo+Yt3
87vd1FfQPwUR2K72A9ltlyBYTejnVMNQkItxkHK4aKKMedLXv15Yyu9mFSH3mvFU
qlenDuvJYdkQ9IAKziRZKycnnqIWNCEmUshkmeB0wIbCwg8adkLQdcqYBR3BUWVA
0/QZYcXE65FpvOchqJgm/umUYr99ufyLcNl/yjxn31/lj1WNoCz9KPKGhDrhRB4r
otILteQoyQ4uSOUbmnQmMtxvapfterQE0nLQDKONxSYwl1YEt4GUHRgq7f38rrq2
rXdTuymlK4gMTF1wJTFyoixOMlCBFt4BZ8irtTBeys7yK9ZGqk06/VDDTu29ObF5
obXpe2oN33D+FbhSIKibUsmtvBuP2FwmrIFVeTbPNxesUhA5JMSfDIW4X9TMJ8C9
uun0Tg6i0H/5mY7wY6gdTubMo35tsH0jBRWphVNgb4F0MZs3y4Ytsi9BK4balJ5N
UeVxrxxct3gaSXcTfxkaMgm19+YLeAHQFeMl0XHj6KoyZIlb3RXMzTtG/svtOAl8
FJpGqD5M9B76/VO/VNDGIimXgz54FktUmJFuzxNRIDbCR8JiqXBMBECX82KM77Hz
HR59hlabZGnAZd+PZyeIX8l0QQsi/VNbRdTYItJHbAgg0QRR4BFtwS9T1kqaByQE
fIwpDha0ML4o7wANWq5Z3N6NzSCO9qz1i+Kbp2Fy6SaLA3zvPAJ+Ageik/JCz2sF
bYPaOhb+CNBQgfeUNrtDpdHSw2/XOaKsg6co2WYG+o9PhzHZjRK/vpW9k3AMLvAP
6dH2dpzFdY25wpLSzwO8crSLj1LJMFXaLNFvoqRVh3V7EgBVGwhanKga4z8dqTQm
z98HUaZ1cNYPhVB3DtorpWuf7zQUQDmtvL4QKIfUi5nRJJPdU999LgmVDvwY0P77
aaS8+rpoeJZYbLASSpIM1yYGLFlJUXJiCNyBF/GCtM0++VY40QPLKG2j3paqanx8
0Iy/EBs1PuLpDCVagLSKQ30AK9NKGoBCYCviggRQto8P9BtSKUCPJgbXnkac/LK1
JawToyQCC2eblF2RxdPXutUbzqQzf/4Vr6WaRw/PXM3LTjoZndm+i1Zvnz900+Au
ejXqT727GP5GoVYt1bYDhsfC0nMttWfVTI+CDctgkqU6JLFWmWYPemMDYPkK0XPe
GKN6VNZesc6XioMTFDVn4c/TGBzHkeerZ0A7OTQZvECbs5TcmZDbuP1kQACN1v74
lpvNJfhRhnSywQ7lsTezygUDla+61ZVG1ugUI6Ji1Mvu62O6eFonJfHt5O0zMnNO
JBdVGQdYurPu5dWicp78Y6RxVGHI7po/ffoNpaVClq9yp8G3TTlrK4evkdxe0SJS
dTXjGQlOP2gYxdENq4PWhTZZqqyoWgdb1lg/UWG05m30Ob6QjQ3KrgAfEZDju1LO
y7uUDy/BhylkvprwMj9QLXxbl/tf4MeAxDUOAEVFMlA+HWC1cXnkhzmm9pfN3BuH
h104TkNLMdRxzW+KpZfurXbVJ3nyK1RTvRrG8vggkgY4RSJw35quiSXC5Lhy3gLG
xkNmrkLCNaMAbfRz/5BDQAjEM+yfCG5OkUyVEhrXUWoL7WFzHtNB1wcKCJMwKeoR
Ba5HIbnSZRR7+L+/ou2WY/S/gNlgedPWMiaR9lu0djGJs3YYCf78onkiE9PmjrXY
CZQsmAmCfslQiU5wg6AQUI4JhUV+v58vqgvEWWt1rcWokDYdQBgRLnSwKikGDiU1
P44d5By3Ghc0yBwKm8iUQPvqZOiql6qZRI7K7pK0Wh/LCwGrLzSyTOZ2b1sPct5x
/SYptVkarTjVmHQV40bOTxTdjWioVnktM2hHpgrhR0v88BLLOYkJv6MKGXDqksNt
5IFcDzCqjjj6BK1TZR/PmkHcHLMgZrOKft9SIz49P5DFITpjA8h1POZ5FL9n3mzk
aKM41QD3mauYzJ2eIVprTYcXWVwtbxxYuPL/IHggqV+GLuhIHaYhTbQsfLsadxPy
NwkRl9fFat80N7ECx1MLrZA3ZxH90k1MLMtkw0bMA/cSNIt4AxTe9aAoShol2XRE
dSWpFgTeKTTTYAqE2WFwT6o3nP805aR/GNBuHJFDemDVyPpFPvXJ9y2say6HcxPL
Iq5DKHV76xX2dheLH7kHeZPGk63uhMpmInh39gKeOAAKhI92gyimnxkhnrw8+nMe
H4cFDH+mXZwLQsOcXjVNBoA/STGGgFk+COtb3l+EcHNp1YP601QsfC+RSSyyg4QE
3X5H4mJNEwJ1qu5rfDVH6ou2D2vYW34kgxYlWDmMCn8OfBBOSfUpF1WnuPwgxXKG
GLmAVs+KQTPuU8GyATRvpbi6pRQK5g3OkaUA8/z0oVVL4iP+FBNKmpY4wbySjRCN
O17KcCrG8Hmi2CTT2Iiw3QEFQ3ggFA6BFrEOM4Q8Vj1hvBzBbXLLQHY6D27ogjtY
oqtarLM3kXgB4izrgQZtOWHdk54IFcqrLpN/nFEBlsZF0P0nEXxQK5gyBZvx2+PS
yBJzIBoca+p5UwgyJEV0IiEWDRNZz1NGzYHaD/JF7zkoUcHCO0Sry5VSFJAYjT+Y
pdVMOeEHjukIlhfHT6qkZZfbHwgkdpiKLTVZGtVhLMovOL8eifzwrC5hYbqSv21n
Dy2ZJnIsyC2SESZ4lahX/T4q80kgs8X7XwimY4KrNMihqeB9ygBJOT0Ry+EC9QI/
jFiNiba5A8lOAqyO8Ae9cZSz1InFW+3zWqExDnvauqcS5UoX+bWydxXAsiva9n/1
6L7EzzAKfdiYDaCquKPfU+3HycJYGJSWTvo0y5j5U0nTdjaCWjbb4IqqZYKyijXe
wXEMaDMbl2CKvn3/2yrWZCCaWwzKXySUff6nCBSHvvyeP5OAw9ruDEmLcTvxhI4N
dVx5/aSgPCSwl3mkDfSXHvD9q+YZkYBF0FkkalperJLIyli2j5hcPUVB1P7ZjCKG
9OS6rXeD75OZWnjxq6g2PsHE6A+D9DCOaOzVVuHuJ8HtcFIkEcS1T3i+xk1A1UZy
Ia6zQSeHb1T2TtdukIk9DbxCEtcH4B2OhlV7NgTC/SMZEEWP6jH/Z+Jn1c2hjKq/
ZzeKxtD7QK+sjnljCCjJh7Rmdbs8t1kED+aZ0LMlQPwI2/Agh6ztp1V4z+erNDXA
4kEygWZJU46LTzc88K0/wB1Lu47CKzuFF40FkOmSchvuXOmPsBKSOwKjytxoGuyg
ih7xZmkP+4UNZJbSAg1B73b4aioAGEomO7QMmEH2ORSVrN8hHdD7H4VeT2kOnoGq
Z+1l+jKQeB4lm2s3t431exSYIRTAMz8O1GfoOcVxISaGCWMJztxHJS8MRqNZzFe2
ams9pe92wmE95s4jiwG/XZ8ping1YDG1R9iLhSKTuS2YcinqDV3gKeierAd0PtSr
NFbXRmO9NaaO0G72j8hHfzKwOvQiR5tjuh78QrYw2Bxp5lQZYl8pH+3XChM/LUdm
9iYHTHawyhaJ1pzkXgk41SzLE8BC8vwDBj4lbP+FxBZ756xirvRB+9EithRav1qC
QLJFQj7iDyaKrqtUGyuZ+yW4LSG3QnYD/ZDVpj7pvV1hWRTnuVBHyvH5QCOF9aPt
+e/nnzvoFH1cjeELpSrHN+5syIwHnCMv+Fo95IFMFAU9p/zAozUAKfas/75WKfCx
FvS7X529SbBIyMVdwCohHGHNcpb49d+TM9yjyazIn8kcVRKHML8qY/HR05CZ+Ot+
ZUC/5BfwPl9sQq69YKoqiglQqndbMellPdWxRp9YRgKWP2USAtuNxSHGvews0Vdt
yn0ddgCf18KESE14gk2180eWbpC4eQg4MwDkgP37A4cGuX7ESQZPKns+mYKNk5Jg
RkDLb+YE0I3q5V4lHTKnaO6JYsrpZN1YQRLvpoJjH92eA8nBg743adeTgHT6rnum
Zb7mPygl4Y/+yqVPDHNZmMv2diSIJqCq5d6pEGoieeKYuhcTeOcl28y+mcp4ulGx
+FHxAGFQv71su/DJtuAjUFJVBta+9XNzMjsUuMJyec+k9Zel3CLug0DunSy+XA2O
iHueQMnjgUmliCrAvPbhc7s8fSo+fm12iYFf+tgO2cuMsrmzDoPs+1br9jS0sqeW
/ZvK684aR+S+KSuwHA0LYbWJreJCJ4Cxq9r7fVFAsINsDXcijuxSIIB0zopultd3
sjEY7+lfhDUix6DRSuussnB05rkPW8jSZ6YV/UXOpsX4JFABxLggINQK6vj16aVu
tRQFhVsUyT8e7Cgb2N16k06AjQVVhMb8qgRLVksrPgDQHyyiLCI1EQUpdjkpiKfH
8Ui9wd5DlNrUi/Ehau3VublFKd/6fJUr4jUKmXvKnnBy/qjKoJHc/XET+8jyRt2c
Atu/xqIw6pqZtz4d8A/7xqGjV7jAqq4yz4RZIJr9346EZfJjmrzga3UIpaCzQ//d
sRNcLpDnLbST1DSv3/jalxnoNA5arFQ6a/McRTuKbsGCW6pPBiPOwPONSp8qmfsE
9dcG6dvvRVNb/Ey8K/kszfR8/j2yp0wP0w2Hn4QEY043ooID7QQmeVgoiQIavQ7N
1YC+zDqxx2nLYKMzFc4f9syy6IWJdrEdfOHFj8tL4BNaENYnOJNI0Ds7hE7QgmGg
R6XBlOYFMJ9/q+7dVks7SwK1XNQEl60HXitkcq7tn62aX6aEtp3FSDnkQoA1zfSF
pjo8+WGBT2Jul08qud8euZJA98Wa3C92awi/rD5rfdBXqVaFklUJIq2ucuWgUbTG
cBSB/nLYot9s072+Ym28ETQh1G6hghE3U6TINNQfJarLfiYC/lB+c9qzG4iy5FMz
CVFeAWgrjOWwnN7aSUcAc1ILuDYgjpyoCW6NXRVkzt9rfK5BqaaY05ixcFJEe16J
kVP50LjXBCkGS2/nMGLFjJUvtW2/gIVMo7pWcsEZ7uKJsTkP3uU8iIsQPRNs4gy0
ym4WaPz/G0hi6frH749HoABKeQ3MnbNlnldqZPIpvv7VDks4+vQchkLND9Swx5i6
vknfxdJmyoWxb0BrAYP7maawb2LTOdzz05iTY8f8UjiTZGQVN/eVsqcqkUOsF4S+
b32I9vsDtO/ZDoo50cwj2sfqLxWepAhtGr8hitfhWDY+1aBmDTWCGp/8Uh7tKYBZ
X5pnP62UgKF/u4JK5BlCz3Ip6o7bzDJ3OZuRtnCSS6s6FfmVhUIEognJPpMHibwo
6WMFyYDLYtFWFR1mDknHzUPdfZCneAa5RPTnVCRWu6NyBQ6c467rx8zOUUz+DZy8
idUZhvHJn9Oc/8eS3LufG+ZY3ejqT3B+BkY1KG3MteIknAlPLV47EC+JTzWQB/bF
JdaW4wM/pOINZhdG7RC9odeIr+QB/PCa9LTa67gNz7IcJ9W/S+dHd3f5mHKLhv3h
PdxPCiLQnfwF9fJ8FW9vcFxn2197esnNCh8wDmhNO9zosDgN9soqv6Y5ESKQ/HD+
JfXdo0sXSJJLvDBhLkmS58Yi1Lk0iWGx8w8+Mx/qAtMJJiY+b4ZcTryk3MvEdCGX
zwMb0dlb9FBdwwSsvSvaQZJLbXZxZPoQPbF+H8IZ/DX1CyLgWGZO66bwLSOexeb2
XxHAnWavwSs+l/0BtSrEx3euZhk3WhirxzKgDEeylQEdIEZgE++5k3QskKGJP5B/
y9By4DvtPQtS5sJMUPgm8WKEMuf3OQ1ddHmK6vEK/GH//eGYgtDvZfyOhm3wbiph
dzcaOd4xL9s2Fd69yejwxiHhVQyb1QooNDgGffUMyja5n+32d53r5CgpbY26ok++
bQf2/xxmB2Gor3z53izNWYiMPwa4NjwOp1s3DRzshpd3q5cNCApGUci4vY1ZMLqA
kdVe+sSLpaQUd45MvQTgFhzjnL+pSsP0IoADe4pa7rR9LE+KEfJm3SYe1gQx8mE0
fw6leiqvBbd2noDMoFxZ4ZJywNPG2OdtJbrrTI+p0G8jTaCP/C1I5pvoj/jw5pxS
+LXV5Ns2a8xs1Nvvm4YyU+zRTPgLRkkpcozS92/xEVISyKhuKtG38mtRUkcnALvO
fhXmTdGbJgYOZB7z49zRB6FVabbVPMfD9DImFxT/heNLHYlUzxAo84WmgoDcmpl9
Df3Uc03KvLUBRXUsNqW9yt38zyxh3BSLKqca7ffTz+oqfPPHb6hJLbG8lp9KD/PN
wvtgQ8J7RNxtSJKIeb5LkkbPIzZ/fcpnesqBbfr8ELzaS8uxV7eA47YONy9zxLSn
K6pM580mDx62vRPDGDU/FiG6tE6mSG49kXyoFWEhz3HPTKgQ5LIQgap3ep7W3Zex
bPEVO2JeB+oS9CG89kvt1PPQR7W99Ti8zWodwLNlgKJyvditFuMEDDx0CLfCD4Jk
w7WEYg8sW8H0kXA2RzrV8Anc1qwiLUZa8y3jQFTOEsgWFPd+isC4K5Q7T8ZSsbti
sv2jdRmftIqSINcGJYiDhCoqArjT0aYOEFdp4vGCr0wkRuCEojkFdPRQApmzHnqo
dbF20662EQyQ4Upp/wLrQcISsqwX76hL+swKOfYvOpIWI18YhfbaZJhYv4b/MNMo
agUGwHx558ikuzaEyL0HB07pFDorvD/QYXVbwzcg5257Ogk56/HyUQInJRAwhL9K
WNmED5bZ0JAolI3EOaHi9aGxXyBrbam7JPhq77cSg30V/T4X3KxbNO8iiVP/zoVZ
P95igSriA7AAyl5TotCPGugf5ZgrJFElSQi38D2aK22cJTaXGy7RJJC4U+Ekur5o
sFwIkE1sI+wgvKImAdqvCz+bczhd5K/lLlcVUZyU5wXmhC0gniuAnzW45teHIFzs
OJeqheYzZv8fM5YOgFpqKNtoNNDSsFnrC8yaGvcm1eRoj7Bhdf7qBB5cSdAljWyf
GhoRPTeksspMEKvt+2PnwWrrxZSnWZt+3Q6o/crSq3MDq2dmgIlOUoo9yJFuQl7W
qRZhex9TOsEmtM+WINVNliOVLFNhZ0FWqtqfPWzfCSw5wdhL/J2/J6yZsWGE8fdr
TtPvzyGVXkPabRE2Oin1stVvpxYtCra5glqDF7TjzXzyX6b4Qv2vf39a5CHW6qBK
Nz4Xj9s+ucwzQhFUTMufXwD4vqbZJIZUq9ktPPM5DA7k+6DISUV5QglUvvid+Qkh
WnSv/5+GU5BjaqfAqdmiaB4XVgMmOfZa94tX3saukR0fKxMAt2dxfOIgmXK9SSHy
ix7pomDR1upXSowRfY8UM3moHAr8+HR5idYMMq+IDeHA/mpSxbIZa9zk3GpzRq9J
qn0rNM2Rss7z4zHQtOjl1TB2EaaPIed9fh/2BiGRCrpXIckPCafKS8MsyNZHm3Lo
6CotnD5PkP+kyyT1pdso54zopj/O4X4MK4o9D2dx1XJmC1zrVagZmF8miRX3HXL4
EFj6tomZLe1ILhkbd0p03KYt7kR60U2qIMWUIM+NcQNd+Q6KxQF7/1ZA/XJpvu4Q
I01K2yI9CfQUbJGLlH6kX+tM/2undSgS8SwUldWVWKb1xrR6t6JQsTC6REPG6NRZ
+dOTdzhE6XfTfgrLnqwldPn3TPr8VrRdxK6mH5oBIBm9+nXnimNqjHBvchrrLPLQ
LyjFc2HgeDHII1jnnW5m/83V4AIzKkvoIaxP3UU8JC0cgQgj2zkqaTEbA4gEmbJm
IpehY8gD1ZyHs/KtN/o6m5VV94OtRqib1n0GqoJDpVl6nIawxUG6UxQ7DOxQV1DE
e6lFMx5r6TJPCurK/AgrRKfVKVHUu6nvhnG0HEmxzUxqgNFOu1rpSr+CWSwAo7sP
4/BOaO0qbsQKohJYuzNvfkmK/XLZseAAgml2WbC/zUph4nmf9K71EDELqWruc0CI
46dfGnrMulKZKBpKVBNVFXidtL3xyflHRIuqoAQIPpl6mP6mkBtVZbCMRhegyyqI
itAtnhzTIj1SgguAAaURoTFzLD8b7Ozdq+7/tRrZv3CK607/di2HPr5hVSl4HUyy
1CNDACOOF93u7nCMObtT3v0TgZGuRc2sHDc8RHQf0mCEqe0yxI7+KJQNiEUOfWVA
XbATPMDI16lZcbuggsUpaZKKlOzgIyO3B15odXlbXCP13tRjvXoaQO5HnP0Y/eaY
bA1eAENnduvBkAb+c4vKEmg37VirrXPYDvZv4LWc4r8lPf/dLGwB5OmY2D5Pf4Tp
PfS/Jnf1i9tTthSxDUV0cerU3YU9qB77p+ALmp2j8SprKP+Vm9DQcazpXldcF/hE
9RdHwkeHAWn3bkcvtZHZOxRQYlsoTcAX97s91RK92escOALMVFfuvlE4XQJf6NY5
gdTgWbjYzPkg3/poDm99wPLcmBMSQyIt7t12dCjBHd/rMxBKqQJasFI0rK/DsKT0
wGVVf8uNQO3ifSp2FSjiO2vxDPsqrckjjrjudr+NK+vnfRG/vmzpIDQv1R+RJe8f
i10Uh+rIVTg7KKpTwHbvl+jG7c+i6mLHFETt3bbbYv9zRVP9ByK4iJHBnrRIkmkx
X3y6A/nloLMp6XoLVf3qA5MwMZ61NVJAvcZ9rnunSeqrL1H2euNOWDmPRaD6RD6I
qT1p68j3ttsapVCredFpWi1r53Gce4N24/UQ9AF1JdbhruhVwB4ryc+nrRSy2z6q
g0xtVbf5AgrlTmSQnmsBjAyrsuM0aOfOViHFKlqW3pYFN2u9TRezTkIque1sPSsW
dKo3ks5O6LKraGcXvpw9ByQ4mKeIukaRTY7CdhJMxGlkVk8XFxDEmXVh0g7CXQDl
gq/mjcakXwrSSm1evxriQ5EVC7T/ctSPEpynMpRL6NEKvXhn+Yw8QVUR73vMdryM
iHELXg30hoxdQqcZpQgyk6OGaoiBoSKLZH4B4nSHMcYDscfnCdm4fAOqY0PYOeFn
oKUNSwFp7iwaefIMViOrk/EyacNtlu0bHlMxxwYydHreSGMi9GEw+KNnErgpnp/4
ZmRD04aLLTbO5aS/cCKLSh9MS7r9o/rPaqGA/I6NKUTs6jjT+v5Q1sI1OM47M2MH
1ZJ/UaaVKkBpv8THz9yrZZwozH2nTJd7OnNn8FVL54hftG5HJPkM2UpSAGEQR+Bh
O15k5EWk4WQNOxFPivba5EDU9woLg7wumUM1+qFzLxUQJf0HEApD6hYetkE6ydjd
YoLkVbWnRfip0F/1Vpec+SIBPK/OaNO4uOw2EFenItD6fWhw88Rx626DyQBj3Xer
SS4YO5DeD3Mswa5iXNoy7oF6JmkvT5lGh3YTY3b5k259nFyMmzSiXdbaAYrB1j7p
NVhziMP3vEvKrf0aYpuMP+dMzELZOw61e2Ee6cnPcYJ6TodTHxQ5emQAx1RBwAIm
awfIdOWYCXm0y98w6+SEkisy10OX7j6Nbw34xslcCOu/MlIfdR/L3/u/e6qk4Ltm
ZfCLh43+24tdSzFBEoa53pHVPZmTClzM/OSDv3jJ4UImsSEfgh6MliBqe1MLmFn0
kGXs9YUbziXJkX6eXwjK1u8dGW1my9Tc1v6JIXhEuyFbcTWVKbqBanhRr25sVre7
hQVI3FLBXEr5adbNEzleax/4K6t7ongqvJaHHTF6vjPCwJ5LZxvxgSR5CE6E7Prq
I1GvjKtU/me/3fIKucmOUObcNeIGq8n+cIH7r7n9RRw1a1KjM8u8hX3Ah9vLRTcC
DBs4V2zfMCTJ/PhZgmmhJf2qvUzE1DhQUMUbba3wvnZMbgxAXryfib8ckNynYkUg
o6bZFfNrS30WjbnzZv09E4mVU9l+iSy6Ne1g9YQJLFxGTN5ZfqqvJfnq5o5kOb9O
1vvSWm0lEJtW8LSTwatZnHYJCH/0cjJQbtehwXFqviyFk81ZP9Nw3FoS/reEsoAm
GawumtUoasASWhfwpriCDox+D7s9cMYXaa79WZ/HgmGB8edkbeXwqsNQCbyhrjkX
EJtN96Xye2yqze2Y9tDUMn+Iy8Tt97ReXN0dEaa+251WniUMT4o6Rno63pr9nGuU
ShzwakY1IxEKgffoasAXxWWR7piBnYEUe30KYeF7qyb9+Tql1Z0qLnEkZhF0neRa
jJhKusj78KNfjUIrvm7cEjoa92NXTG6ntaP3H9gktXwAyX9LFikXSvpLIAGee2Xi
KGrJBGrV432L8SHYA66Z61frXBAtUCXAljOK9zFRnMdKhf8uqCBql+Xb/IiLVdSJ
YabCmaMb49fUuHpyR+dTYa62S2c1e55f9uVBR1Y6DG3x482AtK4Ly8uTgLz42h29
vJRFgFP01CLkE9Gy1x80EObpeq8jha+rHDMkYaGpO28EsPT/m93yczdyLp3kud0O
7CdUFTrLXYcDh2pfJjvv5QwYjVuZeQO+c0sySEvoM6IUXi6sNW6MzXmCtyEZZtLw
jYWYclj1g+KKEdEb1bk0E86Xdv1IJfCzxTuxIWNiQWy4oP2IY9p6S76Xv+0i8F7A
2ypkxrUGLarTrFXXerBHMB+oximgqfEU9FF7scLwInsR9kzRQO9nOjfarq4kWjhs
xwsOVPECR+s9RP02/EuL62OhFNxdueIjDbO2c2b0ACtDfzg83InldOZy/rNs2Aza
GsPevXXhwO5MrfRtjWfuVVPd2MOFJk8ktotqlRYF86U0+c0arJsT40Ms4DY5hA9z
5Hg70fO8xSDwgsg05ErPnKcudhAPNMZOQ1eykfzd0Dqx3MWhDKU4U8IlEwcGqdGU
/VoZ19PJgu53WYtJTVNEVQqLukerHdz9tx/FzKBf01R/HEzcW72vvyFVwFRDq+CD
xqO44b4HN8SnAcgDybJ2EHpENH0C5RkkfVuA2Zdcp3FYLuen2L+rs39+NzQCJ9ao
D7hwsBK4WwL0cCtXOOTJTp3Y0yVd45Dqxo5dlZR2AUC23qaZkj84DFhiEJJB///g
wNIzY7j+Oz1w3jYGzEFyomDTqEWKjzXPftFjO/Ok7hUQ8qWQZ/Zdrq25uHDEaseH
KPh+WOsyXENXmzeKB+O9ABpQzblSidKW39zeTMLTBuckV/QsGxCbl0MMrFw4njRb
grusv6FY4G3N7t0rTJc6geMyNK1sGxju7seh0q3mNFt6xb7C/bSSDr5Db6a4MmKb
Y/uFVY1XdXxTEjlsNSgeecWh1jbWn70PnEmGUn5KwKps+kgCYy5eE7tvVUs3eVzj
MxD9+82sylGJU4en1oV6hPt0638L3lhrnzFOHx5Q2GOTSAS3AfkQQdlHMKFo89mT
n8XC4mzmx9SL9Hz2Z/hNfv0dSkM9q4n00bkGbipQWHnpA2y63zNfUeU22pNQf+eU
a3D46DdtJkhVeDuVmaqKMqNKN7PSlJ2vu3mx0v0EkMRhJEtmPsKV7eQAPt2dnVys
HF/B4A+zWS71zb4Vek6Cagsr9jaReBQECcVr0Td+JJ4Er/TyaHKrQA3o4vNzrtbK
HsnvBFahk+Cshy+f+wyhwWnf5VQejTr+hQBLTZ93rTvZEGHgggz+4+3LmACjWxwU
QsHkxf7qtGfwNWuSfmRITg+nry+6mbVFK5eyrGG1kcbWnIVeGDDD0Ogt/m+4pYon
oqvjkoUSLtX1v3YSxxaq7vJgmgszh3tyb1bwQ2DdBoFOC3bW+77N5ZMnvQec0X7T
mU8d+Wa+brojee5ybN/xwh6qwwwnQDbNNZJCMDxvoTOqhB62LvpcISjfSxSGgHns
f+/sLhiB1npsenKZrGbFTBlQcBU3rwM1lkvuu5cvWWW+o9KJXBvt5nHM3xuBqcvT
X3UYeiwqtUDawCP9spPHt9aPtsS2Ra/Sagddgtlu7Qx+fnX9OdjKfNnN/1yEWg61
XMEYwQZyinLAHOTewvT2y/TalC2JQMlRyX7gmrlmTHY8gYTPjsQlvbeXwn6jxh/Q
f1VwnaP2W7IFs6FzB2HU4lRtPkGoXQk7VL2O9gF7cs8ECkbV4Me3Ktb7B4n/N+nf
KYlQkGAmb1yK9TXrYy2sZv3kbY6P5+rhFsM98yU9HZIboFDWAozY7Vzv4hEupkaN
7YarBuBnK/osH5iyoiMBWFxWAjMgpdIHbmdrVmhiyr8DTiyb6n9/cjYdHENpjBYw
1bXoGCScSIhZd44EWGSu+3r+nSFzu5kiNp8BukUYXOdT5biObwtWHEw14PVr6u/X
IipyIvDrNoaDuiZ4iA6YJIdHdL1hYeZ/e0O2FPDu95jOvjRbN7NzhFK4pNPCzv+1
beG2m9SqOp/MiexpLGYQOWeE1SqEw7dEsAG8+eTOiZDY1MCcR5/XcNTOY39w8Rvg
M7hOLfTC9Qh2nmj++hfspKXBCB6Herc8QUWgL2DazE0Sb+M0SlX9MCoRjoya+rak
X8Cka6Uspc9cYXtEd5OPF6YI2y8Fde60iADza5XZX/Zb0acf62PGmzPOHMitgaRk
3RY7sdifEAzQ5gUEfKulOBKhhfFlluMZfb0NMkpeOkrnIQ9zqpB9zq1Vkk0iI+56
aGFl2zMGwFN8ZX4Qa9IUvLytclFYnmcpqsKh/zNtdx7tsbwO7JuG/9QrJctBmDEg
AunZILycH6qRQo+kJtKE9qtYw24t5XynSus1JiDoFghuC9Zyi28yqJ1w//xDe/44
3/Q6ODOx1nSgEIbXpONkbbOlTuouVHW/3+zn889v1jBbLp5ARYqCKjlY8GXbrgbs
wPmtFO8GJjBA6RgBvxyn8YFSYRlkM2QFIrmQSlxe/HbGwDye5Xd7aMOf8wqmYXoV
srL6QzWA2q6sxaDC5b5Ylrs7j5LxXWS2W5gjac/TQv/z47+o0ogCtyQSkU2XqTzc
q+2t6LJHgK/58UwbXo8elCn7uHuGBDZrhBQMBe9xROmeZtRSQpVLPyWhgHkzBDad
IJFWWuaQBPTWOOJX749JolIrzgq1Jho2Ci7pnE1pjaP9j4c9EHuaiHrdjWyaJbvO
QaI/2Rz7JqyzI0ozcs7mdJpB94jCCj9JMm/+KdEVDF20zkAwyLQuCvKod2nbz2jq
GkRGEnnKziYqFy7hYFW/TnU4Z0YbpsZF+JDaXnecwcYwJFT8HOZ1+J7+T7dI+ctd
DS6TsmcUBp1NFEyOSyMZTsAEgGgPxQFBjd6fRdApBDZlvcEIm/orn4oq6f6rzter
Y6PAaUOZztsjaXn6UX2sC2YdEKfq0fCu5aJVNLEEyMzUWkcFSjfys0QE1+E4qoZK
FzdzpWtSmgCBcaEWKtVL9aG2P0kViF7h8QT3kTtXLq+HkcYYXVmN98GwcIsGgKlt
tIifAVLb6ixyz4UpTOlnbnf0wnt8pEsqdZLbXtOS35x7Q+5SFH5B4MpwbF+bALDH
hPh+KHKuHZo3zqowF6vQgiWCPijb3GlBzplHXzMNhMVhHCR5UJg7gkPRLndrflk0
pubACMqsw1oqII8VdwoZ0Pv/LfSxlPLVQJCurDeqibDvVUqhd/wPGKRMIkfAWfjV
m1Cunk6UTUCE3U0pOe2y31VlWSr6gCEf2DBmm1kB9nmirkF9WA7iH2q69taYDtXg
DB6JoTPBvp998kMQ5xVTEOaRwkRwtVsC50VRbsUbB2I3E/ZSb1pu+gQxWv2uw517
EyVdq3R4p4Yv72CUqdJUliqr4SLmcHp4cniCJu78KyW3SFQ2a8n/2T7TsKKRI1/S
6jCXKiSwlyQgghrG+/swvLuJPVrdKO2tdh1xzB/GJl4/eYWxPdyCqfNs/Xr2xSls
jbYxGb08ZlYkAoKveqG3wFNA9hJosj0fJ8UhnL0tpfkPGdh6DBuHjTVXkoE4eHYJ
4dW5mJvyTuoSuB1r8r7JgYU76892FF4hcDhPi+dY5j1v8Vp+nR6S8el1eD5Ft7za
P7xAzoyvicyILhQ5kXgxZ1C7zmYMJhOtXMZT3Nr6AzHpShNEhPeeoPYAmB5Vv3GA
fejX/+TZA8j2NWRZoyrEhvfAFW6R+zDVDRr170lzWqhrDQjrVyE6ja/dxF2IyQEs
EZwGmk/tC4uieUFm2U7ho3V3sI3Ifh8DR6qhkLJKxlt+7LeLPVARax5M66SZfAOc
1YazKBmkg0EeukUd92tBNvwebbujq4cm3L4JkTSPRduZJDPyHTaug/C4eB8BPA/G
yhwFViIQPMW5EMnMpvB6h7e+Nd/CG5bqjvAibtkBjzys+yM4NLI9bD2M7kWW4aMj
8BkWclU4EDv2vF1tBTBkZaCUI5galv47NcF2QgCVm9pVxB236tsTj0+diKGgpiG/
pbzktUvU0O6pScE00CanvpeH5aLYTSk3B+nCpOHZ+2vxFW/SWcM2eTS2CdG/56Kb
7MaJo3oFzp5ySHrch2UTAXv8ujT8qkbAE03XLXVmoPSgBJn8KDrBNagrFQ+kAl5W
6j1FMcLmC4QOpHUfJKg8BoCothizmIgq5VjBKwxBmyzJa/ph2v6xsLWzAjA65MDq
0e4zZ21ac6+M3GGDLDFbB88Ychq/TVb5li1SzLVa+1NiG+Orbma/yYdjMJTi3tY9
XvlRKLyE6fg/ZQp1d8IODCWRGIJWWJRWyx4vtvh25Rd9KMANsCs3Hv4CTikytfyG
GL8E7UAH2syvuADK0LSlCM9Qb5yZRP6pAfihDM3vs3gGWyvIcix7M+Ha3U3byj7x
nM6fzcvdi6xPhip4GH+KO6eLKa4MH5r34qbxJ8iwg+8QMxWmgo6NVh1vP/lqyfMf
b85yCNrw6onomvXmFw6WBtjKTTUZ0r0IiWAWI4bwDK8F6815BGzpTCgdiTxZTwaf
lIypERsp2GrHzoUvXL3lgUTIz52tYV8ACt8iB30llF3z8zwL9ziaJ/1ZlelFSOLw
ejQAmi0ZSUluDDeLUcMTa/490Lnlv59sy/krz67Gt2IPfwDMWku3eA+fbcL7QtZZ
qAL3U6HHdzu7Yi25F3QFC1RdMn0qb6UhgNlZOuB4RO1w4Q2F0V9TsIlgrcrcRKsf
obxO7CX9+owpmx6pA2tJGQsf4cI976M3TsIVZc92nJF22iTmnEb4tzA57nLkqfUW
jDUpdzCxkzS6h6Sp7MSML9MNC/VPNtluLPt/odi3HV7OhJHzTBgQq1TvYgFZueau
bqVP9B6IWDYK0sy88FgEK/g3O7Ny0pjdzZPefX8JQDODuL0NWoVDiZ5iKA+WPSAm
Wgd7GC5Lm29PQpAn+SJs4kD9oAn6FKSkyLu5geHVsQYUkrdOb51gHV7LdOZ6EeJ6
2jxlQt33qJC0LLrCkDx7Cz/b5WNYwle23jTAMiV8cBSw+ginE9kI7HECoORM2U3L
HgAgIyeICm/jKvZjcdFBA0o2nAf+kPreUXz+lRsNQMg6VFpm4HlN1F++b3sdkHQW
Iln0cYyt4E2IheqVH3cxS8dPolKDAaEZm5WTk0ynu8y7123i0ZoKUz/kz4nikmX4
GAfk4L7KX9yZDEKjbkg0SKxZH5wxqWCd7Opb6Fz6RLJuqwvJwnXKEAKduwKWZM3U
kNr7+txf2flU+PBiAx9BH1gFWXLnFZxabsngjZYs7RQY13whGU3urfei9PLPUtRK
eNHs4v2Q9e/qJd30PNwOBXsstdVzqsfUlJnOdGIDayFw0dpVV05jmeulRN6qRhIN
fe+ebRfOcwiukCQj2t2oo/sUDxU9IA9ZUBXU0sK/3W6PqKcLn8RkWhwzSR6UFJGV
9GNbgBYhZskhrq5EVtOGKhXq65zFnOJvKcFC+eRFELS8wM+oWjAsl+DWiSiJD9Rc
c2/tAOsZvB/2D4fY19+AdFqt+JVaSm9jnI2BCjYxIREu2594oCRJ4viwkmYxvIDu
6S/hurd64u3I7xoxlRL6y0wzZAewtDCbYDofSU2td9kC/i42VFs/FbneRlJky3GA
x7USsxcpaU0TF6BtF790kFdeCGORdmFMa5i+gazYkRlOyj2xmR+AV0G2wl6NpWng
A+0+owrjRNQWJZikmTMLmlc+gHHW/amdjdwORBiIh9+9/F4gyKrW9FKkIv2gt9lo
ca82MPVjTKTuNGczVTKje7oiLUqRHA4a/aFlu5BWpUP/JRxlZcCjPrp3qZkNdn5U
zFY5kkv0aPDRLeXpor0mDz9n1P5RX2yWQEP9UPRKCNDPT4SbOe9oic8ynnlJk4dO
Aq1c275W/lwNIgrKOzOQlvYpueAQF2owP0RhEuzUzlz4cN9jQZqaKRBSeeQyJiNz
1d9KenErJ/THjDd+DP6zWEcWa/xygX+J1ojmDtVNUy9h56wasWHRkE84UKpUUs/c
3BBuHTc/759wnHp/MhZc4iVBuLqZCsP68ZE2+0ZRfMufl0gFJOS6kZMaC+KOGnrj
v16OermYMCZZyFRa2RfR8TKPnwVFZ+BOh1HjrxBi7ExoZ/OlZ54lZFWXgS8DiNJF
gwQiILDpAQN/uUg+n1qJ2dan498AKI2/d81TM+xSjd4usYbO7UDwlC2vw1kMweY3
4DGFpqR1OLeLDJ/haJ0iq3vaAAocH84lshh8I3esW0S7EtBu0T8ObzZrnx1yr/9n
D7Lpt9qsptHxQlY+J9oMossa8J3w1ws4hLIB2p0sraCFy/Q89nKyyLjM3utWphLV
aMtn5a3zOOBGjx0SBndMwWgz3a1WlqIETlyLfAQyrbMDoE/v2XCEhldh2DRNI4eq
erWE8iQp9bdo9IbIgLup03cE2GH0lIPrdLq0PqcxryLhs3IR3mJdTCq8CVI7dKOf
fDrUaSi7NglM/gaDPFB4JdyDiuGrDQC44y8OvVYOqGEEWvLR7tjG3S9rFS0XEjhs
PNgmoU/sts4Qcg4XY8nHwnNtFu4DugWlowztrEEj/6m1/HVPvNFhFfzNBBh8NKh3
4k3H+SraW6GaaVbtdQADTKjAXxNjvEKS8OP0B9/SvjT2ye8hPFw/nLdo8yGecVvY
2iUF5Phw6DOtcdw3HIHZuvFvIDJsTN3AxfA3VCXB3C9erJgojrvmu5utlsuQ0Wlr
5FgY0MpQu9SR2u05UtbxtBBhOjuAJ2MO/jtteQ8YJD05a/PTw4C3lNfwo+tpQInd
c/Xl7Tt8V85EnbpP5x+rKdJTRUAqstKBc5MoAbUwmqlebuVL0hjWTAW4uPASTBeZ
zNM30SYwXSTyUMmLfo/RXMkTTrm+epRgz/AnxtuP4CAUyvLmP71AMxNCNdvNe4A4
+lBi89IKaXcw/EbuxwFsbo1U6EoghEQ0WdANp4KDt0u82ysaTcApn89zhSND8Moq
crJAPEl6jJRLG7zLeENcMzk7bHbQI+Zwc/6qwNwI5FwhGb/4y5rSOfCFBPLd97nr
JTZp7G6YVzzxlsMO26Ewvz2CJc9AQR6lMMtEkFPdqzI4mAIKSUs1mrw6mprtq47r
uL/+fsnLHZMS3vh0oosQIwlSD4xCqIOqc9mRCpDNhcR6zFTzDNmCe1kQmZ/gEe45
k4ZHoA4kbiCb505MROx3ZZi26Ms9IFxo1AGETEyHWOSMXz5eyS1BXQu56fwl/fx+
2T3RFUGbDFxPbAHhpV9HNDN/y29VlYiBIgLft+3bGGf7EcpnY9SHKTiaYf1efi/6
8mWDUc3m/bEO74cezne0vNUC1cb0iKqpiCgih0GH9QcN71QaWpmQSJT5wMqfQa6X
nrALFXXBUJtw9xl7DZFczYJnD9XcY4oUUM5wOB0LOPWRb9CvHX8U5vFAyiPCB3u2
nWgLlC6J9neibVJIX2pGVfaF2p/dMFsVr6nUJ6MOJDGtSVA25zLJCD91HZtBdG5H
wJIeeWf6qf+FLIzVBRMkOWDgoPUweVcPeeH9gqmPMW9AtMLsI8r2RYZh0Qs6YJlo
ZKYcFiRpr85t5fZRf2VGZUEe/wQ2j/ATOQz7PL4TXVjnAWo5GviYshYBXPzDGGMQ
vTyuXgc4NHWAPYR0BpVoH4Y14hmWhTcrwjkbtOw2SeKZ96Fh5DyUMLJXo6ahbaHd
/r8A/7DMc/h77jV0Li8orGprHIAf1AoQ9CgJOL+x0DPYya89pnlWI6O1EoanxflT
ABwcnzRwDT6LWangMdnylDov2GjpSyJPfwjYeZTsIaboSe7x/YRJmOOvAhVZL8zx
EGEE1d+MKfiFVLXOygCp+KqbzRIdQQpSkFQxs0BFHE7gfX4CpRCzvskp8UHyypFz
q5ODEd6pK4AWGJwspZiNWA690t5vt94sCVNj9Nlk1RGJJm6FwuRRNEHf7I/Q4DO8
lvNxX9x8SGwEtB9IuZVGjKO1s1wEq81Yexo0w0H1yVxgbB9wiZ83gCVlM45oomgD
pd+3r8PC6f50d2UJHZ1zrQXFpszsRZ2mpLXTXeWUv33ck9tsJ44m0jtKyqisLr7A
rh7ucbMt0y4o6mvTGaGCXa4aZHGcrdM4Opz2QEcKCS7F/fDXdu7c58WTP2bgNsL1
WrhxB9fWqPX1NXfbcwVzqYu+t66AmXsjYCieKNwAXNDSwSGlqk6ls5Fhfst6isqF
OdtyI7V9XoifBlclsZW3PsZMIucSEFVn0no/9AL4mBEyVN6xpjUiQMQJUZ+Xx3zV
9izgmZSiy/8DbSO6fbjxHxfc9B0dCr2lHE/dkecpVfpszY6wezVPRCnehhyhu+rN
NzxVhsx5CKBJAJ7pi4WYGrKGeTuAgH/0MTr6khpp2KYAzpNJ8Wy5GxkhSYEV7JUP
4EbLvxy1tfpsPavoK1GyD1P2ICXZjvqMWuxb8ULwL3UmWHmsd5Ii/00rSUIb5uab
HEo+EEhqVPCeACB8WfNggnVT7+M7i4oDmVXSfnFwAtRU2M18NennKJ8yc+7xZXBx
OqHGratJywKe7RJca5Uilq4D4giDqRlN3PZ/EaUJD1AX9ZtreMXCLc2clNopy/2/
h2jTaQ9IGwCCjgWlbFrTxMN+a3+4ZFUKnGoNEJTRHkpfo31C6m54M38bl9+2wrxq
mHKKi7/TRinVCanU779A/QcWgI9L0g19/Oq563dgVs+XzWHMkUMsRFvK/MgzM5y4
wQZpetJfNL9lxgn4ZqwPBYzNdU+z2J2mWs7xljQOe1rkF/oa1fObGjR478CbqEJJ
Moz+xMW97ltgf/iW0jI3OXGH1OKk+qyFvBdYRlSfK/P+yuiphmmpMeRzcUIVfsSf
YyxXvY6IGByABIznvYDrVQk++jwOuPidAW3n1LIISFWp9nvjAx8r8LTJCOqjA0UL
FDUUKdFtVOWy13m4vIJ2kcMgELop/fnP4bD1PzOwFApdy4gBVQKK7vUF8hrvccow
08YtR54hxnD04xNbauoP3cBxANAX9TZgFmQ4lGbUUXmwy7+41QLvcS9QtviIsoDy
J7Ke9x1eIOMAd0C0hZTLrX1AIbCHbFFH4Gqxwr29juU3icR8lBY+R6ihTt9D3mVO
JkNa9dAwV4l/Q3iIquxxfr6NbaEkm/bRnO7yW3RTw6Fe/mlfUrr5msf5AAKL6HJy
YxWjk7MM0ND9RE2ysLkZaApTWH6/JHaiIRq76WMiK6uyrin94YWHmS0T9+n4c7PD
bcXrDTCeV4HSCerkje5BTRlEZIVUxk1Mknrg1igx3MlWduskLpQjb94QfpnQiSnX
6VsGcCBnh4vCZ5FA8VaYB/eNez5Cjpn8Kgg+1P7+Znu3UIY6sjqIkG5zPyVj3XZU
BB7XyS2Dtz4DxM84TaMPctl9GLNPrYY3/6F7LK1DIk6QLeJVchHhBpnivTQ2t+vH
6N7GkppgvPHi1sd0pkJwom0Mw4Az81uHyW3YlUwmtJIMHLOvkENjhhz8xx0AQ3Km
xjj4LO3VlzEOezrm7tX2DQYPzk1hOsLUd/jL0BdtrNi5TNsKvbKHjX76Dc0utAJp
9dCu2B2uiFw9v6Lb8osaSS7Df2qbS2GeWE740rMFJK9QGcg73hWk5Cqupd+DS5My
xe2RjDrZry6FcU31ovFvPwJQQ308hC01AxDJcduzaylgu1PLSKnOBXnZmrCDjUrn
3faxmkn2i08E4IX5fTbWg6mSIaAwu8Eq0xTF4o1CU53d7xJCvHcxTnlaP4LuAE+r
51ac0Udb/OY7Ctf4sYL2Jp6gx5ikgFre+l9/HYmQxJvl9pP1R8rdZWRBGBEgV7I7
R5rJwx9B5ROIY8yZCnIZc0obckIQkWPMWah8Vh0AmqH91fVhGPYM/KfhYozDYlUV
tugIsN3yqvkKREFdxfJS7Pxyn7NwpR899FhQtgyLFVFUuKRVrOw/gwJ7wXIQ2dac
BaFKMaxD0FRCxsZOTMHAr9qr088VYoQ+FEMR2XgTn67AAjqHcCLChVdBXNXKljRc
BbIhPwUGpBTGEv3KKetiYmEZQsMQKg5vmhpQwuz8l+mEYGchJKwWwGYX4ZGufzSS
ovvOU3CNnQlDDt8dcpKXaakC0tX+TJ6yL2ECQcZBS8VdDJSs0Wpcaoa6pDuMFq7f
irUGc4+Lch4oRzPx6HNRvaqg6iyGKIg2cocQHEyCEiJfJAHnA3WULXvUXFzzVWxR
+sGy3SzDM9hRs6zMQZdnLfKzCT0IsI22BlsYG4svmKrdZqB+8RKi3OCcIBopnOAy
nxZ8ozPZGFZZbb4jGSlxVahpsujDwWasiV30MLfmtSYIBX7pDBPzNnMaA9TLi4/O
yrulZmuBkIEdQfr0Oks3tU3Ts1eOJOEMMoVRCWY/8QzsEZ6g8XJxj9YV72kcwVcS
lBI8ZW/2FJ9tv+QNzCPF4Arb5vAsAk0GduC9mCMIcudxKTG/k+mNDPV/pOaz5Z4R
g5Czl5kUVtMPNwdFnzQeXHzRQ19mbPDUxaYsWCKB+A3wfPg+iPL/nRVM0xjOv1iX
QreeYgMhbSOfPILPVrdNgsTFJb9jJzTTGs1KLLmAJQmx0RPVCLMXdzG8xs1jXuf+
iUXcDIjHUK39mgdegpPugwlgZPjlXMHBS2+ib4knSQ2IZtvo7B/T2GOH1hZJc0No
JXlxpgntce9nkjL8AuptFYvocHhQgBK7xXWrM6xSO9iBlj4ppcZqMZzqZf9FckNu
BgmEJiqOKis9xlvbXFUJwEAXQHMJlpItvrMdWWBLt7j+oV5/YaNd8JR1MFxRvlA3
wNr2PXmBJp1KuEGMp/2FhMgHmMyVf7O9FRUEUQhN81KMeysTAZi1DoOWSCupgtDx
yMkWukSKS6D4lMg1rpqsEBPgryXhoRxjqH66bfholBxvkX2UA9OMiRFTpFHqPSGV
spvfwscxXhuzSNjd5uuPHSxu+YoP3ZUDIz9YtP4+PgUPpi6aA4UXgutHOnPKqVkO
OTXl4QYjJ6nddvhHFOIBXxT590GHafTbw++TzzhqekFIsx3n6mUgBjBYIGEoVKN+
HdeKGbckTRWwalfdHmDHpTAZ/jvaiA7U5/elfeyHXfIJ3h9nzwwfMqlnQBu5IY/x
q4FgRyuD9/jLKOLamZfUK9/sDo5j0SvOdW2iCPu8riqBMVud1BOUL2BYaR9aSM4y
VbzOAplvXaEGXbO6TPcVm74fACqRZDmpZjJ75iha/Xwq3FpPnyaDlbE0oDub/Ysu
YcYpFQL6ILvQkaYr489NavNjcBtDQBBCVpE1Vw+ilzWGBxhUgkwIpAiq4HhTKLqc
vIHu1VDttpXodKsmtPR8PAeoauRE+YtJAmkvDm32b8kNqGXp7hDjiptKMyxEgerU
S/kFt1/wOobh9KpIQZGkdQrkpxzUe6dvtHEPWHtuI4HYcQmq/bdPm4Of29npPHjL
thqziZsBt42GOb26hfMz7Xj5B4c3YLPzG2nhMmOuFK3KcNc0YhCm49BeTu4WHc3G
eosRpOuhqnEtFnwef94EyzBStq4rY0ncF1OdQ4VIb1WwzAKVvOR9OCpGj0AOGzUX
sogGBT+9/qAv+FMhST4FwBXCe1aP31VFyAvD3/H8cn86Jw/g76ntNJ3eBap+YrHm
6L6ZSvhx0dS+Eo0V/qzlWcV96PbAFnWhhbWd2OdVeuf3fvTIzd1sYf0UZlsG3ehy
zPud1sTxLaxIpWBrm4zmXXdD0SGAJrE4DVoIJCMPTUFyyTI933U5ACc/qnyeSOCL
DtINgtIoOYKhV8+KTDdt5x7tK3cI/euI9HoANfsqy6aOZ7743xKEsCrCBvMPpOQ8
FN+Llofi6kHgDkSUWTNp96UaSqkeQ6gYwThL0udZhjsPmiU+11tqHWzsw9DlyipZ
XPyTSLb2xxaz5aJb2eq+7M4tvtVlsZsc3g8eOq3hIw+l5VprwgGhbyeJzi4D5e8q
xQbddgTAcMZJpeKKgfgta/VUKULxs3f9whl+dsJrodsG/akOOgUvjchOggjKzKsM
K9xx7NFo/h78W29eWZtzEmIPp3kloAK0aeHZfIK+pI3WKfLsrxUbDafZmE7rMu7i
CO+TYUsg+S7wgs2ZHYwxfUcIysbsKOqNq5PEfbAKxTEo1/CkdnPQoY0gCXOKfLHn
y/4BtsVhrwiwuaRDsduOETVlnNrLPPjxKAKwWEUs+zBSGVf43YxW84RHc3hxKHvB
VAHTijrFU4l75CwsWDn+O7jL9x7VeNn1UQwQHwjT1qCdw0mFu4acLXG6t4kMQ0V8
2jSEmw4zFE2HAAlZRZ2fs5Wlv+r0v2qv9VAyZre2GNiHsXc5yVi/aoMxeSWKoAyu
T7TKcxXO7F8zcr9by3SXWQJglH25UaT239fWHc9LMGWog24o4FcEaibgw74X+H5y
jHsdw1wzQoO0GJ9Qr61soeKzyDjI3NAIVCPZPXwObiiHNFbeZFAevlHkh0vqeDO9
2CHR5uGeThaMt/DuzXY+SHOlxgu8xEN6WJtvO094EKUW/aBehJeaX6dmLUqWOIVJ
FjSqBwk612JQWWTg3rjmeGnoKrVTfIHlTdagwKJ5AhALXSGQBB3RJjp2w9SgJyey
28v38yZB6JdykFQAsLI1evZTwsAct/STE2i5mnOXV46w/GJaLXlmw0ngeSyQfTgp
l/IWZ8kikUWpKge7HEMoGIEeWPnVyQav76l/ndrNfaIyJEPzo7CyzB/S+v9+R6qR
xMZ2mEQnUeGVsAkvqVkeuOYPtE6zOY3LaqfHFrBfEh15AgfcR566hyyZVbagdhvN
R5eBVoSG20cuU1v+O0Ylo+S7GyOKiifmQs4hXzStgbeCmrcVTRJ7cquvJSo5Uh8o
xNrcLAShtYKONAmT6lLHRVlL5pP33k+Cc5vaNTt2uWQjQ9hq7JWlrDARs1JEhVVB
Cem0KwZZ1g8JR4guv59zWr4wVxQTp0oJwsCvE72R/khmMwnpNieW4tPPNijaQUc8
d9SczSF8Tqac+DtSAbGWZ2CpvT+Q9aE8pyt4bCDOj2DTbykOdOvsmR21MItf82dP
Ju11jR6bZ3GNPLQOerBLQLV+nEvoG6hg5wZ2FRqy8w0PRhA4XtSkdYK6eI6uRqLf
48yafn1XH/x2E8WwdbFQhFODCoem4MuW3utHRspWT4br9ORVy5bLi6x+8irPw7Np
eg1c4+T5BS55u6PXi3KR+8td7U+7nmKAU9m3ECwyKmptcB8KzWypQ3NfqcHUCznv
nBkqx1FNr1AXm9mgSQv5aNNNYCKJOF+fDoSi783QUWiKqlQzua0w9Od+NQF26blo
om5SRL6k/X/Ts4TieyapMC6++VzxLpcIZW9PNcnLgs0VSLF9btKbavRQ3jlQNfRw
VzY6IcIBYnKmFGmJqS8v6TJM06m+zceE88FzWIfKXgX53I4yz7WXQ2j91yi7jVuS
CxNaiWN8j0HemVEX1LhecHsUxVfSyCm/CqaGZoglPv5KNVyp1FmUTwe5R/oGMsXg
YG3jrooAjEGZgqdEf+U6fByXuPcjXJXOGMb1qNndaHDbyX2yijxDVUavRw89nh4n
Y/ep+nmzM3m8UhyhOvx2DtYCT9oCkXotBqdbUWBN7GcXHukvyecqpmI0nR1aAnh5
sXN9xO4mG0AXvzFgqZIh9ffnCbtvHsYn+fztGVYe2nTCLLNhbtmO+r30a1Ofy94S
vSSeH2RnVHsoKoEkzvH232OBUqBpscscjaOo0KPvTTK7ENMwHGAIYaskU3Sbimxq
f0nUyuDxssMw1mpE6Jsekwyr3xRYGWh8M4nY5yva1Jh4is2c+z77qtSZ7FoAuhez
VM+pw2n2TGIyvG+qsJITPNLSKlORb3lgh7d6eNYs2HCF6lAXIm4Y82rZKyrtCnjL
QWtSjYpYWefFt/oqe9mzQZRs3bT/aWmuVdJl+AC9lTtX7r0bvgUJZIFuLhUIj4pc
OBQFmEDt/RM0puDOOA4YXqdwjyX1z8UEUqG19RfDcIXRj1NuHiRPuhQQh3V41MdI
4sEJSqS+uaYa5dgtLxVsQwpshpyeZhRN1PKiyUOt5Q+zoqacsTmxo31rkkYVbkYg
YhGv1OspHPr0Eh1PeCsPtYGPD0Elzfykh96b67qE+QhPx8klyMOuiHULsY9eHOLA
GCKxv3ajPhRnh0LyZ3LuHo4BcIfEZGG0NDfhvYyZFt7VnguERCGgnQ+JiP6ATZ4t
amGVSIRsU0CAWHJghU2sd5bmnmXuMcGiqk0OC5Pa1SLxxH97Sdia9Rcxllxl+Z03
z7R7WiWJRVac4n/Fo+8ixeBJsmjnSBa6forcX/3RvyNQBQbu2VfB2yK6nfoOcULH
RkFop3rXWTYnTSgWVlLpLbCgTapaUvrzGPu/DLJJDdt6pZOzI19Fii7n7dCJqY8f
zymf6EtsOCamyqmriKXYCFaIacqfvI7cyIQAiqknK9P01lrPbMYQVVTJhJxQKImM
50zJpBeBGggMMUDEi9hRaJJQXX+darwCGkcimQliYaW+snLmekLKTVvRfyGtlmEB
KqX9OtREQ8YfHcLpFd47k8pycM+Oh/sp5TJtIP712uoYCyLB6l/DWS8lT4eRhsLY
M9W/+Sf9CWMn209cZi2NSszSiWbnhPJ1aZ5ZuQvPog7Fg+SgjC2+6Ga4paSwEGA+
mHLAsRARdMrUem0PakfKyoy4D6MidT5MPGy9ylU3WpuxA2eskT1StrPqvtcjMjcH
D9v65cplu8+dp3INoy4Ww+rhTQgroHUe90IOM7EC7xM0qP2wW7+AMof77LsBf+h0
FTDcmFYQy1nTa2MOtXIA735h4O1RiWDbqyFOGwRaJqwOcSfySJ2MycIb7I7xqbSt
kTNbEgcIl4hKYTauqpx8IISUZI814cLdfDh6Zkf3JaOcOdLyNrBU8BfROfhE8U4q
aYm/cGJRqR/NlVBCJ1Q6reQkhOzz/oR4X+4KT+Y3oM5NOK2ZZ61uhfP4i93/Hn/q
KEt2GPMcFn8HVKWOZUllIkcROyglhTV9AO6j4FXLSa3UYzFn5HFQcrrwj4GHJIIy
yEE/grB1lzT+iHDgh8gReTlERu1loZ2wTrXstYUWJegpf5VCM778KjNQm58MlyXI
TsbgL+4jpgqpvpP6nxgpaoAMEL2XohfcxtVUSPm9MKcylBr0QTYsQF845YyaYbZ+
KTnYW2aRhJSnla2cncser7rpKsBps3rC8i769egmDOAqdGtuvujIE7GhMlAk9oiS
MnRaO/TmtIlreUqXtWflGcVS5k4/5Abn3FU9eI1ux2CDvXxYMc8xHZqWV5OifQ43
WoLzswadV5zxihlcv0tSISy0TJEltsbmtaCjcLB1KSUOnD6eGuA2kYVfN4mm1bRy
FnR6LR6yVs6P6CC7JkYph0uCLtc098Q5nl48bMkJUGqUh+Lmfm55hluQIIMsV2vE
u1np6MKPh4Q8+KbqeKOhjiaQ+xeS898UIoPgSOdCLJF2lobgHtQrDAAm3UEtZdA4
POM2p7FW9YGIJXMtEdtY50Ou4v5mgO7Xca/75MfEXh135AFP8gAb5wUAXgQTx1Ir
e/wGjZFYPGfo7FdzsEgakBBWYRVKUGfvcnHc95Q34NqMme/OVa6V8TTaERT0KXC4
iAJFJK5H7LJ/LXuMQM+U2fy4HVFIgk0n9Iyr+tl7CFIW5fbPU2BHVsA6uHOyAkkJ
uhTJl5omEfdOX2VOhWEZ9VcvfWlf9N/mdeTjcPI/ZFEmk9jDQdRIL4HQE2fDT86v
0CMr+mvFN2U7CxTUEr+iqVRRQM6WSwYHE1bQp9PileKSBX5QdIEUVeBinaaUw2BM
dQGlQeyySRfttadrvGdeTosYsgRfGi22xnArVxShLl1zu52aH8/Em+6nU0tdgYRw
Dyc8jkKBhAoMdRgOPLOndVA2Usn+fWAea/oTdNih81jeS/GCtNMzRms4h9IWxjE6
0LfxK61jr6bvMFiPe+QZGlHcUi4lJH/tB21VEVCDMPjn1CUHWYIi4DmZjp7YOecq
h+3LAnas5Q26ERhS5DoeENyS/4wfyofdesQy3594BNGk/aoh8KEB0DgSpOJFYVj8
RhqCHaFnQOoI7KgWfalo+FE1no2R7vvt6vAbFlljutc7VxtrWvzQuejo/TpvyIkI
bBpkoM43kRq9843CEJeI3zxuM6fZQ3jeoz/l9iN0FifrSYaawks95WnF6JgUmr4S
An2z056UyFZXyLRDnEse2Us53wyDNgHYHF/KKta9pBAaM24iKs333596+eD5OHet
BOG7Kdi6YgeUMnu0bZLXn8hXuJNf6itK3FrCcku5nyNwrHyfKWwLZGnSwxHyBGgc
nclAYlrDOVSoI/rmfNbqXSytdeCLHsd5JKBSlyEmKekXDdPvoep6L0XJViMYZ8H5
YVd8qd09aQPenCUpmctR03KYakfhf9kZMF2v3xKU/ABmVk46g1ySWz8Aonp5/bSJ
Z4xFY01dd0/NQzmUDBXTVl8H1/oUiRbsxA11BAlpF8NbTpNFBJvRxywXfZOg0B7K
rqvypoWcUPsAajmDNjdltb9LICL62E3EIaxtWCRQG1IsV++HO/eYp73ntWK6s7H5
Q/j7Ua2qUrH4XUIWDbT8BDAJURYLo4wfd2gGYadKFfZvZI0ddeSnMCScE3DsQOi6
sNTtVvAM+w1QwuAXz3lNZmYJ1NRFOjaPz4haxgyFH3+Qxt2ql1WBoFcgyY8r4KHo
1nmMIDisMiJ/23BWuR0DEjAiRIsWhcZ4m03aL4jlJVZxUsXU6h1yDLDDvBMYV+rD
nFYHz3SFaHFvkzNXnI3Kmuut6AdsxjGnvfmgN7txhGc5rxpDsDN172qUuP/y5ahN
ZKJuG8ADZowirjic/2Ko8Ozgfa9cEJIpsNXRcvmW6bncp5NSIgE7nbeJxDCSWyw5
0kZq6liTxP9B+Kjy1XitPD9unDLFwYbjbPGgOqVFsW+4ukWBe0Q2qgtRJPt9x+tv
GwoInqHW5sSqgS7Mv0cOVPoonrlvts9BCsk+uxj2GZIabztLfW8QMkqiKGn3sNFU
tYdHLuVtmqSwb8pXeDkd/PBDbyreNTH0JvjEDoh8sWLpV5tszhq79I9NOsmK/LTg
8+o76d5rEpYdypzBIz+iiDw06oktPbxJZsOeLsPnJ0xkuGPBccqJhK4DyzdJfY0I
5Q6F0zMT+PN//5rne+0F95DnXIOOoyZ7HIPYGZ+0gsm4xqmRyhfh/kdJ7RrbkAJg
bf1L5o8uUFCBDw5clJhAaaehBPufZ440mDu5B8zvF5R+ksWYoy2kODrGqnxS5wjY
B/SZCvZwj71qMdSzFE6m43N73jhAZvwWyxdihfdgUgwfw2VZEccB1RPqxmIdYjYm
CG7cZ7YKLo2t1eM8qjf8ktNNAZoP2NpAVSpChujdlBipAoFtQVcawRa0eV//F8X2
YhJtwFVWiQV+9Ce8j5cYT37DlIHnGeq6YTnToCFk8glReveiizcPsOVIeZI+i2ao
r1BdKCywXImdptjzTrNZPY+VmOAvt0x5uexNPcKP80EMLPmJezwiDHu4+jM70HpB
YKRRWZo4ON10/ILi7CdcSfFrqEFRyPSNp0W/SRXbnBhYf91qO2bZM+0tREcR3Qvl
U5fM4vdhDESvG9o3cCRKHGExaiyjvgtt+sv5HaB3cvnDLe15uhRveTZY542YNZ7r
3SLXGme5mo05GLugFxsfZglHcQs5bd38TTsB4sJl8gsNvNG51q6y0rcU3QI76qRw
cqU821iC75yknj4M74LWP4WoZsELKnBxuGdaMO2kCodeFU007AtyyFh/hGhPdTCN
gKLAz9bYjmESC7ufmrbpAhUS7/XO8Q0Ul4/OzBi1fH+ZVOTg7Ie24ainiK+RTuLN
XP4qfWjmkmcQRKWyX78d1Q0ZjVJUQEyXhy8xcVcK3DqWWOO+yQhBmPP69gdyrV5K
1eoJD//JzV6So3eStEYvy5DtBOcMwfuxABmVJyjVeoWhfNXb4+5e4Tlg2Qallwn6
PJu/FFm8qNflSe3HeDhB2llFT4TxirI7y/A8c9eEaU9lm7d2TUDSiPP+YI6mkm2y
RmIthn7YHCS/+I5fwWNT2STEYcAt+/tDlyGUlPXqkEAW9iJeTooVFtzGGcUy1a0e
QFGwMaSOa3bw9NY58JsYDNLI+n/JHz927SCEW6UlLgjUt4o/9+0JGiC0rTEhMaMT
QQLgwY4PQCpgd1XyXZrOBYKwEOMnXhohkwQAfhpq4QCqsnwNNnC9qPDQlVpuppwn
NLyJ2EzZIUHfMWN6CiI7byyEATRlXvKyGMySxnNvRB+uXWS/Fr4GFSWzKhCC2tXl
tmMk4lUm/0SW4JSnC4pJko3WMoqKgz1kHeC4AoLTn4Bl/65vuiWXA1fajcrivC+s
V1AXg6rcUmlCCfGDNl/quohLS4Yi32ftpWNVZo9qt44P2qzEh61bFlN5phQt6IKj
GjNA74e02EzmZgEXFF0dbUcBgBNDTjCjbdX8Im6GGEecdTochRxXCtciLVw9kK/8
yP46+04d6MpJXkDk+v8kVKwjLXlYWgCuA/23nlL4fXO9QEwxnKuTWWyZ4F/fqoI0
RnM1cY1PsYQZ4zSzOi/XR1/mzAr8HvBJ39tS5dYEDXplpIzniEQPGHY4BF/1sEEh
fJRfK4mqLE1HZZN0Ro+iRQ7bq4RJkfoUVNeNxarf42NJBJvuXZAa9zIt/EzWvdnA
gmCIzPklm+teCUWsZqvF7dG7QI/orJ1ftifK0vma+2dkM03+A2DJvW0+JE/uFUXZ
LHm4oHc5Xb+hj9TEXD1KjY6mB+WK5u+qm1FgUutpAVRUSbZs5t8hh8qSpHGG6avc
foc7BE5NnUM1a66M2hY9TJuUECDJpgWfCEV1DalO1HkZaFsXlVUCwQkc1vjJZG1S
wu5kKYZ8fKJM9WoSPn9+lKECNlHgVu0KS7EFPh0IQX417FJFmk1R8TC0m8lgsRgQ
e/AVGqCHox40YQHIS/cuNW/n48eY+WybvNqQcfdbAZ5lf0D1N5bIJz0b93Q2KA3G
77BMtCH3x3dpJYhPjRDmWbzDzauFdxv7oFSwXDZiL8YsjqIFcoaEsPyqTfBbidj9
R8MA4SqBHzq3htPTOI+SwcagkcP64Fx8609DGSf24OtX1fZy765mwaQ6aM5P3ykW
rSptkMlBbfa1pQNXcJP1x+2ZWbekU2Hh7Dq7P2keXMECHnqQcHtU+6wZb3QQpg+6
hF6o3rw2o4CkF2bGQ9P6gAiWSy1Z8PQuCutFuaYKme+qFOPv1KD62lfg0m7s14Ue
bqQ17rP9lyw/g1k45TfYUIT+FbVz24b0+SzJ7Gb6dSfdRFrAom8yYPN0KD19kZx2
i9W1R3d1QWicv+MXbtO8Zkm1A5x5BOOr8CrAVvYXHO8VKvywVDhEx8sSvOwRQsS9
KtMmDRN3DzACx6rFf0+EE+kNdcvdGILXKts1R1ySR0l/yVd6+mWmhwP8s97/P41U
PDoZvrepctqD89i9+Dn+FcmOrPo7Tc7gcw1wC0w0cHPgBgkLil+lWuwNyRTT0eQq
u1Oteg3tp4aw6JupVnh7x4MnW/LDruzIEoEN5cjc/FfXblJNIkFJ+xWFOCTw404R
6tTdZHjt4Oc/Vp+W5z0RHLhsyilAYAx0Radw77qs+7AaxkBXKmcMPd0sInPTEQOG
qnXGS4RG8UddmNmT2g2cwNMsOBsmJgYJy1H9Py/7+qPLsYq5H3zDflN/VaYec/Fi
84kXNqFTXpNTJW5Q/avaEqydEsEl4E74jqUI6fVB/zFtSQYl3mHpucDQvrlU+yEt
WKMFZge+yeBDVkWSiDgwX0o2oVTWacgvURAnk1KjEDgZGEMFj53mDucOce7C91cH
vZglngCP1BG/DT6hXl1kImKYyRhh+zLuNCCHsrvZtp0xCuUDhY2YYb7LSU+tc4TI
Qa+1JdEgVM9pDisaGlPR6koQJTwyJyMW0Pu+ilJf4cqKht96JQWVgmAAGd0N0cBb
h+S+2nO1QTuZ/JpcYyS5AhnKC+/xYx+GmQnX/TGcm26+yXEBFMJvbcGFKuiww/vF
Mb11gSZQHwWK0JWm3CqLo2Tvqkj2VYuxzPlGS/9llqEMIkExGBKBy2AsG9kqqYso
JWcI3HZww+rNETzQOMXdU6HTL/VXNk/9m0QE/gx8SZpl/x/EVboH5xh1tbYsckM9
aCcRnzHJDzL2BWVextedq9rKaIJR2Vm9qerTWwswAqvZacMcPSqh18c9QDcC2iXM
/PdZ9phtSO/40ugllLvhOv1tFuY+Wp0WzJGWwIPN8HyM2stKTWB5LecTq5pOPk7q
9QYqjifcgjzfkLv/1bxgRwEhJDI6jJ4BGIbze3XjmOifGY5iu8weO/Su2THrw0Ww
6qGV8rlGOmYl6YhFOmxMWY/oYPq1qbWzLWmy3gQ/3wbBWaQzbg2C8WytzbE/7OG4
1FjvnJBgSiadaxbsAlcVyDtuubfr0ZfHm0Fe5Vzcqw/tRQvwaZgyGspyKfnSSBmM
dPu6qnZ+bkY67XOSngvyvpQCXQ5J2PrWE8UUH6BcMbaiikCzamiGEZ8/j8X3XWf7
x8J1P9NEdtsEUI0cjd6ZB8t/g8rHZoD1zOZwg1PtfzmHhnkiS+Wo2UzSeVY+A7L3
it5HvsdWYjUX8/FBZvL2MZHSKGkFM781pr5Xb3KRM7Lx+tApnEwcNMwEjtaUb1sx
+6l1AdOBqHeSC0AqtoL4nwd2ij7EMG0M/FaNfDfc9r6L2A2BYKoL6Gq+5JYGlssD
GwC8xJyopqZLYu9ip5qiOCTckOz8dr7btfo585KS0JrARvz0EqxRN/3wWFQBiR/C
YgHObnqJXqWYcKYGbpUZ65OWNYEoe38T4MQrZ/te8UhyIpTxZN5i/h9/FcZOI8Ts
9P5oYk1AGgs0MuQ/+769JOc9Xfi43ZCuipIDL5ZZjLjRc2/d9D4wM1R70JOY3Cq+
laSFiEmsFZ6md72bdigJggjBVYna9dI38+/Qslrkeqq/RiI8+v2Cc8yGdTyj0wwb
hfkYseMWW4XeNZOQ21OR4mM+/T0oz0uQeMKPPddLEqkNu7zpQrhpvCtO3EHSmJkb
qM/pTY2yNIGa5Q5rVbo91otsPFtbeSgQ0/bczoHkqx2l1ozq+cWUZlFJjrJmhk/e
2o5jpQey2Dd05VHzHUcySm0IlODxiSopoUno5Kinhjr4aKDaZuvPlC8mp4r5sAz9
VY7lFUrpgCx4RHeO/aFZRvibkn2AFxfCd3t68h9KIw92LbHfmfbJWtATqNBnlH9o
2sV1qV3Qlail4Q+eiJN2BsDqAPbdoxJ2NX8vsKaWZ4ABjOF9SP7MEZm3acj+6z0S
xJULOMUFXB2CgA3gfF2mLMJbBGS4fVtRFugpO72YF1d8BEOV7EXhacKG5unshaea
WdsQVoy5QyWbEe8rG2v+Gpv9felQEQaHEKNREt1g9aU3LDacTqbI2NsPIhp8D97g
l5AOiSM5w2QzLl0jrnNN2oCSDpqDCoQEARTBBMcwHtpaJTekrRs4uejw4QwzjK78
/+zXKE6pompbgKB6fegFrlC/pHnr6mgdAOyNSYeuFNmOyjjvUXEsjkwiy0brnpah
IRiBi5qLqqEKrJ7C3JJ3V69pnjPOl+9LdIozpO5u/JuJessY+UV7dIjGBUpAKRZY
3Ergw6h1G4irOLS1Va9yz3SFq834jz2EwI5cmjSZ6/6lGFz1sHuHw+en1r75zFcm
vmkQ4zaw8eu24VZ23RqkLh9fNX4xg1K1s7TxRa+lU++TNcEVNjjQ9rKP6Sq04G1n
rR0FsUELLHqVA9WsqL9ntSViqQAao0t9hKMdhlNzJSHF9hzomADoORuzQjXBvCNg
UstnnmoEDNl8p1BDoPHXbFaq0prqYmlZD+2W/vej2DFILkjqyW9H7+HXfAdB6u51
uGXflXpQ0UNsjs0EVDMrGJog/h4vLEq4B/u2EbUlh26LDao3PQk/iO+h3+psRgh9
KtY6Zw5V80qNt6dwWPAa7QLM7mbXFdpNOJW8hKCJWEBwD8DkSIcghpjJu5dp53Ux
Rkk3/j4N2BtkjCuk971e/opx02WgRPLqqwUthws4iiDeuZVJEavQWlpMVItAqiDM
+K2dGuwcFGXNJv8QTMGqRcv0Iyp4Xu68C5zNRqGIeho7UCr4Dn6MhQrdMNpoVIrX
N5ltxE/mIcwvAcmywZeLchrlPlMZQ8F+VcguJjWz/dKnncPNdOdvhr4gbHbWWKQl
pGEXlh7QXhMzaaZ9zrDzp74JDB00ZnmAu0TJehwxW/dub0wC28LlHik9z9nWW1ta
7E+vivHJ0j2HnV7hGsW6J7GYcvIkMasHb/FwXYT7AOr/AQdEB0pE2Z9Y16Coxtmd
JEFFWvWHMxAtGsL7HHeAbkfLD++8OcmdHKp9iFq7PPD80b5katghDaEwh4+7iIzX
bS41wxdmwVny3Sikx2JOzzbSSXsuZRWcuPwPj60WDuL/FWBhZCk3PB/sjMsvOFac
q4TiomA+fMxCRPIfoCLdo98pD8vGj4+gtIlDkw/B3g6N0X1H/CRPlIEQdFZKBABF
fp8SLClGl6TZv6J8Si6xmKfhZVVVUjJaUTm5slz7KsSS5d9vfHU6hWSeMV7//MdN
CZlgfYpD4DKvaimOzdUs1506tYPWjH+dKw5EGs2hi20QLNbaGwwVMtXYTHJp6TJX
CTxCfYNU9FwbI9SuXpO+M9C8CuQKtAtDe9pEJkMQloJ7xdnfGmW+RvCM531bkahk
mOshOw7un7luNwC1IOigmh35pZE5H7lSKqr4g3Hm4fKuoaNcS09pMFY3Lo2Kd3vv
4uKOpCnDHoDEWK8N+svwON21N8SFTyM052rrN9jtcy0IaFjpjmbl/8vw1Tqr6Sap
722FE+HVglkvReXKaxNuBBsmJngMK4bfw5Sw1tml65l3sRPEh8OGsXY9B+h4UKmO
9A5vX6YFK63bbmVDanDC/cqmEWseQXStdckKhuIMIEyHPIIvHcrK96IuzjNeUPoV
3c6XBrOS5fPo0WSS0f1u2oX4wV0H118kAXkoxNInsQ8hPEy/Is8nZZjPBk3iaklt
sGzLKezXWv/dSd/AdO9ux4bFsKl/jIGHFG3aQh1Flgi5ueglqw3HJMuvgx02dxyW
hxacyED27/J6eiT819WbP42SIhDul0ZKNS+JLYOqKAxiNThrJMKGeJh0FYNFhuAU
Kmjbxl3gDa0Ia1QtYjDF/nSVCpVHs0IbimsNoRnvMRUUcQjrNK5LitpV+z1w51gM
KDnkVo6y8/Fu37PPRBtD4fqbc1lRxzyho0TOF1zFyb+SVxqHgdX4m+BJ103nCeK1
z/udATn+R1GNl2gBzmqD0UWmOhgI2rg+OZFCs1fB2QDNpmHAsePOQ3Rox4MNIpTS
LCYc07R/L5QYew/daXlVL1A8o1KbFF998UBC1eFLM34PMxwD6sw2kG6WxD6aiap8
QROQp+shL+Rcedityoxs9JYVDTxN0abseI7cQij2fDZ+GVyJT+5EY8hlZDG/tMl5
ww6m0jPdWNpw8OWQikE7N5i64JgFsfXI7XJHYxp4CJqUUtSCpXxJXZvq88jTZWaU
2ndTPaf3eEfx4/qT1TyE8HDy6sw08dtJ58cOAEXq8RqqlHJAcXUZ4x7Ht/MicjOz
Do3m9DjH3xATR98uL/KWmaQF8VqhI5g9up7h9ArSRMQ5REwyxMbj1Sb/EBYYx0Ke
i17d4fMzg61lyK/RmstM0v6xBIyBVQBLpvhhrol7uAiH45SoDPolNxTkZeKiIMmA
INLypmzPFMFG7GsaS/eQpl/3l51KBy+qLzDEMH3+Rzmf9MDPLyniTSGPJvx6vutX
cPV49urpE9gk2JYvhEfaSOjoIMwKbluZuL3EOJ9b/1usNTN46GHvZjHc1GaAeK92
R92qK6CMWUI+JEeXsa88utWH9zXDjIsLIef1iTJa9sTnQ4V1+NNWJX1TNWkwk5b/
Sbc/NPmaPPJa6gPbLSeQbPfE5NRECsiX5KQTKPyhXa0rAykYzUmfXu+DASBie24y
smm1RQ1YtABFqx+jw8hdIPiCAUMzTFue8tR/ORi3UINWY1aBCi8J0huhm5VmObDy
A5YlQpsuKw9WyC82nYKkXSRIn2IAeY84gfn7tDcte4OTQ+6V0mKMqFgmX4gI4Fq7
Rz5bE38CdAXREb/QwI0Q77B+/GiZmfthL2QpDUmhowsGkzEzbZDN71nUlWXN7Jus
JpbSqQ/p1ZqK/ysDI3gq/dcanUtUW3Pa2qN70eqQ/4vz/82j6hDm0QYa/0IkzdNA
v8aVql+CCoizVeT+iELvbsEOg48cL8XQ/Zj0f6WX8GP7KRhZ6cCr1ZvM/uvwoc+b
Vs1XO2W+v17gy7lLcrNtxKta6tjbVZlOGBsWuYZ8EObzC0bv8XShAjEEUiyXpplc
FBCSweH/Q66ToU6B1Z8pexge+w1eipanXhTTGEMkZ7RvbOoI3/M8SnQhCSTIQzfO
c4v466u06cijuE3EkfnT1zo2kxl2ZUGpwyEPla5elX8QtZ1Us5PNdWsIborUNfQZ
SxrR4eMB0yTNsgbthd9YIi3aRv7WyfcUBL5n1+Qg0JarbZWa/2JkvPkDX+HHGHCX
CWoowxjuDsR2jw0wa6XYeol1DoYXdX68jDRjgI9fuFTp7Bco1Q6A8T4pWuAZUlCn
c9COGns14tQ0HbTZlocBQ4Trg0QtVEgoZpH5jac5pGVgsFcjyhF3BNtWF08zd5eT
Wr6YQcZbInC/DVqfpWB38AP31mgLbLqdrrKX01MuP3WKVnojCqMt/Tzr5gATvQnB
Frh5na93uFlAQPz85Z0KvyVvDq8ekSoaJszYtwDHN2j/A4DZv08DH9CzY9A8ArXM
FpLA1c3pinAhy3hVCX2XIVlct/x3Hh9fAqgZ8W4spEXUJ/binXqppQTka3kFfg5R
37vHbNCVH6UfrNxaukB0VQ6ieqemNE3Ym4STpyi5mYCQY92B+vJalsmGmDGmLq/O
M93Zu9uEwDjyw0u2yfgwNS+ZE9154QZ0IVDJHANeYNV1DmUoySY+T/h4wSKGL0zk
5UcdVGzsW7pf28Ycmn4vO+11lH+zvZerjzTZfMjKSq25C3JoAejtr3aRAy8NQm7i
omNJftArrXIhwZ8HRwyQcjzR7PBQYKO80CPKgvjs51JvCkrfUqU8yluROJpRyUs6
JaBl1EX1zreHrv9bkKUDIIgrrLKS5trI0dF39iP4mOD0rEFLHk5vyjr35Vs6mq7a
wcyPMTcoOEKq3sILNgfzXdO1oMxl0iW++7zqnLFECSi8CRAY9GVj3DzpdxB6vqcj
r9dtI5bKs3om3TRmX0Bz3m4/uSqD9ZA1+wQEQ/EPVfGDYPZkl/ZWokFM1dXK6pEv
yGjal/xUX8rej88wKtH2W0A+zPY4Sh+xrFc10LBBz4abNgys3W3abqNXp/plbp9a
1kQF3r5iku/vraToliiEmONna8ErQykg8082dZKxvVWFFlDSK9kmyYCZpr4AnJSa
wXLhKkP4aCAstbkuwvdqQcIFRvFa5FRYTyUN3WEzo6CsgNmJjBQQSDsSE9RbDzuL
aFsd/u7pM31hq8wVLeTXJdWYpulvxlvPUN2npKhUInSpfmq2/PcJ1aiKR3e5+Ksu
FX4LpMwmd5e5hAbYnMMJbEXopB3we3TTrksrLv0tNmJyDs1LHrs9Wg36rbAbPUAB
HtfhkLDvpXlvL5zTki6GI/0N8ZTqt5Wvn8unZqIRtGYSfHgJ0WYylYnC2LVReLOY
zawORGSVp8PdsS+LDhtk/+rZRcD8E+LCA/91yXk+PnuhAQPPxr7cBh614T9uP4/H
eMyx4Tcngd/Akw2peVjw6F7nGDfnrVsotaOGVAe9+YI6hvX8nAzIxmDoilCIrEcw
uqHgw5TLwaq7HMY9X0QAT/63XxEJp6FpTLM5fx45zRENxRe6R5+XcwCqEk2kMFva
f+JBI3Z3CRX+uSyXjiOH/J+8XvAKRimvrm5qklZm6sUiOHKVsH+5aItk79kJSewV
4HHt05zrvuMFzRUvHG5u+Osf4cgpvVzER5O6hm/YcNoqmMXn8W4CZlzLmJUGA2HP
HNweSVpZCOFziM7ZVOZxZgo+IAvvkv4tV+bd7jYyC/68+L3qiWy92F8WLEihqJTI
BlpFJEvkgkthMlM9wEmik5bAy++g4hOZg2EzuRJbw5IjcwqXGa8obPUvb6/ansX2
eH/Y9YlYwBidjQ8m4yhuL3oZcEglS+/2ocmWl03J7fPuGJMDqgNhm+uV4WID8EgH
KhqDjFawYbpp+kkbC932t7Wx2v30rRDbXqqzQiZPPiE7WW0CZA2wXxx8zKXhZY6h
zRPMcQ4SfUC9AL20gAIdaXigQHDbUFT5WadGtnbUMlQTym40YxXJrDdnDcCIpjE4
gHkZvVyIhj91yBvNzm+pIDqrK97eeBcu/WyfUTY5NfbngpHwia3eyVnpVCZxTFOW
gDkuHiZxrMUeni/F31VQed1ZWVHtBUd8KbkFRxy1h4slY4KTazh/wb2rbu/rgdsw
mz7BEudnQ8DqdkEMw3i1GXOFUb0DegrPjMkpVLNa2GoOHCTite9jakAG9WHnDoBz
q/uVfNajyONEAG7zGIk71m5oknmLqNvOnZMswwSDKlWNzwiNhINeXcgRV38ugDIW
apnRP3JJG9tDF5f4iB5fAj0H051+ui9cw9GQ/1nh5bdjWpy3hU3sEVvCFb2qs/X1
B3X92Cn/IfQP2LCOwBa6RhLU7iAnc1gi39+cr2zjJSB2cN2xIfXcop+wdX6TAk1t
Atnqw4csx/lz/jujGvEO8D3YQvRiMzUWFkbr/sZMV/o5UpHS7OhMAIVMGob9B6yh
GXJwngCg4cGWs0V65l9YmgSUa/HQ+x3sgu/jP1rs9p2sgrSm0j1abcLqPQb9Qi0U
ZsaGzZsprj9H+x+nQSfbakn9p7YmtuT21OBKptmVuJi9RY5Rrtxgu0eKd33tqByy
aIX7dfj/fBOHzQKgI+ar8UgbeO94no2HxOARvsiD5jj6kRDmTY8PYQhT3Qo8/qqI
Xf5rpLvaj1G/96VS5xx0GNi+Jx1Jvlt4t+//2FdqLVthrsHTZDlExSPKOq1bDCNv
fityCXtfT9O6yMgWwgt+ksvuT8vXp3i31uIWb26q5DnKv3cTHa97MLX12/qWR1av
TCqMgUUWdB/1ZA6yXa0RurXf4Wiqt4I9Fqs/lzjIlxCoELXdG/4tubIJamsMFNJS
2zeYXNtydEkc4nhOWLZzqb0gy2UC0f19RphQHCwm/UD7WE1JHVhpS1PPeouyc+K+
ykUWjOj/rIRZssu4Q/jBKvfEevqKaYMztIckjZalq94jpV4+EUITuqP2yH96KV+C
1dU8lN2wSiEcNbNHM+ILTsQWzuM5cp68n/5S7Tnilr2a9LR6HLyEgC4iWr2hBcEE
yEqsxrFR3lkWzKIdLmehpEIaHZ8mbWGUKtftICSRtHbbTJrZWtI9cS16jyprXBfd
fmTe+vTe4sgj+mwW+OegOueO8tTBX76BY1wLlU9c5E8zsHSMBEXz7nKfhCvgaAFd
ghJqDrSwNWIsy5145rgvS3BSrqJj1BGQI/hB8594L+W7a1a299eGSkVfiIrAHpi2
Xb4muAWcGzM6pWlnItYRiNQe5rU+/8fvb1jB1jWs8LZDJLG15ntUXmKuUoBzhjg1
pKanndYdtfDfUiyRGoM8jT+EmQFEgbkOpPxP3fXnFz1Wl9InOpYWnYEfXAVLMKg0
PyTWFV0FVrZOZ+aIt13Fw0Yc2I5cN08HVUfZjnhkFO3rfAMRSkAHWvlXdV4nGiGp
qu6gJ+vU63jRfQtFmUeAhkaRxneRM+YUZ/Nj1IaJdZViZ9ED8+lIPq/0CaHjZfw8
jZms5DOBXqPAJpr2Cb/3QG99KQ6ECKpbXORJoV5Dj1IgfX3b5YixYo38cKdqf0jd
FkYF9cTDgknNDnjNf/MW79UAPmgM+qrDYYpRaHjjd8p9tUy+biVvrWndOehUzFRB
gIGr7U6EaNYOsZzYpZFUqJIB3FRQmBtXPXZQGvHmhMClpc000GNIuXhxorr2LBr+
gIbTD6OKAnz8wtowWSuNMuJTZWZEHLF5Hl5/FjHm/2sZ4nyG0Uw1wSOn55qOrP9m
4ONI1ZmGtI/Jhg3MUn7wzb2pGvndg2jkFPrbXbapxQNyLK03YBPiO6GEcdfPaHTU
H4PT5CYXCFYq6pUjQDnDWyBVVCHLhO5rWobN5VVgk0sAzgfkTu6lSlXGE+L0pWv3
T4jtE7YfOVSt6b/mkYbVs+Qtz08CEFJeodnc45TIcmisyPmhufnViPmzpfwBmGlN
20G31ZQqKULKeJtBxlGh5oRGsxwcCZkNXu7zeiKRYbCM5y8r03j8WFHxDYTCofFw
4F4dR9bF+2jncFovOPk1cJ7sNRABg3mC9KA95KTnpjCXnTm1L5Z4quKujonMlpZs
eF/5V32LW/X6hArYEDjlcX1rm0LbWoFwbTjqfMX4ttqRN7KOfNwXYTAm5iVg8gag
jdv8su7KMNgROgUqZz5+K1IhX3Fvz110wE3lSJiveoyktsp99y+hebEA64CJ6Gzj
rtFMTyfncIJSAoOvEIwiGZKI60taru87j4SMfnwktSAWAAORzpa/s2j19+NbmJJF
dFbk3FOryECJBjufBWQJs4KMpO7bGXJ9Q3o36mrhqlv9wmj6Oa6j716gEHprnYs+
G0B6gZXJ2lfJEU8dMapMiB222NHkHRzsGLSeGFH/D8NltgMtT4gN54r+7dwdyiCX
XxSvh7u0HCiBFHm3C6QVU6On4pQVTasG4oR659iby6p7hMvVLRcA2zAI93cjkVFe
hdXtFqFMcFtnFbqFR/WDfOLUCdRsASxQavd6H5kULZQgcGOO4V1A3Dh4KIrs8Q/K
TDbiE4mjMVigtM3Lsz8YiO3z8iQWb6oW28PcFTnihMXQzvvIr6MQDBSh1ZKulE03
A4A3UMmjQ16ZF0k6EKxakg+3ICrPacMfsdWC6gD3+Cin2CII1ISJloIQINSHzlsq
WevCII2Qxxu6992O+MeRjIBnP63OVzfBcoImEd0Q0G4T84g+gMa/SK8bZzKkV9am
n2VxUMp5/V+CoByjoci4YBiryMtRNuyUE4kP/YkgIeJ2Vjw9RXWUTD2V2X0hJN9t
OMsxzFMGpOCqNdT7ObOeWsh39awTO3oKC+3DtfyKU42+XEqMD9m8KlERg0+hKiNe
M6MDbWRo6i/5ttKr8m5ii0a69yEuDD5CvkJHXnAVbi9K1M4/KURiTHYLH16pkfpN
N+WNR/8wyNjjlX9JtN4wHp2puuc7IHxUjVLsWb+5q5vegKV/LEpYMBzrKTz6DNB2
NOTTF8GaT/l/YEvdqH6+hRVMZzERjYXTbKs7qPO+jEGIXaVKqPq6XlkXmlsKUQw4
g65Kq/s6IixSkt5tm8jBxqUc4mDEYnUyIdX8TcDbq7QwZGpbvPjGhSc+2wZ7VIqk
8oVI81r10GT+XNmNsC1IvZAdIQ/0znlgHrNTF8EgrGuz4Pwf0S/6ib76ydYuMYZv
tjpWf8DBMEcz+EkSrjMd8aGVbJzU9Be03pMNyp6V2QUTs7PoovxKgoTc3PhN6Lcx
iZY5xiw3w6ip7kmVVR3yPjveP8V/mnv8YOb/DOfHf7L3qnsvHu1rouNLmlj0dCKa
U8TPO3QpAXjuDoBJq5NOUIpHIZo+36emcnzPK1Dr/+ZaDnD+WSm4eRJtfVPAqm1N
VMSaaaiqdt9rw5Pi5hJw/6si3H99QoB7+e2rbSqZT2T3DLbCWWEe7ZgIYDBbzQFk
ZwCfIZMVNK3zL0NGdcsrmDETWDorc8rzW9QhtBHx37IPa0ftqTYx9Ou74tYirWWU
lyyKu/eM7DLLI/9+jlQo6co4iZGQxwPCb56GJyYkllIkJPhYyHjh+xFldaixkrZH
lQQ39mGu3NwU7T4M7Ap1yQhJgTkQzh3zDT4unLCql0Ix+lC7s7nLK1gIJjNwIS7b
fLc1KkxuFRyOsc67Iia86MuVYLqarIBEzqiGtV6nLCoVlgEAVYsvjkS6g5DZCdjV
qPGWrnOdn03Z8uT1ageWL1eLdhJ3iV/3t85RQHGaWv2z5IgUqm1HTfKAxycDD9zM
yykIOQfTolHDBGmfeXUfGXvuP80YxZT53dpYiLXmOoikq9FFXp8poI7xdENxt9Kq
jKuu3hIKJnrkZR/ESVf8YoWtcqGGRfhrOhNEQr3Ds8ToRxiGL/SfeemvbNRwTkdj
2tYIzydbZw7LnVMlxWLZAhSbnOdkU6UvKXUuJlbc12+mzIjQwpxM1wkNgDqbLmnc
Nsuego7OplKrpHq0fgzWu2TvICZtKF9iiY8//AtygGt+DoI8IbGMWhdY0JHvzX6D
kNWxtX5U76JkCK4/ciPV0YS77ZicpLOmCyYrTOpTR/A6zU01hpwJFf3HIwnrCgoz
NnrLnEBD8EYI0ZAFo+/UBZNUc0YrUtDdQ8knLxEBNke97lWCl8dvGXfoF5zJPF2f
MnJt/ccYaszdO8FhQqWWySoDdG/VhXKO1ENdq+l3FhgyDfFXS74p4tGbY0o4tXSI
g4t4Et5nZwlVIUPEXFmDvpyIdeDFguNA0GbR8cASaBinAcFNVKK7OOq0yKlVnS1J
FgeePGzoJ1sHaCPjWSuX/BTzbFpIHoVBfEK4sS+cWN7vthMKcypUff8ll6dX+wHi
V1BjrMhdGruAk2rnvpBCHVNYJuzlbUtHLvAlNMqEPdvJS4lGkR1vgL+3LksZ+zwV
9zP9md89SmgmyZ0wet1Qn3W7UD5Y+uquZ4okbcfrqGi3BjoEHxL8Vfae92SRCo/y
iSzOhT+G8x3JPz6yAnmvt2fElVQ0mhfjUthMQ/t9EvWGg/a4SMP1AUzHh8MqidSC
NMCHdthfpy+VWcECNCdZ2E/ClqohifKrBGWY8vFmyLAPRb3vF39GykO615mFW57C
5xLBGf2e+5AlvL41qAskcbut4rKEAFu/sZmf4L3SuEuqaJy0yV8g+B2/UaP4G6id
oWZ6kF04wrcjfAmTLMeUAtp6Xo8BUBX9waWfPzwCUgwv4rkzDdK5sKmEnRqvNBik
5BctKLYNj7ZqXnzA9N5naWkHzYMZfB79k6PkFf+lhlMsReupjdqRnfImFEsxjGqA
l6xNHr/BwMdzFk7r/Ab5l4Pu3vT65nu49ZXGrDrYD76EpIsousoAwZB11dsH7jlw
JGxOufqANDHfeBz0gYNqg2vKyRErRtREpoOV4ZwrQaDZfHP3kktPoWeXXkzA9FdP
Oo1XQGJ0olNoU/2KGjfBUUhWZeDtUhkIqnL5MyXl7Fgcp6G+CbM1K3aJtOYLMPcY
q0oUpE56EOzhB+kNsX1EovUqRVWRYy2u8+e/Bc5+9SeLxb/mcCJYZx/cZm15Tbvc
/Cj7UUV5B+wZ0FhkwA+UT6NClV7bgDlShEyRr74cKe3dVJkI+Ui5SOOda5f195Es
Mns7XeISj1aLZaIvf+bvFtMZpGsPzLcaBkuldQyNx38QFvklU+9XoMRJXT8CFQe8
tfUniXcgRQreOCSw5MLoSotXaxTlafn1wbnwe9D2vbzTj4q40Q5o3n5n3QLK7vwr
7Za26XIkB+cr7JTMkvu4GoG48AraqEDvZ1XzlIkeEoxQB4jUN/v8960Oz/N7BJXD
npwkakt7tZZ3nTeIzz/QBJyU4u0IJcZTmZzPNzwqE/+hYkRQvGtoX4XctPFFW3O7
x0KnlDBSIT4wvh0Wr2YBXAjcgPqgFWVQPNt6oa8bperoJjpFH483TYk1smTQFdM+
0ZJJyNP7LsM0M52Yxqigh5OM1ps7E1P57Rs+QaL+HjuJGBKialwE4MO2DqTENqOp
RHHxoOaVAML19SaT47EoerAspZjUNYBtLxCzR3N9grNf9mHP4UEgFHTn1szjQgxn
nnaI7JLTP7M6JVpjfayf9C3L7UGv2UeuGOJ5IcKPiDuCoalwGHQurUVb3JbVkUnX
C1BJTl+0xdHIvJs3Rr0q7rDug3VXKbrCWRyrWsvBCEBi/IyQqmmn8gdNZkJF46xA
wAOBaV9PSS8HQm7/qMGCf7IMhuaNBC2BrpEHNq3cYKnRwqfgdxZXz1s2F96Fex+W
uHJiT5sKKgmgLeh6Xn+KTQHDM/tJ2pU5YE++Z6Q6Sa0VAKI+HuUXu7a22utjZx0X
fXxc9JgNovglRbbyl4nKdEkFAl9kfZ86dABvjeg3W25gMLD00SrVkR1TQwMwexdV
IkVj8dBv42co9bXcaKjXPeBGCQQQ2TQNqIEGoPNFsysG+cpuddm2rhW+/vNkRvN+
EEMUkIUicW1cs2UuCRfTwnpuqI6gO25JUVh40dbFJygNRn4lc3GdS7qwlmxB4IqP
0G6OZS/ODVS9XTkxncdmb0P2MdOKCfJQbGigb468003CV4GfPJ+koCKaiI3zLSsh
oMrx6wmAddtz/1cY2zagQm6LJgwnMIpS4lO4AZMIJOXFC0yviqDikK0/8Zkt2Uvy
pcAz/K+YnmFzgto/EkwNXS4ze3AXbacY2Aj1967ObC5JP2Aj8TO4gYpYrNBjNiai
rrX9QanMwicnMYO2QpVBGjdX32MLYsTIiWcYbLEWbbR0NRs49tS7HB8P62O5aKAn
3gXJn3gOsvYHUR8QJ4mz9ouESwqrdaSd7gvK7spdBc9r04nce0Z5LDM+IxFjj3d2
NiPIeG8cFyeQkDQPp2oY4YtJifDwDRX2QryhtCQ0OZrCBe6edEbPHmlvwomNUwCk
d+GnOBPr+x30ffTU2H5t8O27U1HV0a2tBYeh5HSu+qLRLcWg/07cgeXqjaVDboY3
QuHrMVf09VStf74reBf/a+z1vJzeK/xFK84Lf7amn43Snv1EYHHJoMzbxC08zzNT
GT/Pl2SOLORThnYih6u8uwy0Oz/IjU6Ur30BtfyaddtQD5MmKiP9Ea/L9jjLkE73
z98SET2M/IDYuwiia1+Spub0nxCX51BiQOyK7Cuw+Vdpwm+QF+i5SBxhVm6FBDqD
CwG4hI8sLxC0rHwWQJ2EdZmamWLrUeoeEmb1jeVyZi8UQ4IxbX4U6j/xZfP977Bp
IbmqnPeN/Xml/qoLE9dyVnRItRPsUB3dw70oFQo1VA5RiGjTB5z6hwTQGBqEIYau
4P+C+9JXSCCis2CAMCmzmZJzsE+P2idcW8SqWzwyQnl+DlAoRcpMm9aRQjqCZ3sL
KA392SL/KTzCG21qlKmCVBK6IW0ZGl1bURJzU7c+hNnKeoA/KRRcyjeMgTLu36Gb
KZ0K2O49xJfz1DH6N7fN89fveFv6jCXS8SyduGFIem55In4tZdz+1P6oL/3ZN5QL
RBqDmA1yGPTxJyzrSTpM7yAxt7JT/b3E3RNpu5ClfoAC4XFaZ1nrj6HDmwBqc/Xg
jns4krLn+H41ICPhH1N2x+a8FhgRlnjSZS9TMjXQVSsYEOnNgmTACNcW9PPGS0jC
fPP00WVicvBp5uE9bK7w2Tef6EiwScw33jijF+Mo2APmqkewidNtgziJchrqW6Ow
zo5lGBo7OwQptnqLrECedt5hJRSsC9wu35G3NEUo1B5BGStdaBm+UbZZi5m9uC7B
VoqF4qBp0XAE/m+2F7k54tc8mdhweSduZpLuclzQf11P9etL9Xws8BoQ/OJ+ZKBA
l1/N2lw3vjugcXlzVCjOosgwUALiLsDg2XyR37/alK/y+5W1/+aDu8TODDixwTn7
DQQGNwI4egDPToNBXfdCqMGvBoaeP3O7WVkB7Gq45Japn1myApD58zs1MfgUwZ5+
28LGWvXhPxlAhQP7wuPV14J8lwk/TwQYEYJfND3hvu7HWG8nUNee1M0rXfoOBUBj
ktuf4XKWbVzFQKtWJMSayVL76AGx390HZ89v+5ysoX4yCIehSyl4jVEIuP4PT0u+
nelBAtlshuceXAdabICmFMMegZWUJbT2r4v6+kVyCT3FjWSeDH0BMf7fjNBPJq5e
QMwArcxGIVNvRwkdg5VunYWCwfM+sIDSPAK3/OSqR8+XltYvpBAPfH/c7rpkfPOK
Gbkr2uQlRvFeci7IwqieqGS2r2jaIsyZhzHO1SMy0i8ZLM9AqVgfhypcc6a0zP70
YgDMtYSCLPyy2Sxhw7w8RJls0QIVqanp6ZkQqbZtq8yDoSCpFYKaAEuODu05tvp4
3ZP3+srkejjkamwOEsHnxSCUPgb13VwbKHg4+pq5f8aYxLNpAnOUEvjgTm/2pTaK
iwDW+bvp3jOcBn9ZbBQB0W365lDKnpIcNMRjpmwtMEsjMFDSc+F506hgS26KjWoh
EAWlsLRTkc4MQYhidfeaYO9LSU0uLBDS1/DtTH4ALtzsZ+p1I4BrqlSLjKdw+I7K
zf2pfUQJ5dwrQ8bwxdayPtuRcc2xeLcq20T+hPVrnNi1MdzJYXcXirxcy/AsmyXM
Pil2r/ELQRpNrHjP6t8wxOSKtiWZcW4ELheQCV8oK8l3kgagoKsUMRwwxLVEuIli
hyq2rmjBjzYIpIBAaRXVfBMYr3Gv35bXtcF3mA0FbJLF4GEPfvBjkSFVfnY/3BRq
MhqCn5/iUthf8Za3cxobGD+mFrh3pvic8mdfIcStqqZEixcSrDHRJHVQf8Ddm0bR
VOSSCxreThjDO7zcoQqp8E4MLTrEwdsLERk9uhdFS6G93NpeNeKndQqKZT21RuTO
eFnycJEDILrBGIehPkp5HW2+ICAIDwNrOlUmH4LGEmq8QfGen60XaV0+hVSE3URr
Y09lu8sY0NN54H+S1wVenDgVuwSWTS7gIW73KVZhZAr7eKTQ37HbaJDGQj1HsvUb
jG0715DvP5foQnh4orteuaDVj7RAcwY6JpDr9wHUPWNvJrjXQtJjuvOpYJ2xYY+y
b7Sy6HUl5ywyw1i+RTMYW9JJ78Z4aid96oNLca21LSS2RXzvByEwvVrhP5ZunJzp
meRwuV+lH1pYtXVk1jP86lo27T71P7w/Qp012i0fPGfyAlcpO/YsOahBkAWp0QIf
NqAnVCmsXkZZ2jLaQxe6FtuF10KN4QOXjA//2+TPormDEchQSwmOpFm8qf4NXxsA
9xw03mxgTuSndnlJM8OYgQVfAtJi+ehDEfwkeZqURYNXF33iXjt4KoIxzB0+ZPTg
ZCNDM2VLto7rvN2+PYk4kfVP0DuFQKYPLIzJQedRNP6PqOJcZAYzrc9SNa+yuGos
91npp2TGErTOMJ/kfIOdm01wvFUBTsDxSQ3oRn1algxiNs2xVn2n446r2ouaHp80
35DPTIlpBvTiug9yHHNWshmQQu9MhO7NvJh4bGhiJtNFEBWd+LEBt5ZJF3dM2q9d
R2OaDw3YCRApnQmzJlRretAVr+bCyRntjjyeCCMfHLI69RKTqurmgyWl3Fc6lB9D
umSgSiATXjGtUIiOp1Q1AUuqWd7N8pijFegp6Z+nysycJnh6dQM0zSBH0QdsGPoR
evESpejOc+D/dNWae0p/RSRDi/oOYv050l/zBkVaLs+rC/G3S/iFSi++xQtgBP2W
ykTDhCqZzvPrx3GZ5HYybkpYd79O2tk69eFhoGmL+ivD+4ssiOvY1TkAk8FdYTmV
gIlXkNn+55Ss2z6UOpGTzTs219MsuG6s9kJ3zUz2GvXBgQS+3SIdwTmnlNT3rwMh
9PXIYbgvucAHhqYN139fyae01zXd1QEd5gnJYet9xdTBm9NsqBWZ/RhCl4GPfSmO
RWatJVFAXnj2xKikBgSN1MWA4U05Jr5akrJBB4aYuj214eg227VCW3BVZzURlan+
pexXtzFSy6seWcTSaStU7Ou8RWYAkOmsKKSfPp+18QmFsCP2KPUgltb4LsrLacGL
TeoamfR8ceFVLJ50FRkdLOAa0qIXmmKAyIvF7vGZ8sUabXFFwlIvs/gKwVbJakxb
ysJEfUA/zJfXXDDYZ3PVP8N76vDHl/ZD515kPFFuXZa0vm2XP+RvqqRJoWRJbJ88
aGCYklFJnnIGL1MzXK/JeW7P2Bf+HYAazJPOyPOYpYGOaBTKbOYqeRu7wsBLWYJE
ACpTKWn0Mdyddg1yH0CLeNxwpy/znNl/jJcmEbMAtLsmQJWxw8/YKK0/t7FIiGWl
SFHI44T5Tzx+N3tHPTaIGXYoioS97VJj/Q9Hpd8M3HEHZQMdkrKK7LXYbPzi597E
S15SIFX/2QXOIgNNjlLbAesdit4Eo4FwIX/63e4YE3YTpekmBP+FvYA1GUy7UkYR
ZALrxPN/I5QlL4Ej+IkFj25/9dMRwFdolVgbgnwx4Fp6di162ts5wmm1GvvkAZgQ
GMJb0qhOMvg57VkJO/uh8gknDl9ibghfpLQznHUvgOb2J0RJmneoa7I7dsYkt/rd
myvGFgj5oEcPiCho1o7EPcE/VcsndTX4fylMgy2uwMyrmgb1j36PkRhVDZSHFYkU
vU3KnlTEV4FH9rpXdCIosRU9pbhC8SdLU0+uj+l90mN4jMfdv0o3PZc0EUS7ETxl
UjSKa0aogYixv/md/o2+E0gci4ldDGBKQ4TguOI5rrOxybSGlbBTuaC2dZLhguRn
kuA8wFJ+sCWzIja/AG5LIxd5uE1c+L0OjEa5s0aKbW+4GHHw4aZEdsDX3ORly0hJ
mpY5OeRL6xPIGS6DcTIQmdl+zqM1AM6nknd83MFIv8lC8UkUO+idU6QTVkkBdY2O
OBElpT+5ejqoqYazyA9h2m+/u4Jq3PZlH7SattsbUIcx0S9IZgaL8FYRGjJ8x389
Xqq5mK1/J7Yy9EHo2oh3Yw1dK1YcWFpe3D7fgDLIKOdmL9D98gi+F+jrXae5QGt8
OnL4gIXbEOmUHkRD7Z0lsQI7SvC5AhTQlKkqfisn7Kr9G6Ce9BmWsLHNU3NUUk0G
y1XBYTibF8qCIk2HrcS6l71v0G+ak8fVY5vX3xuw/ti6eoeWb7glNv/fagpIbrnR
M/UXtyCwKNOnkzFlNw6ANhJApj46v8RmgWhD4kgLF/YTXHldTzQ5NDUaYyfkbACB
SqO5fyo0ROtfaPKgrc2dhaH16GyaYwgxKXB3AH+rJW9kTVjv2bPolJjPI7ldFfwa
qW1ZBhTNETaee+0V9EueTm9qewwFNvIWsNIdX84d5zpUTerhNf/6/TE7YnsTYUAV
JBeZeyAoYU46kyJ3WqFHNstgSWsO5Cs/ZWbzdNfpXTx2ZdDlbtsaHt17Jl+nhL3F
5++Di68wRbwhIj8nahI059mQjKEAUSM8l4JNGFRkNFITlrKnoh3rDeVCHt3DIIRH
iHZ+iq0fV8E4h5VYzT3TBwNuVYmIrLQ+6YMlXQuIB4XJgzM8E6+FhlhFWhJ0uCL4
m13tpqbOndB76KSkGSszS9H+spJ4jutBxjamWP2jT7zY6ZF+Hbzye2Ujy2BU5smB
5mTFU+gfn01VsBGgDJ8EgLYiSsoNqvJYN8F2jMjksGyTo55u3Urbj/uTqtCfbsyP
rlTx0O/CC7VqUXWZLNXSw4FiqbIvabbJTJ/k9MIfZAv8U3xE3dB3noItiDV2GRbv
z9TQJ5zRSCpzmw3IbcWigqHEIakesAoz3SvOEh1wM68qysYQB0TwypT+qaEU6a/Q
uUqjdhxr3Lr93o3gwh+Fn7BOEidvEDqtcIGDfm5DKfPDLocrmrXML2US1Bf/LU5w
Zq5pcj81rNZUBvJabxMVqQepIHXNaRCI1mtOSGN4Z6GHCsNIHEj8dy5sN16EqkKJ
yJTG7T8ergeV3RvsGavOrzKJRm1ppHE+T6Ui65trUKP94D+COm8nDD/imowjzfuk
6aDC0Ks7gakQqxGS7i8HNmBK00KLR+eNFmGKUwd1216ijhiBBDAOaBgQpahJEIvm
6SXwjJkkvrl1kCLGKasjJ2dOtbAeTm7ElgysZbGxLd4KMbulCuh9XkijT31Z1IEP
LrmvXUddFs8HvMgV33oHdlbndiOmZgDUl0rBmyP/bDMTEBYAPsE1tCBEnUC2mIeW
J3dtlW2FlB6mKQhASM/wgk6HU3MMNyj827HwmKqvY9+o9EwrkKJzWTWTsX4Yd3OY
dNsVD41t9jE973TZ58f/T6lqVQ7RDXMSe9G1TiCKucecLI60PunKy8fMQasdWg3s
532XntqjNMPIW7o6V+vFoIgcp7/16t78NyU+ODM387BozUNK/bdB9z40VCL+J1xU
Pkpc3rm/F8UTaIeUKl++SX+8j/PLvHEh8Qn1onyOx0+c2sAu8EIG7E1fMsUE+2nd
tVamB8JqTigzqjDSYFDykwVJ4n9UzTtPlIkUiQiAuw6bPD5lxmctcx6mjvRkKc92
pJpE+pvm5M+r4zwsD7WyyONKnGLpTjEFgl7bHr3KVNjw6Q2NkuKYY9clI6rwehpL
dkWHlGyIMpUdaJuMD6VBJ0zkUFCzqZKoLZs7O/ExecFrDBqOfF7Sz8FEza9k82G2
ljlwN6MafcxUPjAbN6BMADKpLJlcNtZWA/nijDZGdP5OXF/erva+T3nP5U3iHBZJ
tmTbSP1UJudEmxYZRj9TvgLiNLBuCMeA+WjOferamIZXAmACJ0gfxJCm89cze12M
C7veLuOHB8OAIGPkx9hikPOygcl30re8SZ1AUlcUbH++msplgvhmfWYXYddVHoPI
y9AezNJw7ZlOyBv7KfiPj/m2l5fam8CAdgI8Lt/9GTRSrzOM6m5eCT9g9wC5rKjc
6EW1P85VPcQh0jfcG9wOeY99ndqxftxhLXm6gFyd+QMAcgbAyZD7mjxlRVem5Gkq
V1QpE5IG5Ed19zphPul4Dql1ap9Mhw8v1xBzRNip/YY5L2ncNX3hWsTz1flsSbxY
UjmQenypz/Qm/U85a92Bcmk7pVAGTHZVt3srRdsD8jPmwHdSbyeqfqTZ2r74+Wgs
+a6HVId2sMkTtYmQS9VjHQqDEPi0PGSji2qksaNFC1yCnVzbkoFQfwe/fsqfTzm9
mglBoYNbptlAUOpXnChF7Ovt3Umbgnvpe4jjkjW12yzES9NCi6zxrvqdc/qPY+wu
1wk6DVRihvbozxd1/BbRhb3U9mgi0nWoOFdDg7j5R+/5HC3U+b8qpvpvlO+Gixc+
6DELxPjuLC92B9Tun6P67P+Y3gZ7qMa+i4ym/q0BfycH+WgetPVqJztFwH5WOacS
SdddZCIXbitqtlFOwZMH56lJFT26ZJUgMSXM6gVFqnYHAcL/+Cs+Fp7J1FkPN8px
0+PeQo18rn4Xc78rUyOfdZfMuGpVkB+GUU5URqHQGDQuI3tPTo7BT396T1r4Uuwj
jXotcnTYx9wYjwnUNfPNjBHPI8bMFGg6PvLpsLB7kworJDb+CQum4Bl/WXBto+36
N3eddNxL47r/KRHfanUD+xPZfFg6+RYK3GhQvahaGdA4/GY6JA8ix/yFBpMiUFGl
m3moFVhJWmJYeMConOXcaTuTv9MUS/qU/tlxNU9ijhZutCHYiR1FxDmxAfKgsChm
UV9qRjiCG+s2WuFAycY4Qu7rSh+WDunxoNrcLVjmxai2Phko8xWrZlM80/i1vXI7
x7HQcTYiYFNqzj51afgsxHhXvKHQdVXeCMrDUaoFhXz7X3U31izKEq4iUanK9Oht
Zuqu9zsJuR6qWQhm+BvNOeBT7elxbrVVDuEbk/UQh+K6BsCM220jTuu9xTCEVWd0
RWv3i/V6OIfXsXFMb9o5SBBcGuq0QfGwEmCLhTrFfPI8OSyo7hNtCXEKXo3iKbyo
ZzGXOzkJIZjH/SsumZKzaQf6GJKAAuYMj+R381HOBKnqaHlrsr+QogP4Zlg0DZB4
cW4xZEV+5ux8ojj5SNX55p0LojSnQinNG/Y2ACu1v7AT0HrpjeVlFN5iFtHS/v4b
QTpqBHV2akfI3VIUpg6MfH79VQ4MQ0PQula1+laGNSBQI6JGDHeee75gVukC04hy
/rx74+8CnMaCxplerMxl8FJ89D2wM813GdmunhQs/iYEGSX1MUP9YYoJ/sD/eaBZ
1Zr4o5kq72VXkus4TNcop0715EJJcHDWiVM2+LYWbh3ca32jWXg/ARbysv5FVN9l
w0Ds/PT/F6q3ma22VS/moMeel1Lx2cxkJYQyIfEKlXlKcLFAa0nljs1enyWvm768
VsXfQ7m85RwY9SzFZpWSwFvcMDv0YhoFBZ4RpIkxg10qiTlEeKdH1DYs23xrnuTh
6LxeEnjL4rlnWV/6Ynv8dSBBDxPy2yGfp83B3yWcAaqEWsoBvN2Gq1dnE5Zw4iMc
j/oqxFbymD941065Va3Xgz8j6DNKUynU9UxCSz4ic8pq/WpLAHGfHJEDg0UdtqIh
bWp3WxniwewaNu5B35wU3g3j6Vvt54MSL4eTTThcufJGP4c04MkSrZa+LsYkwOMg
gsOc4xk9+zwhBeCZFRo5AbrXzikkVWqBLk9tYFeaPYbdx7YBBmx3+ZulY0sY47De
OiL5NWPOalLRB6xpNb49bRFY5nedz02oXx4mPtCH7+gfrOO0RqFiok6IBuG51cpV
ogeq5ppbXg/V7A6bPPxeyUZi2Pf7b0/Gg6fE9hxZxla1A8PoEcD8YDV8NdVS9SWY
gjUlgcRAfvNCynPhTevZHTZiq+u7WlCq1D8cvA+s7Pr8/U0lAEYNVZHbwtl1XoVg
0pkUiW2FA0gxsEE8oHuq5mcrFLcQSGSdZFgDkwOlKFBruLnyvDMvPF1AXlrXkrwK
KZ68Jcbb/xFGcGo0R5JOROu1+eyiL4vs4LI19eL/Y7ppUuxWEBhGAOu+r/1C7/Rj
mKu2UNzoXW2k8VR9EGsRhn2vgfGCZABrLDggqy/4beNz0HvTrsqY3w3Q4EIwICt5
HmpUzWMx6BgksVNEtcZfdwM3FgpXuGLyuB7zLPdkPrHhwjs7D8AeQVvag8lSQJNk
thbEXEqzE7KufDGb+cM6J7rPJlQMIZX/Ay4FhjhGXm+zJr2pBAVWozaaAY9Kq+Ut
+s8YlPh3r0gqfbu/TVLkRDE1ascIX7j4LDor3RNjohsJXdcH6dvxnm/Ph6v1YNg2
7DguBUMgRuLOaAeEXQBcx7GwusI22DPEP+IMdGGCbyeR0liddWdznNQQB06MZYD4
iSPc3BdRJoQ5/tnu9D7S/uGvKardW1n2Eu3ymR+i22Ahn5z/p2+eslihtjQQ5gGV
tLTM5nhp5uwnXMe/MznB551+0uWUZ61A7n0aMlfSm57DvEzHVwQufptOC6hnjU9H
/caCartMAno6y/OdFgY+isApRMSQRJruC1ZbynwB4okd5QN5FTboKUMbTlA3ygc3
4nW89Y0Klj9bVmznJ/+aw/run7zZ4/lM8fA8vMrX+UdiDgBLD0+tlRe2ngk8jq22
tuzWt9qoS9mhnaIkADl0aZR42UdChMtN1mIAOjdzT3R+o/RJ1HeJNykaVZtMAA/1
6rGr9ZZDgkWdo97zCtZLp9Hq23Bixxp6WO5q8PzVUrfJzu3IwjozTyJWSwZSOCiY
avhVEc3Bf8oCS1ynkFHifTJXutpdfoTD+oXREixEG7z8PqzjkIP0tLgPMiwZdsxh
7RFVQozGpnQWkztNfYbg0nulOp5db6hDGwqH4slkJu4i9824aPDPnLtkwLN2TecK
ZJc7leT7mtijvfgWJsitBoV7qi1L7B4EGtbMmX7kePXiJkYiKW46JYOw/twPJa+F
3G5B7h894I6Jret7QWjzwiIYYK34DkgjwpyfbjBLT7oGuHJ6avUdJJw1Ww+BlwLx
IgU2grL0dzuCZWGJPzD8bLNLZqVcJQODexeHvrQ6YVqDTcsasB5Hk7vWMZq/bCTo
Q8i59L7sLjIhTX8jMZVVBcfB5rSEIgBtZTp8g97RtFIvw5LbQYbx5Qh+qXZ4i7H9
R/BDLTUWL7lRua6jzHCGlXLlGzN9wTUUSDpR9hn+5PLP+MO2/75Uj81sk7eAMGqu
MROFtGwP+erAy9wgpO4Fuzs1wtY5x/QTHK4lMyTA6vxJn+WeWtaqYfr4r0PRhpeu
Sbpfe2oesghSayYlkH08bi8hK3dHvza6YnVp1KjTthkVnmxp1OGVELS+Ax5iJzyI
qF0IlGrQZqc4hmyCWGx6gk13zMTVyINCel4zxDxNGx+hYNQdOT+iMINMv1vrKOZJ
qTDro7d0iz/KhFf0RwyMcKRnwUc1xNMtiKouPXjIhQKNv5VuWHlMhIxwL6OFDY2e
SQtI3gl1moPoT1HNzGUtDIfg9mqF4vpi9eWeVLYjbHDVZsfPEVWhOrxBqmM9ztG3
XR5tC3t67VIMdSW2NPyATQXo4lMXP9fz8SW/Ob9AzHWSTKZz8ECm+S9yWaA/tmqL
U314sQ++IQ9qEia+SqFI1A7meK7TkdlQt5O3++nO2ypy/+Fg2k1TDhRM8foJko2w
4687i5NF4hJULRaoWiiGv3pITDrbRDSp6WUbmVkupnGc0do7Q34CLKwGRli6bbhV
9suteZdvkQnuUtbe3SaaTeaDRCjDByzAlNWvsvy4wlBZ16BSa2Y3jnUO3xuxZjBx
vbD348Ojf9cEeBZXKLnRGDmc6w3tJwwtCDxCWpLLd7+87lu/m0UyfFidH+b9LfG8
mzmYFGtqGxnDRKrm0lGefpamCVDyfSc0QTtCVZ6wpL6IA/ZFdlI+xrGvhl/ve4PS
iJyGLbyExHGIEgLM9CPqU5KX/0Dub6K61wkZFF80JBmFzp69NOmSfddzUqG/sT8O
vAOTwI1z/1bCLoYZVVG1NWEg4YAZCe9yHLvIMORnvxvW6b+QvINqELm3bWNqNMzl
IvNlFC2yApCo6m+mLUhLJSLB5Ho6cYNKekIqZw9Mc4Glz27zdOJqnGJq1Y89I/L3
ef/RRTvIJ6bjuFtKsedeO6YD+2c5ZTEXXeoDiy1AfK7lEV8Q0T6DUaaq4nzTk+Dx
r8k3HdEbaVrDV2bp2L/dhIEqdIXfoUE7CP9Hc2P59/LzRW9RTbfudS1ytAk4VgOV
v9mnbaO+Sx79fV7pfBvMDDR9+tBsf7otKGY7R7OWMQD6nKVi0SCiaTWOyM7DLunK
u2A1HlOY+d7eBGZmL+///NK3uHv/8SQwS7zXOmSwvLSYigV1nEdKQ2lfO/11q6sA
23meD/eFjC1TtoKJdU+Rgb3i9AZcSn+LW5Fk4JY0cWDlNC4rD6bWzgPizhD6Kbx3
2mfdnLCVHb+myO4WzEgngpj8KbjIaiYXhGRQ0ckOsOWmkprBvJldzAAAQKuKPWsS
oQgRIKJv1LKuHSgjI353c04OPhVgNRx50oGeWwl3KeJDUsq5o4sgHFXmRzBrc0Xb
//3FAZq48hD8NSSDUZXjdB5o6jJ0CF5IQzxbPyligDYFVUrNEdov3YFo9uU7qJDV
3b/mVhIfiQuNbr8joHwwDVmP+4dr1Zx0fT0ZMC4K5FKpiSzqDafyV9X8SD0CzDEG
m4+z5busrzFIeW3VhiQWJlY7sU3xEg8FQNEAJrqd0wiV5yXJejGUn89BR8LEO9wY
8yBETHGqErj1x42i8w4YlF+px7IgP9LF1HCODOQT0KAn9hdWGW0ob6eB9UxYvRX8
nmpLbU2/5DAUzATHMU8ZKGBeaCiYwj0XncKsqsai3yEeb5EGMSiNBiEhYkQlJWhG
Zop+dzmpfy1HGzh2urpmy+VRw1qZ2YHCcmynz/I/kGEBTqjtN/g9CP5mRu/b3+LJ
+TKCshL/T5bFPOc7ADY4vXTbAMY3GDe/6Tpt6xPAFxZWrQ/kQx0NHEgzblmVkKp/
fSYfQMVCmi1hcx9AR9sM+c4YHGrhtxqic7vVWS648ghDC/MlJjRBhGxQQa7fEI6Y
OrG2YWkN4vc8XI8l4quYQC5FcC5JsUnAIRT2nj+QxQKp+BQsKitYajnLiLnAsJaU
Tk+mGqrfsNNTbkKtmZUNpJvw3yIoAZvAJOEQJc/xEcvd30EBEaORtMn/xxQiyvHE
DsTViXGtwIVYN5chY+plEDE512ZCjBO1emcw+p/dSU6sQ9MT02GNKef0CUwZ4YqV
0g++XPLV0IcukGsZrv7sJOab0WLp8JojdjZ5XNjp4rRItaiicE+lsT6MjgToNVPd
cJj/u6nq4BjnD71o7BOgMSU4oz851ugewHWTYGefOSBqNoy6OQLyq1Ohu9Z0EgBP
G975+Vr/RFgLSF8E21aJF0qlqrw+Fb0+llq8qGC4aPqeeqECYKP/Pa2AoUgiY/Ao
euGjw6LV7AZf1cc9K20DRAq7Vr5JHPEnDV/BzMf2/e4c3pzF4WkOd0QPFALa3EuX
NlOyPAa3+dAo8g+TvGJ64S2e8fiIt3iP+rni7rgzIPqCad/i3MtjPpGd+ptPBQMD
90Vnzh5eOFEJX9Wt9B6C0GyA4yEtaFOt9GWG8O0MGC1lrrRfiyQt+jyjUdpUsS18
dliacY+ksGYH3dV8m2Hn2flKmaq2i2P8w38DQMEEg1tx5M5C+NCG0GFib0hXwKsQ
7JM2eQp7xJpmafAp9tRX0wx4yZdL4LAx1lB6fbwDHtbxiXT/F3bf1fhpy32w20N6
1lahx1scn8F9ZjTQh6uLz9c3c93VUjluaQz4F915aQ+DNk0EK9IAIiI7bOy4mCwn
214CR/ia8a6nz4YIdoScDqWmpL4zzmzxkvpSLSkDBhLCeBNRqnX4os3G9Ny2Xun/
36Duf+JsD77XzhOH5SFtqQr8yrbZ8m5VV9etlfVeT9P783r7wJJy8MTH882weoKn
gAAh+NRbCsvpqx8L+JJEXPyRO5B8NVg8KiDP8q7NCrha8tOpc7vyokVkm0xLLdXr
9NFwrbYwCf/+7ih30S+GPnrYdrE+AyletXbgQYBwcjn+g1ZGEYdV6FyQKWjJoLEw
KRjq2ELxuULcsbfKP8mqr27v47L3RITiG/ZEdxJCSGgwdIdUAVzX9WJ83EsiiSqT
cFK4UkwYmzQp3qENmlXcxtkfXeIFbG7qI3/XvaD8eefWZ104DyI6dZVZhi/h/275
Bs1Nstt7eomrhfXXsK5FNcrsts8oI5Ca5rSio/fL2AVpqLb8wa75SCy3jVV/xMG2
iJ+T8X45K01jcl/zK5m5wVhJ7dYylMX5MysrOTCNMgcw+lRpWbE6yYAhDxqfcUL/
qA24iTWC5gUfv7u5x73b+luyBHpG9cDkNkCaxJVq9OCXfUd4gACM8ufBOQpbYFg5
jd8LcGrZPPO6shUVDu4aS6HoxAG37l3IajMaSOSyiqofbHxOoDOsGvjYNxCGMezy
y0ohKFs8Uweb1v6zXljUF62h+/z34gxdKN8fdQJna2tfvqNWIHOtM5FoQYzDbFoR
LtLOOyn7ywySELyg7DV1Dz4OzfWsjE8+Ah3p2dnN7lykhBLK9ztuI0z/OWYqf4aL
8lqhqeut+k1PJQC5Ue6lsF1eISZRfVWGiD35n5s3J4hwGPDbqA9q2EZSl3dIH//0
WqEI5+bvJFbVyrVPp3ffYWccjOgFAGzOX0d7y1yJu5lN/GAMd97rSX/6qOhZlxsw
T+T+sMWKSysOBTwWtSaQ3rTrfe657pbUhZXo3uUTGtQUoY1/gWjd0B4cJH9TVPat
x2aQqb3mOt9Y0xp7oUZ9prxPlssu9cHt01rrAxkU8xb6oayNVjWcyN6lsZnHtT6u
p+J1J1j9hpmrxD2hk9SUUWYzQMyksFomD2+hQsj0+sQweMPMQeNCKCgWg/1X7epk
c3WE/IjDJp5boPSeU5Lxx+rPCztecnIeS0g0ZfME7bARiIKx2dLq8PEl2U2iTn63
LfnVOLjuGQG+g5iyFjsWjy7lKnRUg4qymSvJj/eu2zqoFBHzzqyzVjFQac6B3MBp
o3834SZI2QZMuS7A6mjQTFGLYAlNrYEUZySuiHDPE8pXhnjh7iNymr3hr/EoyM5D
BT+JrI3uB0VpZff7g90Mi7jfUywkROlPtSokMITI37P7DgoMInEf7JSdZb5ZKUs+
yfXqDbY3hq7ldAlReJj9AVgc/+/gXi/icItgsKFUoQuJfpthzGRhpGDf2zIyVeDc
acHUqn6w82Dvp/UYm6qFVhJ+vFDUVFwx9W0HiCyBVJhHEPbG+T60BIMa1Y00juJH
Vda2jnAgHrPxV98ydfvFUnpfoTbZArx63Qdaztrvs8HAfDBc9EiMewaH5X06CQvo
Wz/XWtnRPsJsgt+WrWgakJngwtIBICzIExpdTnVJ/P/jhn6FD+R6vKQsM+YytYVH
Xes81YrNhUe8FRp0kM/+v5s6C8moUd7am84dX4/SJ/SnvMKdZbJQsB9mr8vFeJpy
XMfruaGw7iH4j0ZsNgMwLMyzzo76cAN13VzBXUgHmYoeyCMfU/9Ta2pHUyf9hX/D
pVTGkgRXrnIyrY5Y+7JqLVCSEfGQyeUG/IAyLSNOmWExwMDnZvLCnu/n0OB5Z3Kw
1Mm1R0giK6neMPxosiRDoNkfuCpor37PqtM+rq10CSvXMIMNCPN6onoYdDDkmvb3
b1Z02+MWJFjY2lNdIv5EA6Oa/8WIifnM6fhtsi/3WiPJSUeY7fFsRfeeX4zQi4O9
vW2NfPGzf/n7HoNxyVKEVJof1kcK3TyJrfgSH04F7mUIiustAroaSGY7EwPjl7y8
whXsDDUmyDlrBMob1X8jIaC1WGaJLVIh9xj+4ubdI77KjZmGEsqkShpeLbufHYVL
nCbsynEDQvzgLexuiQxnaD6QQNmTopUsF+j3LR34P/iJPpDpdjSsrSUqNyYlgJ10
rqT7yP0EgrRgzTgts8k0hT9Zvj8OM192qM8gcIxLpUWjSY8Of6t3Zi4FN614ireY
5CnREaDKjjHnpbaXloVcczV+0+hMNBKFGkiMjG9ufvkZhncLPBJTzL5JBFzrWM7h
3N6YT/7rVavp5+v+k0fXbpLl8tlqO07nn1r2l0Dx+Dw7VMMogKs0jIff49gdcrE4
oQzxuqotwYt7hEmLb6VjcTXt/+J00gjDQg2DpFolvornItqjw1h127ed8v1cZt78
NumrmHo9ntm2GEAp8NQAiSpIA4JGM2Z9uUuPdY3X8Aa4fwsCW3Nn/KgUusKKdq64
06LISJ9N/0obUfjkvmgSrXklLR2VbwFqM8CI/lhAEb9bmcKGWwDVJQ3uqBripT6r
uz/Hz1YUg0u8AH0vk8yRJGwqvgAKEKeasK0NFgkwS8wjd9RnzDY5Q5/aHTx60VMT
aURfbeKjCN0kTJc8Siswr56JRWFawVJ7yi+GNP6rPRkWBeWEsiYnr1982fMnttfj
8XXgB0N/LsEBJ6nDfBaF4MSNGJX6Y+OPGwT+mummOnoYvlBKwfiXM6a8gZMgEjot
kqv88SRu5eh4thQpmpFLkrNLaML321sT+hc/FyosP9BzZcyIA4HBB+oqh1VV3bfM
5YnJFSY3K0Mw+1MHqk7b9t+xwsfabe7GOEgAciCB/ZJ4FIZuysVyEyhZWjXwjT5s
R8IK7+wMv/OQYmTNknSR+ExEwq8UawhKBooMzCVkYCQSVfeUdetvOD0J7GojDPhv
l73xYIbeK/MeJavBmrSOpF8+kSY6q/6lPT1lBCkJu/Hr8h1MeR3HgE3rBvVIH1+V
xbPXY5abG2AVnPb4iUJC3BbkQvU+YvhO8XC2PgmfF5wUQG9AN6Vc65vWKEZcLA1j
n7yDo46VWvdIo74hK7DdLoXXIobC4vOzHovwb8+YnN4Ed7HHGJNdSqBz+9c8zWDO
yUKdE0ZMlYgUxfujyLXeSXh8iiNIYNCXYk+EavmO/Gl9oIZIOJdazPwWHwLisy0t
/0j7h29H7GQI2upi30oc5Y5aWbNzj5RcLQGKpk6hnDPt2JEg5IrvtpzF84rA8o3z
BfN3dSszt0nO8eUnp5Jif3LzLCTVbDk0iwRIxJeN/egaefASNybh9NYsziK4ySDq
UUTy4MGYMWFKx1Ckrn6GVffVSwfgypaGYTXWdyF2rYIZ0B35rJuDKueFEun9FzeV
YnTelKko3mO1CeS3AATQ2DBGB1Regm5WAZ1b7o2nRpUmVUA27NFb0ZFY4h+LcbI/
tsX+ZtGHzNZDMFEGereTMpLkNjfuYlyHEvvxEXVLi6FFnP2JFRmMXz/Oyuay7RZ+
inx6R4Pa1cNOFlJsvbxLcId8jqb0bp2pNhGjM7KWdbLqiIC8mrtvOnhZwrStkcb9
jd7DFtbGOzvgMUzI7zjagBrikh1JTw520hWu5yrNFarbfHEeMsr+bOR5AR1UML4x
mupUj+ffnH3+ig4Ysof4G0P6i2WoIx4v0OrciYX6g/EWiScgLIHW9Jqj+oZJWJi+
8M9CyvEWg9iylEXgKM8uIXgU74pchs1T+IEwNQxJCBaqTLfRLx6PgcwsAKvMFI5o
NBDA3RIzLkCAIjmAp5g5/FB0fy7PhqKyy1f4yxYxcwb82R2OfaAL7Q4217h6ZfIL
ezokEi6Cy1vKjnEkzv0eVLv6+33X+W6DwOPXPF6rcdYXSNjEu0+zCDe86JFygFLZ
4LUrLa6Bu8wOymgj+qsHkBhi75ZOvehPc6VoXB/1oB4B8vn0snxFtJps1qWp5c/i
jljPjulBc1YF+Jnb0Sivr2ZnP0GzslR9CRQPMh0MhurI4ChhgMIxs8jOMJ4YTh4y
E6+JgCdKyUxU0Gqh8N+xX0ng7i169ByM2BFmYVWeGqrU8LPgxyi2FKyjdnJBbFKA
cL/D/TdOseSF552TsotZVf0nAyYq6VSsDXVm2X8ATMMgEa88bHI+dY/UPREa4gkE
blsVC+oVPxewKpQJXFISXZwvcW+KLl4sm+0/QNr/Q46MfvFdx8bBBkPU1FyruEec
gQXg93Su4NO7/RPvmHCLHmcS1tDcqYFUn8xYL6AHlnLmzKsz/N+QiYYOSukSNt68
HtlfdVqvyOxX1w/JWiGSI4U9gnmtr17aPCwL7NJ05yXOPpOr1P/5BmCkOqRdfCty
8ucEhDGlP0NjolUd0QAFfob4p/EfFX1iyio8Xwck3LxMu1gdwA/c8wpLnSGfQWU7
fBACB4T/0Hzq8IJy+zDEHOErqIaYxzxdTPM9BJQygPQfaRRLbvltJQn121A3tPgV
WgyC8vgDiNsOu7zyXKvcqqF2sa7r9CGaYQrYXD65hTeBcfjdJlk3TIocyKJbA7tB
C/35SWNb5EU3uCKtaIfuMXtaAIUg5V3d3xK/tax8LSBsiVAzFuOsCGlPavQOsmaT
jybs8/MDiKRqjCKk7Upp91dIPkVRwPt6Y97lzDIO8+O/ivxS+TOq8P0HvL9qLy4m
ofePK/iIzSkyLaKlgL6G5Uv2yc7zBM2A7wg6vIEg7utZuHYB0nSz5TNdFHo2zWPK
GuyoKQu+i31zNUIF4aj2p5JhBTlf1Krmcw4D/WC7vDQQTYxbFjxnoC5VP8URigd7
FxFhkOsEsjYMtQXxLzr917+hVUNgLbPFrFs1EzOM0N219JxUbcX+Pp4JDDojB3Sk
br65L3hN62WVt6Hs/qklJ6GfTPZkJGBIKq57WudJ9J8Ho9jR87ZFa0hXq7SoCTD4
Y809dIrU1cQJ94WzXHMUJ3UGMzG2qPzK92VdrF3nTjqM3ve2TDOOz/8yTExxnChR
nlfv/gESSBt9dA96uPJl7AAGWUqjI/jeuOgicnfJJxHK/Z/EWdqMz2UNlHynTrR5
BqikP+Wvn1UpbKtIJvjMsqXJSVwZxpXAneMtEWO39/U2V6DJXvgTfLL2yz+TYs9Z
gObGSfRXT8w4uKMmA7Q0hWpMp+HuUzJj4nRGCclpq8udWML9t6l6irvj4pHoiBHz
js9u8iFcQzqwPCq6jSi65ocRsfhRoJKMScL9PRjEdu+NIdfQ6rpSgtEQonpI39lw
uveUfRqZOV4nzbuZWZSyYFNV38IcZpdJBTSDhznvTZMFOzLZK6huq0+UWD7sGyCU
HuQvlxP4f8NLhV9fcQRya/fQOTx/M9PIejtQ8CVTgU904NrFuk064tIWWYK74TEy
io1vyh3GifEU8IE8N5jjleyp7DAjwYysKvb5ohz9CzEHCE851pjIZAFGhI1jMLZs
Z7uqrSlTwy/t/O3Mfa6fA2c+bfFo4M6cQMDCGZ8OQNo4FlePnbG4SroOdL+sVYRB
tfzRJfG7fUZlvrHSNolE4l4AEwDb74TnbfAc4RHM+M9hKM4+cnO7z/cnrFm29YeZ
KPXZeiFs400nbPSTt1R0a/zGbqtnQPbBw7Maoha/ybprqrw8UdgXF2d3hsU9tRMy
WN6WABefTcoiK/uv06ZfmitMEt5tJCejEGZnD5DAzgARWLQefagf510yJaG4wbjM
ZPWuJaf9sMqx5yc6mS353Rzjy2cyeqvLieNlbjX9U6lzmMB08NEoV5oc5zKiZCAM
MxBBAzwkjn6+5txRPJcQmaV5HHIlxaKFaxq2O9an0kLDtR+RwqMd/oNlRNX6MBm1
B2R2fkz+Q+og69vSfPxGRykJvi/PhaCdWF36sStfHJaP7Fh2CNm25dnOWb7Q7Zq5
N8IEtRnDoTy3QySnrUrolXCmLKTcGizAUUt+oPCG1+VlNRqoA9O2Gm9+FLBu3DQo
3RUWqi1aYYjW6hre1uWi+ZXVnm5VX5XVodXiLm1/B81Jdn39rWoPp931n/1OBYWz
FKM77sASkVM0JJt4EVA3qdrQg+NFwZoy9/j1YL6lucIlvOdH0yN3tXJwyvjMKAPI
8rYX9FDQ/mWwwS9NKKAWFFXnP5YoiLwQTEslePwZMEVREtfyNeEOFD315UWkFnLQ
cuXGoNgMPX7jRsG5l4KZ+jGBNud11gQRwMmc7nTLS5RksXynieXwQ0Xh0EdASlHp
VgTSi0TewORMArbuyr/MsmxNno2wpfqyDxuFsPIcZvVF0cZMORKeFZog+2ZHHzth
EOOCRVOKkzNtGnUFur4+PK3o2LgD0yzJSILbkxBjMoz75PUpwYL2YmRkMch9pZfI
lXmUHNWIYo2pbui8tKWn6sKbVAaP/DDXPCMyKZLdIfc12RhUMAQ/q5x+YeJ69wj2
rec9rl4qXswnzcrrsLr9EMkVCQwRXmZOreGXTkyTf7n3g5mOJKzs1XwttCxlzANd
S3FOIngha2Mkga7kKKDoFjNAvlha6sF+1f8ZHR1pZf6llTn/tIwNj9fNjkJNzi9I
0hMSGNS7TVgSIw7//um/A+rhpZx3AVbuisWuA8MwUSbrW6FbOXQjL0Nqb4mW6UMz
wQ0NzBOxAFriDE/Flz5kbwNwhwl4HPzOlVwSVKjreooQevmyEKd+pUhZDAboJD/g
5re/97FivdQHJbvBr0OG4JmOChft4dunQOdzcq29rHNAqezrnet2zzcEQ9NS1D+s
/PBTZ4tdC86n9g6v19Sc7ZSwJ9QbjCTpjaA7EBs/uTODLmm8zkQSPM879fj6GGfk
9+nHo8jzQLMPUvj0yY7O9soyovnAWmquTBpAkJ+b6p7FN23RlCePisNisJD3iplH
/EH+okToPVzvtPdbPbT2zedEskd9atzNMyFdAoD3HKbK88JbFTynT3Lp1b0ckQMZ
fK2enw+7VxbZIlkyt4RsHpQe0Td4zcwo0ZWV2DhSybSlzPhhr10LVtm83yqrOUnK
LlY64F0vxltvk8nR+uDWCIsLTnJG28utHLud+SNZqIOmw3wCmylI/ROzD5+L4DI+
jkUxDHIjJAVTTjHiFlPlCki4srUJQ8ffNXkKDcchaOqJFi6H/elEk3jpj65Rv3Ol
PvgthdMp0y0cSMvayPzKNbINMEuv7b7EAZL8yLgKc6nJeTPVOC7HxKKzKK8eocEm
bHKKH4z1EobENsfMuPxcRkya7VFJmRyrkEstMTCdPBGeL9prGSMqTfau0I6Xp5+l
IA3LqEz8/T0nytx0n+oTn4Rgp8yT/mkE3TqoQy4Qozdw2S1qQCG59n/p1RKKvs5H
U04KqVNPTXTQ0FGA5PAs/t/M2/bEy17lLZ5AKZUxLYOOVgVSc3L5q/OC+yuC6PJI
DKJTKXIqDaUgoqVVY5zKw89Gc1Y3cn7b4JUWPBu2m+fk0TL3VeoDc+539eR/zBwz
PDGRfkHZWnimbEk4gdCCNyQIYFujl5KRTYawqrU3fS7rvF/9F0g81l0UB8GKHTGc
lE07zxkIRNnce2JBfzOadUij3mJktYfShJ/0qH6iTFmOW86fh4sBKXuzJhFbcZBQ
vd5D5tbiOUaY7IojBnf1+OUVClbbOsDFCH2VwrTT4XEhCnArxqorkfNj7+NhPvf2
wpUprj6uY+/zDIu/MG5J4dp1/md8fP5j/zXLHeCV47cDQQt4xo5o2bFJI2gTgnv7
yJJnH+6KxzlVyezNoF7gRAT46D7p9XdTPlK+vHE2uJzYgPqqGS9ixR/HNjxfL34j
hzCWSONxAqFU4zq2ITWOQqTS/gMWliG9i2wuBKO3VcSCUblX8QQ0VnmsG7MvOvCT
ZfhFtD3xUU2qmql9yRCYXTnvu/vWmSH5wWOkp7UC9v7avl56evgnI9dc0lZKIppe
bmGVBkMBjZAPetecZ5n4FyijU6bjRm6e6oKwvamHQrpGAzbmMsk5UMK+y4BB1URA
31YiAetPZ6MpLf3KjJiv2Pyv3mMmw89fSezBzQtbmlNW7bsec/u94StLuiwkgn7h
yelWRERq9J4pidBo+9AACX0XyETtj1ZnMmpfZbEGbWaEZkq+S4A87m9GkluzNZK7
aUnCbCM+Vp+0FIYKm3SeY7NQUKnzQAbLiRXQLFlQ7h2+voNC7pO/MtjeewYAn0RG
EdUYAhUh9icqGBGTic4/dl7/hdEBMRPi/zNtylj6P/kRl+6ny0H6U3aebkpUlmqu
WkrG43B8d6safjoX7LyMGOUU0BLztnCACYhiLLcWLppf9C6GVmB+iYp/QTJCqDze
+YMhllCgZl3UUNf0k/syJxvIP43L4Mn4FjjhbO1ajUDouRvSzYmo9c2wnb20/26T
AzxoQDnbfhb/2kNy8Fiv13bnH04/Xma4SVgsywNRD68yDGolzTtm32S+bEybk7jn
S+nzwkNc5iJBDiq9g5XsGCIQoO1UF1WY0zc/0hN7YmVz3uKjJ4+VAZIKA3A2iiFk
n2RrI6P1HaOcCZXXv+VjOmKosM4U6VrqyVdWf+oK5yU5E6qzFgmoDTCktqXDbRV/
83voW/90a/uuRJS5CPkof0IPSCrgOCUSBZdVku0UOByOs7X8t83RQ2hIt2qrGqV9
c5QxMkSItpKFgl4FNAtBXjnBuT4u3z51W3NbIHIrKaZBolB21aqe8TbNEx6J8YJg
GK0iygRNiHyKLox3SiC1FjfxzdtGs5RV9RmqdBs9Xt589zR8ZyoZexWuol8UV/B/
2u5E7+smsMT7N6iVC+2eElSdBXpxa7d56DXKgWQR/TewF/DExeUt4GiN0TWXNoq7
AP9iBDP7IvpwSrLTI4ImPuwSJpClkNjSNd5iukPXEYZtwR/0m2Sy50V6IRuNugJN
E+XZ0tT4ldcDEeFeqtNK0RlpDkDG8C1vPK4nHCCEzW1v4IW2MhhxHK2zO9SQBMcP
uJA0E/r91ctAnaBMtoWAwUj1UII6wZ3wfI+cPFTwzk/Bu341TKy9wUmNoq4Qfpui
3TCGq19k9QmaYz41P08Tf1UKjfln+f0xJDjRdHUtz881ZiuNKr2Z/YX7iN7EIHe6
+0FRUULh5xnHZro7kyXjHKyU0JB4k2Q09QpTkEFVU+jzSxbvz3uKZMIXFNSAeJTf
GMsLlaI0GFXP+8LKmibRS6Rzt6qzd+Tcau5y2EqQ8vVJkDkm6SojiMoaEChprJF9
CpHlevlZyfWeRG6MGyJrfvVWPcczt4DoIHg7QLT2EL+YhESUnnI8+cJ95g51iLc5
/b4snH5/+T3ENq4G4cjqwchuo15PWXzcx91G0bbpI4HpHigekQ31M4Yhyq0rn4rD
z3JbrNShM/Jed1j2K7PhfyFW2BRwQ1sSKFrM75qgxuF2UYIm25bSiFIfgj+pLBsb
WNy/YV1fVeUBFAOzfcxCwNifrEz9ze3S50e2Pq1Q6FVg3mWdZO+rxsTdbWTvPqCl
50+4+S/sfwbcd44/RCNK0mbG9cJ/+sgE2rRnGPn0fc834YRGlnG3ettjKMpXijdW
3znsUXueSIVBJM61sAeBV6kTk2nw+P/14/ERJAqKaHZnXUWJ7cHNw3dnBmdDI8qe
CQT4Gd/o3WaiGRSr/G0VcmtHNZzqtge4zGY7UFkiAkbMGQzr7BX7vSdvhhV3ZXWE
fEAYkuja1+nTlFCA3OmowscW6tSlWELMRjFOGBiEpWCoGECiJu2Twk94Y9FymDKv
lTrMSNs4umMse5IgLlsWpzw1Je38wzFdGFF04hB8pd5fPPp+M+jpNQ5fTXLkUZNF
YzT2qOyRQlL3fiv9z4SZQE+ST5Qxg373y4tPM5Xlds4ZPEBDu0BtTikk/2ipTPmq
cQgfYyMc3eyclG16exRZvDow6thBjL3hkjkFHx86Q2PghJLgstWmoOD1lFR5zib7
DlnGfDFKksKP0Dr5CRmJLZjaLyEe0eWw8H4LB8Q1aTgo+rzyz78jmnOZFAEygZHv
iRIV0IPOtfCNomdRSqL8MBHgXDu7P8NODoSGXOffrzQyjm29KdaSlgUm5hZji1iS
ZTe2WNaV1zZqCgfAmkmEYR8QeL/0NfMbhLIMOhWvYPJN4S4u3Ru1FplIT1dfu+d6
ZJ/NeUibfNbJoAga94rtwIlZPQXI6etJ9CMiLkrxfHrgNCPsG3tGLZZQ1rMi+usH
9lH0bfDeoUSWjmwDtZTTST6BTb6fbS5ujkeBhi46xa5JyUB21zxSQGLcFFdGSzCM
9Rvf4wUV2lVJpuJ8m2ZV3VB3OOC4NJ8EbYNdYL4qbF3q9FfOKoUHMLeq/16UpAZ9
exscyGo+VcNmNbx7mjEi5Tn5/rJS/XbHdYkx7tGEIZbmf2q55/vxOiOaJ9RgdUUO
f3s3hw7tW7y2vvyh44irH3QXKPEZIp/xaKIIp/hzxtksmfHpSM3UBUhdZ8zHZqn+
7fLz3uMD01YB3YYA0FO1/e9fPaMXKODHNj6ddN2QPL+6ETLQLUpy9HinIpSoxQ6e
NocLz3hTSGy1e12sklL2Pkr8P3P2TXU3aL9WjItFr8kdGtl0QKfvwl4kQonevnFq
0r+nVPrr5yURRucIodpjbHiptcGPBVsrymHK0oAwI8923g7cK9OkYSc8CMt9Sex5
U6R0IX+W0h3PoBTLajOK6Uy/SEZhfTZzWtmXy67RhURrUzM+OPWt0zIMJyBJQNOU
hAUkr9m5nKkZiMFjrxPCniM5h4ka2qWKjEVM36FHW/cEvAuwEiASt6wQ93o1K10J
1u8ktsnfS1uN0aGaDDZbU7XMBYIFzgkFQnXLMH45oFLGgDlRa0dXEv5QyvVKW1Yg
aFzn3Z7TlCEApoq1lu9P9R4VURt4HwisANLVXAsoWYyIr1XDfV7HtN+aFz0VPmq/
VY8mxfLYt+EZrh2k/KAcgK5v6ujq5fiI/WMjLr5+VYTjl4e7RYZWiUeFf6pcvJ0P
mwUePXKnzrNBnqZRiN/HMFLhLIpR0YLqdZmrCjj6dmmZM597/gSJQiYWC8Kgft/g
M6s5RiNKo4rghwXBcszL92tygL75DfWaUlWSGGBHw5P923OrLsdp/R4G85CTxHnl
mrM0z1L3gVP0QVmvUqyJwb6GK6Y0ewNkch8cTtIG/t3O/+0HOLKqukvmWKuQAdfo
MDhYIkrd7C1NZ0g0AovPo75HVy5MR0oAbzxINVqzqXYcItq9oX14kXBHiZHaS4eg
j+39rwAXtLmMnvUgFDGHyiNDI2Xi+tLGoG8XpWo77cxb8q9Jho/JQgGcw11l2Mk8
BJRkeTspQwTfchHhXpnQqkczq3Ut1bMBrgXXCufcALpoSFo9kL+NhbbAru3pYJE3
zB68i58VwXIz8K15OyF0zMwUzmAQEwtE3QSoB0qE5NGYDqhnQFtnUykd7Dbv5E1S
VtYtPA5XDSlSE+VpVlCXmQM5Zv+NHHI/sqY2nTtx1Oo34WATEEOPR8wen/i9R1XF
382nEFRTmr97M5uvSDlVvnDbyYYsrkk3td2jqBRE4/tlhZAqiNSzZ8kQgIzEIxif
VgWSKe65mCSNm33Zuuq1ubDLPQxAWvnGmZK/ASb5Dq9wB0zYzQ/5TBKvchV7DYZA
N+4AM9RbfWy9WpQzakg4qIqR9fsv974puUX5n5mtYP2viFM/Vvcv+vTHtHNCWKOy
sUMRvxiMHxy7uhMzuBhowcJnb33f6GO9EDKSKI9ZV4f8ftIBhKJSga1ND7VSKkVX
uOhG+6wFWSRdedudQOpR4BllR83+0Ony3RJVOgRymsZWU9JJcZb1nURTNhEWhROf
gCWSjfUNxL5JUiDiuj3d0cZTCHKaxzRU1hsoZINArFzrjY4XVBhLhMaBAkwEyK4P
J5eaGkl7I96eXJEEeN5YrnYHBPG1x7EDSY7NjEUnSOl8EaaU/LESI0c03SZeGBXS
PWyBvNISY97Fpg/5Q78ZF1jd3mY1lDPRRVeFFG5bv6Wkd5SWuk81YkkKB4jgziBk
WU3mYTGGJcfD+iehCZeaZ3Zo3PR0d8hI0QyNua/KpaPORsBc1mkM4tO+Itx8m0SQ
xzl1xEKavwVN2KaqvJ8XEalKvucfLgLYfuGYvQEZcfo/RPWrnUhTCKs0FCbD8per
/kTSNdGnP/bOvcaiAKu2jPql7xysembmzLtPdxNYnd4Np4POzGDS1PnGRFDgFfCq
b5yV4/8NuAX6qpF2pXRPh/uuwJoLVThNGarGDsd9RQlDhRUo5fQPCyxOOgBBOqML
PvizQMSg9S/+oLJUk5yB58NG/LGJZnLzahsfChKqgcmsTHiCpsBklUcsHsZ8fDNI
WplQFaMs9SigXll/jBycpGWTfTQdh3367uJKyCA8XG0o3rOcA5g3V8DF0myJ7VT2
HWhHbw1R4Ek4pwAQIu0JqkWTVgPripNs0GRFv70mF+PKItzu5rUgqyUC8swJStdG
OwVGt5pbKnYIMF+OpecSufmnWhT3nde6Jp8n/rt8COela1Rd53Goohc44KynD8IA
bV0Xz/K1rvcH7inbOWqTf2/fz1V6mBtucnFIuebtH1/OZ7g8ztVQEgLLnmO1rJHl
9rwBuQP68z3EZ2UxERQ+Z1HIIWoGPHnpAUVR0l8qrzMaWGjAzwArb4bQnK4/vv5g
iWIVXvmytUym04pTVvuYduRlbRLeynglSoHViVWn0UavSI1Qf1SRrQr2k3aISxCc
uucCkL/esnqxbAJ/fPMcJ/K1m2hNF3c0i02jlfuh1d93o7iK4RUyD/jv2Xp5UDHd
B/WcFTFXGHSPrC6d9H5G5lYcYLT6FJot6gmgBat883AKsBIzf1DzK96ThD1MvcgR
7OQsQ+ferHbNE9JYTq+40ba6NFD+CATXDKDxhcFhPwBRVZ8OxaZxHmJjAK/gEn4m
8S/isBSVMnwrmFd+Daih0N3x5DNTHTGpT61xh167SbYNRahBRURS+scqbQUCtsZG
x9ikTPbo6axODr3LlPtaV5giAENkUBgFFn/AgV4mSDVl6e81yfUJZ5B4awatQACm
NZztUvQWQY+iZYZe1r5lK76FflzsEQBSsfqVKgJKWSIQeqeL+pBd00YrwDEwO1GV
nh5ElIQOrMDXjnAUs1Z8CJ4bwWrM3/0GMBrkKjROrHDe6I/fpo5io51JFAF+LLMU
1QkkVD3slxdU4TjOB8p51cA0d8mFzl9GWgwINm5BZYoxNGFL+q283n+mXvwwjeQj
lF9/dMv3ZB0pYdn4/HuO5TG66D8/8rtG3nZ/FhtL1uUhPpuSU2CGSnLDTH7W417c
Muaba/HZvEcimgOr/ygUE3hueRnEwGU620K7DMrvKt+nMxFdma9r/o23ufCDzGxr
2hUQV/ClyCiOBNKMapYJQx3EAnFyYfnED2ME3uK2PRzcejt7a24V4hYdqkv0GSGo
6HbER8w1sfESBmboEh1DcZQtlOiXdP8XFb/5uRYzU5cs/UKbEw9Z78ctJ8/bmhi9
dt5Z2LW4l3urIlcqRcMCA7JPMu5sIjk/4VdkopsJqmzGGWut8Yn6phrPOEkl+wtT
v8vf5eqvmKggAtRU3zXFhEDdDXlc2iUvcuN7r8QywCmRUC/JVGSTUdY9SM/guAQ8
qMRPlAtUPAxjzLzUy7mPqAzajll0aLSE74K7GWRQUIIqHiiuLkj7/elFzX+FsTtW
xc9cA0y/Dsk1jTtx7US0bwvMDTvkJavj3jFD+gVkLfBgIrW+t0sfzelc6FRg/NAP
2+tdd8vxUM9rA7OTLndsu8uTDRYy8HDhM/Y/Aj65jB6+D52amVsEi1DIdTwqEzlw
zB9A2rp0Wzpwhv+MIDSQrnFnBS2f7EFyRto/4nrOqxmj4/IyYbuczdDIMOpnZ8mi
Jwwbvh6k3CSXtU5mZerJKGQGO+C28fakq4dFitIjxme+9LD+rr7834kL7x0uNTWM
q79omCDcuiYK5OjfC1XwHidzK9eDzb3IfpQqk5Qt/dSw/UeNaKDtuvNYRCiAs/qI
GNXjspGp9WkdwIt1pwz76/dGTpNyOSgYHNboju3MOqHxKxBQJB68W/vKN+k0LH/8
uvEHa6HHIvWlj2kAonfQal+Rd09DcaNj+X/o5R7z92RU2jEZl2uA2oumNu3vf9m+
e4z07NHuuRxVOztVjMbT64cRmzl6Y6+BclPOYudZkOdSUzBwg/8H+mT5bSukDTS8
yWkjIEDlQajiW+5M5vqKh2Z3kc0ExsL9MP3bPs7ibNLA7ePxKIBXfMKjJEFC2bDP
CBvKX+y6GZPJIRVOof2FRQbUMFFbjlIGHfuCbfdXeg7P8HYaKp26qlrLmdypch9X
7Py/B3W86Zx+ATcTCFjg9PlbBMNi6nAyml5wseqe7QG0wF8EJBeiK25kvj8+M65E
KV1SLdi0DmWRHu20C+wFDEa1pKY5ITxLG/VgHaEO+DWABfh67bL9d13Y30CCMC92
l/H40S5MjNwvlDBHyxSsOScFeJc8T2kZ4MoCPXKX31DTfmNGLAjAtSCSojLaoYtm
oBWNnrNvgpMqGk+DERxhEFerLwVyy0VG36rISFHX7xiirrjkUTBXyVy6BuLg7qwT
+tmlgtqetWwGRaAC/KbZTWBuM6JVnp2FvGFOQWNDPg2eTOKWx8xM76BDJ+SnPCy8
cTqAf3mumHThgcBnM9dkbiZy2Ey/RdzQycO+CRKXvAiH11+NHWbKxF2qOniLFy4p
UwYFdG2NmR/2vGHnXRBt1CQVVx1NRh9f/srj1K/yIinJ4GE3RrOcbWkSRyeR/ESe
CZF69dZqoJzvYTwwhjgcD4okxD+lJAtnCofvDkipyOgZOQz5bRVCowLS+4xJjhAN
i++XWQstnaqhFI3wBTs80PvfPUeDEULk0y84U/E4R/JcCYSspXmzmylsmD1IaKoe
kQMmHXmjCq99NmAqZ3QBlzv/sUu6PW31me0LZX0xCke48rQX9VsPU9zIVSONi/kE
z3S8imKqPioExtcFJz641NOAT4XxNTDS7YLlS2IUasJ+k0ysyrZdftv1B9NGkreP
+QXxefSYULQClOqubj3PlY5lrm/CUd5rADUf1vGyu0jdkuWrpg4K0fDKB8DzglES
1EGzVgYNd9D1wWTRDs39QoX8PGTvZhudbFD7dbCxnoD476dvS4z9XJqBxR5LY3xe
3ykv5q8X0yFZDwm1pQh+RcV2mgDfCwb2lwcFF6Bp268Pzg7KYCgakYQMKRVmKsAR
7AzdZylvuB/s7r6HTT+hPICG6eNh3kW1iCgZS346BXJGFq03Ugmvn4Q9dc2oAQfK
gim/yhBOBu3X4rhTcwSJf5vdTmnjxlP4kDugAwglnd9Nl7z1pcZ6Bot5smXAByam
tO3VNEqcoTIn493wFTXK8LOSvfo8HOdXDdQP6On/opQ+HMZnv9cxe8XTu0KTcrFL
DVlXaFH6nVp3tT3ZwURnJc4cOgNkgnejzy4MX5cyuYdI6blqcNoAA5bwnbxSKNja
Hj5D2f7Dsg8orRkJlX1IOb738garctva8GkfmkgErKfXZZD4VqlfBrSlmM8U5CcX
BNNkBbH8z7TCpGyHTuQQm0HF9EGfDLgbm5Zp5keOuzRewf0C36VZ/mnmpuZoRzYu
wgXe8nFwGC167EdeZ2hI8Bv6af9IvPj2f2Ywj3n3jJQNdfACekFH61h6WBSqXHK0
kGkLf7/wv7bFtzNQUIdSwqpb3pFg9ybijDf6kN8P76u6JjhhtDwhdl0ckcS77P4X
dWBMNRfBo0KZPlsrrgIPc0z3fcaMC+4DuJQbWgQQXte1+suy8HmiNDrEx+QYZTug
3vdVG0bVxf93VYKDHvcr4zCnVSeJRqoyAbJSB8WpKh5SgPEB9U3ePdLAsT7M7iph
rdqIh8AcJ/SKODJwWk8e+F/3B5AlYaydiBxNO9b2UW64z/mU2xGkIxPV2icF+rMr
sjRYL5a/fpbLD4CxrJv6wgPW3260rckXMcp8YNJmKrC1hB2Qu9D2AHbMjrTSH9bi
oUo1svxi+CxSuX2eqgVdVpAgDjZW2/1UuSVT0GjdHr0nXx7chux+iytHafa8iXq6
DOJwNM/J1SkBPG+UuLKjN/LUQFtz3qyGr1zhM8UvSdEPnVZL0fn+DpWaGxlwauzA
T8VjKW8JRoaN6XReHgvALHOe6JOZDIbeEtZMHxWGuFfOn2Y4VuXqRQslYfujq5TY
ja/w52+tpw0vmCbXBCK0dwTQfOz1U0UdcH8oPPpaFyih/AP7KQeNzRONM3T8gHYS
/UMtU0lnJGMMtgLFBcTCo2OakAl90UApr76kUS2udck+pOdMXz/Ks7dJ/8a/bqLv
N6dnyMzSLDuCPGUAAsquZwQh/jDZeKuMGSI3wbVN+xUoUkDLz4WdmZeLRw3kzNAP
bKWay+4ZPRYpYml30j1aEmpKAe50PVWer6bLTBx8hPqkbhyy6aIvQ4y4BfY/hQBW
YxJs7zSLX6zHAmeuqNTAhzCtHTjRrppSVHmG6YM/uryPQpFFahxBpinmn+pOM+r3
h0n8A8oFnN0yCad4wOdE6c+R9biU30Eqh1uATSB5dKMNRwyDn4ewmwDkXdoxOPdr
3HJIwJVOQkXgjZrIU3aSB4Evq+Ufp8B9ZxaixMLGlwEkbB9lWAqOSg4dEGCycfTr
3zEnweQq6R6ol3y+8tdwnJn9QQu/cr7U5T1ctJdWvQEa7yf9s6Jy1NPXrk9LlEYK
wuzYDCTJ7A/vh6HstME0e9OJBXa88GjInktbSCxArkK2S6y0CKHPuYGaIYjKhbTx
f4rXHTHLTMNc6rwBeZu9OgG0F47Nz148K4xt4GOLJEUm3Z31FjUQdnq90oAbzNmt
qWTPWeBzCsMuSrqXln6GFE8MkivOVhRMveAZ4wPQid9sjwk11eORebF72q8wHsfO
1lMLdOgC/gUcGOTQ7ePjCxAol/T3kZOT5Lv+7t9L9igMC9debvyGEVJTRDDWM2NT
0qTUKxG//SL8TD0VwRthWqK1rz2maTaZNS66uyfh35PPjO6jauw5hLbv2LCzh4sX
CsG2tqzNhwmGSOBcnfvvv80xj3NmP/oY9h0iahksUyqzLGYjgYauaW605HZ9A8wW
VYtDsoVsckKjJKoZfJ8Muys4RtFsZDrcvpUst5DrCq8Td5jVBjTB3KQQSQPkF52/
imbcgTM4mLXPh8QkUO6NXQ68bUSbxvakwtkVkRySPz9H+Z2hPPWaWC/DsVBjDNBW
mKyubN8nxzbWDCMdaAfpJzLvXgG3IAnwYX2Nu8rInt4C3gZxXLivC9PVznCz3nId
gJTG5h1OHysuGOUFH7V12CS7hxx5iYEuLYyD/428EwxVeARcZC+E3XE4od2aPPtB
eq3mXQ0tz/zsw2OGsW3nL1BR7dlb3qAsiEs56qWGNWxCx/Lxgw2Fn3m8TV9QTjkt
qyGh3wP9I7X9j9pTAjEdVg1AmlkFuyKZwQGh/diLwWOQHfqXA0//uIAqg6hYMJB3
TnO9CV9gdPN+xUGBrOttUQqW2L4OHvdbBv9uih5J6i6AJRLZKzwL/022u0mAX2YH
5asbHR4YRisvFd3t78uVPuv7pubGTln2tGbsaHXE9X/CfgaEKLsWJuasbTVI/SLw
La+Uhj+pFHcP3J20t/j3GKl0iLfrwwUOXec8EZAmt28s8xhqBbIZdXzxaYc4o+U/
Wfhy68+xrGEOkvX+uHxXjwP8K8yiQMCNFD+ijqj1Dgfo57vtsNkr473qRsbhVWvj
HccA3NonJfqe6nYr47YCfe+qu+8SlmeNW1F16rFS1VDOMnpJKbDFM9wRwo1OMuUH
oaQk9MqyUxAVmBRP6HsAF6p2KoIB+rNUtdR0cSuvkwL893xaOHVoERFIOWygRNt/
mmi12d4lTI2qbq6MytukNN2nOfXgnZrlsKZ5Z0AVrT8Brt8f53SKQxfftLoeBHr3
bT83PY6wsL7J0e+9X/FPK+fhTAhHBEzwWT8c18zSd2uBT7rfkLVLjPW1t6d0Sird
G4vBIrw5787NzfbqxeYxJolzba60kC8xKuDddzgMflLDaaHE1BqVvoqxsiD0gzgy
8EtXwgemL/LcbTuF0h0VkDAcATwEEAi4Y3uApqhkCYc2T88RwYCHB7uU1XNIFYa9
81Cc7CYzGEmNmI/G7fWVfuawJkDvk7WhMhDwFjGDUTFa5xxHg4dGj0p8WgfZH6NH
NMNMH9WDTsqg02vmHRZ2bH3v8Pt4YVgufOojV/4c86ixEQ8pkObzYjT3FXRq8Xuj
C1jLyzdo2vhEMKF5aeD+lXiewbXl4FL7YtP0nGzZD2tGJQYk98PlIDfXProE+8tG
YJbdACN0ZdHkKpM9LBlIrwZE1XHjyy5kWQNKkbhThbUXPDrRHxXcfycucOipvdm6
fQrtP8B8wThF1+bx6ArHpK7wp+Edci9IUBDTmIA/aPeDiXEu5d+4J196fEqYd0Hk
ypaLpc42HcfHH/mx9kxZLEA5nUvmPwfHH4NkJlJ2mCvkKdUY9GVPUbI/dMYU5MuY
I0yZMF4PgYO8TK6LF7SRSwbGPaELGKsJZ7mzJ3x8naH7Iox8U658XvTAWEpmP8RN
neLZE3s7HW3UUOdX1rnejYkTDZ9/BxLQS0BXgJoHB9hkKAtrtfaLRJoCYdHwfc0+
IYFJPwDKK+qmsyAk4nFXoVW2qufSUF/uSwhQkOoC5O/nFR9cFSm/5+Om3C52aDzM
LbN3aMb1vaNc0J9chVEAlF+SpLje8zhfYZlDXdi5XKqoboz0utTm3Hyq4qO2F1tA
RBlWv4XNqkxwPdH5HxIZDBMlGXruLJ8p6oHfvPFBgPrxSSxFLvMFAQBJEF184PaV
iNx0TCkxMsg7K+nou8doFbK7SuqLf/zReKr6wnGIGb7YfNs+cOd5wZ5/ckNxzVNT
XZznD+GSzgZhiyY5mZRfkemPXFGmMKtIYaC+wKNUhHx3QR2jD1HxJI/df0VUoTZx
C60blTeLDFpiyOg+SWlcn49CE6KiMZ8hwrls4TLPMMuGIL/PF6IqwaK/DmX5Hivl
8eKaqbClCBEC7cQKeSOzFyGhTaiyeANiXJwncTBNj9SSXD9LicRGUcICGRseUjzY
xLt+OzOlio7e9rNZ2vMRAoxmGiNARsN4rvpE2+zP8ZJnGC7VPkUAE7GmuUz/KbCC
mC1Jc9aL1xyiCi/p/kawNrmPtjbN3v8T2CWgOOKSA8KvznO/+k9AeNydd5ZPSCRW
uRD2oo+GnzITZQYFnfDXvsXFWS3pUydphF6zUQGBCb4CoGhXdIr4F5ByTqyg2/x9
BmdkCUo8JjEQzW9jZddfF6AVUJP8NG1ohR6qi9Zgui6Vqeij3/sKHTLpnzLCXjgB
s12XUlBi8gEfYicGlp1EqK1/JDneWbHphmTDuc4zWuVtwR2seg0GvBph2ruMNv2B
DusiA2KntLtDLTxcJ2Mhf0eRdPBm2elnvnqu9UUoNCQ8uQKPxZtHlUxL2iZqYMaD
M42TKMuWrloGTufvGAeWwRYZK5qeVEZwqsRkol3bVe0Otpl72PcrOq7+4owhukWl
yRg5GcCMb8Hmjqqg19TG7RCcoaL0rm/lgkoQdwVnETd1Nf0qH9YQ5XJqUrdlE1Bc
J5b1DtWrUDvjtHE+Bjo5iD0POD+1w6PlNlUUKqEv8TkE9nEJEdxGZ0G8y9uiYiT6
WLQWXgoiFFyKRYomXo+03ulSBh8Rs8dmshMHHWVjG+XddDPlBUys17NjiN9PQIo4
S4Yo/366WXMOZOtZfJH4KaWoV7bNkNGEIg53QF2lEl4yCoGabpzLKN2XyGDsUieL
zCQ9vkyTLM4nnLoebxMajHT3jZcBRGxA31DBDafYQIcbO4RwUcWV7sf0nT/VnbAs
a8hHYuzButkFRWlG2cpyXblVB68VzxDYD3xx8u3sq9LB1Ny8zPTcBz6snRrEhyaK
mzoTli5G9TSftvQvmYjQ0LlXcGobToNSh9Dlh+jeJTgQUPUmU5FcWAWjwKZ4qeHx
rReV93UI74NbHHv41lAlGY/P1haOdfN9KX/xJje5+M9WzNHPfNtkMbXOKbhcfgp3
qv7exF/bBhLoUEuRkXcAa6bZoynJRBO0y7V7zCEBKrN2s+CFGyAFCG9hUebjin9o
wXrFpZdlSWJcn04VVM2CQ+pyagcZnoiMB6zFDPc/5UawiOAyb7oNQYKbegqgj+s1
ZFxlP1ptAmlmoxHPuEkvq2qYbTyHA7itAA2XC5dHAbwVF34NhwC5hMVu+PO9W9iM
8xK1f+//lIE9BtatF2tqlg9AGfPay9SxlN8Sq4gTHJyqH2exLt8WOMvqkOI+W3Be
cO2Cbfm1QH+c1zkDNofAioYCR3HgDsjxnrIzJ6fREUgbGmgihTCQje2SRUk6/knl
ycSdSFPYaxUWy44KWFKvXH6+1Ntfo9Q3bzrJl3Bfk8dH8jyyl97i1daV8qLEwqmH
WLly8YnOz4eFpnKV39irARCAaH7DT4ohmclERPeGOmvQ+7/ZYFaRyChAmIICaWUh
Bel8ZrUwj3zvOuNBc8ahAY2wzPV3T5ZQTAmmBFto/9Z2TMssG2my1Vjz3x5a2Zyg
1Sz/HBFeocey9XM3tKq0RY0eiF+ixsRY8fIPXD/SbbZN/YQzANXZWDf99y/zoww0
TVvm77xFEgAuOJEnA//tYuDLG/643Ix6Xl9Yp79nnviQ0E3p122MHRsFNZw/dV+D
P0goQ9sKuTIxAkeXFc8UBN6gR65BMAZZOAw/abmHOFnL+sujEuDLMyiPr551qVrN
JW7EP/jM1H5TnVp4rVsbDWWSvbJws0AHcJNvRcIXHelN3euOr9ULAXcsB0JDrP6Z
Me25MrYM4z+SVZ4Z/kP3sgTqDUusUStjxFlnhfh8qqd9U8hFsA7jsmnnMqcs14Ip
zU27LwZHHn93qA/IYzPkNdOSRJNH+jxUzaFlaNKTIXNywPZcMB7nE6vmekR8bfwZ
iGQTseHH6LmmG2O10bXaZAL0zEmKFz4qdnGfM0B7na/D3Up5dXZ5pE/EsDVfzswS
/j4jZT0hLShk5TtzEReE64Zy9eP8LaeeEEIzcf4H9piwo7FwQjc1ev0sLQMAHXpB
LZ4k7kgTb/Xu2i4UnCxAUaQgEz+rsdqNJol9Lq7VX3WlBO6LP9ICaWASYjdCVivP
ssxdijeE69EBi5OzQokB9Dc7kB3q0OdgyM7XkqivXIaqI/JUtce4feJRBSb8RAGq
jahA9ftCsGee9RiWw2Pljxr8pBfCvbfErHh5uTXrk/Qp9mCrEGkh3R+/FcB9ywAv
3K1QEpFWMtWcBL+8xFS/4kZ5nW46gOh52LmnmnZHJUDHmUM1fxHtkNHUoUmloX/c
/Xh9ETqs0tx9IIjs8QnndJ/qZB2b2inJW2sWnYvNBvbj7u5Dbh5WACmiSzDx/Ba9
TcIB2lmj7hiFpmO3wbT+Y+a+Y5HxdYM3NPuObKpB5j4Qw6poiMxpYnnlI1Z2D/Jy
nvEQj177wWGwrOad8whZKZNncR+uamwKitDnSc5fu6/8iYIVuzUp8SQKyKc5DoIl
Pc+8LaeFfMP2JFNqHJ8pinBfUTXPgcpoBp0iYAI0YrjSxJnz4gtJeNCRdyzQR8ZO
6dGMzxQqIpqudVsuxhLFD+O2MjTXrhM604SRgbCBmqZ1+4uswUijAhpY/q0vq+D/
B+YRIbAe5anzH3Tc4cT2yZy442YVuNAHlIF8lwFdvJ8a7EukB/HY4wKO5hwv5UNF
DKmyozVU2OTOfegF11JSMlLbJr4avknHh5ZQe25sJRnmSO8dZ20xyNWMSg5uLoid
x6vn7V+m+vY3MHnhgTVooKwJOVvi3y3o2H5MPZHJEhqWdFBOsn++7h/A2jCv49wX
LxDHcRfPkjgTHO2fP0yLDtxfbHFL+LVbvUW3s3DhFrGN9I3SDNcgwn/r9pid1jsv
bZ1rtAzWmvv8WeJ0arbuRqMlnoC2rx9B9T+r/L8ofuMQpYynCCNIvegLEh1TZRCd
NQjJSjpSwETwrSw9rGP7rpIxijeYujWtc0cfq599kpT5fm08KEXqBqKsqORD2j4C
Xgu4g6Wc/31RKF3CZyw/FI7FvwJfK2SvhqXReUU+iUQ25/2WAOq8ou6bCYDWJeQs
Em1NtSUyu8JYH/RQTKO2oIbnh2w1ukJUNEsEPlSMCVyq0nwf0MGBz8udTJTZuCqB
YQjdswJYv76b/FrwV3iKXWDbzBAuEZ3cKVa2BnLviQnmmyjWleYT9Ld+P55xotUV
6D3oNVfWMFnDmladiB2vA2fzLT2R8GbaEQKBLGKdnZIHOWrQP/6mByyslsisl55b
Uewf3Ii/VGnwnkenhrKL8e/d0JWnW5XwixwT4W7X6SrTcD3IUII5eUkq3CI0x20s
h1zz7+QAH7Fs9S0SywCddudLz1YzOsiooFIHNytFYZnYDPe9vY8TsKqIOYN+dLDo
2uOHGTvSC2REz4pNcW6l7EVj6XqmbR4wZ59uQK+cJMFiu2URGk300kZD/Ag7Htjo
ScnS9eAI5Qvo1W5O9W1PkvxF4PCA9V4aywW9WV+UKS9t9vKm2QEnUw7fHSbsCgq6
pKCxldOzs1AqsoMgbXmQUubGqarmOEewt07MJu8bW4LcqaAM3naDPuUuMO2A5qlh
RK8Ta10S4SiQpOel34ouZWl9WvyRLgwJreMIrMGOdpAFZwc0GLjEDzkarFYmZ9VQ
RqRnG2xt4o57km/yIDkpLEnmd/HBh5IjYgaYB55xEuL6eYh6lvMh7jrfgC042hZE
V4jCbvlMKP0pDwKZFnydqI+hnbY6e4uNJs9pzvLYxMQfDTxF0cBx+A97qVxC/kew
sCTYln38zF5lUc3v0qrPz6xVcDlpT8ZsTvy+3FdGHeTKttSlJzjoS0XKRItXfBeo
0GaCx87iC7yoVQQBv0IHuVPu2TypWcOmX+I8kPQfRW8OReL5YkEhnb74xqMudERx
4D/ELVGMNunK6bVgXV3RgLflZq1ztfRbvOLh+3QMp0IOlO42W2Wy1vFQCwNjghpt
OKzFu4WA85CvcV2U/qsLkx7JmxiLQbJ266QHCbIgIQ3UojJpZIlhzi5QTKooZiXD
Ec0vGjfc2/WdDIUfMsCaArfkWw8gPJ7Nzg+4n/QNsFgaUbXZ3FOpVUfmE7C6huxC
/MQrNmu+jtv0C+M/huDzXYHtq/LdEEW5+6iPaTTGLxqHdIvKyc+bY9matpKhzOT8
ileXx3VSut1mXhcmL4J0QjZMXhhYOVYvxmJignehVdJLdzyRQNX8p1+apRz38vSY
sEhd511fsiNCwAuERiWe2EcdGcxdq4iGV6Js0jknO4GaxFvws3zW3WbtBv2+Oakc
pm6mWBi9Ts4+ucXrUxRrWKWMsnOzFmA98gSk5duUod759s+945UgblIrjHvk9UXY
Zt3AOv2BjGM7NbxWuJRMALRGdf5mE6u2zkz/xOMPmnCJ6DpI+GgOWj185v3wPrVp
joNeiT5EKQ8G+r+EklXwECzVHC8Pab7OZ7JDKChxbcfOsd1FCvRLaDRQkvSbVTKM
LScDaPO1Qkhvtw6UJNJISYRHqr5T9aMVbfyCIPz7rr61UIIlJfgtt6CcyT55c0Y2
PzRMSoZuqWRjuzv1IhTv98ttBqqdZnH9MBL8Sph5U26ciE6c4RxeDk8wOIVRmN4Y
H4B0FqfOTGNfpq0kNDwsMxrLpTZqjgT3udTFqpN35SX7916t7TB/1C0CEDRFRygM
hTJmOWCdT+xXAX8rBrUrgn+GriOZVf6BL1BjigYREHftToaJ02Rf545eZlLJg5X7
KD6DCUTGhgdPdycfn+b08pcU9awuhntj6qTe33/V8PJX51qW/VN+M9CLky4IlgI2
LLQ4v6z9WkOWkJDsHqORQMqghbxnk46TBBWoNUAaK9wd1rlOcpT1FVTvi/DUtCdK
bkM30cikFPBBomLpUchBvkQpP6kuguhGcGVG+ycBNxkcGaUJpBxcgurRTz2MxewA
uWokGnrHNAhx+B014h/IZpdYnvawIRu0ARgOXl9mt6bqC/0g6vjbPv/Zzqt0jRot
Ga/d15mPKkP2+jRwmsvtBN08LKuwUVneSvxg3lOTjhTkg8MBu9xwCydEPQfl5dpo
+Dr3QeB/4DbO7GHmnupPierE2cXpbpp61+N9dAlUjqBT8Ma4cR8PR4m4jPBQmUHo
7FuU7ftKWPhmYKCNBGmvgjG3NYigXejWQOH/EWqhljRcWAQr+cBMH7l1MAZ4Q5K6
cr6yvbCPHXz+o5vXTFX9EZChCzrXJhZniVM2R9LvHDrLLiyctTYSy0UYGreAp0QH
9QcxJ8pZh2K2iHVOWd4h8e2e38q7zi1UkEYZ9aSjzvaHo4Bb9pu9OVpvKY+JuaQa
bYn5xe8Zt8K882nNHhDfS3JLOHa3dP/JzT592sz6w/YFhgJvi4jLdKQ78fkEZjEp
Peez0FMMBlpzOopHPIDjxGQCRoyJNj+ZsNvhir37ZaBKfG4IAu9G97aXsR626KW7
Za6dVsBBaoJHaf8WG70qKQqdcsQam2bq5FJrZLraARcf6qzdVEF2r3Jk3SH4ZirH
1SS5cFCKZXvLxsRbaxL+eKmCWJUMd4eQPq+3WRIC2L+pSFUg78AMtz1syaOTFil8
30NY7y3jumeSIDeHA4ebvEfi+TReiqUZ4Ybbud2Ml5XfSXLq8AoTdNJC6qMMxgRS
XKYkWuY6m3H7gQTBLWbNFUJ2MLGYNyDcBnfMjp15Tj2lhZ2iPYxzywUCO/w4OdRR
e9VBAKFLgBejbSwzC/rPsdwoz4UotF5LjoWWkjOjhSeQkqNp1j3SECKYz7rjb9x0
7WfVLfToVCKHWY/aIOKd/m+ATIhAvBvsOJnS+f6MSWZLTIbWU52tcWZrJfDd///E
EpALaKC2jd4Xhm3VY2y6uHkYQ0kwq9kTD7DU6y8TcmyP5FNqOgz//MM5aTQwhzEy
ZMQ1CCfJYA51wGi6zymcdejDgu/R8KtKH/lrBv96UYko9y/icNQMjiB+S72aYDWq
uwN2UOAILizWDidi1k3KVmdmhq/6PyIXz5btHXmfUO60ThFuHDLrRsGOC0rirllo
Zl1HDQm5V1IRNeb7gQngSUDdHtKiuERnFMxyzK+Yhf58RMLBkMsBgqNOm8kTEoiQ
A8v2+BlmKon3dAoWymnjgnQE8Ybax6cCflpUHWX8vRBqBixEts6kwcdxmqJJ7k0I
lAQyWYEGsiWtZ8LLYy8yTyPAmVCdO8DF/3VJgI3MCuZMI5DqsbiD3ZUGbPWNQPHl
e3Jd7LOyggiahuOxOblKZX429dbaEgdIJEzTclMVX582Ci6/a37uXyy2zF1chLoC
ELjX+GZPB3fbTMaS+dBT18RTT2MneXhg0QTiPg1xaIe3Ma502nUfCWjMRT4lgLDg
KwSfCZtXPC18ReCPpcjRwTMIYMCzY/SmgIAnZlWVdy/Z1nd+vOIYdp6BNvWfMG89
gtxBjWSp+ETwiI3piolrdGTVTQ71mIQsnSmWZSvxZEEJDyCuU7Ux/F0VmNP6zXA6
xGYSi+RyGLS91LPHVKT49dswqysAje0fbEmJmw7WUEEUmRf5vH2aaA9hm04nobvz
lPOmdUZAzKtDRVrP+wbIhNFQdkrIePOxggg+tffgnPPZpiGX2vDkf1FOcCCR04hS
oMV4HLK0MoCYnFGP5Dwf2vlCH17zZzTJDitqD5XpR20vcAilsPWw/E0HMd19xuoA
PIOXMgYiy08q7zIxUvR4N5nA0yqC4aUvyDvXT1GYDeKNqOQ4eR9cAQ0q94baXaBH
peSEPSP53cmM5CvjC6dIXzTrDNHlGHtDey5aOe23O5WqWO3MNUt83H0mu4C4Nj0h
gSp4nOTcWYpVAsscdBzT5RHxKU/lFLh3Dh/qX4OFmo7vMBH4BON6gNE1rQfENpnk
+WhwVGOX5txpHbKUIg73A1SMZhoW+SrNilDjQsqA2XN141qtrCirlsbNdHwnPdsO
NvTSSDsQ4YqGpwMXsa8gL0WQeukbWyANSj+hvweXl0KOJ0SQZuOqDG6gL3FeJvPJ
ZMrc9zpK2UHLw7mEGWDBPcqj205PP9DSfQ5YjjiZaWGuARxhVzxaJ7Jixr3nU2Iy
2I0uzWCbTsIs42EkdySWfqui1/OVyuolIqFR7QXaTq6N07iyW8dxEZVBZuLn7FOJ
YHjGH6xsyRvlaSr2GFZcIDhViSw9uykriNdqBpwb5kdwZmK5hdSsZOBgsAuHtg3S
+GQeaHK88g6DzFjXj95s5xz64RESFf9BvhLK7fKpNzeegO9kjo+mxqWhQRL2PrxA
0Gtjo1Xk6plhKgbP2Smegb57RyjBuZr/Vxy3zA7JSdq4QM8xdywh56DIyPFgty8d
aMQRuhMPl43rnrmC7FK5eLzm/jsSd1OuqrwRXHki5eilOIt0d7VC2WD9IO/vq1qr
YOO1V2DOAEL+zzuifh4s4v1jriTbTS71eGPrQitV3kFE2VUba9zlpWMttt0wS8VT
Z9o7x0v9+J7IZoedp8X//jlQDXExv7Z+zpvNhYpZRXDGwhSqljCVGWQ0ve34MBX6
7iE8Ro3KBEkWWYeBBfgh4Bv7I0+qyZhHhbSchtKcO5rgcQUhKNDrGD4YWbeNaheA
wWt5bpblNjsVwaed4LHr3cVkLRmkILZGhxmAzneBSQbcvHFpQY7zJMd/Je+3aGY2
8np8geKQ+4SFlxZs/9UyQrZOF5/w6JTugKFt14Q/WxSILdRukIPithe3efacMryr
CDvAojrBPadx93zRETkJgYO6cKUQvSxNAIMnhP8hiFRQC3FawcT+NV7yF7ug2kzb
R1lMYceJh8TdBRk9q+Jm6KTLxIYGL3XbT2TSIMOO+iWcjHyQJJkBLpa5qVQ9tBFc
gvamGQVhMK8iLK0ZhyznsKtXOJKnacvKZw4SHM9VXZt+R2WY99bwBFyom5FmGxhb
WDuMbGAcdrBT87LGSqlQ8WmEsB8cIKG7CRLHhhiRBa4VZ5TV/UAJcFkYCpT58qff
HzW68I1FSZjXEgCsf/SyNYOjIhfT9Pck1EVYQ4QXWEik7mHCXeNj+8a0NdrLTrtw
vMmkvVCNlBZ8YYCoaM4UHiYVB6h330WvGDAWryGT07f8z+xrs/R4Hj+frYo7f0EB
RpqNcAmr7c69OeoHl6o0vko4qDScZCp8J3m2wag8Yj+t/8oHYiihVHc9T4BoJHsb
bE2N9JKGPIwhxXDsw6E/CHfrzxOFHM/O3U1Sv09Fem/lcr3WHs7LDcvlxniwausm
rBObTL0TnET5E+l6n4xeC2oc/7fuUbq9E2cGSzwxPQpRclCpAHIn9jW7YaGa6Xuo
+QTActiC3kijb9yUK4UPYP2AveybkHf9VeJfs30ZKdyEtdshLDwOJ0jsbQhETxus
wbMo7zrV0RGlwi1Gs7Kda/N+6f3fCLH4iHAE8brUclQltApWnJAFzQDcMzaCx+Ue
swWtfPnHWVNE8njDaG+RT3oIfpBJnaMvWnG8xxzY/ZOrpT46QOEPghEsc7wNB4XH
AXI+YRGgjXhSOHgGf9XA0DtePZ3F4CrNc35tJol/HmwuYj5tNTpQrUV0mWFfa41l
VJsfDxrbDed7+zJDkI28zs1hzAhEenBkeaN9KDr5LXK3gR+7EwJ1RMxmNZAH6ba2
1fVypuauI0Cp02hXw5s3/YxBMdroxreiy6cFQobLZpvM79rV+85e0sgqlIoQTwRJ
EjIwthT3LwddOpChuYnctqHl970cXHgh790y81dOaCyIbgpgSorxCgkppL0TQmgq
6Wgr6tN3KQC3YAkAkwn6OJ2MKMfKJ1glzdJMAz8N3klFcy0TpVY95DvaqN1a7FAL
T0+6YmcrtORdTuaMbVJFjQhjsU8N719jMv01nD+aSdJORwRra5CwuazbU5a74VXX
GN8cXm1KYOCPdBvKYUl911An2qR79EIvdlA2J5+8xLI77a1vksn8NYa10EOu3qVG
7xqdpKan1Rc39WeSwq/nUEGdxSApiJmlrzRKARXJSja78OFUlJuhZ1fHFPQ4GNls
Y12YqKjuxe1V2Euyc0bl1NVbWWu4e91dAM40+1LCMilzvfuAK7d7pq7BXTbk9tBK
qALzFqinsu1fajO9ZNjryaH7rwJkZaI5l0R900H8eL5Lc6BSw+f4jcRVNQd+vrz6
lu+Xsvn1Tn8wZPGwfrDCyyBIsMdZTKLKJhfITs9MH1pHE2UGNjb/hBNt0CEKma1P
zkW6FrXf6GjV4VsJ4ExV/vdKHfwuIL38dV4tfjs2oLDCh/1FuT9bVjP0esxuS43q
afM0m9UMe8Tb+YveDZfo3yxbnSCBsJTyrorfMTv4iBwdu7ffHlBciaB+ODqSGUoE
ZRRfvQtsE5++FU3skey7KsuC+JDL7tlT5b/pWdqr64HDRtg/5V91/37a/EfiDawe
ulR7ahD2xzw3pypQcpfx8+gZyWcr/KAjMMN0fnGWPOdloqZlk721enQGhFV/3Nhs
H8yw/4d2rWyr9eG3DO+68d257VEMcgWucU535kYh7bPB1MB06hftgDP4pnIv+l76
UMgjrS2qQWHCn+a49/9XzcseyRjluDw5y0uDKbdy/oJWvlt6WbaO+rGnTjnVQ2Mj
LVyDxP9SGx6KKoQKhaKL2jGvN9arfYnv/Xy2dDrjYzUUmtIrD4MsnIqLuDrMRxm0
hzBc7UMFTQJ4y8047aFevwYYG+tACZGa/keYUhiAGrtkCcz6/c5D2ayJrC01W2ET
nH65B08wjnNJwSGAONRUJTqlhhdCfQNfYetEadsX8+glwdTVDb7lsmQ/vaclm4YH
3I19Kye4mcFmAej7I1+z3NqdR+nw1NLa6IYw2alaHaGH2oniUmmh/UzRsdRs+g/S
Ob2Hm+yQbSZbML65xpzYjv/8a1OHfENJdboGhZXb8fdRu9zgXAmqgMUH+6bu/0O3
gb282DaHqtnrpA4/eofKteDD0tT3yF8M9Fcp+YYCDaLn8o5qt9UMKXa7xhDXI+x5
Yd1x9wtL9VKhHf/QfvQhSyxGMqE3P97sKCJZahLXvK7ZJybAccbRovaiS6fO3A3S
BTBKpsRyTH3NvxUkuWSBEIyoyGCYd3hvoqV6FfrXQuq1kozaDH6LvdzK1+EldoIV
RH6c/vrYSeKXqtjOm+5LVzHB69++WI2ajnFZiRvcorcj3xRTxSOqYpHjKqERSlQs
dXid8Wbz+OXTrCCY1f+SL0sGBAzfdNiz45uaPSC31lA1OtjbzClrtxUUCfeOT6JV
BHBNwLMaVTz2P3/PZ9CQ4QXOLJuz9S5kC6uuum34CZ7FEXVXCnwysPUP4lszaTEi
QiETpHtRFkI2J17Fv1x1ONc/prgoqlw3rZ098obgr1HFL4sYpBKTVYEYrfGPPbef
ffVeopD0BYdsE7JbqI2W8uTw4nhsUXz6u7pvc09httjQADaKQULs8KHPAdQUQgPc
bSHi2lBDWX7qxysJi9gHJ/9QiBg0xSYDqe806SM7tXVCBwNKR7ZloAz7Lft1Bo7t
lp+2IQZzB2o2SVHsuWBUwQebiNlKYaTaQOTu8Ep9NxlMZZUa3RBHKa2aPVrDBtOz
5HiezAcngwYbyds7v/JPzfgb+WZu/1UufxuNXlzyUh9kQRBiKZD10ZIXeSIx5yOB
Cld/03IbWZVZfTlFZznHUVqDc/VnmxDteMOlZJYcA+H8drb5uDdQqPBcUKRd8ntN
dTDVgyeuXPdP7honXODWGBaZDTyAmokEuOxHzt4Pq5TxDm+Ec+lDtOGqPCCE35N/
5BVE63ZHftbmCR5zwdj4KeLeJr2Rpn1nidTUBLyqrBkGmTvNWCisItKewlUhadX9
7uTtjqb+DbBpEg4Tkn9AlurqzliXMhc7NFzYGirnTyE+evWjaJ4DVmA1utKJ6dzH
T7MX71mtI7rnWbdWLmX8HFeVlgAvKg7pnEhst4UbFzdJW/lSvf95Tn+ZBRNdFrJ4
Ac6HCTt8PQbB9lfRyaJFJKlLvTnNzJsYbk5RvrH24UDp2R7dO6zfQo5QsIB+e99S
FmYrptlKIIqgiLq4ftbo9+Npnvqs1q46cjgs2fhDcedWLLbDMVctS8ut4JLXf1uj
rcAdWBKbQVUZOO/SdAKGy2/qK1MyrmEpGit5pYkOvuZ3M7Q5zpTM5ud3JnX5LNao
KFDNsm/Oti9L/45bqYiZPUYZzCa7+kYOK2VUr+vYHDDfRy/VzuvqTq4/eQvcjPFs
OWPYrXyRO+NzHsa9KKOxWw8Rbs370Ulpo7P1cevGLndvsI+n2C1YIUjdv24bUjne
ST7a/bUMkVj1uwJgABv7J8aGkeA2X1ZRujx6QieJ6xDwsFHmphxPKbmY8TR/KhnA
pjgUf63XyM+WXzycUA61Dki1dHVP1buYWOIzIyGQsCKzLD/j27q+gULdrQPJdbDG
wSi7llP2ZfW65don2Lm1ooN2jjIvxJmZhu3H6FmyrKT4diE0DZeb9HYh0eJph6Tb
pIVAW7U8hIjJ5obH9ImWR9aLktgoHchSdOvlNqQBYOhy1GYCvyFKIyzEek/4FV97
3w7GUvuqmaYfQ6yKiUrxDG2H++mgt4lzudRDQeR2bTz1LDFgyAtutV5uQMDKmLsi
IfwWu9tFSnAeYG0bq9SieFOWWLNifaktFEYWSpLJfRwe6lX4Ox6nhZKa1oL5HLrO
J92LcCfcBYvoJHCsB5WkTnIUQ6fB5+Y8mSqoPquF3/33juArv/nJlBdTzX2Jnh+q
ObvfRe12CL27LEfgu3DFNWfhZz+QY5yZVRB4eTKholbANoNEeNq9oRrs1O8vDT4Y
d3Jz8KcqUlC+qX1hwZpISudxQhlfwFwkHrpaQWXO9i/TNeJVDn9cIAVEZyH0E/m/
KV3wDbzLcRQLxY0lLf5B4L1DGjYC2WxHD7HBo/uot6QZIv3clRqWEBeVzIZaNhO2
WnA30cmRl/VFVsXIBeV1WmGpG0K8SXdXatPyZU3a25yMiSiKY5U9jIUKkSlFzN44
mB6MJIB00OIrRZaf50vRsuUSDiTpKS9WnsK6F+PC5A1P/gSl1zsaGhU+GNyK9eVu
V+a+fkwZ7ZTy3xHHM9Oq6zF/7K3AF+4RBSpYIonTVm0lnUKUzHsYeyTQtiHx8NkH
JGGwYqm8t2PjNoQAdE4/EzssJp3xI/gvwJ3TspV+2jPhEsHd30y1SeES7aUSTA5I
nAVnX4nmRc92ctxaVegDjk4vItAr//yt3dbf1OqY3Qf7/9B1bvdRNP3L2+XiPJ/R
n4CMR6WEte20+Rj10T5LYZ69v7lGuG2tuK0nCcU0m+jzQU801DL0Im+3fNqBGZe/
meNhVu9xdpf2DWC1MJTr2QSwax3D26GZ5jOqUwz8XQJbW5X7xnhGkFvZDPN+w0PP
8iFgNQg4Ayzw7U03mRy/9fdx3v1zI7JRME5kceQVr1jAV2uGDEmsulxBAak6g8Yk
bKLQQbp9L2ItyYyfIcyGg3++keezOTp9giPzhZxnoRYSOuCtdUSKN0Rve2FGNFXQ
S/9v6Nlq9303+o/NQ13kQruSu7QbIi+aFFXcE37KRqdGXlDevhxldUFUe/L3pHZS
7cSrWmN8gvvSV9UGsQGLF4VYohz48cw36HYvrqDFBbvhLkdpUdD5540LVpCEU81Y
z9uDx7zcZ7/mtPOjv6c2XAjfj3cg86tZTxNAxlF9/4PFWyxBKpTRtnUbU5QKWeLf
2ZXMbqX1G8q5nG4417sfWmlR9oXuz08DXT242n0nSpxMdYCPgSFbdxhaIuFmTzo4
pUiStVDI3JYdzwAOs3aYtGKb3qNvAadWAN/Y5+LX8sNpcZPwfsgD0ht2SS14HPli
I2phKXWIzkm6F/3x92ow2/qouiWFhx6ikUuRf2GIY09kdRGkBc2l4AcxMsUUguDy
8NUZH5ItNYnl9b1P57ZnJpP9oclfvxFP8ni9Y+PoTKFLamBjGX18LTX4bRAR9h4u
PTIK0Eh/loUZ7S6BJbWFt//MzN8Ow5ntS9/KSFw49Eg7MXtArzmPNtODDrtnm8yD
3LWnfdvYTplcchCVBIm7ia5YYVy1LqTrkfXR05CHPJeZy4KtaQ782N5FAXBrC36A
pmzwKU+jNIDEHTnZjaXA/5l0RKoJvC8U1bh1mEuIwVHn93Ets60KwTThXvvKDhF9
i31P22YqsUz0dKap1s2y0p12TG5u28nz0+2/DPxBSuRnP0pnMrfCxzI/DTZjs/zr
bEotyZwhOrwwPYOeXPAL34jFtrJmmn0Gi2Ce2EK11CdJOaXqgH5nxhb/G6ooWyuZ
1WqTtbO4w5VCF1t8kViJjyNviTjsDB9ttCQwIwfygLWJl4zIX9XJNFk7r3XJo1jY
3lY7twq3CXiyIB1bt0vEeWWssmvqofa2kxOT0rKpyu75jOb3IjzUTdxanlRnQfwP
EKo2FioilBnhWSqvEdN/lILjJWuz/2x4mN042q0qmug/l7XkWSkdTLNbQek4U+0W
vIMHD4c8IOdvZxMLx5W/KgDvJCQF8m3Ir7tEfGucDyu2VXVa7znu/esQ12KixQkO
FXxVGQHA3EQLTGHiubs0bzUzWx3aSjiIT8TsrgdA7KptmmlnSgYnf77/PmHj4ZHw
XPx2cle0mADbcxf+w8XLGwvNVFN6WgCmRkQzjf+VgUy2tcTegTri53JvnqSn6qzC
vOJ8k8h8l7EE/tvAXmmtcTyND71VbuJwL49Q8rU9OXr0U26ciTjiIyfKAopO8N4G
xA5ZawkmbA6/t2ld87fKvwAoOvIW6dInISW7DBWk3WohbhrcqFZuCvS22dJMmHk8
rGHfZvTdUqtkhBzC+jejqPTKq6cm+ZqW4h4BGS/Lm4GZwHvMJhMNn33r2P6RY46V
RPDv7GY1WPz16q/Gptn5wqvLMbYlZ0Qz6tjByJK8b/kMK8H2EgVzfrRT91ea2mQc
I7faWTeqMZaHwUpBySIbogbcKjBjopPDFgOW6BaMyrNt2WJdyvTD0fm2Tfv1O5kW
VdQlvIqDSBqUqlHVKSvPHf4PVL83l56laQPzO878RdHaJQBykOqEhnhJiedkUfHJ
PzyEG12we5q+UBk06rkvQydQRglNZVDuz0YHywnH+453vnY6O5qSyWRBdWboycxX
+nDXoFxX7NrHEGn9R0gLopD3Y1XR7Ma52MC6dGZx41Ob+OsFZqgoiC9kD36ehRp2
wz4MhWqrHXf/5WxpUzq7e0Idx+aneZncWWfBssHiSKgkQEPzxvoQNh0NUvGwQ0ZM
PJHuLZRF+2hSynUT2R43tLdnRag/XBShirnrKM2Ill98wqvSx9XJo/a1EI3RRAlj
lCT9pU31yODshKrYC6Ejgc2001LvBHr6dOJAFtWf8i7uf0jn3mIaga4EhE7ePS4X
mTaMlL4c1xCDdzfQelHVxnh3SgaAA9kAo2Y0Lm1cOFy5+PGN3ftXIlsaUHq5ZS7N
H0R4sbgroYMDU6fuG2rE4/E8QhPShgwX55b9JpNG8CBZDeT9g3qUsLpnAcpSabdo
nhNyMwkesssosoTPGjHnhn1tAerQvnxiVPdZVwFDDHBCvIkS9EgqVKwBen34+Sue
5Urn+sCYv//G6w6ZeWP1Of2ZDkvCjG/jAk3jJxElyokZe/j00c2Ips/1UwUNtO8f
Ifex7pFLAEs5iSSeordUcwJc3BnX8opy7uW0UgM5Jfwq48ZjdvkVJOzGESyILzGh
mOLL6iOqRK8RV0lvm15tNcRK74ejRM9b49dc6KOBRSMbUrseqImgQ3wEC1d93jnv
sKzpxztfitqV2P67tKLtOrvG55+WmlvdeIS96vDByHbfsalpwoAk8B4NDqkVHQH8
QlTQBTMgXwahy7dqBN7OXN8b3hyqjbHm/zcGy+ff98C9p9VO381+2mukqWgXWvAt
D5Sl+t+jP9oHqHv3ZV5f+M/x/K1QRcIvyoLAm1iFVPGUwxDJAooXwZKGt7oDn7mv
uVa6FhnhdV5uijrctdHAhHtT1yGCSSF7SSnsaVMiWO/sEcdvOGlR4aISdsjwDPFh
MFVqzMfJUS0R6i2753fsvaJgNmOKJquunmst6soqJYpri6FBFzTf6y8zdUUJpuYt
87hUcHa+TGs7WZRe9MkGxI2GKCsHEgAsgCNXIa39BbRupQRVbulpC8qruGMO4YK/
ZmHsamkxlSfBo/xo85S0BFhDFpztDdrhLBqhVcxPE7eiU3W4VyfFEteXxET+T/jq
vJOMCQmur9EhCsOVZa3rlSz+ATWbnfkzmMmVwbRUQzKnf7gMXr2P0cu7g34aUD9M
yxVCfx4PBuHE4ULJHrCkIfS138OaNSBecmpa17JZbvBvt2w9d1rTiue04J3S5Kkp
rAjs1a1ntuTLofVrJ4h2eSf+YTw843FNKGXLg7/8udRebKcZ+nCXwpyyYSdtPw8d
464DjRhhyxSPa4ooTROs60KngIJ3g6iNl0L8gb3W4WP6wZgQWSSX63VI1sgkyDqN
etUWnrJTwxoKx+GxIRDacPc6cSF3iW5cTREuXo5TQtfNHeR0kgHlVTjfaqSPBzJ1
CE28DFk89t56jhsoLOpwyPnhRUdy9jkFR0eRDr2BLY+1kVFOfawey8t3WhD54haI
GVLCPMkSSjixArlJwMYqcOf7PQQ5B7UR2NLaOKF+QELjKSkWFRn9k5aTfcW/vqr+
BqCxK38n61r5d/WR2NvwM2MkwSIkArM6Mefo9vk4szcQUeAJxLosEbXV2htT076u
aUkYzTawN5m5YmknB3Sx+KgMua9ZQy7h3woumzCsPcFfQ25EV6VTfkgvtECBLUNf
CIU594ncgkw3V+KhGrjExddcK1RGwXgOWL7Zoqmw8kOk/w3+69CyzZO8VYTaeCkE
/YpL5AdoTCPl/ySWHBPhiRdQfoacOnfIQunxWdqZ4TZ4AptXdSTLtFhgGU6g+pQe
7Pmoih2DjINZe9nI2q+nl63/BJo8mP4dKGVdKWZhusuBSsABsuQCd5tXqeEGfjpk
8wJ/MmKl06B7QKaiPCjiaSqw4OYnl5Z+OHVwOmZ+i/W9INhQuAz3DMvEvXk+LXYR
cotv/v7rJY04kxVkULNmFzvo1wxxmvyW8ga+rACLSpQ6ogGUw9amEdYYTP537sy8
cM4OPgTho+t9izrSvYOpVmrIqJ6FwkaGDZcf2Ct1m5VDXmv/ZJvFBY8qQEs9X1WK
mV+e6qYo20FXoLq/l+xkx5ExW3O9RTq1tYm+lrEphYBiI713CW4corEYfvwSR0rN
2TqQdqmxtqavMCJpnz7n9kDDTchaB53eUxa8YXKfQ1Ygx6HIR/xVvQGctVvITS2f
y9VYPUB6zTpkyfJUMzkqTTdldYB40vHzNcng5+7q6sKUh5fmYJRO80YQISaCFpsA
l8dd8szH90Ze44Sx91cnq6NRUPX4RC2NldEt6dlFfARx43W9fW2bWc48yFywHXSq
jwErAxcPKi1QpjShTZ2ubV1mq1MveiqvU+ccYSZkL3rEdmPrh8avZl1nqUGBt7je
e9hZ4p/gwFMr1fNApNF9uDYEDpyIld9TLa1sEgtQJgiqX5nTr1Ug6NFiWzaDnk9C
TuqnDPbeiftm0N6CjR/UNRSe5Zxbi9iM6unQQqfQfCp7AQ2UDhb789nnfFc6I4wG
62r5O7DTjES+9YeX1Tt3lZPoGtAyawsqQ0Nf8OdLB1DKRUbVEOvSSSajCBoCW5mw
cfeL2+pklw0P1lmx2Htc2SjYpfEt6Xz/N6/sCPsA8rLrUXR4jmM4U0/liEVng5Se
BD9wm4GMO7lrnPMdq1mfJSNQ1NTNwGPBM0hy11ACi5dwfCqj4ponjmm2jRkkjN97
H2mxAn4rhatWQX3LQWnw0k2ANEJ5oL1ClKra1MvUgaSoeLbaiQrTh9e46ke9iS6e
AfYKbMOPhhF1/JP62T80EgFNNSFWO3iyl3ptGbIN0Fh86AO+YLd0xRYdstTDY/1o
jjQanC0YR0pL0EGjafmXbg3+ItIzsd7CwWiedVnBSdKKPmDSQQQBZn+lll5qH2F+
HpFYf+FT4TbQl3RPAGqMgHoQIjToss/8ntU4IkWYMUxT/K7egJoFeEacXXpxP7+6
5mhCjc5QbMeQ+8JyN0TMsaW6Ax+aCOYifRSazfD+fQmAoecTb7vHcTuBUj9LJ9pS
YgBDvjmPWOfOX9tdarOvXioTU7vXtewEcocTMx14nD8S9dVZ49v0Mbdc9cxukwwT
uIHoHxOpDALjn2CVMBoi17zamB7kQ0SDz+3Gf+D5IYwrt1f5RpK9Bmk98hJ+Yjc0
0ga7Zt/8ImAqLJwdDCkjYmNHYJF/xNM8EQWQdBEhRuppAut03SzQgi3MCPGZXWUf
Kq9OFRakyyGk+gNuTiB0XKyxOESE7uR191EgQc+9h71Wf1p5JwxVqxBQ1f+eUogF
SoTicdpkM0hcFxwTAEWZ8oWi/oi2Olg+RIpN91wDa6K5AFXi5tAMFEULGiF/ZDGo
zjMgZN25QDWo0rbToZlC2Z9H9oy5BEu7/M3WhSC9qrnxT59mD0p3d1RMMcvVO1WZ
c/6+ecvJb3wTw5piusg7GAKxm3eugTwY/VjhmMybiHnj0BL0BhWYUWOpdyoSdr15
dr/9g5GwdfIxHmdu6JDan/mutTNA0YDZ8j4UOGpfzf3PVh46A2NkBboD6Iz9aVxC
hrgS0fOFBT0XfKdo1bMYLmUw+aflO/xZrYMws5pMYVuqRgq5jDHFSbufJCnD+wbX
0r1k7kgDYB8sdM/DieBOkjvVeQS80L+4wd7Z6Fzy+9do9Dmvb7M6lk6/eMQcnN86
OjGC5X9WZ+v5qWOm7wbUm0yN+KGiLHxAllc42tC7MIVNufHSCjy5wpFUpDEZOjKD
YzgIk4JVos37hlR2BCfmtF/JNUWAjo+fSvQhLq7UGdzLO+RRgNRB9Gjicuetw0LP
KeTHxWh12WQtgNSKsPxkzxIUYkKEKCpkvaUTvHQ+kuRXqwG25WA2Ht1eFPiqwlo+
9P71WzDP/E3Jo22VOqkxYILIxa8TU6TAp8pmxVFP53FRag6bl7qLtLvGq6Ocf1Be
Mup2u+P+ZJT1uw5DPTKUjhHJWXpiRZrwAPSZKAnI6u5PDluAo7tH/nCeKTUxs2lj
RZsc9bfnp5zLaJQYRGIPoFHEdp0JM5DhcOEbS1hxMZM/N3dwZgHSOQ9mRWhqgCEN
jPQt/gTNZTtSmq1FezdlesMuV+N5KZyeTJd9YoYOQPEcVxZC7BW7Ujt/oy+Ep2D2
+W17fYaLCwpS6cjXyfL/mJChsJLjb4GEtq7cjxu3OxmtG6e9Y77UWWYMWR6X2Mo/
LQhw5/Uy9hfzKdopMJ2COYG3cvqL6/Li8fBF1uJFQFUpbwNO6sR6z/RLZnVtPJxT
TW87H/X91l7/48GdUfppTeDT5UYm+ZIp55QuOawA9mg4YDAXXvlGACJbJD0SSlGZ
UihAknLPD4BUXQiAwKNJA7yw/xOSfux9vvn2jDM5et6cWUOr/IrRdULH/pm5rMl6
m1UoyWYbuHyXX2A4G4DAJiCj/BPZeAtr061R4Q15XPyIClG06xW4nmn9+HY3StmM
X8xfaAHzyNltaouFXHhMPxSU+2aJ/17cojG1vGrNJqkHDDxIHwzOHk7n8MYNOmDo
+KHKQ66hXybheDH42ojBC97kRxa2T8zULF2YF8jpKeK6dHag3ZwVvrP0bXxyNtJk
uq9dZKm/2kOLe4P5h7LV/FHoSDZ7x3E4FASxy2mRfAOrZ1JOiDcZBDvYUGU5ughD
s+wVs/3SE9rpCrA8Ro4eil2SUd8l6ZxQu79qn7LKiEIMxha9vuykEKGZ+z5qLYr7
A/z/TiL/eM3Dytk9orW//uDpi3S81Sa73fmjJ2KXaPyIgJ717rJR+wSfBVp26CMe
gf9GIeM1lGPC9c7IpPCloj1/H0DKs9vR5K3z5nby2Iyz6Iwiz2H+96RqiaeyrYcz
JqYat48kr9oZEU6I39EmZQm+snfGXjUfS0BnAixUCcfkAIR4/bKkq/IcfGbCOk+d
as3mINL4lUY4XHyiD68q1qknpJVgKtqJpANvI3WdMjlgsUWcf9rS6lcgklHKRyZa
ObaaT0YDNoLyelOLQNBJxr6pbJIndxRb+i6G9IKaRdRffz2WRVNvV1mNpUXCa2yt
g0FbvPWWOESj3VQbUJrqnihEC0revOa1/jKKlgdDbInLyPV7MZUXb4EQjsIfeiu5
3ARB0Lzej/sLI0LZWTxLIMYc7/+0eqNK+jGKaB4/Yy6MV87YCsdMB+LC5jXHN8yw
ed4P0CW0SViCPM7BordWCpjVR4VFIKoHDM4KWF6fMB60x6G0lFZJ5tfdvjhWRwgv
ualoIMskYtHGG5zFWOGGHZJqGkOONVLhcyalTvYBv10K1rhWTQVBi4SR/WV+P4uH
Bb8e+s8/czXaaIg7Jv3BrLALOPT/r8TTrmgLSplJueG6BzPbae7ufS7Hwnw9IgDO
m1aYolGvhFH3UN/f0UCOnFt8MWM9ZhiOdec0zgfMRkHYZQPH7yT+XwzfU+s7MUtB
KN7PxXIJktw1uAZiMCZOJ6lliyjBuJImP+LXZop7pT/2lnwCI7jZ15LgAnWJypeD
Yio3mg2ZG1vDqQklk2VABf+nbW/hkYKjrBOAcoYo+dqGu3fAymWy/xWtOWcjuO/L
f7+TwYNgLgZC/skL8ytk/OdOXRZ2vAWL9Pb+FmS9lr3xdGVJwF36B6oaL4VyTfhT
YpIViaPPKjPMI31sgdCmtfsDH7QSjaaikNZ2XdVCCC6ekIVwbjW41FD1hkT5dCw5
O03jLhN1sHqUy76gd/fYKxIJZ7mxlQO4aBapm0MksbTY3TtJdoCaJGA6JgZPtLvO
Lvsk+yIwbZOYjS6x2iToaiU7NDqfaX0dgv+LW2KmFmX6ckYDuip/iC0Y+ZNXqC1g
6dPVarWN/f0j7NpCsGohKw0BRZxpm1You1IvCZbY92iiCQm+PJrDJt4716k+d7Bm
Mkd4knYa+8WfSOrKrSqViyTDlJgZ3a1GSzSUoFUQpu774NxfuejZ0d3kGZp/g7CP
Qvuq2f/pOmUCazq2vw26zwaveuwE6BIrze66Y3qbfe9y4XgEQO2oFfpW+jxH51Ik
1DPU5WqHd6tqX+fbiAnpC7SEc7binxu9g6WG58+Jt+V4NkCx5CWSh4KsTfCt9w33
aEJvYQqyWWgNrFqg6VlDFLtMEwg9lFDvgvdmDwhWF9pCq5BX8YmUUs81ZqEGKWIR
0OpzkFiefi1AndOOoiYY89M+3/lmoSamjyFotV2CesCABtORpiJFOEBgUJAOoMI7
/PhCeccq2YoZDgrqELPw7RkccPoNEebzddeQyF2NSfcMS+vvkWCI057tSkMdw+dh
gny4ybud7ClVPTADsDFjpJQ4foHcLOEAnMTjpicxsRR8PTLaEws4y1+UV/gRJOcd
cA0KUIqohnSB837UJs5HfzG5+fJz/xcO+o9qx3dSmaXwmuXZr3bUFhMisJE9z0nS
2yni/TpscULRA3ewfIdJOGxVRjrbev8rBYiWTIN1cVwbPiobpYFfUFe2FfuCUo45
hs4kfkgMJ/hn+nHC1M6lsaLLfaaLYKidu9zDoCVG0NCtFINU6DEvKSWT1wdJC+H0
5v5l17b8g7+oB9J0HfvcAmJTtMEoytSqqCZVRBLuOeftFSHr4NirqG15YpzKIlEA
PlCVXQfF0QlKTOnsWGIPqTdBIeOd0Mpzl1XKYSShnYZh/+EjAenvkmoLxNJMgGJG
9MiYYovjZnwZ1LU5oru0K4Yz3dpx/UUb28ZLa6g82/IIjxPVoFLnvwm2Gdm+o9Kb
LhUV+aglHJx/diBJ9OHyq4lQBiUC9Wfxrk7hZCHRd1EJUVguk5pForBF2SScp3GB
ufyrLvvBsfdiXHW+fLF2VFWYIEanhpUQCUtv2EOM52EhOl6d6ZsELrA6f2iTPgp+
jORK3RTX27MqSdlJGhVtszr4xCc7tU5F6BFjo8R8/+86WTK6bg6YaCX6jk7WWAnA
wkwuM2sI7lrymMa1zE7PUZhD8n5NpEvnCURnkjaJAsv+HIgN+WWyob+tgvvrgC+L
yZF1/Bu1h8btflbgBPVhaIhgw25MCe0Lo6lTX0jtiCu6tlh2G828KKZKUa8gGEzk
nM6hDYw7P5Tr4DjCBp0X+EE1cwFqWfWUjC/tZ3zC3WdmkbWncuM43SZqY+4aq3ZR
tYVRZRRfEI439r9/EMAOgN3BdkrANsAChDAIcn0juhXah2EMVRkMfI1yQrj0x9XW
OBbhcGhP/B3/Iv30W+H1rjHlKJbbvB40paH9y2EaBrxr6JZU5BXfDczhXGRdxhwU
QylxuKFy7C6T3fzUFwAtDdcWFmTrxKvVoMCz2ytpH79W0XfVF/b6wvUdSX1pVT+j
H3IKVlYi+A8rR8ZwEKG+kxWNkvTIpA77JPweT7slx6+qFVQV4S6CSKXzg0Y1OY+s
VKavRtWLewBYwrI0FD5MofF+rLWvsofflHzo+nOHWbMonOQXnYza4OKzJhQIRJKd
UAwWTcQ0do+TZgEd8UcGrAcetA6rJoTopiaoIOsIQK9wy/0PKlgHsowQBtTJHkOm
6YEbrZp1W9RBb8g4iXaAcZsDvQoI8YksTSeTWjhlimB50y9ZViFhstkdNvl/GIqO
JddXZd5D8QgFDt9fRCC9WN5NxuBjHpOhFLIB9XfZg6w4zFYEU9DLCCyRNyUo9kfy
S81A5DyYkueTrKHc5k2MzxkxIZ8e0VIraI144IiHXjtxUFoaA9QKYUislG2Iv6gz
6RHcJNO7+jvzn8DvTKQlzgAHuOspGrMDdH/13GtEbn4VfrILfiV2MDJAPYwDMda5
YYRl+ZX2vR93Af4J90P0580J5hW2Gb/rH7+xUztE+sMND9J95w/Bq09zjOlMVb7a
HQzmqIa2QfOZmLUJBe6xCaKowDOAFAPEVGKvkgPznd/znzfz1QUvmL30/wjcyqZ3
c8w1VpqcFSLYUaIbzRCYboBTzdpH/e7RKh8KoFPWF1PWSAPdywk1ceb3APda+XuR
gP5xPa/NeD5YhsDVzrm+Y2G1vSmqVHZpai0kGg1yX1dxExe8hrrEwsfgBpR+FhYQ
26cW2jbTZALVUg+2WYn0u1ZpEVR4CRyJXSUHgy4AoSxbqyYx04nOPXlJ+5o79FFP
3EcxN8CTy+39MiuICbOrb3AovhZHIykyrwtRf8kYB06Qd58q8Q8pNmEnVb19JfMy
UmkC3iR1sVlp6D8sJSKcETeGdbh6TJ+2aphNkJoWL6uTirWpNp7PCQXqWlXQ5O6a
zSz8uVdYXaSKXkri03xExpnAvlINSOQrsaqEo7zF5KUiYtjjk7tIffrAsYRUSxyH
mo/OsvVDcU1+vLNnxwnHNOXhMUmtQ0F1LYgeZuBDKiW/morVbfHwu5hdvpe+lAfw
IZOGVzw6j6aqZu7MrZOCDOjiG4TwlxwNnhuMjMth5T0Q5j6n7s8nU4bdsSD35won
wwzM74IMkWud0ZaQ4vN2v8tehxthlMODgnDFynOuuoe7WGGCrjAlwezC2PG/nXI2
Th8NzQLSOljn0dkAijhsA6YkLagHciLTxMwtO+ADqupjv/p+IXtQ1K3liH6YsILW
c68+bDOnvrET0+pY/HaTQd0dcXpByA0wDDvhnqdpw3kBvjgh7kPuHSctA1raQlxN
oAu+wZUcMJXO4rIxlyQ71nzAy0tIEpHZ7nmVSNCXP+S4HWLa/JMehuwObyEvXM0C
ukQC807PBD0KcOdqeuGiSzI5lJoda57Yx/a/yeljH7Ax2KhDT+gjpG8Q5m+NDwFY
kQSTl1+Rv502e4LrSCo8E29xWsRcrJcOqtGfjR0/Sjdxsm/r62O5/GOa/hOnjoFg
2usiqNA/DruEqsiwZfv1xgZw6mcZYfruWuIh4aGWbj/xC5FxQZNcxnB4uqAf8lsn
8ustGgCO+xNT6xiNIcXeu9NZFbSGiAYzyEKturnfqq0wTPAuxH0NSIO2EkaHhIc7
m+4JvAj2j9sU3DfFBNNv2inVAYATj/zuQl1NFVyQHf0X871rOEDn5BOotAZXJTo6
U5HPplqvR01QU9EXYx6kSZycdouyNdZ1xuWnc7bpCKg2YkvftXwBPeLHVG6ZbVrQ
DDTqh6tF8uCvGlSAXhXrO7AjgqQAbfDLtIVELsy3piHYK91wgkgYXzjC9g4k83Nh
zqJhGGVjbCS2LioDJ25X/VWvlLZqtSzkDZe2qTfUIIY7cvNL2WsHeKPVrNdjQ5Ef
wCiGLanmfc0ONl7Zvm+zsUb7hsoj/1SCzso7CuAg5wuQbzyj2tmyel+TN5fbLkWP
Qh2wwEQi16mY15mIRUziqM7R58OA8OIhhExzs2qK189dhlvFxorEfvdHENRQQWG2
Pvu0Gz2lmtUf3W6YhPLm4JvYqkzserIP0iWJGRApbLFNkTKET/NA2TVpwwnXk0zK
7UGfPioEbmgzxI239t0+jrhLphvP/FV1B7WQ5/uqEu1BEeafkM+ksIQhrp/hch9u
K2bGcoPMQZ3B6h77TcmTqBXVZ6uqudJ79vFi4xywXFK7VaLuFoGaBkqFgxRGKueZ
O89rjqiohbo0dvG+DUThceR/GastjzbZS+iYfmYnqY/Le4Au5htLQZZCsr97VOtI
Gyfar4csJ7clseE+yq3WVm0zIURGAsDI9W3XcIMv3UzmSzGKKWiIuoaWSLE6AuLw
HyeMpm6bpqWH/h1MiiwoMH+G4ygHslW2ZR+Ur/b8o7YXz8DdXmdjR8Ka8eyHyE6P
Pufrd0TcghTFkqpr6yVufhU4QwS3r7FfZxIiWNQUJV7L6e7greOfD7Tc44dExAIR
IeOt8sEeAGS+9S4XSw9uubrthDpqX6kRs6nm/isxCGRyQNxc/NkVXM2hBls1M17s
VPi4y/YFXk1UGPxW9o2lmdfoQ0MSx07wLS6wtBZOifaqOTYYHItah6h/57c3aKp3
hCiDMMiF1Zf30+gHqwyP53GSkTXTKRCF+rj3+U0FZK9PlBSxild3erlDSc1Y2FVR
vnlwXD8zTKaNndpTxDpVymsCYYNPEbsC2Iks8Q8Ku5TwdbpyHH6OPwoetkF9B+pN
cFOPl6qFIvUmLLfCAt26RUlKov7dW4JHkxMVfl78/OhJP3mjN3nG/tazaa7amdon
4pSDWGqlfzdtIYSC/qqLVR377xyLftvls90nVRUUyKRr7IIwvYeUFUeAUSI7HE/V
NzP6hk9ItpBEzbkMdrL69zR2JaInxWiCBBcUjivwltNMRli8gUkJ413/g5vXBXlT
wkv+2IS3pA0zt+ufIV0Hy9AhRsxTnuYS0zdb31HqY5LhpFjn2UH3ioAwsHO676rl
8SoXSVzyXKmltQ9xzEiwvYgQkj7KJE/DjXr3w8EIsu6MK+3Mc7gMQbuh/mmrHXQU
bVQuzOVrUJOQe4YH1zljftqt82Mtm+V10RMWRjwbRZXGvhGFuZRItmr61iUVSCmr
zIyqCNv7sNrmLVEQ5xVHuDKnUU4y+a+2eeJUUAGPHMFc3KgOqRa4Ftw40NoJy+LV
Bzenq/hddcbTBeuG7LIYXEZz26d7I3U5mhtfCk+DRfrUjiAnxnY6AhNTn/Xs/4/M
E6SG0+qOSXi8LBvXrceM79PwuE11SZpnYG/rgMId9PinnkE6Elt1st9jn3b/OyZ+
V9KL/qtqmWKTow3QcfypVie+/vvHDdd2YrHmmlCrGFhFAiXJedM12ps16Gs7x9Ct
jfLPhBx/23WcLJjgBsFJ+7Z0y2k0wZvhtcPDz5AZ0Ec3tCjJa30xbaeCztODsM0R
z6zjIkdLKCVqiG6Rmtk0BzMdwkXX2HLU5Dy+VG4O5uZsR6XchmUeLF3huSZPO8eS
Q3gOqGdOSQedFDO6UUBntK0tTT2oUdx13MBbyF4l8HYcvR8xC9MsC7Bjefiu0WqI
NatOSk0ipROLnyG9ZTVeQo59JuEwX/t16PF9dY0jY758XI4DlOADfvT41Mw8vUgA
8SVKECppAqLwleBBP7r+qP0tDN83sLWcC0jma08dmlShxrZXS7NkIHtls7C81TdJ
SOJSVNntmjjMCb1ztdyXJIS8uAvvBkNM9uydERo4thrG8rj3ZA74EEM9GP1J8EB3
WB19kJGbAQei4tlTq2RNqfV4lmCh0WC8ExyTYp6QlxhNiLCjbC9FRHkhpFLMmu1h
J6GZs5UQV4IMiILJZDpcMCecipbwkC/cqKTYsW7xd4qd50JH1yxI7jNPRjG78p+g
L3g+GQLPdV+2MbX8jPIXYzdjc4qHZXSZrtr3oNNTvW8ytuWTObXID+aeihT6mcbq
TjUxuNRPnTO/kPCDL812jeqE5GXQZvnz+whHYhVXdCbtyJdHwd2YqcNgMx7ES402
Nevj25uQpjBR8BSCGckepETNeb3XCzm6UhSuBjepYL2hst5XAEOP3BUUCrHTqAVB
tORJPmOFWLl9yWjnV8x7avc0+vA7WyHg9X7GMXsDRJeRVJ5F4IqTOQJQdh5/ZCjf
T6R6qjJpopvsbXlBdzo7vmjpJrImlMMW+Up5VzWJHJiMC3xs5PdPRPwWvNuVcERl
o3mcIuc75RS20Tb7v2zdJZGgYJ7Humm+DrwJ0eUARw1XhQ17HT2b7RW9len+9sZR
yjsYMIVYTC0w7JspJ7sMZ5mYknkpt8XOdXMrTim+PLek9roBy7ZBSZsIjqT+lyjh
DmKJ3vlCyS3DOPjoxYruf6tOr5omgn+5cJO0YmUiIlh755JsYlVddBdXIwmmwni+
2l1CyNQNliCYGZ6CeHNtDCATOjZ5KPm4yLrh5hUJA8ar9QdQWw5E10e+d1CEABNf
0lrs3BTqhuwymqb/E+gR//6hqYGSaJq1DpHEbU5YovTj90BBqVtY5blO4mCi5T0m
83DaPOMkjR1b4UtneIfVO5uC5CI7/TTN3TYh06AjEh7H11/GQvwSnlEGr4FUih5f
4IezwRzElJoUNOvxGrINMwsDkbiwtg25aboqDhOb1yg9dmr69jLUpPdFUa8wWDTr
AGLUW4IGTGJ2G0VGvPbQppeApc4YNFaYh7nzlET8lg6ABHgikhk3cz7dew95+1rD
StP3AsuOVXX+ii8n5AjT4mIc19lgt8IwFMEf27kE9D5sA6vJTVU3yu+z+PIb84jO
bZKwMcXPZLHbwg/p7caPeCWq8xiDS2qtu3nMg12wS43TIYP/UEMsRtP5xObZhvBq
+xJNBnL8S5gSUnrrH9foDTXzrKTSewk8nYhLc4cz5wGgOebuiArJOr3O77QMGEcs
XxR1d49X2j0/vARPhPagMxq5ikGiNU7yJAYMzLgkC56XSpJSs0Lpjy/Xp0MPIeoC
X1pBYWmKkoaV5Fm0Ppfu6EU1j9GdXQUmPT1Kjdvnpb7yADYZzbZWI3F8yp6YC3FB
1lsUMHFN5+y3tHKRusor9E9FhpN58uhQ3DRyfFWBuGtjy+YwXeMysU+4vaTdpEqD
8JAStRYEYI3zh/LeZJSyYQjesPUHO8H2ebqgxsISyWJq6/5CfuRTwLoCObh9Q2Gx
kFrYS81Z8YaXBSVtAYERms1RjjDQCCmnWy3n9cs6kAzvH8Gv+cqABOf9sIAFCS3b
3r5QocaIk08FSAGIiswUsxtWe2USCvXT2nT+0yh66dXNksKhqKFBej7GfPwUi5J7
7zVlmT+fUNI4jNCJyDyOoihHaznbNrizfKXM2RE4qgrY7ikO7uHapg0kVqf2hkJI
d+73TJtj8odw/h0F8H75cTJo0xC/YTiKVCO76xgZobEUafLc2rpYJqD30QEHtTEL
ZGAOnsyTaxhvTX4eKa0KvcaOETmDsycfwUpA4iIF+rr1Gfg3l82BZHNWH+mnF+eH
kahokerx5WqHVMb/jtG1ujpE7AVV1BSPqSO0HBqOlKzhyIvzKtWH+Bcqr1p+7ri6
Np/rUSs2znHtSigN2gFzNIMCNTXHluTL5X5LgzaazWbNQeZupkGPa/hBv9QR1cJF
SOZerEeNdUGwYmcWDZBFDSLQuA/eHgou40ekBcZxkPhaM+OM9ec0AElVokx5keVr
sC/GiPdSvCTpMHHO57vukLiYeCMhpvR3Xdc9UYTabTn9difMX88hPp0wTuVGWVmG
TiJUf46VwbfBvn2IwURXbp3kfo/lR5bjumF/SWhK7Ino+QxgVZh5u4nnYPWgkWv7
L3pPgYDC6FTGskcPdt4sD56SNTvOaA401ceZIyHW3+aXxoVQYZQhQRt5+Xj/K3+M
442W6+/YiSgdqMX4Z3fHYsj0BYnXuuDuDK3jj9Koogh/VFxRzQDOn/rg/4Nvw2mP
wQZiMXES40U+7fKUsDb/nl36Eitx+eRPIs0EH02Ngq7qNtPeEGBywLOL6XM4XnYw
oV6L+LR34vv8b6abi3HNmrR/9NhmvO4q9Aklvggcuuc2Z8YjkcP8aaoNBSkHoWsB
xMNWzifdL+Hx4xHrD1INH2x0H514kM6EUFgc+Rs+jbk/4mySD44W/f7fXAITZUhx
HkU5eF+jLC0XfDaWnhgfcxPgfyQDt7M5W9B82+5fBINq8IlyYvYACvtvBnFRBYdN
xhBjVGB+T8axIBRkYvu2A3ngTb0u7q9PUOSzW48NlpDnGxQJdrXma0NdYX8r0RXr
9YIf51AVKqSRrt0I7d5FgLswnSDbaTV+QH3A49Gsq5SwmdvYi21H9TNKMOc5px5Z
WOewSINARu6fBvlisaqk0SQKw5kdqzdjyjiFhENY4CbDlYksnMTQYpTtfDkz2I2e
jgrcD/J7rv8AMiNFC47TEbIbTiJOC1OD7mF8+LJwsqEQRmDOOfbjoUWErlj8HVF9
rirXSRk5eesW3yUUFwLDg2PgLWcWQ88Z8IvMqeiN3YwICtArFcE2HONKRU3GN0L7
Mv9H8Og6MGcFnzGbvuGbuE2i++etVpHPcOirrLTdWDjazb2p/9cRBozqmxQsQ3ZT
OeS0NjGulHLXzUTq491RZrVY1iXJ8jKS2LgfIoMpzTvfSRHW0VplZh3AXQ7Vr24a
+WFxdWq4bGElaiDZC2AYF3EShmfFHU4MmiATiszd7C+jeLJ1B+jqt+z0ASrD7i5l
GeBz+sw5dCUMwi20Or7uyMxHHElf/XpnMYl9WMXxY03uw7IuhAeYPLxA74vVV4tH
ExTTFuaaZxIGIzDEXyiCWvMDgj75hHbBDPIL1w1e/LFb2cNwrBNjQ4265fDeAc+K
Ks6MD/GL5ah+zgNsnqTb2F3lO+bA8StgGescTtL9H0CSYyvKHnQWmKgPBUo0UpGJ
usj0yTZG0LwkJDzaIV4jEZ61TWb5YlNdzPf6TlHV6Q11yGTXOMOc5MCY8vcIySED
Vdaw9f3UkUmV6Us7g3sKZ0GiQ29jZlF4ekb8v//iBcya2uhM8JRZEwX2pDNO6oNE
q5KNAAu1nOulkbBl9Sin3ItZnjGir544j5k7wEkTSxVbv401v6m/ggPx/WT75s74
AZEw3/lx/G3BwAke2Zf4kQG0DM82ABGjmJ/tvpPw51KYtdoaixl1TZMrBp9bjtEY
GKK9E6wHDSTpMR8X/lWjvSHqzAy93EGnkKLAATM8Cw49m0l5cwG959K5cCZ/rSPR
XQ0NHGvOwUcH3VW9To3CZiA7k+k8lsIqJ7Ts3wIkeIIpcYD892ozDlhZfVJ/Qy9e
81m6oWbX5CwipkaNDMUH2WXChfV3BKhDEy+u2rlQDLtHaEZMHgpWr8seXpP3hENy
HeO0nfQt6vEVSSO5hN2CaZt5k1t35lTNIC05Zhpvg03HTA7xwxekbEkPI0I6Y6bY
EVcaHaxJMzSITgVWraNXbHD8ReOBLBhbs6EiE7TtdOvjOsTe0N5umVpTVyAx/m5j
/hZSGH6pa7udA9yKGMBUSMd3O/O3/n2CE0AUEHE3U9k4cjRqiurAfhMakZkJPF/U
s6OGJf/NPk0e3wu05/VZnfhd3ynN9JluLGm679dVRW6trM9wta8eH4cmZkiQUqeN
I9Fw3BuHh1PZSAR1G+BkrarLx2aKi9w5Bg58odXrXqKbziZsWmEC/7P8Gfe/fRmG
GPUi66hbV+7pUtoZKw9OTL2pZLX/Q6Aor36SMgfGRewgMwRFPB2XTyMBARc5Wcul
thGKwAkai///4h2SWn9ICGV316RCEYfHoMBT6eLkQRgUhGJAHAMyveZ4GO0qK8dW
J72ziepv7h6Ms2KCCDKPtnoB94uGRXotoUNwb2v4hO9N/iVU0bf2YWydnSvOGM4K
VrfkYj7EcsWjqD2W1Ewi2mwLfWnPPXwKYNlfb7LASXg3dV4LhSaSbB8QvwptxbIw
nFiukSyN3G/bQGo61mNt4tXtnAdneA792UWFbz/ZKIYAxos0gcnk8JvPYH1Iiq49
la4kJshIVzheBS13s2LbuvK+/es5TiuHwrSbtk8YRa9LfogZU9HGkv59vp2fnNtN
/f7XSeikrYrDdyxgJbZjtEFBGFE0naZBUhLK/Kzfw0dgWGqg4vXTAdz66wMV9f65
rDRkSiOIOgM3H4loaxm9UEvrZIjF6SYq6S4fbLzXPhUdJutxmBvOYDS54LQjW872
+VKZh1Zwcr8IaxN9uFeK5MAu7aeTiqkFlkkmqZGt0sH7nmajof+ypTy1a7sONjd4
zJdJm0aGDMXIe4OjVFDfTLdyc/apldPXcR8IpCR7pS9epxQQeAifH/QikGB7Fb8e
MLB2VT+7myAEtAE3numUwBKhpTztbsNeQDshcts9TiOKjwjoo+bO+HKeBuW1If/t
vpIH/hTMphldmi3oDO2O+Vzm9p1U3YagYldxeGFjfLExA1mWUMY7YetTgviuB9H3
tLCaHAGm5I9EyEWVmHvwsicrlUDr7EHBcftixu6YPs4xD4QuHDX/j6JYcAi/6jd7
37RaGVVip0Ao01rzLpYFbadRic5+u3tPI7rlp/BrUucibJQ7O/UNuRyf5Eh/0+Zw
zzgh2avEnbNNyX5nfGjqo9ad4eqSUcxn39wlFG42TWYPKMOgHpkRUwLkJANl47UI
ppr/xkWhuq90ULKSxFiKY82wJF/T+i1PdPqZrctlwGMNqWMg/J/wpETeS4hCYRmw
LN+chNJj7FclcZWdiUOlxsDuXpQz4dklc3fqzOQK+T+7zRIYgzs31ORAWOsxxJO+
Pu3c5wwYPWWKWdvBUHNMscOtrNqONsGtLI0sjZYQZIgvcs4Ry6J6UNN3mT/6lJaa
gr/l9kXz7j1e+xPL/d4yJAYOCte31evaJiWskyChfHxj56E1amDyBHvkULMdtK2T
ijgwLwtHolEanpl624jiuHBGbDr4ZUhhccS7v+E75yU0idxmsqCRh0NWXtry14yu
2BOfB7xYkSEPt5rtxWNfKuBIsNRnaGJsLpW8KcAoB9qYrABdXftvBA3H9i/+gtv+
Op1c1XrK2NMXhwbXbWH5uJae49GFWt5LQO9I3oK1n/xjgvexVuthr6yv1tX0AIOn
AOTenXXbXdcpCbXIZTx9MfhoHALISiPl3Ua7XTxS7WC0OgX696OBh4SHm3QqDms+
6szywIDJnFtsSb7Q6c7QIEsugjsB4vJuWVpWQxNs14Z4P4H6gDciT4oPuqoqL5JN
PVTYu6h27Cg0dY4Lbc0e40xCgGOObSaRpKrwWaoDfcHE05NFKU+NqYN5kV2/2zG3
xoba9cfUyx3Svk+wtqQ73SeX4owTSg5D3RUsWDCBpl2pZ9VqgrZoIa41YpWJKEQN
VtxNqTt+/c7a2b+04gu1HaBL0jubIWNOPKBbJDtV9IJihtcbFBtm05WyxYHQbiDQ
phfzNbkhEjmIyHJiEIgLOgx2cPn984H5UWCgNkXoiAAp2Brluu7HOja6+sUnH9vB
ZDePlPf//EkFsmRBvRxCwUFJzjeJe9Ghpai2FVty5soWfdYis1bXu8rcvRA8RGQs
X/hWps80m7rWY14V1OkTbuucJo1swNvZHhKCCt2OXN6DlsGZoEDuQFrHGyczaDNT
0D5bU0Lt10NrGjR585vVBeoOgjxDpO4Qr1MOiRqp6721NEBVuajLjSpjibCDrO2P
eqlQ/YAnUAoggTx0tvtI/lndRNgkkQkop+5rEUhZYxsnpqm7CfyieNa7jTgR0yjy
7QaafuPeF+fKMmAb7aYS1a8Q3UyF1Q3phqVd/Y54NCB4bRc+nAIwGyKANU8MbtNt
rw6YJHs0IJowNZeYlUp5bA0ibzeYEzgflwgtjdt+ZwhKuzRhuTh2dQOpURPHK1fB
UIcUDHuAD2B40M4Sfg6jikll6mdLtWpsHcvU0ygu9svGGmSaNQLD0ZhpDUkHGz8j
Omhf9WT16YbSg6VX9siO9d3J64pkX9wSrd6LRdLFfNCSFK+BGvswvRZOjBqAN7eG
IZSyufLrA2eHKrXTFElnqffkcazYa9dg5hzlgCOV3su9PbecHg4EoozPKiRmG7v6
1+9PCeTBsehYyRu/uTw5W1N/fXehTrVjryTRPr/bPVCWkZ8Q0ORtLIYrKBJdZKRZ
kOQhTgWAvnn88xUXjRn0IfsXCpPxNgF7DesEm5UqizPvZicXvpWQJvT0m0y9queW
3mJxVa/3a8NwA103ijOheeXwG0Gmn7+pvoIwWYxft63h/Ph+ACxL3LqUWOwq0kwb
lG66K7+wU+NdJxDwbCRQgUYw4UDRQSHKEsukaeVQ6ielli+ysDjzj7Q+fQ98g9tX
EeSgH/AHFhgPInAcr9/87ObF+D6ev8kXsFOFLWR7clDqhl7K0hDtAB5ZfSNlrHw/
UfLVUrduto6ZSK4iR+bY1MWDXW6dl5ATFMxDsW8hoxJlVe4iunmBNvBhHVmFAaHN
FUX8R4RcGczhJ3K9itgbd3yz5f5yf6Ko9udOYq0+W13z92glcL6SyTP1ww+V6FHr
PtnPe3MNDKx1aPhg/xo77+GaMhvPNNzVDjN04IkscoU+knhYezWvmvFUtCn4X1SF
ru7i4leo+zJYz9OEIooYuvgnS7mfdCWD6eCMsSrJjK6Vnfg4k9PvqcZ7F77vN55l
Hq3/N/lccVDgwFi8s7Oww23jZAakRb0pMVI0sUkrxI4OrUO5Ea/ktjn0HRLkgAOs
uTTdMIMIuo64nYTB513WAc1qiOoJdZSnGDGoaAK9xBlKa4ZP8EbzzSPmKe1BPj3P
WeEWIijJMXUL8q9FWQRNrzWFPWI4HArUj0F+IHtjNMrMtwfCx8iK30Fq4P0JveWr
4zmjNhaovV+PCx5WKSqezM9wMHK+IfIypkuF6nt/vKQKEAG7pPofg/satn+IW999
SzIW4Jn+fivTQ2SF4TFZ5aJYzCxESI4BOMH9gwz8Owx+dNXK3diSNpOlMzwQ0CmO
RmdqP/r7AvHNmBASiGKZDXynaGy1xZngYfgIRIP81Hjf7fjtEyS/mjdz7TBIBjH8
K9HSFL4nGZhXmi/VnVX7fc8QV5K6kNuGVuJOR/vWq6wxUGzttcn9PWKx8oQU1vW/
KhBz9cxYFQUvMCERmtyAOLgf17tlKc4QtRzaBbxsVbPK/HZJ4WPzeE2Lnzbe0eDm
R8zZFzyHjXuFMNWa4maD0mBZm1ivKqNyYKOOx3zn/3UzBJF2ndjrJ8Rz3mgMePz1
VtdrERJW1f5LFQifTJRsSuOIrfCIP4S/MNn4TsWbO+IA3KPO0fbWEBgKL2C73jAl
aaV47wIwWYh7FFDNf5sbRID/TZB76VUxKVSloERIq6IVuTWRRvB0231xjKcv1S+L
b0QTabF/T7J9X+qvgrieSX4AlQ+f5WLELtckQTBWqV4GobaBjuLwANlqDij5BCKj
lHfzOgPJLCWc5JWAI316MMLXwP2U0vj4vgTHXUP4d/CARH9eH9evRqXfYZ8MRJyD
W07cq+I0cNufqc84t3RpyTC82X7DQyhZrC5ro6LtPzG/wX91CFTBffg4zkco+xtF
aQQDNoIb1qlzGZUFZLWxWxNk+AmXAhB8axKAVULb0u57lf5CTLe8pVUyco3oLXId
PFUxasoJ3DlJnA+Gpd0/9lPe7ML+WdDN+bW6CYuvwBAZ3dy61PgqU1ph4eFjprU1
i+GQBv5AFh0zvVGT0MbGei0d3UuNqe+8uo0aNj8QiLYIk73lXqof+F0O6d/Nq6Lj
V0br/SRXspYjR6y0NjW/BJU0oAudzAW9MUzPV4PB2+oavV7FTHjP0D7+oVik0XG4
LpLGwY7Id3Y5JimW/ZdbYUIKfy3A1/XWylZtxzh+ATxJw5/gUqLR0lKih6J6p6yQ
mmKKOua9BAZhGJfGDVS6oC0XyW8eRgWxlRRQm1jT3U8qVxoATV2Yxx+f+U1xGjDi
kkUWyn/3H05M0Zs9V2LSX2RsFMWgvXDmXLCOCQx1OAAFIqjuX6T4VnjcR/3mqg48
R/CzylR4DzflzJFaK/KkQpZFvrIBsyhDDu2L5v77ZNqw4KY+6vteGjRO3iQcLJFy
IS0NexeK2ZT1Po9nB4hejdof4JF5E0Gj7N2Fcb3HruJPpSGQf6RIscjmsrtIOxKU
UonlZiw5hqSAqf3YAdbSqDOY6TJRcxZGGG9Schgy+Key7qO9fnGiMvPT+rIwgG8U
Bon9UWCpBVinGPnNS3mHjEmUdUIslhdagLvu+vrKGN33ooG2GDtHL69qQSsoOgop
hQdMR5VGujdfVjupecKWcVPdK0ERUy+aSvmCbIggpsP4vSDJ0U4ls4y0lldtl7wE
/T5xe1NdGEKwDnVwOw9zWbSrCJpqZXwtBeSY0HyMqMhkN7ZgVvcT3+VLrUtsGisP
yaRXwDKg0whyeqPowd9LAJEMovIIFza3gdapEk3veB1gg1+x+oFog3/rpE0S9cJX
ALpwLY5F67V3DQqbKtJyFnlrcNqQ8404feFIuovu1dKX0bYCX9p3y3RDtuFH6AtG
S0Zqcjm4NU40pwwDtjKd6rfvEyUrTKhaxc5xPgFteVQosoDmm8eymMz3gYy2u/lv
yg5KPcZAXBVAhgtM2wyv2sMuH0K+Gl4H+aXeIqW+VW/0GnYt1GE9LoMRD2xBxKDL
vc4FmJJ9Hh7ip6XfUXu5w4ZssqOyoY7/w2Fe+ZHI68zkeWjBC4Ihf8dlefdCHqxj
hB0ab4FLdfqKcAi1YUFa9BAWwfwP3MS7W8CRyvPmYVjhYv+EcTTjBLPgu2UYPHFN
VD3xuqdpD8tN72rUNj7heMrCFwTRwXLRsse+oV5IndQR1vp9hzIdx5uLOhNdPqOo
ATFiC6AFzmmttDRwBv5uRXpYYQUGcTNWUyVEk7zRAdFNwFKkgFnG6iDJZUwt3sPj
5OmQQDtEo9J2DrXAortCCGOuQKUXpBmTVPfrmEhiT6+uRozQkHvy/eaEZ5E89Z5N
1aoahQk+1Jz97TnY0J2OH7VqyZWCLg/yZDXM00PB/JsTukZEzPu1NLOT9kr4tjwC
kqrUR3KmxHyagwUvNAKGABgw/RMU8qJwQjmpHb5pg0kDqHs70j23M7BEtNa1Z6f7
efwsvnRkuqJXJ7s0Wr9IMqiltlLP3pbO6fWrWVShucNcRkeRWWVoItlXiUg4LLVA
Kf/ugT48lucyP0c0MEmtQNSmiWW8uI7X9F+dg1TFcQocv/Ip9g6Z9qBIqTDIXchk
+thJ1aT6IpGYzTTq0izoNLo67pITh4fzR8Xx9Pk+6VgRCywfu1fsD4Ho2NShsmfW
9F80onThmh2pnSGZEAN70gi1v2SB+P99vqbIxDBD405Yu75Bg+y0WnAelvq6wcUN
3IhV/cMNxKJ/MMnPu3pop9jQaGLCRt4ewmrD9TG9s/VyzkvRIGOQVo7/yh7NffeA
v5E0LuoERjMsXGPbt6wxofxjuAmAI1yOCjBpl6Gq/VTpzimbqdeYAldD4BxSNnbD
UoD3DLwk8xfK+lvZbKIpfD9MiFnMa2IaY2WirahTqfUI3XEvt0M5PCOwPXYsqsBB
eWJ5S5ow6WhKWKtMYxK1Z+ek8PkahegS0M2fFkw5gyx52eAosAo+e4kkjIKfDotL
rbi0jS12DJTu8i5izz4aAd0EISPsKWGABBVwwWcQVLih5xhP7XW1c8C4BIYwGuYv
nueElXJIRL043KE5L00DE5pKtrNJs9paG/vI1cde4L2zedtff3wwXHzs889zWSID
MWBIqBXBNQqSje3a0Py1owY09AYOSgIaePJT+BmKvn2UHXqD9rLthUnZbQSE5CSi
oYa356k59PwgS9Piyit7LyKd/w6WgyUOIhjbUD9wfb1E1p55HB0cpqoJzuoQ6p8Q
BaEvK76y8vsXTSyfNkwYaeNaRn3sTCM/n1BuhnaCjVFUANKkBOD4DelOax3BNU9P
Ux6jQXiaxWVhBIc29KDqqmOGdKsAdxEvWV67jUb9Q8k2kr7dAEgq7dtcAHyJcJGM
23yQ/klSz2aA0/eQYgH1Ao82h8qICSFoReQgDTB9nZphaKxRVPHFbN3Ou44qvCMu
Lg00hOj+rAvqYvkk0yG2io0t+/6/oo1ffzZkyDEFQuInSvOh4aJy+zdkIxQ/kq4K
upD3KB156xfgQX+Eh1/oVJPLpA9f3DGq55LeYhDAIX1rlZVBO/fIBhMmmPsj0fuO
TMTNlWXfandbEQCnbklqPGz0oKdTAEM2FtLrU2w134TOFibyYh0Su3D63ypPGVVF
EdxstCy+9/S3Y7aH7GfdNathE3sAZPv5CkNVGjTSINydAuAilNimiyx0o+ZZUasn
5OL/Juy6/SBxB3LXx6X3GlNPnuYefi+ZgawXWcez3rRvHuAQ/7FrhIT/9+qgsyzr
zuqHIA30nZuikLiJPxSJzxwnjwPUiMlug7ViFtH1MggjC+LwYAvnEEFmQc+3v1bg
unevl6Y7+mFalFjeuh0P96fF4deci6HWzQIxULCqKtX85DMB/I16mulhlxg9efzk
HOnhm+iJpe40WO23GPLkl6cOtPbl5W2UUOq2/rDmW50GiHshK0Ud4BiC8DJhZUEM
uUqoBD4nTyssTiZHf6fEwljAKK1ZP/Ujzp00T3manDJvEknXJnPi/at52xPYfmMR
T+S8iViCtBNqXr7Mn4OLs5I9mX2DBJELt7qF3sAz8yBgwq9aOg+1yRRdsuspYljO
yvaHmSmUu5juL+4JQlXcjlC7YcQsJBqI5Ej0Sy2VN8JO+4pArhohBhjZd/QwIUE3
mZO+NWFxDz6pYvTmRtLPb9B/+1ScH6EwAYosI/ez04A7nmVhdUKCkaLIPOysqVKy
fDR1EPqdlM9S58G7a6wSeqXFyfUbD6pWWff4qMYFH1bBZCA330EUJZiscOlKdba+
Tb0go0cHy9qJxEOujaqv+JWU9v4drPI7uaMnQlVYBAqCsrFy0LeYlHMs+QI3+olo
kO0S/J4u/NP0y5XrwfYvGmQYeW4Yp1O1bdPhmKiAOg2AgRBt/6rsj0c4gWnBPChu
dg36ay7XPnuBo9N9FqYt4tkAZgqUbXqoWL9KAz3L6GX0bawrei1dAHtGWJaehbj3
G7rebbQfqGv0DvYb8lDi8mhH/Xmsx7hg/1FH4pUAts3SmYSAFhUMRkhtPENmzcEA
4CioFly0ZemOsy+HFAv0iSJLVioM/zg4pErsh72ayKEtYYeAjoscSitzcY3433HQ
cX5HsYewXUhE8biO2EwUzNtQ397bZPDEUOWGH46uBd1WznC0ZWZLjy4gpzpU3bxY
gwykcLzs5VZ4Me89kBO4UQUBqK0dCrDaYZ6+vc3tdDOWmV+q07qXOgd4rQyIJF+P
OESl3g0kScJguaaOQ2PFx85K5NLrjtUgG8D336eBjEupGoBf1Oh8gSAZ7jcAwq5b
6Q5AZXBn9lxd5LNms6FF1BkVbmLvNZpN7Q2mcrBghspRgzZ4W0XIBgLmWwYlGdyc
4nlzznDEaPt9j2tFyqORRFkJu/6/TitXyL5PgoLNLTRqAtthbvSFdkYNz8PBb2f7
6DYEIU+KOP8QuHlm2aynANe1SEW//NKHEn0kaNOQBrDvxkVQfH95XVtG9SKCP+PY
GPmX0IEY9aK8aJAv/iYN//c3ZIi83FIuQx9oHMgMbVGH+UBDmuOnje0AIX4JwUoC
yJTw9W7Q8oKdT8UbFvNsi5Hr91wIgM9EuhEzYQYaAwOuAJxw1HT0UCH+51+gtyCL
gtGsxv2tXxdqAhSuYtUsaHsB/zQTghnEzgiNlEwxTQZU2aLcPnGApKPLnKHNLGnl
2cvC5iR32n3I2w3VHt5cIFyoziwRLYvnAWYv6wsEP0fDJ2Bfs7UmKdCAC4VzbIG5
8WEb7dGXwO8VIguoWfhsdBI0Veg0Ii6REm787PaLspsxsPIqOGwMLKkjTl6Ek47H
A9ap+XYPCdK8pkgPeYD6fFawdp1AJ2srtiKWpIJMlSLQlRx98ljm/Qyydmtt6lia
1DTti3h+5FF4AgYxZnPK55na8ejb2a1Cuv6vPYv3YW5d19kVVQXIcwQ14m17xC/b
cWs34oMIrTjesElM/YE/B6lqW3azrlkl7FC7Ksci9AnA3h3s321O4P6heT6M4FiD
sFTGD+vSPeat5YeAGH8/QJbLKWHlFuTnLxd1nZH5Iuq+5cCTcyv5OEQRt2buoEJO
cUnHu0VicJdM2iSQsPX9mSUy5LLWCOL+A4XO4ZhMJkDrwGKSSjoUk919Ry+rMubH
GL1ExolFhsA+emb0QB14mDCyzdrhxK6X4VbB9/1H8m8VmPUfALYBb1b4pz+Oo3rE
N5YCys33pNBPyNojI4M1jEIcI17b0OusdJ+bKbIB59VqNH+FABfv3t65ZRKP5GY/
7Z0zPY2KXJJCX9XqFFyfNCspeGcqn/4V9+FDQ6ZzlURnUIMGOIkih5g9EUFMIoPq
XcavdVPi4IJ7uno76K14Vf7E2gosvTJ8K/CRC0FP7QZ2eJ55dLwC2xqJRHJzeCjW
y1U5XvCfoYJYF0iEm/PaPCB0clHTG2PQh5STmu3tjWUWd/3K+e/zxYHMUehRTIIt
CxV1GA+20IlumvO2VceNunPuZJ9/n9nC4O86TXjE4wyHmN/1Dsa+nFGyjX1fcMAO
lKdw49jBEQV8L620wcS5UB1BWtYK/sOuIyaSBjHBqDFtDAmhKJSjtul3YUnQy63s
wzMc5aznNF7YNEKqQkr/a0YZW/odBEpmTQP+hnUJ7c3LvEqaGm7+IXk8meAW/RsI
l3+71Onit3Q4k/OtElP3laFxggJZu7+S1TUTVgYjGUj8BoCKb+/QrBBD9nzmsghg
cY+lN9+8t+YtDKnUGz3cTXHl/x4rmCcbGNtejcZc98L6ewh3LOX1zBLun+wYgOkv
M1lgOcfLk1SGd/ZNJ1b15dSCqKbz7dBACBc9B2AwoDv/Mt1mHqdDOIaoUNcYNhmG
wyENyPlo0KplG4knSn4Llw5f66NGEEOclF6zaSSgQYo1GVUo/fhV5DP9YNCtkSRc
9/ZnB/Dp0PBV6MIkNiutDqfWFKzc6I1sC7G8yTQOiIisat7pJv1Gh2jM8d5+hglw
gsLok0eOUzHoSKtI+rcs9+so4j2O6654cp4ZBeVtr/Na86P8jjeZj3YZWJjxb7xC
NxwA1/okaTFGPqVLI/8yd12AKmdFvB0pcPVN3z8pwu0I4oyzlCJ8S0PVXd49LxtD
FhIM/9/surS984BXfpH9NOXEPlDzOH4JkYz+x6AOzJShJ+CPYxLZzoNsezmo1ROy
pl2rQvvCe8ozv6zySj/oT9znwvIr4GFqEbUW8xKdTq3c0MwPZm5NwsLPDB5UfcCy
T+QdhQc9/rSG+QjWLlV2mYe8QT3o0anVUHDi8HT9H+DDPTilhPUeVYddsVCkahRW
CAHFVp4YSxhM4kF4G8BViRmGh6bZF4Vl5A0HD1UBE0ei7ZvMp3HuM67i136nbeLO
dZusvLxQ+N7llivhBdRM96cR3fZR1eeOwT3w6nqEVADuGQnFyzQ9GJsC4Sg1Y+nd
uNf1p0asNd9Kf+LXAjCYg3kchVojxzbbh/6IdoCcqbkfvWZDWkG4L52RwnJEwa+5
IG6oHgBy8HP+yUmyK0GQZ2XFkbqdQmw5gvcj4aCchhOsjGBkQokaqa1QQxctqcZ5
5z7LWWBPBxHZHWx1YfMkbG29GBqgWxj3q+esjLdTtUJ71BKAbtPJY8NCfllPRIeI
eQi6J4360ijkSibEwt/3HM/YK2pVtIwny29Ime1YrI91nprPdIskgoeN+W2aKFRC
hbInzF9iNFD8HZgH7Itiw8JM7c/Jv3K/riq6fmC7NX0BrYHsAGHp4AIQhoSA0jxC
Rscba86qDZo6dKG+Wkrt/IEmf1qKxadtUrT4vnFqod8vckx4ZxshcqSj+ISD4NEm
KNDCfDb5j/jNjJmAiEIwr17YD5RFI8PJERpsDA4jb5ZA/n1Avb3XWqraP71sRwoK
A7XhEeZoJTPK+5qj971QHT4uT/uCnkSfxqrwVhLK9g0ntc14eibzd9Y+4SSPrtI5
6N3DzgfH6M9jL2Y5icuGAzJrvvoDYFEowM6F+LnZPTmn9F9yrKANO1fllttBJllC
kD8e8gsXK6qWhR53w4d75EZhLUTM3pnnlyi5iHTstwb0I/l+gnLq0OKVoVt2AvJO
oadh2lkH277mKnMZZl6BX/yR8FbuYO5fkSROzLFxTpVlZOh6MLX0bNfaqx9qXDHD
soCa8bQAmNdT0mVawq5DCLRBfdKRVgTLSWsUn7TG3xQCzSdClN5VSzH/ojtqbSuO
sz+FVj7KWj2FByYOJMCwfmGmV8Yp0WPQkEQfKFYE9SA0r24v3Z6BrWa0JjiuUlGj
TvPNCgSyRbzsdixxwgMxqQYs9BXr2Mh2CXu/GwnTMjWf0mTlGKlrsb/UC+bQJRkj
6AkGB4tAn0P4NQsVNpidsVImwpKVASZb+rd2Nl6xFzeejuPagXqNBePoI0uanPaD
1T904B3AzeKS0xrl249wDSZB4+MT3T8TYJqwUJGeLR7Lha0793Iixw7zm9cMuDo6
NYE+qQx2a/eNQwjVpL1pWnl3P8F6HodpZPOxGn48ZlLgvbWUnauujcinTQ+V8sJb
uReqMnwz9k3eBzsrJxyMwiCZIMwXUPdC+psoNWOrojmmgKSGW5xqirV/Kvxdikoh
nS7BojGMsqptNabpHokUNh+SDdRF4vb1uVc1iJAQw8d4ietPlujl8hUyrQ3aPIUD
QT6HeVTYDEJAVhvgy1DIAhx8oD/+bFUhG0pV9Yt+rS9zIiGXg9CRkIDBUNk1s/Qz
lZqIWVpJJJjzyo4x/MN7CuREytU0Iqtro6YyHASkRr6aFtne3ciTI9ZvEY0TfyXO
iPuSmWcEGicsY7oUxXW1pFZuUU9zBpLHK881SILTJ6ajfKdlIBlVIuWoxooxOisz
G3r1waX9gSMBxn10n2dTaz82GImuGYaQyaWJsxonmvBmdUeBIbuhTo7e81INjdvD
lvQMZ/UVATGacLeQz79seUAF5I/5mbrgzgJnaaj3j5ZL+IYKItL6lH51m0hfmY50
DaRX391japZk4982XBQvs6iktJiIlGEE67nKDAjXpSjnylHFM5Txo9IpOezx+2C0
Mc+sCD1QvKUCWVKC/VLKdCjKhKPOgCPgO7+yozB0KgshCqzdPxfePyL5O44z9f99
D4VHPePTEez5WuKm734WzVorZ8aKoGZoKGetC479j0sGpKvw4WXeVl4Yd4eeswie
oonfrVrvjtc7rXIEXW1cpjmMSzGrTGcujC0Cu2Sr4OfEO2NesI209J7vAzx7mE/q
hoMYt0/ZtKgIqZEI22wCYybfO7rBgkcX/3OXQ56MpIDfTJseWVei7hHODxurnEWB
rPyhKvIl5i5qRPQH40KbH2bP0hxL2ve9yUgJwy1LuccJli49C0OrRh0/D0NZWApn
IEKA8VZo3SkAMANjTHvvS2dghTteSO3dmQKgUcrl6jL/Ia0Y/GKoZzfgzTQnRh2C
kvcc9w/iwl0ORBFdJsUCrOmz8QR4KvJAXr/sRv7PpxcBvhz5nwevAb+Lr4OHf6Xa
GCk6O6lVH05pn+kIRcHs6vJidYe8vKXibuzMH+uweJxY0pevPHd9M06VDDl346hH
1rFlQyaGGr4oHNUsqzgtOB0hWRGLyEcfvc4kZFFNIQS6H1hNokoOLgUQWBM2k04f
fpa0bzM4zGAlFx6zy1KlEavgKpxz+DyxL9m5KZO9BFkiT/Fa4RTq6mEir/Lkz/qZ
dsGNeRJ8XkB7G19BfrZnK+RyMG8jgFDh4VR94I9d8U35mOB223NiuIVs9WiTHste
62eP3CyrmIpJrkr4IiFowMHOo/3tsQjBwCQOsuqOIYJN+Ee7jBzsmtIRdvjExrV3
XJ/CcG45h1QbdKCxrs4opJaCovqle0eOEbpERyGN77jYjBzhK+WjNZYbTM3cKHZf
D0SyHwpkXOWurOuSzpcs0WymgK9bADDj26b/uWQ1KLHooFxAwhoAJQmuF8IbsjbS
Ny904RA4f2i9pJWp7tcqoEceSdrGEbblSaIwIIqptoTIK3H9QQkNwVHlGrZE8G60
5zQCPwNvRwszA5A6tGkM9QCvMnCeFmxBg7orZ1PIb+WEsqYMwUcIeR0fkRGLHdGp
Ck9c+SQLt7btoyQvVj3nuaEHbfhsh8p8j5tNFiFSDaLDw9qIuMu/BB1YEB/t/hhw
j8dFFZZxGL4LzhxKBCEWMTCZgZdTHSf/jDct8pKXTqvg1ShqNN4Yb514ccDycylP
efgbKnbNMuOzg4zzklKSCvzHC1xQZo6JR5fIMUqJycQdPsTK1u+fS856xtpHxRRu
bu7hzgsscAAkfVKC4u5CdAdVKjmPc4XStrDzXHCuF6uWLkuA+KB1T2HDm8aGvfaj
XvYhxLTDm/WUIwqUUhNl3sAmcRwn5VDBiLgzK6VPyqSZ1a0VGpElW3nuaDVjs8P9
Qldicl2cHs+fzkeDd9kzbo9QSXw6vMS2s47Gd6iQbGNTqftYdFDw+hr1f+7ddc8+
MScgno8a/OM4KCGWZfETQidNogdCFVMIqgnFwcSILlo54Pqd0560gUgsVFMOcFrC
49InHFcts2aipTlIvW6KifDx3Alo2iEFhX+zJmK/E7/PyYrYyEaPTwTJlB4djc7x
KVi2YkWSJZPWeK9sizpCMINZUh/EwjMfRPc2aT80rPYKVUvI9s/mKAMF7uoWIlUF
IBN7VpMdM/ojTyVznxfjKrecrpMJYNgWax4uCBpczXTVFZFIj1hqkjOnoFMzs84H
gVnwMS4swLahX7feW/lfDMR7gjVjRr+BL9b5Ong03ueZ2NZDEdqXQWCB6PQE8Kg/
fCOtzmP1PYKbts/69rqjCHR8tiE5jTZGhQsKeB0cJ638jey9/VLB74r6WZbDHdbj
aC5x70rylZdmYCNeWaViEg3hkftNPnX1B1t2xXgkYo3qcdeIXtzP83Cr7MjWiipq
p5O9YWSQC/KuAR3mNh9IMFMLpI/LSEE7FrYMJYOplFalyrmuHTJVE277MzLfdqsQ
eoOgxx+kimaT4eSdA/hKWjgf0S6B+VOCSguAlDX6I40gVN840ZT2VgjhiSMHZQ4w
Z3fYrX9TOqcT6/KNrFQnvttxmbQ22i0SRlg6lLxE4Q1ffjY2k40VckyKC1wipL3H
qdGKRVOckRgThU3iGy6RTSsVz67qq9IpYiazDmhWULdG9NVxK6wMwsx1u4thuhv1
y7jqwDdFE0kaDvqbeqC0P2fSjVWIPKVLfFcVeAksJxquPzXLz35KHzWnoRq7CI8d
raG7zfbgu9c139rDRYyXgTpTUMMXezigEd5jO+UHg1pU2Vwal/XW/sH0vus2r8cu
MctyKa4S5VAUPhiCJUzmSgXAUkt6jD0OHlRtZIanbxQd+rw1gc7TDa3Fx5yg1woG
UALpTbRxQiDZMrfRXnhNZHFt87APXkNRUBT+rt0etj2BZrwBo8Mdur8stwRdybiw
F5Vp3RBBe/4/MbP/Dy2GTGooAWEdG0jHbVd9vTczSUyQN1HYs0lZQda1qSCvAt0i
+Nl5+V6GnNMQJQI+DP4BBCCNVBnNQeM/c9VieYRQsqQPaDBoQObunxi6Ox/Xj+hQ
EMv7DNPae1Zb3bjfVIDEUfbX2iWmSViiqFbO2ywJlHFTydvK3ZKi3QfLqsLlVtk6
gKG1vN1Hft3kpXSclalnpiXGY+vB8+zNdvQf00noVfDbHamI58ZT0qjlBW89iZv3
QhomeZpv19zi38cacoG0OTIP9NNZe5GoRWCaMLjA7QYJjYtK3SWPWubCtBCljC6I
CiUPZb+++i+E7LHiaFNUBv4pQOxMZClej5RH/Z8FTwbIFTfupiuQEGXoaD50W0Hp
AJennqreRobFnrf0QL0bgUwzRk7bX7lMhu0RV2J5QehE3AN669xxXcmZNjbQtjMN
pZKgrYckctmtVL5E0pKY8MFBBFUQCwzYbqfftmzt4clfnlHTHyyAfRSr04TaIz7Y
R0A3j1x/qVbBbRgUelI6ra6qcUSyvFIq6QynlcH4IiiYRwFA1BZMwv8cPJRKYHGI
YkC+CplF4koG9qAefLnCE0yuqdJJ3E/cpliPlRa0aqKmqY7cmjNItsoO3eBmRp0q
XXsUTJuhYPSyu9SvTE1PjXlWKUrF8R9Z7/7I3xLN70UdvpCFTH/8WbKQwQh9sKjr
PdkgjCQjTT0Ku0HzRqGU6ApOqBolAa0qT4+WbmGX5xzadewTjmTIHYfQj9kgAUMc
RL+3qtcEKCoZzhbg23JOLhAbv0LYqr4xMP+tuH01QyEwiF9NEMxJZZhYeJprCS7Y
Pm2xBwme2aOQYgrbngcmwRAXdvQFWBByIsm9USBLwDA3inMkNu0CcPiOPYvPXw2L
L5KxPwMGcBHqR8QeeSzUOiERIHHeoFpYlUnEaHVUDtoVvwnic5EbH/30Skp1pnZT
sRy1FcW11vgR/iIF7qMlMa6glBZtAy8J4+aK3gEwKs6KQbKChJEWBxjG5myrdRv4
xTHi9j1RQmnDNKs1NoqzNa2N3ksj6rcULp79kDrqV1+Wqt2wDYfH9t0RwhEI5D5I
ShuxmxPpdLd3Xh6jpICGWfvLDX2gKEZJshnOedXUzaMOErqLxEJTJ4PrS7Y2u/jE
b63SM8Rn8CvGUWDP5Q9UWLgkeNNHHi7gxJZ5dD/A7WZrNLogWdgPyklcALYstw1E
qDRSnqszenNWYg/CB8wB3DarhNfcR9TiFYCyUAK96BOTc+1B+zyq4Ohkj09i62KU
L8QfJ+0Z3X6WqMinMBGfPQ+u0WraOB1dprfxYyPqGsdj8ayL0t9v3P5Su4Gdv1zQ
UmoLTxT2pSRvKkuzSpGsAKQsYG1vHvURdiy8PwOXCVPMo5iM38BeSnTtE0HPuT65
Dnij1f2tiByjygY69moqvVQc1JJHdfYkToFHTmJFrKebCWKvxkNh3vZu+NTwjLAX
6964pSLMJZE8nyXppjfUSB9tKGXyW3K2dtUzyo8l5QVJ3/nONyYUz0HuMqf+3Ke/
dkdYDNN6RjcSeb7DKwKJCpFFPnZ4d3QiH1kamgJpRrCkvBo6+RvSrQjjUO780pLL
6hqS/JXCuu4iwQXnrwMvWFaObwRSrS+9L/RHtQycTOvdxct5Sa6yAf1Xryk2MJ15
AzoXjw/Ixk+SOM0chHRbYCpjFE/gt+jP14gX14pr8TzNqFF1U/kXPdzKySkwbn3n
aP+o4Pj9HoBYSqlHf8LRQzUGzkH/UrXikIwsuQPxY/TqzsS+BOKBlMl2juxyna3F
cvZ0hr4Kks+gb5KeaJVu9CLX/YP4z4Z8Pf3JI+NhGdjJ1J741sea9fW0wOw/86uV
uwh+lXDwfDWzW+6iHF5NXKbZUAaXaY+PnZsJe+ViaYCSK8kq3kKhGTvE2w4OWrik
9uxHrz8J21gxEUyWh3w9Ymt1hFIKJRHrVhvA/7/u23QyKwK4lMdqwC/CZ3iwfXHy
XFaQ6o+gGKvUtjnJ5f6+V/3eyTTYnSayqkjDfgexcWXSNCabgMJSJHjqATsmN1Zf
NpxAz2/CJKeAnAWgrsdq0RiwJM0f3y/0doMHvh/My12O7wEvKoDEWBJ8ThcsttHa
JGF9tpoBnJBOWtgxZZ/+BEPxA2jkjAg+ZlULX5gRXEjpUPNMgha6a0wGeeoA9yfL
PxY5c2C9gTZlgMQu/La9gASGRWII6l1z1NvKOlWJ9sYvVvWixHKiGkSG97h5BYR9
huwF0h4oOmFPhXN3qVZ2riOTl8GNQZmSXVoId0nNLuJwKYWWjkt5etF37pI47x+o
4bjYRwZwZmV5i2zZgooNiKsDKWOxiNioBkbJXaIlPGg1VXpveeMV9ikxWR1a8Zoh
DrUVBG1ryaRpTEcKdrl3eg2JBm4yx6mnPygoNt/lC+NiUojFmJP6DjFMTbnf2LVT
+RLUJ9h5CYd2XQ9fg4tbmgkhpxVjJ5/KpisL2d8oihbENbkjHCAYNWpYYe35la5e
TDO1nqFDa294SeIu68PDr8KONEnm1CdlrM6aEisaWoNi44WJpTVkQJhfEaV/Kjhu
fkkm9s75uWk4sLRDv+MM/t7Sdx8MfriikGrAUOcEvixHc32yqgDPFZFqxA05j1KH
aXsjj1ZrtQPUxjx86vO9t1CXazqVfI6D5uIqgk1lJGgUq8zx+STSr/C/nrNrcIdt
3BKUw8yz31h/bX1fXUpA8plfTq0+nZs11NVIIqPWo3thw/79dm8Xdhl76G+Rmyyu
/Y1JnsIbL8ylhUV/Oadu3itWUKhylmGWDhBxkFK2ufd7eoXESjiUVP8//EUCKb1I
5sqXJR825wuPsj1Iop+gQpNnPfFR092wqy65xeUuWx+sCzo25ZKlIwr3P/LzTXGV
CDfagAuin+uhYBJm7MsWmtqYsIIHZOB6UGMnUpJqNL04COLaWwRbNiGnAf1WBFAG
ClUgxC0wOPqz/PKOhXV70V9jduOrBeDaCO30SAqWKhGhY0m9sfWn4n73Bj4Q93R5
5Y/U3d9m7mxGB3Co0HAaqEGMc+kbpjo+HJTjwPzcV1kWPv7J4GnGwuPH70i+NCad
UN2yAHjE7tC8hAmdMWkXyRefjI9Q+7DfB5XkkyS6KPtyqezPbogTAkRlRULvv1qX
njFzycEvNU0/19FN9omduyw4SPOEHIZz3S0ZspBeW4AzmpB6I/zMFsyDNp4ECa/7
KIrU+ya34FYOW2NSqlJOTNEkLDH3IIof/ddClS/zvsB2fHg6iJODT0i80mJ+AKJQ
vzJqoYiffeyA6xP58/JWEYkzBpZGpwj9YmgvHzOA6SCwypOp2/Ctg198GLGz9r9/
9yojxqjKIMRuwoas31tjnFrVq4jRqbVLSXRBeC+jTCrqe4C9mTFj47QzcnH73YT1
zz9OGWzEqDYMXRFEe7wFXChuF1wRY7VAPf+XAF0/zm23vluxEGKezdi5kb5aplmI
EWzqxcCHbXWIHOvfsPXTbIm7CSLMFneb0pLV/vO/LA7sZMwmdUFQdSXqVz818L2M
hoEDFBD7W+L+BZAevijiYKmGqpdPyFvU0Pede99slYIxQLQ5i72E0szncSFuJ4H0
YgDFhqvKIWMvQIcQYQolFCT+PI1FCbbBlbSdZxlXPpniVMOtCOoeiQEdmrBFKkl/
i/V3M4rwhBFUujSZeHI+TJC6U2AahyTCtNePum+SO63DY0YtptWelpFbSogOCDyW
ech+QVN4ZawyU9vt31yujUMFV2HM+SuCfTTO7C1Rbrdq8Xb0dCT4p9za+dzPU0Ri
RYKJiRRHUP7EiDOQ0umFVuquTYFE8nX+I/fUa8XbhHuaqcBNQzsd0CW6MJxfgxmQ
V2StUcIrVpgFPO8UF2D0Lq8YxtLsOkcG1GIqbGdETLV8eCYA2Y9sCuMkFyAnpGzU
J30mrwAnMvIbPSx1gAmJes+cLLU+qVjsDZ/MiMctWPi4dZ/SxJ44e+3d3lzst73z
u4mNdSiMeLnKlAf3kNAghT88lmsPzh7Lka0ycgTSGwW1hxVYR0yIv3smZ9y8nxX7
aWqXQn7BkxrxJWsOXa4OxB14xp5i+YoEtoMsjYfQ0spOXmlFdAz9cufCGN8G2KXq
xhnon3nRfJ5w254R16SJMOnVSitI7bR16BV2N8G7QsckgPOaeS/iLPOkqVe7k1N6
2o6sioAdgPChePcJ0Gmf27vC4W8qHJUbOUxK3RRtIekkwtgv8Q4EJmBsaF6c3oUl
YAVOssipa5z0vn2Xcne9BHbFqvvXOyU96veUHsnw/ZhGHtbZLLpB+FhhWug/tmDJ
ndrWJhg7hx0S18tRQA+81lmUp1tYir2h11NbMwNOtlGbudZoxlFT3//2znnxlt3M
OFkM23B+vowop89EUeAWhSGygTIonKNMPiBDejxK07n8k9rr0eykqCtYr/UaLRpT
D0sSaQuio0VqR3Bdi9F3usPKhodQZVg8rzOUBgHYSD0jLmmtcWpM8Smu6zUAZxkf
JOGmRsGYpP+WhvZNJDhVGcrvc7NHytgTA/ZBVr1Su6brX5zyQbUnKx+P0SyrUKUY
cIQAPfKssIAxd5GcH4tAlLqD7z6/weTSj0NmoTz9KtvkLCAQgUjq7xTeCSE0ntDG
f4O/p/moFtmz+HYO1i3ynewjPBH8+ty8ZWxD/cjmChV+9twhNjyKRauQPUeL/KqX
O9Cl0gp2NsAfcDaSXEH6UcwbZY7VWxmqdaQdav2Ianp9/p/0kWXfPMBPlBLaIgtj
rkZr9A2bt/iznRYcgLHr4C2oM9krXRDek7Te5vGH8py1BiHfDo9BmxCEcSC9t+Us
yofPAIl8U603KzxUHSZlPWvKsC7snkpEBvSJwl9vqjI8RULkgzFNO7a1Lub//euN
iUq1h98XCcG4rBfdf1YErrujtf0jqs14Aibn7wwW9dvUbpzbUF2ReRJmHc3dyNVE
7iLn/9P5C38AJHvpEh2H+7krVdS0mO/pIfIgseJfe7QyLs+CLyM+FDP0F5yL7fWz
/7tBBCxZdAV2p8cDkC19PHRj3X56KMNO91UXeUKtqY3US35V5hE6I3wRIUXhKmrd
BolU+2ClBfQpW0ncUq16Ihn6C3OjGLzIbppuncmVFqzvEkBq+u51pZ6H82mMEfAB
2OPUbjcA9kQyR8tc/6mUanz+f1VBUUZ43BulSSEuyo3yg7LAyVH5N7HH/Fn9EKmL
l4VlHQCiNuiEpxiXBzmzrMod4rmTMzcEaj6NW9akT7q15Zpnxpmf2xZANRr7+1sm
5Pska4d8SVnu2hhLK3zaqhb7oru08oeYJcE5L3pGi1oPFg4Ecpsa1s3GFPUttpcg
unRCNbFkAb21r4N8sXsDM2FFLZiW2Mpq0UfDGw+zQwbuchCFhnWcmFeXKqUvEf5O
FeV1balghadFnNL+WeV4qnA3jk/sm0jJgT+d/GPMwf1Szjyw0J941/UpFMPaP+j4
9NCIrhsrcOaiXVvO+8D95TskDLEXTj8+4g9BK0DPoLL/GZQh1Wa4bTzSxpKTOLPb
l1RW4UA1f1ljXdFDoQ0VRpUhC6fFJXBexYsVd1VF6INteAJYbqFKzEct5J7WyA6u
XbUx8MdrjjJtwUq+SSkrZUurFU2otDC9aqCHXH/7KTW4CrUSz49wUbv9Mt3Puatb
P/SgQgFfclKHYX2KcdXq6DFDjodAOvTGUMN9sdex90vwhlBh14P6U2sJpvVuu8nk
A3PlmOJtg7Aho7bQMrn0IA5PDT2HBDxMukalDxPWFmVfw7eI2vuJC9m7l4RKB8+V
O7ZexOb6QGVrqxGxDgDtRYdaZsVabPlQ3m8HzGB4p4GhtT2RACgS9z3NwBSkhYZW
6Q30LhRAeGdQFPZM4Pyk/trvyhb05n4wlPhT8hM/Qwsuz1Pn3VRa8fuxn7Qe2PrY
FCAiodFYLdEOya0bPbL2J8H+7eiJHr72QWRDTi8MSr9RrWfHZ5SfNM46eN5LAsu2
nHHMXvd33zrq9KDX87uASKuKpvWMLneyTtMYNLcYY+AaTA4YEi8OxhkNecQSsAAM
q9ODPf+M+uvPiIjnhuU4qmqE2JeMnFkiYPrgZDP2L4vCcemSr7hhQoPZHf3/caQW
hYqF3mUIyIXYJ8z5JsRlciF9uQ9ryoDGAGzUrZf1DBdb9p/X3N6l0ug/ciXu9/CS
dIeJF3gW82k9Vx2eazjvdUoWx7aNRqq77PUX4wpOsbauJcMhGXtmJI+AgcM7l+UK
cI/isrwTZeTydGtEr4A1+yv5MlU8vdTbbNfITvGljKpl6H/JtN4a8qolIG7xkJsA
jUnSGVjh5bkkkScgZ4wFB6/W7OvYPtyQfn3nHXYrDBEcid7vpzNN8OayYP0j7SgZ
jG2NAhoAhVJr4tEps3pjDLfWrf2dheY+6jzmCs7dXWk6D0MmjxClo/7dbTmtQbuf
6gSCPxBXJr6Zod5edZqgxciNxZdfQMzw+KlRMdlD9QvO7KMQek6CkQ05t0N6BmjV
Y4DG8UC2lQZXPa3k7zCjEMg/FRCzsrUzxqv9oUp8ZeVddBxTvWAsHtiDQY5aw6RY
epljXFzIqca1MUqcaSbGXxjl2DTmzXFkPebrv/pXLL1cf27MP2olDEWnWtnxBTfV
ZhmpG90s3knpDGq+TzzvigoWgbLVZn8l3mjq3G8p4JXwTpYP3RuBPtqXfKj36KPe
+oXq5ErUVtbG5JK22wcRFG2EisgW3C9jpeFAzSgQf7vQ6OYXRxABVO3hFNItXIRw
tOUptfqDq2WGgG8NCQMttFDynvTf9uhkkXibwJ7wNSxuxjy1Mu3uCzMiBTtW5IDV
tey7hEyCncIfLl5rWpAN0NwxTqycvPudUnUf0AHKJdbNmLI/aHrfXjYQCwcZ1xrv
nrWh2I4T4RuxP4C+hWCNPlTxky+D0LqzzYFsF9rFEyEW7AV6fCpyHXSpI/GtKqM4
lVccaBnp0T4VWZKRkAokUuXiKrhXC+Kd2w4XmdrDQTsjX9wC6CsdIyj8H4TnoaBY
Rw8UpnyK8VSOKxA8d6NUBkhPFXbcgFWBWvr+6Ur1p0dQlnwa1Vb9dxtkUGAXq5bv
Wfxfdsul6BYT4zMOiaN7tBjfB2MR7m0FSr5vvq/tU6lG3PqvaxOMS+h7aPDUmX0v
Up0VzMZvOGlEPApqzQGZsAZSBHH8j6yzqsNv3WHS7m4PczYJu1e2SSVv84IITNPc
GEKn+g9AMSu3VuMRv3VF+CTesddqJ+UjyBeryZ+eiDWHFnngZt2P0F2S4sv3CElc
uVSicXK2spEh7vhtxF7Iux7P1vUA21C3vrSJZusgEd3Z/L84+7WxaRDAQ/pa9z5B
rJbxiCLGxwLy46fmAzHw5KoCiig9aWUuU81luhNHuKAdOSar1t6SsAStg/TP4ChP
HqJMKdYfFrVFXPW6+Zg6kc041DC626ODvE7xIpdrdh9n6Yfkg3siUijKb+qN58In
8yiLq7sl5hEzN6tmmITSKoPGMmEbAaNIBkOKJwAu6cJ8j8TtDrykY06whaaQp4cY
N+PUofjzJzijEEUqlOqBGogWB3OiQrEWa32IeBzGXBvUUTrprzCEMHHu+gFo8XFY
HI7GQWxhBb0v9RIcaQwpS89K3M/M5Kml6nWBC1lAuBBHPQQnyGL+YLa3Z3WNOGdn
wG+6whWqNpjayn4Jxrt6vaPOqcm9YK5wu9ZUmD6l8Ib2JrUkPXLdyD1zByZqICl8
3H1a+aWr1cdXbdxl3+OVh4DcfD6jogydd+hzGbzrwju4c4VfPuY2+yTX4p5nQS6L
FDlfcEdyUsSQLjX8Ocypurdsu94zPpHoz8kVXt/ukr938IZOdvIgDw+YLO0PuYAs
lSjNlDRQ+XNvjhs5weLp9IPw/9hIzds0KNpNFCQPabJZl8o0Ky7RYDH10C+hB4rn
9vWFOceaN9+SB1f8Sk3g6BNkvDB1GlBalwKyfyI1IEl4uCM3WbidCqKd6yKeNlye
wJv1f+LcjofZfxb0INv1HorhhjhKgCYsq+9YAz0v4QLIGnCOcPd7KwpXbjbH3BOg
v3yaSKvRAuyHu8fu7jBxZCYkZy+TwYpD48SX8Y/xJRo0kF0Fs7NxUvrSeK0hWkPi
uNitW3LbNgymB9XVRC6mpy+gmWop7T8ws9Tud7rvuTSU99a1g6zSKAgWqXtNbaCd
IfWW3cPTwFd88L8GtLN6vZOv33jthZU49RSuJMzQeclgeX8VfikYzc2t0Gud517K
NZQNrZ1sfEXDcgE6gRgR7E5nByLxp7Ng7AN1IDFmGwGwIEZPM68iIuNuB77iJVhw
kdUfDKHH3nCYlHysAgOCaUPzC0M24jyclZUfu4jWzSLEnnV6DsBLFrXIR2BuW9uH
G0tzxTNOh8Et5IDAhSiJsYgtNRkfF4N3PPtsiaG2X9d5vGfGI9WiGJmtFVf2tZWf
sAaa7LO/hFgElXp8SEk1AxW8BT+ycryp0sE91H+gjk3wUY8815p75PcEug0jZ3mg
/2wqQN91WrNfgxYhxnZxUE8dGNKYVNWRWiqfidEP6NZeyOy5jGt0jk+SpNSX9d3s
wgxh1tj1ptfCnS52T/cTz5nPfKtUoWmoJXtMjtWeElqaugEP6FrYrT7u6Ll+F3tT
gDzynvFoNoq25Nfiyddk2jDuRhMwh73rPHkMdZPP4lpLSvLbMxW7VH3yedJBLsc2
zIi+O9laVjZKn4SQ3AD6WLlU6LK5M/rqj8HRS1eJNOxvs4rdSn2esvtCJLOoELGp
ccTQIubXeYHvmrorF5SS5CGusMT2A5xdCSvvUUiUzdSe6zd1odOewB4BI8eH1NLl
KroUTcMJBpSB9Vf2A227+8JaWvsoeqPvGDEHYOTkKTiULKUjWVJN0mmbRKmpVfCf
YYwC9B2Kw0Yfv69SZI+3pjJa9sOc61/gglcAk0tJov7NDb0uHgcrAa0hqOfdeg0w
jRKd7Q8WGX4kQgOIydNbKHTrH4HE+3bySW4Ny+S3UPam5KLsr0ZrnNDnN/e68OEH
Q2aWpjkatYb/d1xq1WKPyG5h4GU4Dxj3RO1cUXAEghbsFmgVmAOyyF3spXkGVwOB
g7jILHEEvJmcPOilZQSUZDIzm1hd63HtCDgoJVA1xveUoNySiuABpVKg+1ikToJF
/JBkYz6Q9K0gu4NMpjFwihcLpLczas1taZOcJ9f5j8yvDYIXuHgJbtjQx+s2BUtE
0X40Bt7Jb0YBMmHjhZFF9r4D7n1r4qoJI/gwuUSDlH2Jx5ZCIWrI4mEculMOkUKr
qj9FnMRQ6HgdAnScVFRMbAWkghm9G9/VjqHdlxfRHaLwVWp2N2XwDXf26x53jEh5
X7WDU6aOorsjq8PFpV2Rl/Xwji/260wnSFlvw5TwMS10E8/kz0ehmH033N6O39C8
t1lJjuoH9it8roHz+XWfAT493/2L/6rMqMM6CbPVR55vT1w6aGw5HPE3uqO8NjqP
hwEwYKGUiF05jHCLlxgY0G+UdMjsadM+GgTE2l/hyiemV9qsU0aTv5bkjKDTmbz7
Vhk1paU0P9PsFwNJ3BD8rFj11l+J5oxbqrLLLICSHjxoiXLVBXd4nSypFWxQIViP
ewU25kDzVX8n8FeP9LLaixmfYaXFJCzfWWDmpXCWNfWpm5FGUeEVa2EnwxpPn2Pi
Cn8/hz9QilM3e+yVZEPU51DT5zRxc001EaPMA9y+IJAYIXX8R1cm6HSnNHv392eo
kqQ7Bha2Py6aXqKTpCUichWMuCdTn0k5Ht5Qe+hsVpab2yHNwAVDpAQOOmFxoujk
8UmfUTJRi6J+0Fb4lsDVzdRkdgTDKWgivAsUGE08Z9QNVPGFA1JyOif9665PKYXj
r9Zybw7vDnGH8lJOcuFX2T+aLFUEn99M7mVUDHhXO9VbMhsI5Ek0H1zUfuqt23Ku
U0JCttyC9CsBVSPYxkeQbcgI59TEIsVnM1+4xofyAdjndX8eJTguz52i5LFFcU1x
UIM/7OfnYiPV/BTSvFLHw50VIpWN1OwVP6M0waU/9dhN5/Pcav/A+/DuezK8Aik2
JPA3xEK9b5ihfbv+v1kb0D2376xvY0yJ2lAEcYfSjNOEmBwQGqE5ZevtZVDJADRX
epiq7dhhjgK7bHxRAm4l6mobRyqUEh/mpBeBamVaGwtpLwvMTGpcTDPSIhL0qb5c
t7zJHW8VdOXTmoicZmMgUyjBtFgRAiMZAVMNX48JS9IDKgybypYZxbU28lZJZbxO
t4FhpwOQ0v/VCZUvDGBrOEzFa7B7zEXjR67Yn6WvM1n0jggNrJbPnL7ZdVfU/Lsc
mDidZ8x3GC4rcrOchn0m1FA3QEugXgitC/zipZI9LB9gF1r9P+HtlqR+oXXAJ7v7
LIaJBdxqDSETZlqRt4aBlWap3s5TEBC1dgIL8yhScLJOHITwTtEBRELPUEUEFq5O
capcMcw3rUaSbiYukr3gkbG31yoKmbrZrz1/72aNCFtQuSOsW3N/daT5lXrSlVaU
zClQuEOCObfRpeANSes++GKVja5KMc9hweEFfsrhoTUxXw5NGWd2HXUEw1ei6uKr
YtEmrEJ6ns4yYUJyKgQIl58go8dwD4W+tnxJa65YSPseuccD4RShT8etp34koGf1
LgcbFmjXrkxEHSZU2ZE9XcerOSAlvY79NJfQ80feRN1Ys8pB7ycZXtaI+CkSVjdi
xQFb1SjWDeHbPU/QeHikrDx5h/5yqISQrb1EdXWOCZHtHwtSn7ssFxfOQUU9fkd2
YvmXumtxrDx4xENHUPsMHq7m2oM8iDFRyvUx/IsIdmmf/fGO+Ml7d2WicTKL5B7h
Uw/0HZTsyyb8prdSkjSJCcGqhb3StVuH6yQgM1njgJLlYoAZkS8xHmM3uIBQbSc+
xId8bylvfBGs/OPDMTY9U/EgLPds5TqOfKdHf1/GZV7dRLaTxWzGX1rtx2ROfK6/
CivIHB5QSeMfm/Sp77Z63QqRAGMjkPoa3g+FUfOBjasv+qvbipnq17+5Fgn9nmkz
I0I0djfW6VnA1wi1LogneXkEA9KUuCok0XGgbXxv+JLjlDeZf8ID7Erp5A/aEm26
I/VhOojJDHhF1GWdOH3O7rsVk4RsTLvEtZty9z8bI6hy/2IHg9Th73ZFM2ydPHHA
0EUS49FUieqmZkJW9peqhsLlMCECscSiimllBIJVrzBao2mBPL0jLDqJqkobfRYF
Hgz7Hx+biwHcdIIyCFffaMO3McMIOBuVZXlKF68Wg+BWWmKX4aard73PJERivNW7
wd+jlS1X/7d8I44bF3mgq8Cx3rv5AN5PCv2pKn5viMsqPvjs0xpNi5+Inkv9Yug/
8HzeCDJcDNgvFrD2WQIPIabJACwimuGpaYg0qcSfFhVz2sQlVa2Xy+9UFpttCfxc
7IMIDYOuRcY6iV4Ter2/MnauRE6bpyGdJIHuvPoI8/a/WsNTUFZLuQ5FnW/w3Pey
LiORXWBpNgEg28zJCafm6DD/1jRzZ/9jv0PKsBKfNJsUMGNrcEj6hUcSB6IympCt
w+XQFOR6DYEKhc6mU4MEiXoripd5GVINKZALW7FOFpqQxctwmaJKWDHrXPLPqLWI
Mcr2lp9TfULfbHyfB/PIgIebFyLEfaE/5QqdOWq6IYjGFg5gqIwEFoYGRYxc0Ij3
EiJGIgiZEgrQtVNVYlwMDDY6OYCEH20167FHFRTcPMNHT8XlpaWSEEhggGo2ngU7
gXXm3G1Ah6jOIp79AUXHxRQcewUn7e+CSh1nEinJ8huIReO26eZUfug+ziKr6Q6s
lJqbi6nfvKP666lkTaO/uA6ldStXah1GSeTDrSTuOY2d7yKR15u0c7woHAYfTExt
ybnscmtjNlQK/+xkNHyD685sbbXj6gu/Ib3RU8UrrA/Vtpqv15E2J7/3ZkPlQ+FO
G1pwGhUDloZY4w0xX4pkcaCOvBSdsiApIdnabnj/OTGP8L5tf6ZCmaLYb41NrLo4
JSHB0jQxPAnX2SRXDUx1+GyQ7BI32wXdXCvki6FP2ntqc55GtJdfi2kXOnXBu87S
KROLbFOFlarEYTNwP6DJBBa/wyLHZXbomo6ybtkqV7LmeXuHU89/fK3OIpEUwPkz
w70p3gvVCsNhbrUEX8LhaEqa4B1+GzGXY2IIBkkBgSTxMWJ8/DhfTrOBRiO+sUmq
pp7PYA6yUNeTQv08cmAE/D2IEXgbj7bkBQqQBZgEt2pF9ToDwKug1P05PZ4H0OB8
ZD3gecvH3yT4u/My+eNOyOFkeynlrs23b/gj76F9pBCFEVB5f/I97OpfrfADDKKT
a4epbnqxyEUExJtgtcdn3hSzkF1sRK/TDT95XCnMkbKTk4LT0ktvS4fg/Lcgx3dO
NBnx7UAwm9Lz4fL2BrI55p5kCMt7u8kGL3mFxA5JnIFrRNZlIofs1FkKtR07qWIV
K1QVUODyNbU5w2NaxMQWq7KyyhynagSjoPIEXSfVhdV35cf2APQGpElWeCHzU0sX
DIAbWGhEnL/oNg1O15VInsDLaS/ebagQzW8ce27SB/swd0wR+SWZcsbxqt8GCAy/
2m6HHKorVFO+3tWS7IcgcGVhYa1Qnp/aEZZQLrfmwMfl+Nn72QthC8GUkjgb+xFB
3li/kz5lOugeTtLTaqWpfZ5GvpwuIKHAE4vqDy5PQg9MEC2ax4G1JL3vJi2plL43
BHC1IU0Ch+B01tVTp6qiwrrb0Pdds+CRzGN4eDcgk1VfBvfrFXli0RCWcqWf9eU3
Cw+1q/GRCYtos/kXCrTCgTjskfnqJGGI18cHWqXnLfUWwffCSwhu0aZYQ9tKWes5
G1XXfEYKwFqcwfG9MpQnZTGBwRbp9WRNQ0QhmzrhCx8CjSCAd07AnMkyNWJsAX0n
/mvbvAWjGWDQU89xNmrmnjBX3+GboYyXrCrl9UqoCCfHe4uJV9Ge2RYd9NQf8mTt
zkcfoZWU+T4nD7nILYvAmJnLBX6tjVNh13+y+X1VdXNR2GaeCBHQRxtdkwLfAvmD
f2WjDuk7eCKMul0Pf0WaCCe+Z0pSKukolFxfJFGrZRAWLemA4uXDXCaD3zQSCMCk
CkR5/IUkITojVen1pFPDG+Git5RP5462iQdQsn08+w2F83DE2DRAvO0WwE9exNRy
2FpDEYKicP2vRATJB6BWR6EtCe2RrD7+EZ6tnsxK5n/JSy4MiBqoQSGghlgWkIix
nSH5moblLbj1ZiF7ZONxi/CdSzBsWodDY9IHM5q78v7SVyX2+R+p57qsRiogq6G/
UnivU+6HF8k63khKFvaO38CyhelphPGE9ZU33tE0W1rAFXGdH3rx8CRsVPUXvWmK
cUx0vprwxZI9aOIATfLj6K/jihhS3UdXunTKO80rDI2gzASiVd3hzpLZA3MokeDG
69VVUP9qBEYCECy8kNUb7plugnPQwbSLtSXaNOZlah5rCUHp/k2nUAxayyxZ6Cg3
SHMiFPYyJigNP+ORdDgq2353NLSeDKXGptcn+aXi07zTp/IqYNEfndwaXpRcAV9h
w7LxmODcvrdCA4/inCDjEqdkmAhgZ7PHlcwWYdWqo73xoNJLrPRwDk4MNnZStHVd
9ebMm/YBbl/nxV/xNtmp+4pOSExVR8GZL75ePUFy494nMZI+W3M4M1glWIBbUHxE
c/+phKUDbeQrVUAsehPaY5A36pyeCtgQkXujhoVw5OnOonxfc3u82HwmbE2nJG0Z
qilMyNDo2ouVksPR5GVvcMQ4nBws2c63fNouDQ6c0CvASwyqgVjLknZJmMo2z09z
l4yN8k4Yhiqwvf3Y1Es4ic3g6fAkUbFMIMtJweYB3Gm90xYpqLUP1zEMdUWTVfdB
PxL0CYp8eVZT1OQGCsBmDVvtG3Wc0fo5WpsiWMraSOez8X9iQwKVjQ0nqtBRrgBE
8eWUaCpZU/pi1NSoJ7ZLm/DUDsWxioHjMaz6jVK2dUy+BU4IPw2AWVbybJEDGXDF
RFXBtYX18t/KYgkuunzQzphQyddoNgxDlKoMtUub/PentqqUX9/jZWIFxDZMObhT
g/c6IwlFfFdjTWomf8Cm395tjyUJBF/sMzl4EISfBZ4wAMWEJ3sx70JS1nvvwBua
qkO7z2xXgTXiMMIoS7iizTecYe4uvWfbYGPTYRLPLR5ee4tneSgbo1R8y8+/evw/
8U2f7MX/pLR6isMykricEIwO5U8RlGgxjSLXfv4Og8YN/c1qHuYQjvLEKHFZ5S9d
gQwoniA1Zyq3tX+QbKHuaJyVLFhCdbRUTOa7YK8nWlXV7FJZ2KGSn5k7yVmyTdNe
JaxCZ4qd0Z9itQBj1lhDZ/VB5u0ybxuVpV3N8If9Pzou/WaXCJrMbc2SG8KWd5g9
lLSJc6v0ddSLe2IA4asc+aoQdK9UuFjOSFZM6sVaGagzWk/Ue3zcNWXfhN0hIg0a
GRDMR5H8NIme0Wu0tD3v1bsL/8gKS28HvDB4H+iw80OeO5Lbr/WRsHvwHqcsg/RQ
sM6JjLSMxC6p1UuEKekSUUiZK7b9yzTbyuyumC3uqSlSXQvHEYYKaAG+ldXTa6Ky
AJDn6OMs1Hxv4YtwAhcX0Z2jIKyr/mQfWA3ns1bIwC55Z92eCmGkry9jRiR7i96B
Jt5G9h4Q0jV3jwBJX5bPbUG6mwmk6HBCWJnLD36goRuf7AvykqWMuW6pCIvFPM73
hEaatVT9FfPs5xT3zWkDsmx+4i7OZnOmlMJa9xr7ebSSR9mz/fIP/wsDgC7wM6A2
AtIdWcDNhz6sld63LZ+G2yRJ8p/6Pxr86FEsk8Eu128OtwlKgT53woOCQ9DNz39S
mismYG26Ph8VTp7JuUeDYtUb+Ck3fKiJc0dgE6vHzjCLwyly2zVsWz/q+xEER6C3
jmkspenYGDVnvCwJd4g6nfTz1JpIMrzxTL6AjJJfCsjAnkqSeCK9g7Uu3QfhPqGb
97hQcrLXOAccPoW/ZXHkUsgiEk0go3Lca47P9Lbomh4kGf+KdFf9b/D7foETnJaD
AoWV7fVW3XKhNI5baSGn+pVipfX7DHrnlpQvklXdwx8Dh2u/KHZZ1ISde5hdhcDx
Jp1V4zPPukfzmrEEifx/auWaTWfUmIW4J/6yxUoCJAA/3Zdjy06lgZ6PW+VNNKEe
UnzqkmIr5aDNlJ6Fsd5zMdAebfFAZgGizX+KgB0zPcykzEkVXek2ATBIsqiTyUBL
Q/lVGGUajzDnLyDMAdaOagQrYTMAKtoDyN7tyRR1DnDGYtp35gej3u99mKDTPniK
HlYl6LjnOauYQrQblPIptGnaCGvZrspThx6stxYLm4OJsrvdZxw6anATPtBM//Tr
6FQCl2uxKTBLRQDQ7uBlWI0MNqi1rsj7tYLniDHocL2UQGbTi6pjQmrdUqXSte/a
W9xtwJ2ITicT9ZhLP2uTyYDtuy3ft3HkVQyRPNtVtxGHikRmKhT3V2yuBSqU7W+F
E4M8yQWX+Z/5Gk2fM2+yxOzjM2ziX/92HnfAh20sfcW+2byakWlbd57M1HdGMjMC
cRj3KxXJ/QzVnaDx41XkTPbFShtEPxVCLmVU7mWRD2V8X+IjYeNTgafKa5f0L2Pq
C0s9EwWHWuZvkyaDfpxAWu1f8NyHfretxUroOik0NMnpwj6U1JNpnbgar3qjxybf
3WqW539aG5OsF/0CxGs5AGP7jb5/hm2eeZZMVaHX7e9wRW+nWPWE8YTLjDf15qD0
oEkEwHM1RBL6w0rhjw2uNQ5FanPfv+DYKWY/ryt2A7hkJBg/0bJvuonIgIU1WgWh
09sYehRbu4L1cxJukzL/jNzZXreLE4R2XRISpHMPzuMu4D+j8PlXIp6eSNiAjP1V
zuBZyQ3ma0GCIDsaq1VcxARQgQ9JJ4GUz1KRWmnMFwEmNarQyy+r31uxEN6d7m4M
YEwxS+fWs2vhD433qKvX9B1HWSGN+25uNyrrhHNRqNMdMvP9vSf/iC9Zsnh3GuWI
YjVj24h6e7LheGgNIem+mYj7uPLgVpLh+1LoNdmSsDJJVUAQTFcG/AJrPPdbuUpg
VQgNwUE5ezf2Y4iMU9rDTb6fT4PJH9lzxh3aMzYS+19zul2DzXpA6VlQ7m0weXS1
VIe3JREHWjWfq6HAVQJZVJe5IHdhhMdNq68HSgc8O8sNfaiXfMugbYKPy8DKWzLA
5Pt19qP89YL0XVuqQ9BWz2G371DIpv9kiLqU04U4bOQKRqTDjTErKpe6vnP7+ouf
C1R9Rc7nWO9mh+EwNV20KP0j9UH5KsLA3NaCTYlLK+nM20gFzcfLV35M2WaAQmqq
rcqJ6H8Ut+E9zkcJkaMEl31yVY56x1ZE7sdbNVegMhWt/GLs2BsjV4w7cwyCzr0d
XZiGvpihl2j7Z3OTwJHtdTTkrOd6+zK10t9Fd7m3wddTFH194LS0UqyLeOuOnk+D
5kTWC4DMug7cViinaK74HjaaaFRmIqEZLHKgbUXI/XHWcubA/T6WWKtclFOgpScH
BfAE/R8B9++DoWVtfJrJ8o7MDt+/j4E8dNSAYZYlZAdj22wtSsdqnYerEPREgVyh
rIV6SOP+3/WCRJ/efktu1aoqpINulZRA/mU6knzm3yVT+hW46/A73d30YvqUnG5s
KTzK4Dxgv/Akbex2yiivmfBq4TOcy/aixVlvr9yPVsxwxIBhDio2k9/7F+o4xbJq
0kQx/6a6M67P3bZvGHFjs9FfOzLEk4LOY6xHhZI33OZkvnO6szHFlU02Z0/6KXfb
pjOIaFxa1fFhlXOmScClMzLewF/+bJlqpJ9yOfrgprMLsxYV6zEz4/AkLOgkodo/
hED9kY/3/LLRamjvEmIUBbI/N/OJk/fN7GHgtneCeDLBwCao7AIi+8/8IcQqHOjP
glp1efYTxSHVUMgvi8cRufShQSHtDB1ghaCsr+77Hl55u9vhAIzr2v7Hgosvj3fY
W0vldMkZ70mM3/01q3FrXs5xzFZK8CBUUZlY4W/nF3EutDFHFSJTMEix8mZPef8U
D7U4DwvJeVw6yD7GyjoMHD0rccrFQHApRHlX/BLevme3R4JfRSs9qFX7/XqMZDB+
3NWw3Wtcb5PrKxx+goHsvdqrkZsblaXP4wRJrL4byrKNLOmXbuuoXJ7RI/zHu6o7
252hebgljc7NYkc+cEJoRsbE9UYe+j4l7cOvB0QrMBFogfsWGkLOGFepBaQpWv1L
MP3Bk786k32hXCXv1WlyTLXIxqmGbtXD0Pcjk++YjvnZjLvdlvuNu/nLDW/cCNYc
XwdaYwIMLXiMDfBNzZbH2tb3MU2FVkQkjwBOLbZHQiUGrn+NdyEH3MQEdR0HjSXr
RYgtx+8XttHMnCY8QBfo2KXzhBVoaT6+fZ5qS4GZqHPZEgSRcsF1PjKzDzBQ1xc5
bFyUHpYA52zTiST4hpSrlgMXIC9EHF7mE//7TLQ3bn9+pEEfA5KWCfJpfqbKtYV3
iMOs9jrXvhZ4/Q+UYgnBBRrnaYD7YpfZE8ou3FCGLDhg6+gcDIZabzRbhLKQmusB
sGLvctcOFQtp25oDgMQhE16uTTGyehEcwK1aWgUbRmESKTeu1MTxsg97GoJnrrlj
YzIRlVAeWSvxWJ+NPPfx4IEeK23DE5INyFzLQvUH643P6ErcTirdCCfKhj0QUtRj
5U01AzFD00Rrmx+1IHO9wg5vQFKNJxeb96qaX+m2sb6a/432RQ8xWD+8kJzlZfEu
AGBkNsm1LfOPSKhNsZjpXoFlHbnNdBXqWi8OhWA4Q9F8YArFRifs8cfdbLbnnoSn
/iV2bec5Ses0sOAmap8R46663JamNMSn7EZ4q1OuKgK37OD1r5zWZcEBpYkav2WZ
eVwc2jIgc3h8zG841Nvng2ApYyrMBuA4LKLK4ANTgMel+Rf34CWYBOPn9S1kdFu6
OjxN2x+wVceKOERjZUI2+5Gwfesy6dEcZW+Go32jgNE1xQiIuE9fevYX4s5kjJYO
qWUj/9tiHtKN7zyVDtAVe+lCY8tnefu23Yaml/4AWvNiEL08uWwHciaJrv1E5UBD
VWWJDVZX5wf2CuHT4pZWYj2RtklubCfoy8Hnkx6x5SDxheoMFu0yLbz9V8mL4ahf
mzjNUqDFcJYBnWiP3a2Oqi8guWZdzk+XanW/VFK144rOIrc9Z137WvhNyrQqlEP+
ADJ5Ez0X0dYWPavG3nS4tAIhqXQ8UwJN0oR+txl1mAE5qnhHheg+tynmPIpk2opK
NVV6PkfEo2SFCzR3C4XESrg6BElmh13UZ2F+vu/5B/meCMLobMMf1izAw3kqDbNZ
eHygBmxEQxGCDINq1EvTjVL9KyWeSD0oFqF/fP2olGgffNlxPJ+dP2OHUVime/pH
HpI+1wmojgPrZPVbQB6B7svhArVehM9h75CcyrwBESWt6feAw/QVkP2juDN/NvgJ
AD5GIEXnc64C/SnB+7iy15rebU00cBomllxYiXsRfPb0vkIg0lpitrgVBBDcG6ng
mDMu+hvNNbe7DF+UHZFPN5B09ZmO+QriwKTFFUvGFCoQtYdZxcosaurlRIdn3zgJ
//kfTVqOB6JHVT9WfZgqsYRATVmM4ZWLe6N/BeNVGKpb6U0A+3Iaf4H03J/y03Rx
Vv/9oG8uL8YFh3crrVszTmJFk/DkkPjYcQv9S7c2cxz7nBVHNLXVgx5RHutsyOya
TwaTYUSZu0ZPFkEe/7GkS1jZzaqX3PdtY+xWjeW3g4eulNX1DWZyk4iRwF2K9Ei4
TrmAd9ab0QSlVxIijxJ/wwI5IgJYh2WI+IFa/uwNUBspRHROtGZYgUh7MQ/ioV0T
cD9MjcEDkWjf9phMj+K4jmPgJ42DZbOwpIb7X4rauyoPOamA+oRehU25oeiI3GuG
kFFVbIha51J6LFj8290ckzR4Aucq1SDOgnOrfXhi/jfEZgXHjDYNipFUUYicB3BY
fXvjmf9eB9W8YPi94eNgFJJnqoxXj+7fa/AC4rh0FGImJBGuctKaLzVeT4n7D8rr
ymGp99/lYB/na+kKnwFDOFGsj9yKQfxl6zxDoRpM5X2vvwnBWdD7VOL7ONHDjaIo
0b/m+pllI5evDKlllURvlxxbyiBg654XaTMsOOc0YlR9vnmhVfSIj0Ixv9i9H6PM
bxAwjYX7Cv1iDst9GFh5C0wcdEBm6koPzrTSHfAdXyDeO38kIq2wgTCscLqqRkve
EH0YUmtjAgUXdTgSFRuNK4HbFExl+PvOumvSJitU4cb0KNcFvlspBY27r3Rm/SIX
oj5brVH8sq/QUybvBAdCA3mVB1KovwW/+PHEikg+20BXLS1hiVKtklzdSD+xHRaS
kqHUipRRAlNWA1Op+DYP65AGRny2d6vasRi9cmFl2rONQjJzAbVFrSpOvPuW3D6F
CoXDqcN54QqdlPJBLkFXLxRh48r+TSSkLc4agJdk6Hhe3zaL3+2NTrptrul+gG/+
HMN+uM/a9uzOerAz/KTDx7bSfX2q7MMRnRvqrExUgcw/QSv07jHCHQXL+xL0JREg
/RyNsm9UwCHpTcxLWiwXLiHFw2k6VFYq5NlaetgG88AKQHFriShbJurWForyuTPN
TPe+9VLzpLcby7WrXyDIh64mHQ2GvIlNCoM98emiGBwrtq/ETRWi+RiSg9QyQP8y
At2vnDsS9n8UcicYMcZDEdtZ6ngTHizhF7hmmvIDTpFhOr81oZhpaHeZLBrict+j
Q1m76YDRLKdwXfBFQTQFIoVEY3TrcwcR1bp8YoxYAkTMJC1CeQqKXjzuYCwxlJED
PhUvW3EEZ/7hQS7tzS4KTgPZFLq8mU21gHzcFCAGpwoazRhxF/boHaRYeJkxiaPg
VmPte1m5ulNtXu2gRcV5rOQKfT0e9AauaxfY7dNLGY9hpBrmmUzBTetS/6aIP6p4
RNluo9yWdJn6VagU1H7Y10094dwYobQSHDYkjtmWBv5caUlGn5mKmecxRSzuE2vP
+2BGDLxVQCfvCEM/7GjJEBYjPqpy0sgDw9wPpcOmecY51uhEaJaCWV2SET0J4sBZ
y8BESc6xCi3ROcM1BGQG/APal5eMzK1PsNvnv5Sm3r8ZKYthFxmx9j30fskjfxnM
grlSGS8/swg+TuV3gjXGG79oj2bfcO8Wf++RYpT6t3uxRCFA5JOv7NEDNiugFjLC
Y2I2R/s/OHVTbv34eS4bGCCmSkKIxZKJB1W84ceDN7CmE9zNrhMtNJpDmhZOr9/C
+O3xjXeY70xZjEmu9wt2RaFq8bLv7rZ3KYLqBtz9UFoxCHJoZLxWTSSGJvsgBmeP
SJ2+of7BZUhsmW0w3MzBw36Tn2Ptp1HQR5yZyXCinpY6OkdkSq3+KpCMZumqS1Cg
j0/pk4+OAzeIwK656o3d3Pka7gc30xX3aiolQ7bVkIbvIfPsBwM6Ot0GPHvCFgjd
WVWuza0nMuTyMY6wgI8ngWLktgEhrnJqbjZvsGq8LqK2NwEc9q6UXZhh9kr2YdkB
gwdL2Wwmjbqq4g0BGuBmm8ABj5LqpTIf8IUfA2wD0QK3DMqVh1sEIisl66PDmcNv
uvXOn1utKiDGnKypvk0Edm2CPoB8LbIrXlkfcQQ8HhfCA/qqVaEcVSg2x9E8H8Ug
RbkTK3gfF7aXcYa859zzuv2/7c/lVsneCdTTT2hoehVf5aXYciN+RR0kqUs+BXhV
F1vyNSslojeKhUcCJ02vYdZzqyc4wjZdwh5e9B7Z+HWMeBIvXBN7BR9CeUusSotp
AvVgLVrv+8ErVbODEBvDK/E+hMKOKm5aSoAelQ47LD21wTykymkOcb43u5AhUdg+
5agobzw+a/wauX7fmJcrLN8On6vWuZFbe9cMLEAE6tNaiLCyFQftkppCiUAVUuzx
rtjX+NgnHZBGXrgCkPq2i9H/HZYMuRFbWSpliWmT64eqmQxqtkxRcK9QLcMOqkJ9
N866k5epSch13LCO/9ALgWEDJG0DyOtQuw5ePosKzNRsq6TGAOACGjIBmEuaru/K
c//oLCit2Hg9pyIcfDLUn+v63jbwvPVdIaDTIXBO8Dyv8edAjtbi3by+P9hcbDY8
Z3/LNJ+SnTkOv4xbK1Pzj7knLM34hHNLGg2x5CV4tAAW5D4jGWbcyg5eMUHwwCso
8DxCS09av+2lzDy3xDrzwiCvAxbRl1yWl+YEom0OwOmTuJfKOAUIt0hQUmX0eT6b
KkB8GOA1OEj2AarvoLm7wLXVJVpYXDH83YBUwxxx88LXH9/B7JDkChOg2b2RaRsG
aI+M9Fh+bPL7Tf+P+MMws3D3kI0mFHlNXX7WrXIZC4MaVATzRDtRWFz3GCDQMlIy
pfAG3stUnsi19hXdD6REgxe/IFvSaYTAfW9eib5/RBERC6pfDSSoSXHUmEZvRjn/
VgUWre/G+YBql7fB5v1Fr5l57v/5zQNSnN5DnyREh9ehxhpc65qJH1epxQN1it71
GmHrAJ2rdkXKenQIvtWuDBUYMUSTlbbpIyun0XNioMWA2Thtw/etkcj1BD7oaCN+
tHsDLbIujIc7eMEOs/zRT0LY3XMDEtz4YcoPbBH+7QnwsDf6CGCGrWrn2PYkad+m
RImriBvVj8lK7D+f4/7qa3msfWen6wtguN/GLjHh+gPr3bYt2rDVSCtWUUyFu2j8
Io7ZZhElhyHsp8rPkO92IQaqZlGHL25P4BErsdQW+vkzIKpE8HA35PyLHcay4qKM
nOsMIuZR7jybLxJzwurW5wtD1nMS0W1JgzjV0IkV0amV40n2xRI63admx/W2Lo66
3oZL1K60NVXrRSfhglGmscM+6Z7qLBgdsLaGSHwIKTPSjbC/MVI3PrsT1+TXok8g
ML0V2i1oRBVxoM3LwkfPTizCJEQY+MYyvA5YwvOPkbOoHIEghg3WhQ0vfQnCufd1
HBUT1jBGZOh+7Kw2O8xjH1pcLJ0iNMaB9Dqe7Wc2Y5X/8Zzo26M48mPHq3v3pOLD
V807rZob/g+/gv7l7wbuK4OAF4A6nHP4D36vGvlwZZD2HdezLc60jkuaz8hTkX1r
PnNdcNQredfpIYS03LUWgMGajKegdcTQApsNkWXGke6l/9W4yooANG7gFXZ8zJbE
FqZ25EVJacbzAx4ODYpQXGAkIqNuoRgXn1POFJ6ZqEoK5w6P3BDEPxH04gqXN379
uW1uI5y5N30sRhskkobXFxkCT2JwBgwS6QBp2vylervGiiGBjBSR9YRK3t9AGi3o
0woGSp7X1ffE01ehmJTd1HWsWuRlaLoS/D5Nlrc0rE8w/fXQJD6grQGbEf7ULw4X
QtIQpzzFwl8+vYr2As8gRaMzYQYUDs+kLebHnJ3loHJN16BGTYYe3Yca/v2VHHUM
rEyVgbqHv/a4di17+QDTsbM1wJUcvbrMnSWACkUT5jdwTf7tw3cUaoqvLT7LgCC+
Tfk4osfxNYDxp8Lf4bNdQ7g01+OhVJdQ1uWlbxqnhaHq2uqxdFdsbM5KTbrvYrSh
zesimh1t2BNW+nV5Mwikmf3aPjvNRHAHei07Eq3vBKCn+coAz2nVKb0Vaq+UXQNM
8FbUH9zraDnIfYrpeHVanrBFjB+5cj0G+8iEfpV6dbhXEwrG8wJT1NcKLDQ/KcbV
xqY7tjUj74DxveUqPFemAOTRwFplS4YURDgQipQU5kirFMcT57MvNC5OXw0gOIjl
oNRInjVL3NGEDCyWveLFQazEd0vrCyhSpF8rvoiOs5zwBKQ3eBa7P/jwX7cXP+pC
V2lwNByHloeAmwm3vr3ZKRMjFbBiKYjCsFkaNVaQOlGqxPz2El4R/nCfiVG6Fjoy
ocNoS4RK97DX1TuIIBBbyCba6TGm9sEUAqVgY8y3Jg7Wu0XcB+XfcVvh+Ffatbvn
97c/7afPMUYsy+1bf1Pjzp++ekqUITaoqBSPhLj4kuNdoxNYbGy5FlJVVnTJZbm/
MqbKMq4nSVOr/rsCZMoItShE72/0SWFchfcNcwyEd437flzrZ5svWCPprpG7tZZK
pm5/6JKKU7WgRRulwrfCCoPoFZi9ajIRLkQYwxNBlQFkjfp3sw4NALJQa33LHCkh
vGBO+OEPEWBsWxXClIpCOhJPvUu7x3e5C1BBcFVhTq1LuGUPrtiwjjECPt+au8ih
ixPXF0WfSOoFp/A7X+N9npCMP4avN5XntajJFGGg1MatL3hn9Jkwy1Qne5Lplf0S
LQW0Nu/7X+ZQQoxLhYN2ieoooZI0UgCyeyEuyiApa/wEIKjzahHeAa/o6QX/b3BK
7EfxCOPjECrnDbzCJyEuAWU5dHLlpTVU02t6MqMsg2OZi8kG+a2TjuFZ7AHwMmU8
M0W0nJjvJJpXJpzzJAxo89khxcQHfp5/Jjs7wZheg7zMB40Edcq8mFfxAPmh282Y
m24vZrVJzSn1djp9r88rBNk1S0+FZ8Y5/Ezhr8BSDBPlWYKVAki7H9RMsoR5MK9W
JilgfZO1V6iEAPjTBaV8iTcj/ybDQhbheOVjV7SzozPBU5nwlzZnz4LyIPKCV4zN
2bobVmP0/OTzegTAlFpb7fQxNzFvqONbJWR2b2aret2eWdL6ypwBOfXju1CedKYi
7T7Kg9ewSacOtiduYj3usuw1mqWhwaURRE4cT7oeQwxkMpV3A/4bN57i0JX74LDj
33MYJwAUGdvOrJkn2c7iXsdOOhzXGLrERRwkgrkcSD57RdoucGYt7rIDQpjWc96M
7rCxK0UIs5GL9U/Pfb1dADzlN65Y9YcmomsqQYISW0Sd+vpftXq4IpYTgR90PmR8
5XjtzlnvGlMbgvUMv00koOAXvwj3iqPBYD+xNYAqoti+c31uNc/QLqMwiUmUSuX+
hHBzBfOkweA18gs9agzOjOCP+0ee2kqpb8NI+YnD/cSt/rbT7WkVrUNGu2i0DAXG
VMvjKEFRIbM4A6jhFgEPQmu5YVdS2dRG6IKseMywVCB0nLEgwlOXHhhD57/yGGyx
ZXK4aPrj0egMW36Z1Mv5hljrzEWyuPE3GH6RoMDCc0a7MPp3r+gCh9DyiMwWXLRL
xABjbRrYcFyBeCn7hLMwiWCiAM/5kOFNkkwLwvFoHNomSwVA3VjcBELErR6lRYQH
qHR/etRdxo3fgElNtA7qFXah/OfA2kWBjcE3nNfo75CoUf7l+s5/W7ESsYtx/PLI
z+F8jeilTt4YOFYGY28LposlUHqYopQ85ZVsNO6g37g2nUk5/fGB50Fxd+Q5pFzx
QRtHxKSDm2jkrT8siMYrc40Rc6fE4TGxpmLipASikgV8t0x3kWL14HPqcpYWGzq4
FnuswaRaN4aMepwg593JBXDpTQVtZZEbnPzocP9of5tk/0BtaaSHNoEaX4Qqb1Ht
+Y2WBbJP/MLL74keQ9KTVo+OZpox/GPusHWGj/ro3CpledA7lU6sqVSVYHLZ4yQh
x4dAOzT7Ua+rOCHNWTe/E3oyc3y4+EyzZJw0GuKPPLEx2Hkv3XYo7Spz9YjGnpb1
0cLjrKtw4umDf3W0tP8rQUaotUzF4itfKcdxc8PD8ikxO1WJIfZ3SzFqOHLFQVod
yX3W3Eo7dRBDfefoYu0gbgPBYl9ZgobdICHRhPw0D0Ge5MB1K49n1NdRbu9vZV9S
jgkZKFHok3oC838wY+Ej5bK7oFZsDY6EcRzeAOqqFlbZMtTz5XnPj6vbeBCeOL3y
hq53i16cr+V3JXiEeTJMlEvSccTRu7T4nF6C+W9at6Wh3fPmeYaheUmwmAUtQfTg
yBzjOqUtDbQNAgXNvY+9eiKXBRmo0PZMizLv8HzDu85ZC/C0vkdzF+wiWLBOpgC3
cIkaChriyb9WN7eFwKKg9XM9FfAEQFaKr+VAB+9b948lwjdaIC+8hZleaDyOJj6F
RH+uDsJw8/oaIog0abXTnOxML/DCjMIgP7h/s0QJaL1yVH82KurGdiFqWzrecRED
U99k3/j90khMp75kvY2bI9uwkNQAV4xli+zU6P+YBxl8dFqiCvylg4j5uVSfXCn6
apBxZM0sjAQ6A21uqIkXDuKQmaD/nteBNiKF2EAeZu90cdOVMjdErHeau5A1V1b6
Fqn3kbJut8u+gAaT/5OZ4bFkWATaxvhcuUt3+iZKu2FcKBf44sLScnyJDb2rY81u
QzMz5hgTMDFSaCYVXwb9Ndw6rPfYaasUPCOf9Vhvc5KQuyfO7mHxQ53kYJkjZ4SX
+feussXWMo9EBPWiJ86L+3nTE6UOgdQvOp9cPSvBhmfmcCd2Lk8aLMJstVDxXxaq
wQUpJBGkuw88BGwDMvABbVby3aauwUvVQ53RLqET4tKA+3vyLIslboHiwtpcf+Hl
94mnuAiSbEQ2ED90YG2yx9Pa45dwagERDqE8p9O3aqyNJVffUTyB2BTRJJRCGV6p
DaraUcwYmT7LJjcRnJNkdPcgdm5KX0+myZuEjypF8KqL76Xfkm09InsFF5onK3fx
nTko5u1mnnqT484wc2Ac+NIAM9ahiFVAxeAySU/ow1nb5f+jouObwHDMUe8vqptm
ntRwYoBzZI9EmcRwh3vAG3bSZ7381ZhkbGlogK0KCIgZAi9kWDaHafy/s2IhgUXl
1acAt4qqXJRdnU02SjbUNw4zL7mZunmBgyOVzG2Tf6gvM7rSkXGI1JfL9wGr7JJH
J11RAgvO42A0GtYRDOvAOGGbJJ7jYSkYnx/dAde1uIn1z884FUsTI40wbzNQUaVa
zlNZkn88yPcxSEnFWrbGoVQbA0yWULhEvDiffZnDmnx+Sjb7xvS+ktTjizCEFEwV
OV44SpbsYliblaogoVmsVBeWP0vRNHPhGm04qv7PkWre2xYwTB/53BhWf2K42ESL
+ch7B46r+qcRkxyWxH5b1DiTysdq6C84XU5eg3xUyQqnMKlPlyN9jA+1+zH4nCL5
cspABWlcvyNkn4bs76Xgf69oWVupOnX7ilbnt+ljy9nfbtKD8XYoWlrZ762Zs3CV
8ym8tuaTeJi7PEel5xDyGReLsnUjtdRb/K/a5HbFoYAK/PsyWBQ9vLdBu06/AV2X
ZmmmEh4IDiIEMbhk8vlJjvH2dJGlJkYqPk55BHEWTcrGZng4/9mK4W7SS6jT2HTk
ut+hbZvifIY2IoEfv3C2TXa6R83Qp70GKnQ810GlHyntJgs6P+wh9vIuZ9POvJPE
fWaBwZAUtFZPTPT6ZNHK07MI9/RD+STGJnm7fp7MAn1LsqJwbVCvSsANtnToo/d1
GdlJspDp/uujCtFXnx87nP7zp/NgEBBH1IOoc3rEvLypg+PZitxitfWwKkVT5lge
4deaIj97SdFxlCZPWikdgdxiqTxQQAdA4pcOpu9bGJgeZYBFq+35CwQvAtY4qE7R
s6D/YWcJUP63lfFAKVI/EkZhjuCDn3Wl8zty/IkMx+66moF740NF9U4nGftRh+lw
oLG7uxb1/GpbWvWgoXbsyJQ0LDOpDLN6bqGFzGfzh7kobeZU/ux3OQdi8fAkRoyD
t0xpJZWvEUlX7Q6OmpiYM/CHkRt8P/f9x1w5XzyQxjonMFHmEwDE1gJQRuYrm8Xm
nzqz0dw0O/BRZZgTEfJSvNnjWIPhaPdnggJl1CLZkiy6M6yJFCp6BB/88Fq7QZjp
m6VHastYAAFIezxIU6/YaAoVxUuyTWvWQeh6UEWewqhbkilPjjMgBFQrZZfMOAA0
LFZf/T7UqM1OkSpqDSU0KDnzxZkmQ34AtIwtAhpemdibDTtZoVc0dhiG49+YwOQJ
BTJo7xNay2CySxbHTSoqbJoS4I0O4Lyyevj3Lc5vDk4rFqM8uF+m9IsheVI+cDQm
xPSrafBAc80H/jhZWanoV6XcdGRvJRhTPOzko99k8rkcX5b3lD2jQg5Zwu/AQ0c2
vg8ze6mI8tTaK2QtBKP2pdfwS4wsN+fS0/RQO3iXQiGz6Jufeb04wi05zkV3GB3O
CeolRLNNuWUS65m5eTLcwSWYbKjVPmelG7UivxaK45At+GRbuJv5MX9b2vAvISiK
vJw81fxk+scGLBexKhDeaN9wm4yvG49UmT9vMr1VV3Mtc+GJ8yRdztJWqTZdxodF
jgrr5uVnEXt7ET7cxUMCYutCrzFlGat88I0oFOb3IJWaiY8WJL9bzNM9GPEiCK0B
ZgVeXzO14yeDHnnstyWE98GXJqEwq9+o1QuN4Wv1bSafrNHtqoW3el+nDXgEMQt7
UtwJjAxot/B0LR3Ev0f0s0pHCEXIQNM/xTeICxJl2xIwDdbZtVvkr9U8vF7GgZuO
4lnoFR8j9Mnr71EHjDVyNKd7HfWU74uBO6WWuZzSHwFcz/pKiTgXVEi103G+JIN8
Qj+UOW27CJgGJ91UXCbu/AjNYBFuZVlCD/HIj7Q1ap81zHx7bvBqR2/DtGYa0KJZ
rQclksJWVUu2zNL7PxNsJoaXv0uk6s3hkNX/qxJcL7hwnvB1ZzyU0VmYDwALIVaR
s9E7EJ+fR5v+wFAm+AG/HokBlmaCfXE22KdMgsKFVZgegwAt0ON1hLRU6AZjaKAm
NS3vonz7i2DK4ftnzGozRMAKxzBEmWLn9CiQqYh+JQbocSxKhUqKN7I4tFQBMzgj
ZwdUNEVdZoZecaCX1CF2FfV7fZ6/FxJ4kdzkI8ZNIJsxW29QAjEjzRpWB8uhYcU+
NZB89rBKf8SO4yiEYCq5LRNsfOO3SJ9rmKEJRpa1fBTC0/mg3SrtUy5b1ZKbOtHw
XTojT3hGpIDwBhtYHxB6hGxaXK/7iwhzbIv8E5kKS4dQLGeYJszooCREOPv24OWq
QgBWlosfY7k5UunfeisorVKpckbOUSvx+SEND6KWP4AzV6nHZ+RqGFw1S13H85xs
mbJlNj4AT/aqNvVAHpvIM+c+KeiRhGUmRXtpSXUUri0ppYthjZoMf27SoNMW8Nvg
LJ7/anuAoRJ8YVVXq2sR3RnZ6IoYptFARfzfr9Y0utKWQGhAxaxLut1jaVSwT7io
uSZYuvs1D+lg5dRcpHqzxW7NOV+AEPyd/bciyQ5bZO4X7DOYuMb6fjLDidY7Uya+
d5vVdJDiGQarNb5qwblnI2oA8AsOoMWYE5TzAYmgqmW8zFel4RmP/OyUTHh3+fmh
rE0pfc30jP3mIc9S3VP1qVQmatsqjIWcsJVaQ2Twg8Q3Rb1ZujYM1qHkDmZWhhCs
rGAToYu00eDooPPJnZmlnxs87EbEZWEvhG1znmWS4etw1NULJMkAAMBxUL99t41k
HPG86EqbMkLI7LyTWvMRXSu9LlAghA0wPAAATlz8HA3pxdyazDqUMrSPHax/jzE3
fGlH70YUk6XKxP+KPmAT19UqMUVo6WfWuWxUdHBUx0XbmHEitD/uYTdgV7X7oe/N
YlK7SvKOAf4n0gdVD/4j3toyISZ2srN6nQZMAp2qd1iFdED1iJasnLGRjmRhuesB
qm9GaNKboHyzoXQRgLLap8dPw75gRDh2B8P8x+Jk+1VuP2IOEtWn5ZC3J/oK/L+H
Jom5qYmCEarAwYqgy0D8HShfv3tjPXuM+B9uYyYIuZdjID/C+PnioH+XrNZNPqkQ
aQh0ij08X46V4DSHV0e1Ep7XL24aV3dhED/KHrX1Tub82zOPJLVao/inHeBwRknH
DMdeLIMn9+/AI7CvMUTNZHAOsO698JoVOE8szaXidDEEW4juwQtNWcIxNrPdbbqF
dNInSWkSz/MARzf/03dYp5qnvSnQ7wBQwuhTXd2nDh5OSbVaA8Cwb4KOJtFJkdDR
Rk3P0CXKkR7z1/r6RbLEbc/OpVk/pcLEjMYM2O9MEUi9YdeC4f4J8GkWx5T9/bH0
Uej0Be4SKALJrkj1nHZfmRtv05dFryoXDk5n3bdGJSsQoeoy58hR/MzW/qqJsuiY
XMR2is3xgaEEOZ8iFKFqKWVoX1eaNPJP8C6J/3m+QwkAEkambaAO+iLFO+ESzPCQ
DmbKwkxui9rh/yUHlYuy4W1ITEscYAIvwp9++A7ci4BBV5hRsG0S1bdnSg027zht
5PR2FMGKhe6HXf5QUNJbKf6a3StWhhZx04N4YjbEIyVckh/QuGxuHR3SINhT6ORR
TLzy4pV/mjs41HovFUGxTjkjI/ar9pDIg9QhnMp7HC8dMj/gBQMtO2viDnSAcNZX
7ChKB7ZfXeG2PoqQPoWKV4vKe3VQcIJ7xGgPlCRS7orbE4KUL1Hcjvks+q20Aav5
LHauhpwmol1wrC3WavBwugbTLL0V7gxyibe9dH2Vwzeii4nbwITWPIRb1XcnEdAz
J/ZpUWqS3kn7eWhbKcYdxlvsgNS23A4PSZx5uVBf/3PMM1l1VUmLD23m+UHoyL9j
yRbnoLeiJOyEFxdF1GX5ym/xrDaQFUMjFZKlppdFJWKyRZQgjmETKImU5RBO/4Iz
/PIWBQpYnEqcdQtp3fZ4h4mj/6Xvn2OcRWyqBGKqDBlCNcKEKP4XcO82LpHTAFTD
cnOXZ88oaQwVOkA6zxgXBk/omDgU98X/YGNtbkJhLtrNlsF1qoR7p9xOUDH9scvZ
VsFrKwJNGW3fy6zUcB73BTJGpu6Q0xdlfBC55xJtQ+muZ9nQCEGU4F5stVtR68Vp
ZZgrBBQjIYYFTnujZfqM8ipiUj6pKYEXYJ/WRrNfOAM+K7E3w46wq1K19m6YowJB
QfMCr6/YtC/SXRpo37QA348nmBCoXSI8wdWa5TkEw8ATVuVFcOqDyG4d3COH8N3m
LydsG/cAd8+4EVFWODClXXfnuPVK7P9a1A7g7jfaT5tBioQQYqdt9v5h0L62evkM
KtPFSP5GohE6UOwgpjWWtGmOGZZwvB/P2rLJg8awkk1tCqSz86C0uBFUEgTEkNUQ
vy2LE2q93HUQyRAJYrnMpzRKV4PIaqL5gJUUeAL2avOHmCSIPgeGbFHphwnhDh8/
HhbpLjsHa1Qeqr1Fcyq7xz9xL+pQuFhfm15LCZm78O01dhPShBFZNOCZttlfUB0S
bjJZcozj660im5rJa4C/+03lQz3dtQgOYxTJH9c+Mffaz+Ccqu3uEmaajb4r5Wzr
uPBZuk1DkMWPGAGZVq5gM4Ulm80/kmvj8YcMqg6/YwpTcMNPTOGJaUAto4P56HNQ
ymS/3rxNJ4/EI0gcWVxb+IVCKR0tjojvPqBJ2ph7RJkuYENSUFW0OEiFnS3Rd3sz
ve1sDV6WSOxvXYphPzyaw4hXUy2+dSdCh5ZWY8sqjYTa7FRCvCRQUmHLOhqNE3P1
CgHxLzep5byN9YzoBPlYQ/f60/SDBMMFkybh6UKDGE6ADIF4UWKqwXoHh8NqSAks
y1oGV2RbvDzGZDyYOJ/rtEDNycFchmrMiJc3dYfxDKNTp7eVK8d2EzrGoKpTFQrp
uZBgwukG9pH453KpuHNITCC0hdGnSCkl4S4dogKCPRqc4cDTo3RvG8q5yv9tRtOk
UYZ1DDOfrZxVWVuJcveHZw68JtiNN0+HvPosoiuulv7XH7SPFVw1ynGAmQvYbWrD
ZOo4z3n2iaXQnMkvIStXwm9l44Q9aB8MdQARIx3GOIzXJbnncxgP/7gcAPUrObSg
RFQVkEZ+BhIRk/AYKGh0dokBAeGsIeXQ3d7ilWy1Ntp/6x+uqfkX6hABQqKKTmKo
k/aEPOU6uoUEnNQHJ8Uy950aBgr/M0OT5ZNz9bZ4exS+3VtCUEu8y9/AHiXfOlFz
WyaAUNRL7bkINviHHCKIbGHjruIjTWZ21qPLoye35aTJwUum7iZKLjy2x3J23X/9
QyFj+Yp8F4UP9mSKk5sRuJbkdfOT0yRe3qWsmsjiT01lh59/hEKMjoHH2uxpOV7L
/XePQAk5M3BwozpL3tucOLGCvr5AiQ+VjV8hnZKLhouvZmfKOOl6gl7mKHA0XWWv
2ocGOEWwtADCodNNLRhoRnxIppnKW9i/AAdudEsswMNmCdSyd5Ekl9lsCRbq2fiA
5K7ASC4H60bBBVEmfRoMkuTwXnyqTfqFrl3fXWOQzwyFncn+wJ8B4JvcAuwjzxX3
YllL3Sjy1iudgAQUQRZTJtg4hYn3WfhWEDyisnoqL6TEzX9F70QL145hft7qDIEJ
8H4E8I9nLbUcq4tJdylmgdteQPzspS/mLp8CuIDTfLSZqCGpxpixIabeJjxMzz/U
sA6CbPh84MJOJVLxckbEq/nR8r5Z3VDSzGaC38f8Mq2wNQwFJt4q2HBdgsZll/5J
YAb32BFA2vQgbSkFOrdsHdoN3kjHEAY8De75N3Ak6ZChs9OHHOYgFUm9Rx4uvm53
XE6Gbemr/htdC8jwYEehhShs+4ZNphTcWftKpu9sFDbt9Ts9WB3BSYsr6Nf9jm1F
rxxWIAs6ph7qH197Q18a35xNe1XQk+0VVUP7DLi8tFn/jS3/CHLOU8Xz/gcvaZei
cUMcSfDW8zWvP3bC/4dp5xoVVNCN7MqBkCLifgnCkJOIUeMHbAxdv+BGQWs4jJG7
oSYg23Lj9h9iZbvnYZ5hVH02MPPgy0tNVYOVtwmepZThrSpaA5OXUOF5PlaQGWYc
5IQ4jPgp8g67APlAHtX9fEONKEKQrVXdhY8wDnX6SVEMEuygpdwI8aMlR/CeSFwU
uTzAqBfXx8sionkJ5+sC66emMKoXpecS+VEz6mRaAnL5fqZOYKai8BosXweOski4
f2lBarR7D/5Sk5eAIn7iHz1kDOQi1aMNJykZrZdIWMHQ18FgXaR0GtDCM4dNI0l9
y0j52WvY2ISN27+gJ42INcotfCjpIRJbVmN4VwiNteF5NAq3tmd08bBHzYxxaNaY
znNEDsJRW7AnQFVZhCAVkcJ9LVuAOASAtftQurtWF1cZLPuOlqi42iAWPV5ycZMz
WeNSnARDerO2BueiJE5UB2LWP1fHIUdf1CpPSoq2GqtOo0v9nl4uCf06fIPmvIwj
K3PTh19sq1A0dYo108ZeM3mVTwe77hki5hlJepwFcalrhE5wLKUZEIhyFHzDZB5E
1vKSIMiEMVjyNUVu/41It9nrOqlE5b0Lo6RFjK2JvbbGnPXYluRVa26g3FThPsiI
y7sIfErMBcLN+O5eLyyVLmcfsRskP4DQrymju02pX8A84jv98tCN2IbGvQRXdN1b
Dv3c+V9oT4LJu8rd8cQ4zzkVi8TP3xRKIVNDjtoLSoLO60xNRllVGFnKr6t5kP85
wCfLZ886tKTsLizRH9ZqrcGIabCD7NcK79fqsX8drlO2Kr8LATDWaSJEuSxYp0qF
6uc7smhU9zRIGyZEDTvb9kDHs6luYKDJGEg0ZiTgZoAA5asJ4RKdKK9yv/h012/y
qjqGobcPcg+JLJ/J12xHRjJ57P/ByaIGr0KIPCWgZvVPOLmDIgiaVaDMlc74r1DH
2mglp9yTHrAXVtA94h3VdsTNHbYpy0OZrRoWU75BvJKxM2LJRVVn0Ov+vy0wWbGH
e23+c3fhySdOEiTt1htTS8d4eYKV7U4ogNe10IRl/GincYTNwADbZi6K9/o1kOj0
XWQ+aZhb4RTvH9tRqT2cV7y4ZTfXgPyTPSedGgLFXXyWo7+oez6OXFXgZ7kNaY7M
OWIDhrMbW9IyPuhbD9scUJf0685jzlYspci0n/FRQq74OKctfbO5bKbUQC2vBrwN
jvpAp7TQAqFSnNjbK1yjL0fq/bDHRhfkE2hKVQEi5O7+UK8r9a+Z/WvdNNtw7ytl
CZE/VEjTXQ2CWI43998vEletsKQpEKfhejxQto+qXybyGL/q3+TLyPDEmzvHFVdN
w7k+jDWNYivA2ddKNLurtHt6jrN1JiZakr8ZdgZBZNs/Yw/PtUttA4PpG7Z8KEAn
8QXOiyr7gOBFKZJaeDbwFHPoK7AXafB6WHMYdkXKtcMkw/WDgWbaizjTpayx9M+T
5PRs8GNV4Gm6vPJw9EO4HwWLhmIJsEKAuTSH8kdw1sdJr6li2m34cIAXljUdLFDa
uN1pQMoa+RvBwp1bQba8srBiGl7rFnxxK3NDfpcAZEZSwzbaMiT2SjGvLXFcNnug
ePvYbOZmr3KpVz2OBOryW+CUX2fxInQYHAf6cq+kiX2zykM9j6gMftsfsrMf8W39
/8Q0VQOR8qq1w+gpxkL806kT0KH+CmNDX/didKw8dT+Gxzmf4Swym/J4ajSDn/LP
Sdgj80o5/sLT1MTqMYnAVa+mmcWhqAvkozvJf1UlXDAJ00uHXxG52h9+wSOMemc8
5Fczwav7H+DbhMlyoUBa50auXGw6pX7ueKbqgA0e+MBToOC0ZbiaUiSdK38EyDnN
lVvOvPYxu5v3wt+MknmUJpqgbZ6t25uFgwR3vkZzf7WqnOUQcyzAz5QzsLHMsCgA
S9wzHKrhdBjoCX3TfQfmZL6Rq6PjXESSzRbST/KC9NtyQMjWmbdWGWctjNKVzGmM
eSL5neaVJRxpGn2QgpOW2l94eX2R6kHJLSM4JqbC3LF9r4RqZLsLhezFwt3Sq/E5
2A1Cr0D3C/NDcCWI4DgrbMpeLQTbLiyVzDE+pu0G6xoW2V2hEtXbiXvSel9N0USw
WJEeUQb36V+vW+ldI/suYKJTQefnAau/Q0KYxl1w8D6HIh5ByPuukYPVOAlZbMzH
L65tU7iwb4wNOd6bQXlQmaDKYmBWgKiayPcreIgvEKoVLcu7ET8jniKySxak6j1p
swdhsklCzMPmlFE4zgTr/9lyBMdUzO5QMVBDnjAa0moqOIUdhxfmjMA/kRxKsPWx
Vw43EiIev9Ov+Dg8WFtCBhyesOWt7CN39HT+bhBzYL5hqsT/I6DSJFxg5a+jaKi4
x0ViL4fGrttS+eB5dTxidIWZ0UB3O8dNyX1j0a6KJR/EwQ0vYRB83pIhktDfllJh
5vZqx+Pw9T7sGrJtsE7Ngj5k+zd5BIsaZnYxAZjLtOScwoHAOtCd5chMhr6zgvT2
fEbFO1oBU5HvWQAVywrYmvKosFQQD/89M+EZoqTLaYWQc57g8nbLWnZmiWZ8uG4M
oIn4P4mmkMKkA3NbZhfTlwTQcV7jykMQpr9KlSamrTEpcGMi4xMN4Km9hT3HauPU
ERMEf8cOzwAzGsso2+U5i2m61ZCzotblFVlS5sFGiFZOWd9q4JWQxHnPdNslBqva
2DG/0QZ0FCfdpku5uOy15LB33OerR0e+dZoqVlhbKksID8Mg9ZKcAXJTKILAa9Vv
4uL0FmQcSA8XjRGwE843kjkRDL0EMSD2Zvq6VYgHsOjKs2zdsCl0hZEus6ue30zZ
wCzv1OqlCHwEaa8IcFw7NU0Kg90ZPGbZo+oitG0/oCuZZCEhuHtUxET3pA7T+Yqd
B3MTGKtOLKaZ1buesXfRkLI4NzmM9Tnp6m5hMxMAQqUqtTBytwCOrhU7xq5HJfXf
PpY759SSyBPNs5d/lENHLdmDJMT5NDFqHbp7WG7B80bCWOfQoOSi6PlLzHZalMha
TdPyxpwUTGBlBJuW7ESAJO19DrrQQ//A4x2LQGIMS3urBS+J+ngoHVmnFLD+9ejM
XrZ9PtbzVoQW7iFe0NeDraDap6PBS5FdNt/skl3Y9K/SvGUuoVdz+4jxDPjr2DZg
5uxPDCba/E9oiihG5VY5170d6VMh2tM2cRROHItbIKtP3cxfCnbndoXkYWRvq+Nt
yVkChvxhKVTVNd2xIqkf/Us2ELoogEhnTqJOuwMIQIdhs16qwBSnffKlkQmF1L4T
bh6KpZGeq9S5SsaSU6cHZX8xXXPZEOkNOfpOtMC6/rQX9zjYXQeg97Xgsp16jBQj
090005ThEs7+d6DW+OCfTzTMUhlRMi3nSdJoaRrNn7AoZ0ci60C3xdKMbnfLRYuP
hgEWIlMlkAB2mZJqAEpFajk1LPa3MWqPnF1UN8rxN/HDjPxo5kHI8HyiLxFTcX9Y
9bqkbKdAdrfSQD74WpfC9x50f0rMG20R6lMnPllvZySRA540RgZRngebwA1sNLID
FRtA6qDXXwMj9HFaN1xs39EF7GzvH34AjhKw4xM2X/XnxBACUCmKnSH3rbbMwcUu
hq0yqqPpPvdb14R0l3x3tdS1mhWn4qFDWjE/qoAdpJgTZmsaWtETi7mKIoQhrPBM
AAcocv6rRdD1SmSdUThvkJFcH3+e8QZlGtQa7haHhkavhcF7EpMIS8Sh67JRZ2ng
tcXaKofqAWOj8KgHPsHnDE8ssyTfqGIHlf0x60+muKaiOcNqFLV4mdbbvwOv3tO3
imFqiMUAd3/ajLC0pKjyYfW8KuHlNGv3V5+wBV/Z1ZdQEhXWpcQQO/eRilveNuBx
D/rxXS20Es8ObocSzMuPfdWblz8913hHozHf/u7ZIfEoEELddcH/a1OzzsPEn+vj
PdcuS+QdbFmgsrsX4l+GyFAaUlioyq7gQEo7bXT7SDu3Bm9Gavb4JfJc7TemGF0r
+bipAErlnyJwyqjSZN2Wr3HT54U1AHTze3XgI5lJpdTLjaERbM0hwnP4XW3JScSn
SdiAM0w187uRZgIzRyBEJdYSKqhMTfZpDMWdWtpwrKdpRFxw+AbwrFGleiiYZt8U
N6URIOEgfMLfwsB2ebBDmuu2spakh0ZwEnfrZykTV05dFyWnz+di2YdBSlWoQR4/
mS/NaR6S36iOOdxpHoMDlOntiFUTsPg23HWvl8B1Ca+C673dH7xzh42jpz54wzfp
/Enx8lHPbq56drTMoZ+JYK4IKoYWWEULTHXbJM0Cptg//V6N5RMAp70dUYtJJTIm
whHd5z/JZrfe8Uk+lTDOzrigrDkp4ZudQvJVqoduNohoDHjArogybMdgStsfxOxy
6SJkeh7HHmse0gJQ7BU68QLeYxXY7IhrA9CUo6uX7Zby/8R82P+4dE9825DNE+Dg
t2M1u/N2IqALvUGv5RWaZ3VP8zaEx7y1pNOZII1MsMxW7TPmVOvMAoxcP9d/sptp
lVWO8dDgqsolf50w4qnHcs7yIbeiSG79zQOvQPuSYB7AedCrDWTPyz8iN0hYIGn8
B6ENZME43kabHgCMD9L/+bP4WlY4Q7rt822jIYbK9F/ZQK/5btG5ooEF+HOLUYVR
pvJ9JiR2BtYjyCTj0zWwKnvNINQz7z47NW0y47T6pjxbnVe1V3JOgF4ehpLocrCO
PqXQzRnpw2RZkfHxE0drYJwBqATDPCpwj5wnf3WyoHPK6tNWv3NsUmsawvvFhhks
Gcp631llKYEsjRaJZr3a3yLNjp0AnVBkcHWSRnXQhxMNjjDW+RUMI96j0nWd6pGN
/rKWfZgVB7+gqHr6g9n9N6+QWFQlqalD7zK5pJLiGNKWwX9/qnTD6fXgxcxpnB00
EXqQVztrMuZ2rhPFDp5Z6RVpF0BJIK5CwooKL+p0zpVH/ZqeNIreC+ypy5qtlTn3
3SFii/P4QWe4sqFVIeBhQv/lPxNTwMJRvsq5a5xm9bML3iq5CxLGcsoVNvW5/B4K
Th6zTjlI2cMnv8h8ShouVtIjSgx5QUzU/gDhWHxAM9IYLvGvUwMIKO8MMigmL6V6
xywy7QmTS1OYNI8pe4hOIZuhhfwcNfqYNSlTp/vq81YUWNga1624YYcJQbS+VvU5
ONVqyi5grP4o2Y0URI8wU2Yd3WwJ9L5qleTR4/1VFNPXDsuoYINtrE/4NXFV5RpU
dyT/fXhHiMUSWZEmiSPm2l+aQPbulhshdT9dyUYMoDEFbcCDKiEUp9Ko+QDKECow
/ZOyCtYmG9b2Rdg4hgPHSW4gEdfNn9qYLlQdICppomkcqUEoK4D142lHIWP5B61C
UK3EIIFTDlyXeKANdcJgM4cpO28mmhBDJP5/Fkueo83EmKikIgLfigf996ahMq73
rhKMCJEvO80iNpf6T5x8W2NgdWVTrAgrgZ6jEs1x8g0CpImYNXCaiQeyVmq4WdZe
gTZOqgRcKsoFlZt1NBHXnOdNLG330oBfyWNUkUlZFYVewQDNEsmi6o8AscUOfwFM
ji6Ho9LNrqrls7u24SimI/qhWjB68t8L1O0AcW266AEpiyXm9iXa2giCoteKO4gA
ZV0lZXyqJRt0RvBSDezfewyvWzwr4WzY+iCIlBzc4ajCOuqrTKpQpGpfcMcFotY8
mQF/hO2cLnQ+D7s20O6i6hib5VXHfH+ti9h/6mb0AZUopL2S0xabOCUUsTBOLMHI
8ut/5jdafPGS3C2NayWKn+S1SM7tqJ4ZMwvFRAyMk6I3KhVJAj7St/l6EoGKyVYQ
HiErgj7sYKHBOBuNNPSbQYyD1MFlXUhp+hhgFOdjTO1bqjxwTutnW7JxncrJu445
CQrpbdCIT+p4RVvQNNN8MB94js8dh6Y1qYqKEpA70adnwI31VFP3X028vtC376nA
5hATfuesXTZaRmFqoFYtq9xM6+UJs9vxf55q3hSWEE5Tbe95VulwQqkU68wL03sd
7bxrimUMfwlRpYmvHKVX3bHjgDVoRWYW//S2BkSq2+ZISy0baPjGiYWILN5oNr50
KByvewfKiUcY1J3if+lMrwR7/gbLaPeLbGdXNJYwJzvqR9dpu60KONqprvoTB/ia
jsOjMZzSNTWVUiBKsaTHQLeEmlMrlTwGf9NE03XsGkHc7L9PHJBuTgCN5WxRfuK5
2wCFb48lYtz/Syzb79/OqXDkn1d5rdZexz6nEkmirbnMQHfaFE2eTh1Lg6hcZjru
68b5rBnEJvBO9TTlMBTcL6iYEHzrszC+ZwwdIxEOTcjCgLx6/qgJAuxHhIKp3OMZ
Ez4xag/9CmYuxnFysbKnQqWsm4VKW86LWbJI89HKSfXIuOhUPOmfvS9QHToUO0Ar
HgkETiR2fgSE9Xt9/0BiToyYhtXe8nRkFOJEjHciKCRjzCnQk5Q0iOo1wAe31NJg
W/ScxWtQMJOrffBu/IsKvXCv+a/02kf3HCcCcu0O2q3bKp9m3pPFBbQ7nVmDY0rf
ZVH8igZhsBD4tG7egn3YR1pQ81P1dD5VAAD8R1DavlcjhNhF86zDo2TVJ0fuCdzW
KIXu/0wrPJ2jvBebw3R0CyBfbX3tVq6DNkz49iCawdq1XUiTihZtFe9FP3wh1LTH
arkaauej/WSryJM7GLyKKdDgUzc4vD9AhYG1YargndymFUEW2KLJB5RC8IB0pUZl
fML1nXS8GjhocC392uR0J2KH3tpBw6xfpcwUNkdpVLLAunRtX7tmUEzeNe5KVX02
GduX1fp+VCGleUiXEg+o7u5a6ZW7RQmtBKeu1S7cabAnk5ZXj7nXwjMoFCSVqRr4
6mA4JajroWI8JtQz0UXz42kPTsXLCiXLzHjcLlYXYAN9XIygVnxkOxqzlKYIpQew
QoVFW9EpjG+eIvwCRPby7fQj7XOv/lJymkmOtU8/JK+KV/j62FncdpG4wxrLe2nf
ARoKToGYobWliu5kyyBNkHppcFYqfTXrKoVg6H5ERzN1VLg5TIxA8Wl8z65uSH4U
wHsBzADNlLsg1L6ulE/10s9RThev5uuetGwLx834ixqUjdrr2hxo4G+6uwYBhara
KWQKisKrjjO9fNnEKFN3TXQh7Fjzyka/J6eqZ128oN8r/teFBb2IxFGTxW5czGy4
ojkNuJ3FaIu19zQhOFuiDZxhpFV9c9dYlgGPFl4rX4uL2kZgbM1WlM64au5zc/V2
+Jh5E9+69o7OPwbS4D9K5UwPhvweeKKi2tUZV7wjSOIhB27Oom837pCYhDRoF4rx
zZXqPy2aqm3P4d/qECaYW6Mxf8akxCtnls+qvaqQn69VjccTdkhTRIIoa54s0pad
hOUrdTs1KWq7fWjNW7InRZAXmNakW1CP+jQqMisdSNq2tLyiVh/hIMmCSz9NmCup
k/yewaJXpf56CGnOEBZAen6XoVnCVoiF7GSrE4CyNqBOMhp7b1k3eh7ATYuz/Brg
kLXO2G+bnR7URppzzJaupOB4jn0UD9x6zcgMc73j9B7mulFETy8LrDBy7BXwFApN
U9BPXBcoSymKtKkurSIg2LbwabTQhBSca20S2z3E0S7T7lJuVD3Y0yz3tjLTADa+
TqKsS/p5kgAp0lQmnQEgECum3gyLA//t2kILUuQvCjG3COfJgxQcQ0cBwBPns3sS
hdm3z3I+FyZ2rtLfIu+vmdKM658MX2R+YiKElaBZDKCoJ+ICIDfy6CclT5K6zWkn
szgyqT5+ExBbTKpMZ3Un159Qq0aAcO8SeX/MzU4+o6NC5nNbHo8ZMAcOeJD7WB+k
FVprbJ6oxf2FzlOV18BTHnSftqwdPR35wfUQ3jOeiU1m64xH5AqA8vNhA2/EtpXX
q0tyQTQPNdCa2H8H3Zf+QHfcK4lOYr3qucXuce76XfX0DDz7PrwNQbHyTY84zve1
KIdGJkD/Ag6qX7h9c838J1E9zW4CdM5wIbFi7lOhMGjUvtTzZyFlhnd0m7ZwIp1p
sKhdYqNblawTJIh4hA4uXtBIRmmliPHStgo+mtgwgM/edw0IKejO+ldrDvhsdwQM
DTXrrwA2Fb4BmDpUmvnCy8/y/Cf/tGnP52+DZl8NsY2A5CWbqkv0XVsrzGFcxcPn
t0NISCuTDd3CfJbT2YS48Cf0zg3Ot4Lbp1G/T1ohVwB3Rc8B7FCb3pta9zofeRjy
KpeJs+1RmXlzBi6zvfBo+X6RpF4sQQUTWC8MDJBNbeMh9/15QFY7B3sbz+/qBNlV
xVIXU3ZH42G5GIAeRX5oJ3MdeCUQMKA2p4bGJWKBwzgXrpxNJprMLoHNznCkXWIv
MDYmTIxUJrsI7NWtCx0Fm/LCDx4tGE6k8Dq5JrgM+9xbJ9SWQ6L43Jx6gAYclaai
d4lTDGHDx4aOFs1BjgA2XrhPuqHEaQ7/pKc7/gv8Z08tFlIYGIdSrF4eM0XFRo57
OxdoRtwt9GdxqP5nJDWKKonsIXLvFjRqgimW1+Dj7lnrzgXtD+5ANPNhqsFx9gnj
nU0CuS/zC0sPf5az224ymEyxYuTBBd8fOHFVrxRed63qf2jjo+Bda6rsEQ7e4o68
EfCUa9uz9JW3Bj9xSrzWnxpN43t8rjHtp36X6IrNkBw99bgd4K2UQKqefCpWu7No
KDES08KwJ2MhMpQD0cKY29P1yNiZkW9/TjcCFZEF7322GiFNQBeNxu2U7S16IsAM
jUAPQ1STSgnhl8wKZajQjkikzuX+JxeyNGWXxf150qb9jBtul+UutLAQ0yOAqZjt
92FW6eka4JIH/tOMYBCCCD4fbMGDpmJtQg9KVmkOijtvRxEXzQpcd39Y5dvAkx7f
LD6sPz+uZenrelFHrGQSxvt8dGaEBoLCCEo0rmYhUxNMw9Yly4Y+JVVk2ZvzeQLd
5S1kyreJQkJMGniKgvCv51R0vLZAjACaiQyBFP4RaWbtTRnvJ/BDAYP+p2VK9E/S
KLftiNa6L9ctSNMQjnzlh+WvKU7m1ngPDTUJMUg7qE7MD8qA9VmM74TFsKVpbu3c
p9ox1ies2FejvaEIPY5K4ZnAWBL7Mzlp49uCwHBSvaopx0CuT3sourfi7rG9ULP7
D7aDFkAC2WspfaF/J3ZrRmSbhvMHQy1R42AThr7jbI9dI7LBXLpDvFku1k1qpMPm
ZZmCQvBaE3WpqKbiRuL1COZhYJ4gn8B70uDntezeiZzSrRJLT0N8smaZdOX7Adeb
qR/f8b49B5l3By6Q3w2h1LrwMYSZfMR2lvKwSepkeOwTwRRxwrk38zhwQksaIgM3
WFXkxZs/O5pCJo2+lw5HwSQghADRvsH7GY+zgio7Vduyktr/HLHoqZ/LrUz7pQ5R
gowyhI+aR/VuF18m1JUDR7rK5ilnlWTUkIfK26o0dxVCvptNCRJjgoBJjM/hK8pE
RbLqxrzVCeuBnbDdFDIWJWLIbqdaEwnvIMHVsRZLDVq19x1ldGKB6yPfMFMZqt8a
UefDdVuxKt5S4gYq60G7pbe/8TJMnF9UbMGjnLNCOm60Ale6Eg7iddhd9TIjbLPM
op9QayJU3DXNOH3G+I49RWUIxytvtdWxVFsxVcZw8hwuddFJGNu7rNrdahh2dIp6
Z59yY9NAYSz+PIfdnzLanDiHUg+lunPh/g/WRfCwSuRkN0fkKXIJxvzqcACRu+b4
lb80dWeKxcN6f8bwtSX6DOBVe5wYGIxc0rn37oSvD6VCtk4qncKiuZVnQEldrNjz
MiawT2P3BXhieEbCmvIlR49L5XEFJWgnKZDOnb+8s+Lhsfvxl6/SV8sBCKiNPrN6
BaZvFdt+CQZGeovUESB8FKxTQcHFPmEaT8Ly7oNHffL28dMIYbi0NHV2osXTOpC1
B1ZUzd4RFdwjQRmX06ZSuyiix3VLH5doeTju0YtAG5JWs+qWa+USrf4GZPoVrA9o
Bg5j6jWik+fk4SzxSjvhzvrBLDd0vaGv8d6CFPUrLrWm4qp6JsUlv0MeLi83wdyf
MTUeTV9SpqkqcbnmZcHBsBRlITf6EiDlw7WFpMG7sLpx9wjSrGkt+nlJXAwMUDlS
fcG0VlEZlKwV+YUoaS3PDCAd6bjniF+ca8wuaWgWJiw1mYCJTFc0zFpk6e7TJKtY
RW8oi1894l7R2vDdZoWCARhBmWPQSrtvch0Gr+V+OmB73FMYMMNi7VFoMzvEazTG
w4gwxENbDa7YA5Tph6u8ZqckMyQhThfNHKSyrUt38aeyE6C0Nx1NnlIrOR7IQbNa
QVActFG5kFHAHV0Nji/XB477t0VBpKCIjZm741l4LK96K6jTE2DZTOu01udT3OA0
DppIvTlkvqztkMS8YcKQ5Mc/5ytP4UkBLfzRc7ez4S50bMPvlnkGJeojkpteJRyT
aa49J9CzoV4FnMULx4zfNcoAWk0jJZQ7ENfaPxGodmCnIIsMEKOuJ8jmj5aK21GK
Pbvhikjbr704JhmS5w3kAHUw5I6uu8FsN20p87mQfsfILtcB/261qHwZi6i8bGTK
WguTsRtCAkYu40A2jnpTCxK3iY3CylI1R+efh4bQhuDwPEFM8UMuFFnSBxvfNEzF
t/Vgi68PJw06Z7AT0ZtZvoifn3Xnp/J9tJ+H54ZQ2hgvdrxrGGZgzPyyDuJp3wyJ
GmubOFUnYn+8zEFqIQ04y+3B3fWg/P19hWd4P/ZGWN53mDYWBKdt2AHKiYgOGJOJ
N7CMIl4FLZwSlcu3ZkEYsCoC+WXexpF2pdnaKVkfiLRysQaWFyeroiwVQQsBLhGs
frLO+E0gjK/KH1btVvpHNYWifS53Ir9crWl7taLDcplacBnquf5hodpK6Pt1PCgC
C9a0FKCJFUzzhxTf1GCyzaco12VNJ1cFmNALHnffOVLAcyDx1Jx+7IkTIMNt1xkX
NaFwxeCPPgVj9bmDj+SfWO/lg0AMP8qrXJSIF2I2SkD2NXO+q4n8HMIUona1OSXQ
dc7lUP5VvxPzUpiuwOpD3Wsw5GbjtiCtJwnvfogaeztCsVMdj6yn8Xql4Lw054yR
r9kbuZl1DeFJfFMgRS0YvypefEgLhTdY5VfZBgHm4Hl/MQBsFV7AAKFRRmARxhIG
p4oBoAM0XZ/a/pAcUIT+iOnWLTBJxAKzPmxBSos99bCePY8Mma2c67/PFHXyaTLR
MZwGT0H1a15jvRniQ+MreUuCtXhU+MFXEQ7pkIAXZMHtHnmL6SKi7r6lsWpPwHGI
6RDeF4giB3zpn2NUkwHKbRVaJroSeooZ2IYVXdrKVdy9LXBRaXEdshmO8bb44jgu
05kYFWyY7EeLwSzuL01GImKAkw7gaT9scaIJEUu0IsPUiEze3jK+93UVuae5/LSt
A5zBqTA3WT3DOfgR8TdHbWz+r7qa+wl850fEHNuij4jg+NBXejeXeKLZjxcNnngO
v/rRa74KrckMuIVVeoAofOr7eG5ePwWscia3Y7U06xmJrrPnVsZnhkNdlRZ16SxW
sj3u4lZfyhLNaHdwKoI7az+WNMH9Cj7leGuhVc8qoAaiVXXHvDVSRRpHk0VFQXKG
YFVRf1/61rkozz3tuEb0QggZI5V0ArAZmmYe/tmJ7vYCAGz/woWBsc6if2Qrk6uo
8rxDaw9/kOMWWXxze3RcDHJs4/mdOhIVB1cLVF5RkoqvL6pS7lJ5o8KotSQ1Z5qF
Jr6IZspHQpqhlFt9/PRigr/WRM3qF2FceiZefhj0EL1csm+Kx/Z0UwA0yWB65ilJ
yRZ0riLYCPpfrnLBZYjHt4MlFsBOqPFhRigKgXOP7itSnfm0/viP3GV7IcWsSFgw
/rxfbaD3exeBwY/wszGt4Q/q/FZ5ZPZQcGCZtqLb4SN/3ZRSkcfKXP/uL6DFJ/Kw
Ht8J2+F1roHSedn/1NDW218XCHPuM4W02MTtIOXnsAlJXQVxgB6AzMRrWDBx0Qx7
0EfGUw6w6wllQ+7GBb09vK7g+olzFudop2toy9TvStpCs+qqO0PmjVM7zyn32+aC
z68iVwcdiyCmUhu39iSK8Ur/09Mf5HHdU3fbbtPcBT9TveZ6WZRzAbQ72Tkl4LZO
0lMJLOvi2pzI0ZAoZ1vivdRDIGBr7aJE5jLlq6rzW5XZRH9AHaCtTa/hmzvB4baT
gUAdKP9BXaW0aCQL9Dn8MCz6O5xsuKywh4ehNGnpea49k9hAWiO2tqss2E6D0be8
9a+t2reo7wCUgshYb0VEKqprXM5BFM6Hd9iP1lWJKjWmvx42qBA9A+jYhH8Rbp2s
ySEdK2TXC7VT+qy0i0VD1ttrn8K0A/Utc+qm385hsAU6IQoaLHlSJORv1tmvei/J
vKq7lyWzWO5bO2oEnKXlhHAQcGq7oYC3sOErS3pCQi7YGxr9tlsKo+WB35HcFQj/
qojoRBMCypcUyUHGOoShpJpsNxLYY8U72R2PXFuxFo9PF9RKo6Idp09HWTytcwkF
C7vCpZN4GunMsXyK1nuRhPI68NE+sViJpLp2C1MRtg35Z276HYnkjJXOC77WHsXx
Qqun0fneeZQM54kzAXZyRNGatzJoQlm2d5GpRhsUope2AoMZjeYFvNhXRjt8fjBN
Egq67Cunl2SDOIBS7qPSuNEMdZpRbiWE5IEqJN3hUwT4cxW0SCdVpc1ow+KAqG73
iiYDjsCD1ohEN4ft2U8eXcPFMDMgqSH/MH6r32wtz3Wa6IssRz4/XKkWpxoH0B3A
vGiY3vOpSBcx+CxRunf+/DdzhZeCMXVkM4ZeEY0FTnPB+aKvuQCM5iQrPDYDoB/Y
g1j1iFCJACWoikFqWWGPBw0l0x7H4N0X683SdTHZr6y7kbrFVUYodqVwsAKAgclu
M7fD7NPNRkSWze6TE9DY2Mat8+Q6Csh6Nx4GtVRGPXCrdy+hUYYGcA4XKlmuY3k0
hJLES6umkJBkLkw7oTwqMinCJSXuCOEDtr74niP2mYuxtWgOtL3Q1lZdBAzLc8Tw
Aza7b1Lzk3r6QE5HyKdUc6APv1XPmsL9JorrsOjmZpfhSzk13kI8nUT5Zoxf1jQA
7N5PnNlECaOK/uIXEQEgbKnfh/vowoxYJKV0mCPzuc8LA+/qZQgmgrX//Rg+j6OX
R5AtEDYoDudkNqkoF14rebt65irVJy0AMuZcqSF1lDWboQVsxlkgls9jmBBEPlM/
r3dCiDy8se61cwXNHq4TQ8Ed6TJMArCXavz/Bf+eAS+vwcpnGMjOdUpKPknIB/Ty
gX8JWiS68HxywIxvEyHVamSYIsNADXYpy9B4UQOe1PrgzEA4S5B8kl/RVKmyrc9p
GdTlewlKi136Pp2fsguxwWedTRkTWDrpKNtdrtojAM98HmIyBUtU0yAUpfd9w199
vn6oYwuGW9XEaJRw666twV9BA1aIrY35J989MQvbueJHh3YJxubKB5WUgaJ5hf8g
gvmPGvGKOeORt0Wd9w7YXK4PFubeukBaCjbcXRWWTnZ9+eR3PyoBKS/lP5r9qNvs
5Q8FbDccEH3+tTvFw5Y6U9SwkUDMrT29NGIJsIX2Y2a7tLAMz+DTQLNW7xUDfCEQ
kTnqljBcH/s/dyvfr7nXGS/FhIat1sNWjmjqRhNNe68mGVl8lO7RYsrOq3T5p3ui
TKJUQM4t84pcdozrt199HraoYh/GH14iGYM26btYqK4Wd9fgmQOOth/9MiRycXeH
4UNw6NKW+l+QhhHg4f7jvBfLCK0Y1EflVj8gRXsrwTVLcRn5PpZoauoCzRpoy9dZ
0u1PIe5lSdp/lTGQ2FSqBi9limPvlSU1w5eGrh2ww0KAjjTz0GLondgOsPHjl3db
xjCz0lHMJFcc4iButq/ngbLZJTQKdPQz5jhgxVcaoFHF6+9rUwvQih5HLpKOdYAn
FyHDIrJwLSirg/AUfiQm0/xfkV35BpB68fkrb4bstspFJI6L31m3qY+YD557HsUW
XHsbDMGMMqOpIIbMnBatbHRZaKnSBaAGQsDNwOaJkxPIlJbZbS2a7wmQSme30srv
5ipH7BQ3Lm2A9XTBHjga/ioxqIqVonJ1+QU7C6cIOJNiJmmvGdRL68teUNNMU9Wd
IWoHT28xdTBwQtS8iWmhh5o0wBE/DgG6f2Ujpgsa7BX9QyFBdGPueHUAjoM/rmdx
V1B8T+JQ3/2YsJsCgxehyxrZW4qBwJsJTg8yOryuOA8v/VGXhj7qawd4JNavR6do
8bCPTp2/MnAA6JBCLro3GSHGTx7uztLPXzMK0/3j4j8jFjg5djSiFBBoguUk4Une
M/JtaSgcjoDmI2RZd0C517w3LygTTSgMz8he8Qpd6lNQ3i4BIXNgFRD2nvJIK+z/
CY/ejoqhkjsAEaS/FNGMbeW/uoAsBeAAfbOGX+cUzaBr5OniWDbsUum3VitneVMk
ls4N2IO5QJGnFJwu0OvhfWYzfLHxuYKwIb/kGo2h4BOgFMgWegxqYLG4JrxjmJcx
dgZLu1uPs7Nw/houudRPaH2aKvd3LOgv/zUxO6+V/iE/CYFaAYwTUKaPAtRsdJvk
LOyhf6B38ntlqbO28LpRx6tMWlj7dKXX7jYsoFlxV3ROw6IgTJH4M2xRhcJf7eCH
qxFO6vDmLfofAHJLS7VO2SVmJWYjb+cB3AGlU4KKCZZIr3U2NrelGMt1uH4V7gXQ
jhZ25SPPDOkXuD+sG0TL+qy110CoXstnJUiYFrpioHW4y6UEJ48S8vdCmM46HWh6
maKsBp2BlHko1km5jKbkfMKyeTXJk8qd3Q+mfos7DpRwp00cKdFtGSdoSXOBOMAB
4cSJrbNFwzpFsm2Ku/hq2ZCviForqgSAuUVRReiO/Rl+34MVGEpQy5IuW9y6fSfy
LclOkDHBfyVtCeObV/JBqgF/UkY6ZMx/hoyqExtWLGhfgdPmbBcYEkG6bNiVrDa6
FTOCQj3Uy+GuPggM6i6uATtYohmkyLiMXwO/qxY3KZiTiJUH/bmaZrc/2BrvCqqu
20wRkrhCXQGmET2cpj9h2YWGEGcuhmvoAe0hP7aV6ce1xXYiGxiD/+8ZHE9spRm6
3FmPt6X6O2baT8LHj0jqDzyzSvZOXkcZq/ovx0IHwNohqsLRVUQyAwZ+xFJp1seg
MMLqic97NT8IO1VQJsH6I/ZovphhKYB1oWnf5AM/j+DdfwB2mZdtEhMdHSPLqOXC
vyLuS67ggEQIJwOhphlgxEzHyg7K3KkEc480mkSvdFvzbWn0zh6K2LnrygweFHOx
62eU23W1wQSXTwcqcAdyQzGLkFTVrMwQabEgkIF6savv47WkeHwWEBsy6iZEpawG
lCdlq2tWIVMIW3iPRxeum4xEJhDdPEL93++nDgPRg3lu0D3vQaSyTI5S7AyQ/f1d
KcoBtgtpjaMKb7zQ5RTIjLiqDQxWV4gt6wL17fgQdbU/NqzOV1RbecKqgkmy/lcf
GjuH83aNys+6JKZUb6kiDUHuUjt2PcjGTnP26YiAegDXWJKWCVqXgk0b2cgP0NCG
hrMzoNXV1ks7fAF7AlqSJ3buEjnM2shrXeB0s60VmRLqqXj5qCWZuwnV/Tconr+C
Hhxhf3t1TBEtKeIavY+nqXp5Y9h4/sg3Vv9uPCPgyEv7Er5zeCgm0L9IW7vZ2apM
6O9BMTwyHh2cdIi8LnMKBa7DU3o9rbTRgL9NrjnmVDPmHQ4i/7H4cGy2sMwhfI9/
6oavJMRbUfWxKkqDYMqFScnVxOSs7g8lIPxCCuqAEOnhvkDAE0KcOQ+Qm2x3l+YC
3nyLPC8JwUHsVSIfSt16PGmBKRvbUCR/jvMQA4TVCMrHScPaTiSXppBJ5LyPCEQ4
npjes8WYggGl3Quh8kxSe7VqtMkkvDBezdOHUfCyt4r5LcFCPaDeVCgleyBeuRWf
7j1yA8PL4jJbjD2bEo1HT7aWJd/BeyZHouY55oTMsL/FaBKat125vPfCO54VKpW6
YPl8IXi3DWOhXLukzzLIH1lwYPS9BJcDbwfnxuArDu+V3CVe614dfvsyMzQT9AGl
ZTZtnS4+RKnkg2od2gUtGrq93/U01hcRgxvRxW4wrIOwsO/Eo2v7lg0jdMZ7ibmq
GjlH2NHj+NzgcGLdzcNMpggZS6XI5oXIFESWbGo6/mAMpghyVt0Ps8Me86xN7meR
MuzmgccUNWOK7fjT2OCDOSa0UzxpQ1bEd5wtm+1fydOjHenStz/Faubec8KHTQSs
uWZzUVzz4oTgfiCShD3hDbfECEIEWou6QrObN3hMPdrSR6xvVWFoKPu95DW+pZEA
EYLTDjvbS7uBSmpdyomkjrlMgmQpr6epzXfqoAcqJn95XreHAQDGU2PCn4FdcPbv
sxYNXIdi4Lk5zs4W40Qhu482Bng08PFgxINEffxp9jbifLO60Q0EMT/f8pnxJ3C4
pK8Cs6JrlhwOsIEukiLktoLnQcMbTKQ/XHq1foe62fnhpLw2PK5UrGWOejpf3Uf/
KHqLviZgmdWdqhSQU31dVufbnDciYS2sw/vyCjju2rPYj6FaruEIQznTVYbobd6Y
NMZ96Y9NGepzEZwhBbx8k37UXrhh9Sy+U9DMEFWwQAnd8DHgK3VL9ShKW3YxyDGS
+wuwb0/1ZPpn6t4wDpkv4hmtPhutVnKGVElHehqTqz+lQYZK9Ws5SLg3iQCZpY/y
JVU3gsO93LXq9vOrYOCkQszzv0GODAoRZ21LqEqDYCkdmSCOChDnJJK+wD6Jk/yO
Zz/KjCNIOqRIpxlVqBXnmpFSsjoXz3UT83F/5y0g33GlBZruw3wOz76jN7zy7L6T
CezODJnr6wXEA4JW8vMYEGYWQ+1kPuF39EEKf5KqiUmf5wL71HA2WUKOuopx8iRs
SotuUGJMKAvvIubN06msBhMcrvaAFA+apeUh5VwD98qbs7siGUjG9N6q8iDmHh6Y
MovsslOGnj7nNsQuYqP6BfBnSl/0wSUtAWtlWXZeD1st4UYLyNTqvE86kUx0Xp06
plLZgHc8MO0GNhQxaI3ouMabcWO6Vy2XXw1ry586HAVijBrjhJs9MWwv6pok71Le
plGx0M47yGmkIwtuPgUbwBZ8mvxrQwv5kcK3loZi87rWSqy1rOU7Xol9o0UEsWVC
9FrxZZHm0c/pa58iHvg0D50mcEbhS6S6+CMOynlas8nXDyr3fMY/4iXqDCeqTmLa
pjuozTVFZAesoEofs+JJ8bGw7Z9UbomyTwSsmK0r3uMnN6nAk+WbXg7rAWmPzu/4
wvE3NSbBq8W4LZz8U9F8WdFeHm+GvyLV19cKF6hhvK0Ry5uKfED2ILeYHd3kFpDP
D0379v8qLmfNmpy1CTM/IsIrwPisT2E4CgbQOYDnp4CTqPNrb1WU4/RnORmiO1/Z
L2QgEwZhpaIm45hDu68bJtDTTVSOHgED/6HJ/0R0pMSStRdDoTYfSzzk3gXftjVp
c2hn/80ydYEsQ+8L6PP8TucnTiw80GtVu2l1HoWjkSHfsrXwNXLmViZNKSY374rv
fsIuu+f//C7S/zDXZ6APfmEedjRiUbt1Nvy9IysomWPer9xlVqymiyPmi9wl75KU
x4UnFoSW4WPRej0qIGqsUBwvWaW/VSmNBwRqaM5js5nDCdQle+zYRDxBPYvTBlDb
kzd34n1/QQ1G9wLI3CikZ51wEg0UnpNr8fYgCou1gHmQvq14BCz3Ht5kCKkq4G0Q
/3ozIfmd3RsXW8pLbax7KxRo+D92xQjqbhgdcIrbm7lSIP9FZ4qdfQmv2gTfG4xG
pPDbk0VBE/Lvled31imGZKFlNNcRD/QMD0I9aNjmkWLHoB7BrWB0gIB2bKY72ttT
t1ysNIPRrvDiE0eEmZy8EYGUIuU4mpqt20IGl3eoXvcXsQ93JE1S6Sxr1psi5zcW
VvNFRyqY1pVCz3Ez3Dbj5DkI6nm+GT7/wijr1V8zK8snuK+JqtPErUQvYaFKB+qT
3gHtPvPke8gybXdE1dcFl/fklZUR2K8rrP1W4UbjvGFD+xsYpOqK5Xc/jtGIo+tQ
SHSqiHQWpsk9HbSMzJJiEGJ5xw6eo7Wuzi95Fx3CY6OY7NMYZDSvzeg9VS7BlzCY
/cvvmGAaTYe5NTqkFKM+OaTWf77gTt20oP98td3zaMKVYUlOgLnHxQHqAh2eRYk6
k5YaZC9iIl0k2EupcyOP9nxY6xjw3HaSmwE5kN2TNaQ5vjt93ugzKI8eIdR5jBOp
ah4KOPPPatppAgGRtDCkt7gOhOGLyPQcBpm0nmgVPvk1vOtBL9DBTgjbMqrp5g2q
d14QGGr9vneiWSu9zZyYH8QsTL/xR8OY98t4SjFBSM68D137MdTuamdoiO9Sw7bz
48V+wo7e52SBFQ6y/InF4KtYfp0QTNO4B105YaNU0aNXihHjCyUdbQUh3s4sjLUt
xpGkfFL39XSuGpVXp6gZFZKBHfwMKVL2KjObcw6WyjF1ffR8J0nCsaSsqjBFQegY
IK9viJY6QqBJsRV1TO4CO3vJ5oa4ZaEWKLHvm+NuEtnVx/Kb1P4aecjUMACUcDMD
ONtl18WV/DxO1FgGTaRmlendO5daqC8xuw3rWFi5zlWgR0nZgpLLr7+6DHJpC7Uv
983AJ3d4NfZAvjDQQmbMimy1Opvp3PxNsO5fFSSlVzcDW72BS3u3xWvEZJ/RThiO
qIpD45g/e39bZwvGqVsBw3MRYLdrUgGZlBIVVOI4HORTkplPar0h0a5s0TbWlNHW
tjnTkXWKfr3n9hgex1L24gIXDErQoE4d4pkfgcy7hv5ZsfnxuUupK6zjk6V8Uqjv
CdzLXGUXPVk+j+ncYDRSCDQcRPpvq7D82PhYTQ+r2mUNlyH/ZdIzH3uegJ8HaqYx
uNQMq1WJzmSXIr5f2wOu947v5Petop7F6urGIODNSrhwptuQlVDai3EanR7/tLDL
+Fjijg/URhi7p60lUi/LF4+oDFJVEON40x9JpeozPfJYoxto3t/CrGRmGc+o7X83
VVCMthJXFVAeIwn+1zfz0gi2CIQVILnqepy8lpzXATjCkB42TD5voIOUlzEdeHwI
PM6S9GpIxIhNVc/j3Z5TIKH/FCbOTrU0WRsJCKcA+oWOF7jNKGyIWON+4YaFbhoI
LKFDRpkfi+xJlwnaE3sFwjqgJm1sx398MpxRiviLNxKXC31A5wiVpqi075oRYzQI
MLzEk6XGttbLlfJdXG2qJSuqMFmpqqJfyY0kPnAm9Ehxq3SwRelIr4KPhfreg9+2
xjGQgLZTicKOrh7/vNGJ4eR2quRdQwKwfUfIVwdOXdWsdH/dEva6fLX5UT1s7fQF
bChabQm2y4PmxsOGWKrHaNhUt1BYkXiS2GgF36RKq2/J0nxQIJzsXQyz60/6U9Qc
VRvRBL1+I35uloMyDt0tuomG99+C+yIBHR4H9MSPgk9CDmQ2Xzx8+ldr8og6WDBH
VKIRq72GPNM0okJoOoGrrWP/fLyx8xDQ8dszRXidbucoJ4t5USRNQi/fXCCIi0y2
9joVgIJOz/Z5m+LDlgqwtikT0zYvINwFW9fFVhCGOCYJAR8KcsPjLs6DOMtlKEmg
uA/T83zEdkhiz16R4oGzWF7qNFvd7b2Tr0InEJpxnhMwB6lu/4cmoBHinl0saWRl
e3qEbYkxoz1X8pRNw3pzizCTb6Ck8u2Qr3FtsXeJQirIJzJd3Fvljj4Ze4QZsOL7
U3LoJ5BUNx3hM6jbqETjdN/kBtTEh6aRz4j4mHm/xBq7AcddCzat7yslfxaU1MvN
ubk4lwsdCTwdqSluWU7CGL9yUPt5Fmn5+c7+GH8OGiGkTyXlp9NFqB6nlnDzMZSV
Jod3/lzLQwDGwUSbHJ+3nHc8m0uKKYk0OMicoOtaYLSZ79q5ZoTAl0ZZis+viY+k
DoEzri6SLUZPWgNjTK0y+w8F5Db+xbEyGsEqhP/ecUO5M22AumpjHkoSyzyD18k/
YUe6eLcDeHzaNSLAmZtT3m0rodnKSgisNiD2US7UzZSRsq4pelLnbL7DJFCZTBD+
iDNF3Ghd3lz9DeG8n4KsuqDfeDjpoT+/GhoXvQnPFSSeIEffCDgG8byhatc4UMqg
weZlEB6fMEO6QB8T3BYBssj9AGRDZyxBi86L1TN2Rj8haIdiLxgovo82LugDPnuS
eewoJlbkE1B5UM36B6NU6YEm2cLgfv8oUMKw/YBeUOG39MMmk1PLMjkrbIkVDhRo
gHzEQb29SiFS/CiiY9UOtzg4rhxcM4teKNU2m1nDhxCGBxGszPRqhnn6TbxLfADL
0EK9l0lbINrAcP/2/XBozJax6obAQEWvZyhAF0Dj2I+aZ/dWDa2WeHPXUgjF7Lhf
xk6EE2bMTbxTV1P77r9SfoSdsQfDM+tH7QywdgDzOuc9pxrQju7mF1VGv621JKEM
2ikjv/lgBEb88P2aKjDezayXyt+9foSL+NEuYIaH9hnlZXOvX1Vn4ZFwW5kmYZtI
xQDqEt/6ETrGMEqpOgWvUgyc7Ua7d0AiIvM9mkO5yYWiPjb6VhrwtQqYuG0rQfJZ
hcXBQabAngjJ9DlWM+EZoauhxIbPzMdJ+F1PViXgsaP4lcOZNT08WHwXD2FpN1rS
y55cZnnXdGOE7U/pS3AiPUY/vaOOuEJwa27gC/f/gMWlaWd0IZ0zjB75xv331BCG
JVdGn/8SO+3dxQ/JHXsyBpFn6IjBPoHKFXkXZlZfBERlrovaAg0TY0DDZ4EfQwsE
yVn4USFX62EldnJdL0UZdh540xHX96ThHMI/XenD9ij94DLUEzOc2ICHGgM/0Mop
6ZEDOhzK3jP6z2GBK9S0hn5cs0dwRSKxDV56tDHjEwHuTrKkVTDo3ZkrK5t5xxAE
eUhR1lPbnPqvt2HNnjG4JJh8OaZp5AKPYM3Ms9kEe1ds61JD5zB41K4tLcbkzNN7
94k6+EDKGTrAlHVvHHEvOmiRGlVLWYaOWuS7bwXbfSumhAj95PWbRFOyw3qnGa5p
AkwX1rzIRtWCikVftWT+PJZZy7EIuAOkcLs3M/cLtShpRDk+YP/AZFMuMfz9nHKk
tLPr6zmaHMzlFFqlw42+rtyFqvauPOshWvf8BelgbNhlc952ts/y+0cdJb+9dDpm
b119uRMbAwgCiuhONB2UwtMQ6Nby6QQafOYPkjpjqx+5NdITQaaAKjhf11svFWQk
Cr7xMjW2B6WRnmlS1tbXExXOudDGHL6g+2ytTb99ViRUkoNFW+E6H3xCe9SgAIvV
fFmCmpNVz8ug6u/rK2rnNF89NQ9WfW4DrNeJelIaOKDBjGYGwutNFjdgBmozCG8/
zB1lRWUK+a1A9+uR19aLEaMmwg86wcxtAcF8W6rDsrqg0oB1Ix9RMnv6RV80a1VA
ztev0xnrLZBY3IVxxWBw1wX/cy8ECu1BaBgaOK+mtWwv+YmZ7F9iPeFVBPAn858E
7g7OVdJVIQkKIX/lT0ZWVUM6zyZI5OHKPrh4lU+uBE0Jv2YzYIZ5koc0iYeNidzQ
3wqSRqZM4rfljSPf9rcPPFAuWgnDVvwAiQZyl8cUSu9MTNCgNegCI9H9gAONfeZH
5wiJSt/P14Oni1fRQkQXq3RorDC0GevTVTnXFq+fbUz74tVARriBK1utHQhVlF/r
WUGlbBfmVzioX9ExB3tLWt49+zWfQDX9SBYCvjDZ91hR13hA/HsOx01X1P8iWnSY
AEcZZtMQDc4YkbL4FdQAJvwWhmXTuV9o05DHc9eNEtllfL6drKLEUTRRxh+ikKhL
Tm1JApoVF4ePAVfwoGm5r9saxfTUfg3kSjA26/UMLWfZoYZE1ldrhONB7wjbBNkk
V5evoFiZcum0mI1lqWK5fybrdDBRWeTxNV96+zdZXQonew6UlNxZHTLvEyFslyZK
3AflUL+S+lnu3NtGt1/Mb6EJz0fsr/z7z5+RBzKmvZThLfP1VPsrJyHe0yVazNef
w5Jns3NDFhlw5fy3cfupaQy+H4EXLQjgBfqXyCYr4MBzN6jerNpwAlMT31TAZZ3t
Ew0CerVlmvbFmMTJfP01uIE038dVT4C98EAM5FQ38rulrQWvW9zo7HAGPGw/dEFq
nDrdFRyaUTPg0GQUxQoFxhEpwUj7Y4v6VSB9HW5dtUPER5OuykfxHwFpoJC2US1e
KVHdx/LidMIAR5MROUVR8mXC4aw/JNjH8WSmAM2dKBN2MX20Kjdk3/Bkb9D+QsZ8
AAdYuQnM4Nvxx6erDBJa6sT438yp56kHVHWeTRkWknvaTbyk7ijzBf0NhDuvjSVN
UUYB48KtA5BWYyU8OE7PawyM8Jo2wGkyUojxvXKe1158qu2vEgraZ3IGHjrGmk3i
KivvMRNc3msPWlKXnG8hkuWFxig/X+Y4XUrcKRMS5Bfxberdp7DZF6BwfRVls05r
jBiKJV6m/1q7tdZNYWAJHqVbn/zkCT7lVVnAbxUktfjTeQMcUCG9RkB/e4v6tFW5
KU326TsxRnW83ApkLUKRuyJBB9P/ij3ZaMlJUpsEWrLiKW6jvvJRTyTmJSn4Jz9z
JVpzXc5mOwYZmBHyzF8e9qWXsY4O9t8Viuy3sMSFlLhitaMJ0azhuXT1kDYQurPQ
U1icORoHUgoV1v0mAmNOvE1jGi7ZxfRBLJu4KhEaXkEJdbbysHUPxpbQ7eOzOYxb
ZYi5eqjNIw3SukYyaYHEzyU1w7z8bXc1/dD/iFxSBNZ5+Adox5HGIWEkpkXIRQi6
aF0SgLWmbM5yDmg3KDwmJZFNeqcIzcmA3nbWxQ9E2nL7IRSPDUG77KhgGH37WkuT
CdRudEwl9eDV/HfoAIJXf61c9pFm3gkaIFCZdoGqWNGzI/TB7jn5QSp43IPQfFjx
7rJ8H0Hc1uBwCZDo4qe+38vFbJJlTRLjet66+Ray6l/l5dUu4oL/+WWIKYGw1Lbp
IS9Lilnsvi8MsSAMSjol66qfIW8f7TcSbeMTyIw6XuUW/u/8XSqBluZEkvJq5r5/
L5SpgQMxIzn1+PrLjt/29EbQS3eevPICSOKNgLd07zgsHw5n+MeWnzDbZPymEivw
oFKg7BdqhxRbHwaNIP3KY75PAWVg1UQ+4RswNY7vdIl6JLWh9NRQCAohfUYhW+TO
OSuYl3rV55ubZSoOUDeYG72wi5/a9WGtPj3HxzkHsiVFF8tTNPa1Dt016Y7w2xJ3
vU8gJeS7qrmnju93CDEVpc/JCWrlpjEMllBM5b/LS7R6DtoORFNjZOTUO9viOtvZ
P2pfTQFy/CL/LJFFdTlX25dLkYTv9JKL4iGXUyrWv+SmulUdlzqYdqkwNgXZO4jq
XM1zVxtT8Z5PZlslkfB4cdUCRYfj07nA/JMursU8v6yQFYD4WkkLJl3AbyLjf70X
1cu+FTL5desimQjnUkIfk+QolSKKqmS5OnfGgvob2korLZhQ9CvQrBVMoh3u3jJ4
vVPkssKjQyGVg0ivSTTZIKGKMqOggw9uLnJtvZnSEqbml5UXnWvC/8IjmvRi6P6o
zj2wVOQbJba0MkD8Fc12kyNF9wA8YAq/mlRLq2qkyXbuQN+tQ+xIAooVHDj6is5M
j182ZTE5eaHpu+jn2l2GGM5wmVvXx0qZslxyN2TeOIJpynvaI5ilrBhBJmXnkgME
9KVrDtqKBDecw7tEoMsaNcbrGRxfg8VN2h9T2E+1jyKBC4wpZwO5Y4Q2hWExPzwO
ZaZf5ueg/u04JcaqxtUuRRPMY/RqH2RWDUXUI2ogC+ROr3/ffqBIGaxhpxz9fvhB
FLXugAz2n9Gnlrrq9JdmpuXu1fO35VPKZuCOHNG/VSVw1sofHrHPEsPre4yp3D0l
Po8eUGnWp5HX47NpBD7Q43xQSsvuGos31HYRFInxz/okebrMNtvO8BHnNu3H+1Jy
uwTlBK10whPMHHSyYClSLS/viC+mrhng33zrhpt+uCLcQZfKSFeVjydrqq0dPPcn
9CQOdX/IC7wVOcR/in6FvNdrZzpJp/nt8Zhjk1abr8uJWz+kO4cQiymCabunqZHY
+rHRejLke8tTWHdRWreHPYDzXgXM0HpK0IFpGuSf4PRqrr2F2Xs2t8TRIsYAqzjS
rZOHzeOUV5J+CTf1ViITNYZ0kphg+YJVJjSr5zL+uuM6gPKSmjAN40jLHW3+rYta
+mYFPhkAv4B16U55WJZNpBtTPfNnbVNkquiR7oo3Jbp9Hsa4n8kKILa5aH8NUpZN
sKpdP9PObF+cdkN/jAbpyKbUAO1iQK6sJt7glW2IQlJNYhz0puM2SQ+WQNS0iHgY
BD7YRxQ5ithDgIS8o+7pd0mMyVM++BqV5b5guw+yGxw2MM91/I4FNDtQ6dpoIlwd
JtoL8cz1E9AiNHiiZmy1seXTHXVHNh9GYVulpK3s1agjTIv12EoI6xj/vlgDFnwW
K6wZpkPnVhtlEDdJ0zUHi6x4X8WuFv0Rv229O9sOgWfHKAa/3isjz044qVcPZvs3
xP5zKJEu7pvVX81mSUq7zgOT+z3QHD0ve7j5xmkQlPnB3Pb3xMJwRstyDVWVx4rV
ERkl56gRXEkruhq6g2S2LFcgZjaM61LzqGEBfB5CrD849AIXsRJXVTTWt3cVhZmJ
55q6VqZAwC+hr6tDEnDBA16CKQXsjfbqoZTXAZVNFE6oU7kqz4VGjWdf+6l1CYtw
voKztZS/QVWbCvjK68nlsQzVO7ks+xrQqd91+1CVZgYdy8XzKC4ptX4BmSpu9DxT
49Z8wEH6i0z3AG06jKh3yD0O4cjz70XwiYFljy/T7FYVF2Oeqq7TZNgvQQMyikGf
AAjq4/sdf2suBxidibWUKKINH2P9LNI4Si31bf+EgkMtGZtDAj7Cg+PvlGuDZvC4
uQPu4TfzPe5yZCLTwvLbqA2vTQ0CHD/E1+e6P6f5Es74L5mwkHBTOC0gUJVIghgF
yOK2PxUGznHCCorfVVbNAcRPy2/NpFHFFaaiX2oaUnvkOwDIZiHIX1OWwf1+ImfQ
3HZRir5+BluYe0wdUOcO4qekaiKs0hff15wfOzQpvM+pBEVg1q5wl24dwpmNZt6H
6ACigMCLFwZ1IwZRdxe9/X9dPqm5E/CTzNMcKGR1OaYpxG0FI1cjmzUE0iHOPVTN
abKXaYmQ81IiDvmzHG6Af27u6Fpe26DjXgef+aTGfeCKjLMMFXCZ1oe/sZoEkjQv
0rtvVRNg+p5IxMNcEa9aA34n5YyUW3XLBhOXRHY0Hb5sj7Q3hGwcWxEln4fjznD/
YAGk0N/YSsfRbhqoB92jF0pM5jGMhDp9PyPDjauheg2XL1LVi6JFE0lISwifEIWm
2ik9G4BYm9hsQZM3cGU+TSPuYU7vhcVyzsboYw5UPtF9NR5m+sewQZuc2kN7jsSY
+CLqbiclPNmCWG63TFtIgN1lDBgtB0fmlre62NPkys2fvTM26S2b20p1iSOOulmd
X3gzy7aQKQW07HUhO/P79UstrRTKModjv3qTLF+WL9bWo0sPHSqZj33X83tRkKtY
v8VL7gKkWodTHWS335O4rS5n9L6Dvc7jgMY3PrAnMO/3v9uay0WiUD/SImcj+//R
B8gKX4dOQoaLSraD+LqI5wA7EoasV0yvOaPM2KfIbfbQRQEhV92dpeAIcAiczedc
vaUab0t+nBS/OosyX55W32UMmNiaQr0PcQiu3s7ajBHlC+13Fwgh2EDMC4Fz8eiu
I/yuWoQNzOpqRwm2BMGxIidyv6ZbQGJ0VpZ4L7DK52RsZet0vJUPrAbZA3gMPbN3
jhdqK2op+6kyHHu3jEaflKNhF8qODsQ5+R9aNwdK3/1weCcJ4Cb+iuoMqms7/zPb
TksmE6uvlUVKwls/CPRYhRxay6RyULuu4TDDe/aNYFYzMrieg6YJ/iHiX87/Xpdi
HbssJmE0Hbt0htQkdMgi5YMpaf/Z1dAePyJ2auFI/4bOSYzqO7Jm/i6mz6YJ51RN
EJtPn6oRfUvA17V1c/D20h04vFHMbxPpSX6tKw0kwymHGxHK7GbQaRc+r8aMPtuW
hzV7M5ARE5ljrUss3o2xBsOu+QywWW3Ppb5v+B2+QPE2Kdq78MBJXWZn+ddCITCl
017gqlm+k8EsmAhYD+3xyvYKx4DbkmlIN1HvKjRIbTo0I64B2g7vLM1c/FRDdtCF
UQTTa69SNo4YQhmc7FeU3hGpp7BBShqsemdwVt3lsj4pZVVZXNLCXS/chf7d3kH2
mgY3HQnVGseW4i8Zp+BJP1L5tPPHPJPwhoNZ+TZqwbiQa7upP3GpdqBG6gKeWPhL
A9x87IMrfyQdowJMRLB4JJ6jxOKwhsv4Yfda46ckFU8U8dqEakFoo6O+w9BvTOom
LdP7TXx2WmC3QCD3O0GNMmYrL7gzeE0SAh+Ae8QymbnT6pzA9Bx2N3P01brAIaBb
E4LfmyhJLt+9eo2j+uoumKy0NNDIoCa5wU3w4Qr1JxUDO2rDpk295JZO5WEfMJum
GVeBGsn4z4r2AOlPjS7XzSZj9T1Ch7WeHPL7/z89GrwTIh8GXhaD60RAzGjZavft
r8v89+pLQF6pX4cVdzG7WZPLgmJno10pBwR+I96AOAxCn0IQu0OKuO9CV2FNo4II
MSKsTJvPyQI0KU18KjRjUECQCDOqQWw1aCwFtwmScQMgsH/VHTFakNG0UPK+Fgop
IMKPzc5ptHpyycaoPsjww4kH7S+F09OxKQiRf7WA2fSTFJ8Ouf5fNyuvMgXi/h5f
ddffSosuNbXXZWRGBfnon8PqS2F8o/RFQs7Iq6ISuk71fhKiJsKiSgEhSrrGyBEm
aCtjEjGXC+zDI+1CYwZQUaXbPiqWWdsV+uTaUknmhoJaNbYg8PgR+CPSCF0eUW6Z
iWY59fHFQWJXuAdJh2J0wnFACLwSdNvajPD/wltytG4c7bwlXxrcph6xZJAS9+AF
vvnwlyWopJwV5/eVdGqAQld8eR9I7cGyGUBv/yO8BL6wE4PEO4jH3qJEusCMM/f9
c/fGBttAJ54eNFXjCqSVZbEWy8FGt32aU51c+AwKBEmnFvuy4AA9GtOCMmufrVOa
wNCrYR3cJNPVpR7aZW6bOBIkwsKO4/JTl8r9+7eGhTg1JhQCHwNMOEwoxkSVKyHd
cD+a9+9Q2nWjFaPwzSCkGC7KClCXB3SFQcnWN3ju6JuDDZemvJspiy1qLCokL7eY
8cBG3za6CveyTwCJX4s2gGzalLIJvXHKbV0mxxaGTPUUoy9GiExCA/ZmrLo7do2o
vBoT+ZPppsRUkuKQ6kjT1TuwXWOZffTCKF/zxAuDdLPTjPELTtiBN60IRZJjM2vn
GkgpmCSsjF+8xHSISkkIrwjHSIxBTPLy+nulhyBWx8RAVNLmXPJ9KJXMS+aRZ7tT
hDMJYsxEuX62RWIsjzh/b5sCoUo68Mtrit+kUWRpak2ephieEdEyOdSMftygUoP0
uwamOtyhZqe9UBIdUCp4Kf/uMbh3ET60by3ZpOwaqHKoHE4Yrbgy+HWMtwia4mMK
C5zbrP0rcBIdP+PXWvHhNyDp5va2/hj/rBu1NFNgvqdbS+EKvoF1iZRjaMbKcNvJ
kFX0srIvRQENEeigxgN/M057VYZl/hzAOfVsV+VABOZwUMMt3Z0i6NNVfynZePpO
7P2zdrVZFjeNzLz9MYkecqcr/UR/pVTopV3AvxiYruDwnLLT8P89gu/YlvIJa/Ha
BBNBWyzFNv6kZe3u4zpGYqepsr2NclqCbGqM6gIgf/qvO+JasXZD3prXmeNCWPzG
4IlQc3NS+bE1hQ2f7A+aXOLJD2tw/Bf/9mHyMoSt1HatlTOvisR5m+6yxiXVyi9v
CQqYINOZeWO3U+5K4CyFFJjjBLMWrUuQUoTJHvhubz+Yhogs6WratS0W5xW58Qjf
+0EiaohwRuKMcibt9VfFPFye++duh57cTU+JjOLdii12OpX6ygPdsiMaDlDev68N
pk7b/5c8cr6NpMNSwOoNlI2vZso9txmXC5XD6NbLOv/xwe8oleQ/A2hD0Rz04SHp
ML0CsNLv5df8gHBbWwF18eg5RETfdb+pMqETC2b5QLN2IPd/1Pl2y3FO2p2aUSj/
ZfHEe01ST/7acBEv8Vxx0u5GAA1F8HsHuE2M9Bz+vqbmJiRwOvXksdjaGCd3VltV
MjinPTFJ7ANZIeJcnMLlh8HuQ4cUnKH+ZHh/gz5kWqYtt8LSCsPlwJrIQbZKahrZ
r/0+omnTerddW2aV/hr3gloS2Zs7JKkad59CCjipdacclUzQL6ToUsCA8zugqidk
9g2Fx3BIjxENT0iJ9WEA1B/1TCfTUVT2nuUKoIlUC1yynauNr1VvyhWtMp1QURdi
mgPCkhGhsjehYpcbCmtAd5BYsJh6aDrxyj6Zv8jCpKbIQGuO+sC5ind+BAcCDbp3
Y4OD1tqt+nW/Xlsr9Fl0poEtHeVntvXzJ+n5Kd7U0rEuRS5zHX921u8cQCqvcJ3B
NPoQ1IDH82fiottHmT1+sQ7ZUn7t+MkojaGK+2Pp8CS7inakKalJurfi7CLC9rL/
Y6W1OlthAELi+d30zVsWDAkTyPnlXVLrmcc9x4IPpGmJc+OQ0JGF9JU/8AFQ1KFI
JwQu3H3XeHLoTwXaUBum79VhpPSLsccTsQ5pKQ5gyXmv1ToDcPxjBJufZPMNLD9C
0wYKpAU3N6gbOOmTwONx7zvzfvolNQuBTkgEDhw7sqYS4+kavF7NjCrIHgS4J8xf
irGNXL0iB+ERgMTkeh6aoHfWGzZ94/UOf2sDX+IiWon1kK+NnYYappxMlSn5yo1R
C9kqZKkZWwuDflPD/8ICsFIqNphk9K+7ZUyo6FqiiaiLq9Z3DA/7cqakpawkJlCB
1G9cjcn506MGJeOs55quOl3lzQX3QTpSjLY3q3LSBiKWPkevnV0sGAdJReuoAZSM
N2RF7YqTBwqPoqQySUSqjYEmYFuuvDCU+327agWtZAZTdkKhMgXVt/R7gasqco7H
I5nlmX+BvUQFsw4d1zbhPNZmc9osGM7E1OuSFoy8CRw8aqXE/xLAzXUheHoz5LTh
/EARflHP1S0dfBaeRI0ARja33nTTCQ2kDsOGcD/igEeMeTzycmhZq23U4CzfzneU
Kc84SVz9we8FfNVEiFpjyz4zK56DKjzNxyVyCQwQjzKW+P8ryqdO+3Zyo5kpcqiT
efI9HgMsj6c03CUXRunHx6GQEd02B/cTbqNnVQGAF82LkMbrFn0YB3O//Swlx9KQ
l0K3L3Bdpa5OFkxqWJuYsF3vM43w9Ik46atRjZmjoKHAImle5KpqvsZnxlV+d0kV
XiPaZnrXUaOrBb3fO1y8oD0yHIpmBd/7Lbea1gIdr+LzU8OSKAGQ4FuojRMg6TL3
Gngwpo2zhN6ge9MIA8ZPLMyjOagf+l/PvUIk+JgH/Lu5XU6GxyS6Vi7i6gFxtwB4
3sL5NuagH7dAm3yuC6STgMDcdF5RqzJgFoaNTLh4dg1h0aUsl4QQyy7WUTvJJC/Z
mw2Jt51uij6RnOPpYl+qQYjbdLczg7JtQzxuarWrA+UzY+M+81zqDWz1FczUsY4+
8NCAcpFUp/Bhul60hq4xDgnS1Z02LaC9X/uOP2Abbt47FOSKX8fu/Jj0L3OKjNZW
oWrmZMt4H4ABZQngJJn7j3q4Oko4OkwJJ1tSgsm0POCUP3c7qSgLbn92yyX1Qki6
pavu6xKOPHOpjRFhCSGQevl45CIX3W40UpgGZ9ZIbbi05pVCYnaujmkMz2+cdSZe
DN255SedT4/xYZszeRRyj3/d+ZRL0PQoUus+Cm3vD4pCIakKlWLLEKVyJ+p8qL5U
nOmJ5giVHYa432dsrIJZVbicQM5ZPllbzrZJ0aTqL1VPx/EBOZ6cSugdattUuHlB
MIN0tEwIspAfAOGhhFiXXIYt2weJ8j5SFHeCthxOfPnNrig0jf5k9++MVIBu9HNL
acGo1XnO3LKyhDwU/NPgGXKQMX6tJUyg5NvGodaWcfuIOHKgxjU8l3D8S4tkMd9A
Je17fwDs3I5EiHcckTGixtCfO/7efVDZ7AMTodw4jJlcUeocXHiyBUnn1jQkQcRL
PXr3TUcf+4AOzHZy4jeS/ToHQHdmEjkivJCgAkU3u2hUmaylf2uySpZbgSU8hm3o
0VckIP9cw2R8LTFkWUg7xkMEkJe0UtNu42g97JowRq/P55Tjv+fNPvB20pzoLg/1
u4BFB2duP1Uvw9qevFeq7BP/qNlKAisPAixXv8YHw+Ri1cts6ot08ABSIzu/pqKs
uPEgthDoggkhxfhzC2Z89YjJRFhvqdKEzGMMz8ks9jmu0nKaIg46J4mi8EmbnPJ9
2Hme3+H1zLxLPFH49dCU3ByAuElzn3dN3xxY2pkp1wr0DHQmrCWrsfJrQnv/eXQ4
r6qs1yilI/dvDWK320oDN2sQN70MoFdkdEjcS5wCyABgEkb/ljTrj15OpkIobYZU
olttBGQ4Gv2yBuUxu7AM6KgwBWV8V8ueBi7/ESLuxA3zD9LXmlNwtVWjpwhS7kGE
Wv1bmm9/e/VCpnz5lJGO8r5n4vAs7GaCO/NpObGNW+JzhFQmIMnsoaeNaIvoC0D+
hMS/P24H9ciXg1vV6uMhMNxI/dPCjA/SyDslYn/Xjk0IQ0IoXW0f2JYDQhkofTI6
WfEZ394I/tjhfhNWfOoutt7Pp3Nyn178ecFTqbYPaiOoTqET9pIL3WRvRMH/8h0h
/09yhL5vLrmZixqr8ZrZCFI3pZ/4FwzWaeKiXv4T0H07otC5GVIUa4UfqWAq2vP3
w1T5ndbs2Bn+6CZ62uqkYePtVtX9BE8ELSaSfgBNE3LuYx1mZpJ6XDN3pjnVPhMa
VUx/me6tJCY2+6c7pm8QzhRelElefJhsVDg7/e60YfsLIq0fq7bgFSp/a+mSf5S1
uOpW+caNQQgYjDRaHIy6qGbq9/y0SVyKuGf0z24lY9HNi3DYh7Luc4SfNipX/jAh
0gdC08Yy4M6G7oWVa0qN0pP+nroeysUQBV8nMtB4XE5YHg2szF2ccNVClHKrzKme
KmZIJ+cqlWf5/se1kDH7RZWit7I9+aYbdS+YD+q9v4bGrkCc4W8He8sdf9RNkiLq
O7v7bOcMyRQwox5MT/HdliHAEU9bk7vtS3DlDQJnEQ7ci/yYy/m5CYp/7ezZypmc
xZZF7IMhywUbm55O841y7MwilDh7ZBi9QUSKLVVRTu3tL7wQGsEP0fcjLmitoIcz
Ks9qMwdS7fjt8s3I0h1xJ0cXX3AVz+l2nS5uXvE7mQ37I6U0gdnTsLeCZMNn9qoI
9xNunOTByP11dbMTQhGNMLo6diGt/fGf+tfBpVmgLVAlJropEqMgoqdPO0zEUQxT
sbI68uZcFBoG8Si2b3o1PnnelWMoc9zLHBvNN/rtnP0THmyc8KuF4ZGVxIZ60BWc
NS4EPeksMdvmcPnqwwI6NkFrYLKzv2j/TVR1SO6KOGI6RGQ1w2d6cFHgsbfPAGLj
hRSLVISiuHuG3/YtymPke378nPDao7zXlqXbtzw+1PEdP9SGC8nALHSI6EWxz935
qkIDGR4ynQwYRKibeGR65h4JzgMyXDWPeX0BL8dFynfPXf9EJvqD4gSfjz3PAl/B
oNSH2OkjBN/lMjqQ+2MxB23Z6HXZVXFVf41s3MiE26DPQJc43Jf2SNsRzsvr8rHy
YJSZF4Evchv/vIzehC/tQDTS4KWU/Liox5WXWaKA6+v4nXKKn35cdg54PbFTqV9n
NywFgQK50j3Qx4gRL+0qF5iViMSrUZv6Nu8J3v/N9NQ9oDG0Gy53mEaN8/I8JwRI
Qv1PtGyrqqL7zhLPvxFSCyAuRMujxfMnpq9bR8ZSWpRrXBHZOO7NvZVWDOdvmpBV
xyDk9h6kur1crHx25sw1qxwTyNaOEwb32zhj9nBkxh4GblFMy2wTdZGtIhr5mZCe
toC+tPO/Tu+FesPQSGxP0hCA+MHt1MZJ3TO7NHpq+T+5DmQSefaGrKNa6N4w898F
0TKocHm57N8QSxxe4pErxVQkj5lcYKbHqAn2WPUhfdx3tlyWNw06MZriNwrbGUQd
SbgEqhsHLyHvntnMX9BA1Iguy1zg8dFGM1I4rXr/Sg4iofLQYlukWskyEsYcs+P1
ihze/zhgarikoGrlKC7XoSkzx+4gZvunLtoM43kHL6hmUsMgOJjAqB/XDtPAiKGt
pf0qUc4KKuQ5uPdzA+UrffyZQEpvRWXLa9etR4PFRRyr2woblxbX5IyUKhbqoyrQ
JmAQu6a57J34oTf29aGltz5xKnK06hCaND1R+P9iHfXF37mGX8iHrPuQnRayWyrf
8BHc+UEk8XnHqe3PVhF0P88S7DB5QQ/wRHAwgLpMapOeN0Bb9gVJh9Zea7u501jq
4fluqyP0wugUNVlpRyInBUl2WuRJJZo8O21LdlJp0I58I1BoBqfZKz/PZxgVCgmZ
mAtwqhQ6kuIwVonHqzPTS88dStCESv+6Pj6nfOJgRuJeDRZmiR1BU6OGPaTZQaCH
B/lfwXwl/CTf0D+Ao6QTDVdY+AWizrjsa4Uci+BV8jVY77jPIapOguGbpknWw9vx
MiehJvFmT2C5I8+3+Z0miF3ImKdTQJ5f8r9bLtyNwzMSawVdGHPHdwGxImxkM89Q
Bwu5rW/+u7iFDFUxcgoyPk6l5iwxXXeyFdb4I6KBYW/WosRa3KH0TU9iHA5aqSPg
SrOZx5sglN/9/KZkMTppWGCLcm17Jgwpun6D4VvRVbW1dSB4YHn1xHpmjOgxt/3e
KruadYrwNrZuQch9nezoccSpG25qBEr1jEGBRuWFGGvTgk+cs4+9pYszSPlE14dD
g3umYJadUzTd5TEF3iZOj6T2LPEEY8LjV9YueZ9uOkBC3e+qKfvAj6Hr6iBgm+Qv
lwXv2ixg7TGUCc0U1s15bqhus9bJW9sT4wZEGn0ZHc39nR6s5mBwHuLVjLJ1lpGD
Ni12E7T2VRxlJtnLKK9bc516x6aFN0/+I63ot34Xvcy2IX7MXfjwFc9CpBzcW3Mg
+nCBL/cLFx0a71jgtn3TqGTV2pqAYMVqg52U2zxyZNpi14zGyEX4Je3eouqu13GA
bPhLlFUK057V0ApJPJjODZw2uMKaDbGrPUEdiyGoHNAQmA4DEtDhpPQ0Ju/+Ar4w
NcmsSIngEJ8eqv49XEHWkOVouFh+Pv7XjqoD1xj7XdBZtt33NTsIFnsmR/fKqypk
9ohQCyjynwRSWz9O8MjVzSAY/ZVSdqnffdWMe9xUgidfiPqrD12sz1a/N3wzUI+y
vEqpo7IybRJrmAY7g3kIzw+EaP71cTmif6kDMkPxRydJQsMiyYKfhXrXMrh6KfLf
zdGSuN9+YBXbAVc6n/YlriS/6I7Z1kNQujkgOd9JiPOtYRJp82t4L3uyInBP9Wye
tfe9QnPsHk9VKsU9ZyWAKiX+gXrCZoLAVofsWMJZ+AeKVVvDsff30c/JE/HN0aWe
ylfgsHOx2mygXAjt1T8Vh2gUUIMA+23i+95vFnzVj0OeP2xTQjyvaLcM2UuiBhJY
nWvEkmKOdQqL8lJQvseESlumazsZlaU4jZpBFxk1fteTs9R0l00ogDYjDDgxF9Tn
+Z4vMjhawUGNfh7X/zd3BwQ/FnkgnQ4AUyohBK0ufO8QGCZVvsIXLT8h7hSKWXNA
DSyHQW6u7pj/8lJ7RvUm0k8pyn0DeEuwf5bqcdPHoT9oAK09u+7zEgkdijuE9dwL
GJaOesU6AyfxYiIQnl7wZjepAI20fDqyZI45Uc3ax0UZ0VuH/cTFI3vNdl4oktcC
fEf4yVIyW+dnuncYnB9Yvcvc7FV/bePP6yqf8Wz11rkfo0mbBrb1NLtbhoPSjlMr
QQVAPUHHPX4TeFlMDqRUIuMwaqDZSeh+zBTSnRIWt9uh6HhDKRQDC5p/SQyFf3cZ
wXuiCKo7o28V1xcb93kkfh765a85fMpJiiOfoNgcIdTd3VS8kvL5pDWKiO7yMrlw
ue6kb8LoQoSbNrvzV1Mga9N1tkaoOpX0yApN65PlLf7VxacH84Db6wb9WLAl1RTI
lXhQJ28ql0xgu1CErZpqRuIMRYukIyaR8unaxHUF7a7nGw5qNY1QoNBp8IemVFBs
EFVi54/vvbM71T9ikDHI6HmttvNdcjnhqGDNUMuuEml14OoDs2IIEYMX4rr72Rrc
xHRVVifmGBGz82xUJ2rYSMBJVDLHxhI6gp1D2/FFCQc7tYAahwp4eyBJnUIcxEnP
dACc1ptAU1wbM8s4ZlhMvtwv8lrVBzTQPfFECoxp1gupc5yIDTpj84AlFc+zTVdM
Eb0k9TwylvJwZXh1UbJIogKgovc133YWKradABvCrEa8I7CS3HF/QIwpGI+r3J2Y
o5tCJVrlmV6X4HzslFQhVTTt1DH3V0oKzp4evfzyRlpA0PSBkVAK1jcQPQWTYB6+
+Ef8WAPOJOdyR/l3z+e2kkl7TkzriANcXDq+UPaU27QoCsQYwUvMpHaniqqtxTnc
D9KQpP02wg4VxmLwlTrzaG9CUd99ECXAEtuAtBUpLBH/+Cx8M5FThAxeR7Af5yA6
Iqu2FquJhnxP1m6p6s3Isoi5hJ/y/iPy+Sx36sJI1icNV2FgzVxeUpyRGSKZzBNc
U6RV4dNt3fIW3hLnkguB6KSayJKE1O0qG9x81dfmiZdXjKPvgSM6BXZDZQecHk1G
hCi4iXytobyGe2I5ZA4DgAqJnw2ySQfKawm1jSW+lbOR8YbEDE2Ov6es91yoLgt0
Edx9hRNxZvJ1z8+3Xub9ualwJcxXD9bDFZ2YVt66CjUb8taw6z+TdyGroCXzfNqs
CMyhOKzcFnYMZ2JRpJZqg9LZvA2PT5K5/iXVpnZFh6J8Wb+l+Y06tMboqkc+vS0+
uYoDm3ER87CnWUgX6LezWwIzEWybexP12mS8qUUe6Ix1WlOE4H8zSQQ+6WEYM6GD
DuRxsoGL/xx1rXbMZqrOjDVURtAPOy0NfVqTvtmsnSdF9I3wzzTK0mqnI3je/k9w
CxKRoHVnnd4tHlDIG2hk5Epld2Ywk5k47g7hPmVnhFcuds6shdoqtMpvkaBO8+OL
PhqinYLe7UIrawzGAd/p0W210WNRd1RPh74BnJ7KVxgLBYBm+oJttmFlYBrxSh3Q
aFn+eoYknFMW0sw4mXHAGICV4i+mvRbXIloNGZjd3G9MWttCCo84Le//rRNhEDBm
v27qBH3UCxyBfxo4QhU5bkueULlFcQn6vGw6UOTYLzPfU2wxerN/vIxypA/J7Ang
knqzg5JlDmcd1YNYUSJM7QAWEIMF6diI6KpyQJKTOrgizrXSChEIDwyjREoGNUAe
sbVJWiGRHepiv7qBQ68dcqDbbHSIcu46fAlo6pqtZ948bW+w4pRwVr7iqGpDYX2v
rs8keYw9qufo6pjRO/294PKzC6CsPhIFc0CYVvmCu6KtN3K9zj+mj98zV5JT41S5
ZX9I/4+HaRb6eoT640zauSGwZu9Ppw3/f3iVGOKoJEBgBAZPnOKGX7Fm0CNyJzwc
NDj4ch01erUg+M6CwH8lVxR3szpyGGFUhXzkw2bR9HewtjYgDBRLSiL1sJkz1REV
IP0/5bVlOrM4Wmiun+aKXu/Y4Eaury9tZjT8nc08T61TPAmlB91Al9wbmf0O2px8
t9FqPlzLevFIOw8fcmaP+a7L3leqT/V4RC/ctHRdz+m/H/JeVOnFhPVCtz2lZHT1
C4EN6rdow9v04wsG6KOiwBYZQt3qh+uGPtmIerW1Wym8b3Blz6LW8FqXwjJVc2SM
itZFC8BtsETECDKDJbZGbSLgBiHoGTdrL1PqZMWs9xYeXw4g5qu/U+WrdZUMTNgK
5F5L3JkRODXl8mlgYNGfLGpNzdRMYUsqn0NxFsvC42GpJ93QVwC3MUBEOcr4MUFQ
ibqzPiBH+AjRvnA8Z4mmUZVx0mqdpmT0syn/pqOyAFtok+x/bhD/6aXKByCeTVqV
K351tP+nONW8D6H1c8isv1xBfkA5Qn/FmmrfIxZ6GkeTkj+X3U5+lZ6U945UcugT
nlQ7jkVMoryevJ7c4vK0O4tZSINuZPiVZJ7mv17oSIqFQQzqHavcGxbONQPc2S3x
Kv+YxTvpSDG13Kb6vzqUKWTZgKlccI+m9nM9QG85n0/TlgcnyBzVv3uIuda54Om2
HHpCGspnHzNF2lhqyABB/xWtGU3E62lNiy2TDC7a0Lru/Rms7u33+i7mi5lloUXP
qWUeJ/JSzMFJO14d+XpSSxOIRsWCvujH1Lil91Ij1AZmeuC+/pQtPUGEbddTmTIr
BYZ9zsAli7wnCd3O2EA2o/k1yllPk1IdY5etlmNkb3sTt8fwbWp6BvG8w9wVUw8w
NXm9zQc9Ww2TCf8SZYO9/ovkr5nVA5FcU/1sEpHkUutK0FvxJhZOsHPxwHFRv6pF
NI0x7uGHrCxaEv3hGeMgLLFnbEwUP3nDYwrQqx73yobY8nYFJskIHvlPk8gcMIYU
XKH7P4dzD6c6vvc8+ZYPZ9kNuNIsFEsdvm37bbdAT55L2YquY+NPidcl9QPxBhnr
xSOC+vP0bEiCHtpuHlh+aXo8sJWfzO00zihEzax+zPOGcdHgVqFndnFpMukJZ7BU
JJscjEKg6wd10oF9QcbQDERsEQj7Q0KiR2BupH5nGKINtfA0yXzRGW6PXrbI2B4z
xhDc/M1xRn+GMhSSr1f2n+oxiW28/KJ4TH6zgmv3gAjsQLwwgk+YrDgMpf5Sn+F6
1NDV4L2gc2RK0YK07nVZYWHmJ0nvYQw613bcafwO/uyNmrv5wbg9dGDwLSwuAuCc
LRRIW1En5Eiq1MplqH11W8gT1CXpiUt7m9is894cIXobxdXu4Zt8S3DqdeoXQHUr
CSdZN9cz6FRebGHUKL+FykqXa/VCmj8Xrm2oU2AbnxHmupKrVVUkLcVMnsafFD8x
cdN9GdKAjvIUO7U0uEzz+LoQIqz7lheG9yEGUeW5lS7TZwaJKLDbyjB/bkwUCk0j
7cQ/MeTIuYl3UiejXu1kzxbfex5PUszUMgSqLdWHxCQMvcI8TpURdIUdXy26whuc
MrZFkwmJ+YpN82mCMqVEJ/IQS2i71vSgMmuwAFZ3xxk86aIxtK2o+G71xqDno+uw
f+pgy4pRlOB45iPdvHjl7BhTUZF3UL3p2gd8i3Io/57EGvU9Tx2OlxKl7BlPbchj
7i3BXescDGBedeeMeAJOZ3C8b7DQqJFUVF0NfTSLg8HwOAAPRgK4nliqn6PXbD3/
LPF/xYrkGyRMS5NDgTIUKhinFlMSasgZhhZGbwCb3mphuyjLct4ByG62LYi80Es/
XYcNPqHQJwRRQPbqmCJs2LwfRglj4PWLd2VBIvWa5iPeklDqOvqtHWl/T9XzrDiU
+wEJlBCx5M8B/y9lqp5aAWF3zrQ/Zk1R7dFdLqYJCMdlj25OPjLCwHdoYePmkzYx
d0B9OldpNbHwy8ZnWTDtfuplBLjD6rHZgkKqWN5aFsIRrpO5nky2TXM15UWaouPM
eOEVN1PiWYfGqXSZzWcgIR8gUmORkGiURYGNDaEk0diaVflO+JDVK1lTTlXUGb0c
wzemHYzHikdr0mZZ/k6oR8tprADSZ0R+bcHEHTIXaXphMh3cULUMJXjvii9rc57l
4Rj4VZBWc2+rzkGzardTw9qRBIOZs61YGzOToZvFHOzIeICUZcP3mhwIeOrqDH/H
9+6jy8UTrTiWphIcwAN1DprcWJlXyvO2XSPhDDl0bUJZDHl6MgcsCN0wwRtfEaSt
alRp592S/2Fn4Ika02dbG5BQw6uTGTtR14DF8RgaMBDqL9WKpIjMPgj8QsqCU8Ov
ZXZ4FQND6g12GLmbkVcgMJH2ymfsxgOURHafRvZZ1NY8Mgo/0hn+F2IZrrhS/Q1S
qk4O9lIT36h3I4D4DUgVyAQfYdFmt8NxylzfMDBArTA7agWs5MKib/G889MFFQbL
oObS0+QZ+Fta89dm8bTdHm+gnHWjRex51QAL9Q2kXwlCrNXzWXaZhEpLkUWOWDog
LNtOVM1GPdJT0WkBu8A2vTvIs1xOwam+H6/GdU6u+RTMkXOhgasHDB+HbQ7vUTBo
lJRMUrWGYPltIaLk60UwyqAkIn9288r0W9XCZfbgIPUTCw8la0FehF8tF/H4uc7i
bihLMIqXID5aa2P/8bwGLEwGdaduVR+WxBkOtA/JAPFBAeju41Eqjv2UTRVvH2K7
GCZfwYZE2UhA/4PeUUajnIA+DuGc0RO6YPc2bW9gyqgnunayjLPAt2FirRymHfe7
QYhF3KFWsHcKuet1R0MVKDaBsBCL7tjGCkhSHl2fkrRbP5q6wQmQIIj/fcvUXfAC
Laae3cgHrKrvFxJCmtXJv/12Jian3xhoLuyurKvsmaIrdG0239N366tH2pMRT4Zz
LLb6GT+LXt3N98d+uoC0oo9S4DH2buG8bDcCv6xxZO0lhYrTwnjRCWvkad9LcACZ
uDNkHTSf9+63ujEQUylCqvPA+xVynvoaSnWg5fE9h/MG/SGqgKGnteJZ2mr0xSLo
L9VuuUb2a5jwsqtbhgUo4ZTt5AaX4XGMHq0fP5BmTmfGCO6/smEkayhB5NbzTJP8
0nJJ2EcKe5WDlvC806VsCaVo23NDfnVXbB+oUsKEN2T2VZAy9Dt/0LqaAYdxRAQZ
rykx/h1zVjXa4lHR+crj/hLwSf9Nakny32WHHqAsCgTM3ijmsn98gNk+YBdPnQfl
pcRR/EeTIkg4C7CsEPMBiaL/OMZrrqaslzqzG+108e5R8EIO/gfY/SajrNw57qCN
8V6KRHWSl4FVTrVuT7DfEnGex971MxAn1IH6WgYet/Dr25nEF1qqF4+tO2ZyQ0M1
ZHfLYG1FMx0U3gzcrUhVeNRs7MHFehewhXBV8nE+4chf8w806Hmhe7cQT418KUyx
CH3cM3a+WqRpsjBkdBgdpgRxNylBHSPvYl9BnLRiXvCfCYq0Y/psKn2os996NuZk
zLTAitfnyV3iZgU0qzN0F6IYzdInsmEZBb+VW8K133hButPBIchu0a+Da3ClVkLG
VM8f/qeC9Uaim7eP7f4RnIppjo7bnAGS43zyB3gAt5DZpmTnfVLL4eryNfSINCxt
kRax9gfm441cQmCSanYmJYrP70eR1LlsDJ5i29OH0wyN4J9W7ojW+iX3Y/UYV1/L
UEJBn/QgqijqocwgUtDeVWRl8wxOoNB02UJ7EcV+wOETNXm3RWOH9yyjj113xEVJ
uvF0DtciVmFpJPYjFusfqkKuVnhnHtouI+tdLSOx8ba7ASvrpaCHKxYb/FIj+0qi
5Ss+Fjd/i8yqVbdF8OxEWNlcsAI5AO7njpsLbayWvqEHM3y/B+lxUOimTV7wUhYi
Hut5zH1bt4C5z9QTP7YokoXsnbxz8/9EH34mw9ojsRg6umG+7+Uz7rvTmqowkd8F
nGgeO4zqtHLLOdC837cgUzHIgYxY+lK6n7pdLYiRovqBy8LtG0hCC9ryacsGSDDg
TJyDvg3/TOtVafx4Vd4MALW2carBlAKaTK/DWApY+VkUQkszANh5KME7TXT8r3BI
Ugs919tYdZb8x6IDtIQhr1YOkGCrWkKKFLGqn3neZzn3T240fiA9MBRu/DH3QZtM
pLHXWD4b7Wdp/2XRFOQXCH1VoMBeilRnh5LCOQrwaQ3eE4fobEf3XbSSWCZ8lRru
c4VhNbwov+psdi95jjL+6ovC6+jdebXisk/3/ML8nqJC6HN2RV2f+N1AXuCgSl3D
+wYJTR5P59AnJeChPKqtsHlLOgYAukPvvS+/UTOm1UQdel45NNOSorsUMyeiWj5b
uKVNAdTFLWi1OS0hzKWrlrkeoQ7BeoIHHW1mfXYhkQ6pDSqlRfHKl201w86xk90/
Y07N6Ymtbc0kJAH7uLzC2U4aKzdo0hMbKDVe6cLhcCBhEIu7pVtTGRXr+RqZwOSd
Tc9TDtcFfzN+Lq/Aq7j/VOmdpJMoDtmH0YbZpHDj8TAgzrMjn7R6LFjTw9WkgVmz
QtkjY2Q3AK02eR7x8arcznLoxo9ExyAsqb9ZJ+wyoPuIZ/i7T9MdARqnP21pdDuF
JVIAFfF6VX37k2e7w3xUUu9nS0tzr/VCzhRjHgRmP/KsvdYW1qW03YoulWAU44LY
t2DYmC0BpkvkfK/STOc5oscj2hbHcmbv7UUDri3shRpPMrz7uWHaXZUJfxJbv91q
id1dAjg+rLblJM1h8qEEffvQrb8hY7yAPlAB92yIVdUohm8ioNZLe6C+ae0zFpf8
bTkAGVjuWvP0FCyxaEiOnzdVgkIYiV6LbggTbg8gQTgZ/OSz5DZie9g1eh/i5xDD
qc8ZsHcSaBBpCIxhPPRggPDnUuPi+ux2KjXPZlfr+LBbvpKhWmGpNswV/rrZRHz5
ztfTlUyeBYQxskzFDDQl6SaaAZx+Fhp0Mac9MsT8YJ/NxS6azP5iUWxnB/8axwNF
LeK2mQC3Esj+DDzvyCB3ZUMPzay+PIPUsB9e5AVo030GWx6elNsKriGdvInh5TVb
Oc/wzALvmjvgh3l1kZ3/L5AswQd4gNL4EZeobz0DnMDsXuT+e/WOgMXJUakuK9Qh
F3gUwfR4BUHkGGeeMIshSGYSTXGHxwMwwVi4SGCRWtPSX+baoyGUu4Z80htqUh43
YZTEITGxq4hcfgZR+WEvVO/FiOygQFx9/R/acIupUGEZCJ0Q0MW04+7Gst1e9bva
Zc8ndtVPvRHTm+MTzpEbIBY5aK+Vi8FN1PXKQ+Gx0j2bkI8PcCzAdu2iRt9B1Lhl
mfwnqIOX3zKxE9ZRv/Sr2dfvQYkvCxNBAg5hE/Rn4avnD1+XCR8WllqHq8pBFFBt
kzNBghX/zlHlVnHqTK/xirp7VzzU5qSvOwJnX3GA9KIJ3K338P01TVM/iobNOiOU
nN/THKKa1e0EDNwMYD91KhyyqU1GQQXirA689oHN6xN3SG3EVG8HvO6lJNZBM9mO
C+kJg39xNGwF2m2PQ1kAduFEfdscJgNiMJpyYprkVuHfM9/l8rJitBW87KBPkp7b
9ZQ6+4W0opdbQVBMCIT6lugCBW3eajxcHcP+rUGSJNCwYUUj5vjy4Noe5HRWJAvP
teUjfzojS6a94xp/9QA5f1yipfsP0KuNbMXnTaxUMdxNbudr0DxQtHVEQ8gORYbb
Fio4MM0wLFmqNy1+5YNizZUnmSlhnoPBPJFTXg87NbH1iv+//AyQ7LjDf/cgXEGl
lNnqL9sSdzU7qF+Z7whFdDLZ7age6fWFNb+/oE443lMTFi65r41C8h4cfKLhs+1Q
zNoZFv4MQtePmxG+f+YYi2Q312az2eT59wwZsdpXo18JUcadAzg6N7Fx8j9vFfzp
tLrtZuVv0MWxace+NY+bVQ4rKhmtpR9AXqWFOdvVZw69uGazKOhK5i9b2uvi2U5X
RyAWF5eAmJww68g7jBz9bAnB8agGuAwb1vGHLv8EDXqmJZqiA5UkZV2WO+psvKG+
5SWcK6r4FIK9M6O+ESHNkg9BI+1qCJ/zLR5PpKV4/3wCrqgDZoy4uv7iUO5hUOPd
5OV8DNGWm7Gk6f5o45u83fiINqhiMT40C4wCBTtdSVUV6QxFgtgSR2X9kIjzmpbZ
oXrmAwrMdpZHoc7V1B9Fdlm5c3QXTYtNHI4BORGJKX2dc+XEmAGVMAM9UdvJpGhT
QPEY9v69+YbQ/UKtgYQj+a1aQOqKTnV/wsVnWsbjoc+40N5HB6nq6wwC9pPr+Mbz
njEecrgU1p9GUCuHPYBcJXs+XS8oQDWXevdxIXZRYz+eY1ttyoxc+73NVK3wGD1w
+U8EdYgAJg8dc5NOUULhiuQE3fUConPou56op10mZdqUOmOP3JmkkiTwEnrflJYd
a+q+JqtUXpYaRTcTKc2+mVo820QQdqcr6lQ2nBpCu1/zghHvB+sZH8nGBcE4ff1s
yAFsoxs5Yy4QLKy6pJAIZpi1S3O0dTHqKuhYLnKgXWVkjn313cYnY9XeAogHgLr6
aH9hevucYM4jp4o2yOXqwA/771khkp+0uEH8i+g5DRNPk9rcCC5m1zVFto/pxJQM
ntfIUe8eBoBF2MrTvkUA8DhBcuZQ4IxpwztAs1Yl+vAx/611ohH8I8nVFgmKsAy3
td5wB9VhZZNn1DUV65BbkmIEz1K3WmAySn4LlKYwu7vG2Dz2LBIsNu1MGMdQ2SGi
NijyALUhwfWyP+WYaDD++8VCMtvAUNj5HrdnUtZgcOFQBBv6sxy8ufXCK7P0FQyv
jvIlKQpX2HLEnZsyaEnBP6AvJ4punl6/1sBltQUJxfv/P+wvhPxw8IsMeAKnDZfY
9J50Ot2iE7wonMhcVnXlLElC/vM+RezYRjkvcQzj+gcglzRnpxWqjMvNbNAcvT2H
tqTZAZDdRUT08ywxCAs4hHYBoi3H4EOnZ6wJhpUr+XNvuAMGV+R1ya/pPF+RIkPf
vYInpUFFV5QmtmlyN/oa0Yj0KTDtZHIWVJ2fXU8siW+sSFprcZGgXYMqDMHmiwuU
WnYDdIZBbb5I3cDH4aQDn5arBH/sDVKIN4Xid5Fc/qMmsUPNEXWB901WQ4sDjVW1
uP3Cj0MVTmiMCC/UhxdKj1VWLymYKBgHD/3mgg5NKd0XZaM5Mueuzwd1sOqNSA1L
lvAAGHOfNP7DZTFXXApd+2Y5WlimSRZDjLqxcRmoNMuLnFQnYVKI04Ltaij+89mj
uxV8P9NJwyvM7lQbLUZuQuHESzSsbJ7j/tTK5sRrIEPYGvqFLxiyzlag5ebYnTZC
2Ks92LVzEP/cqR3j5Vrp4AapUVbW9WjOxuIWvKZBwHZGGJFjBT6dUgUqUT7CfDPY
901GkGVEqK+Zs37QJuftlxB4LNDBL8I+hncaSt+MnkUORHeS4VZbe+ti0zPrsogx
L3FTwOrEohHcZzZH+tjjYA3Y+m8C+cBGSMMy1cl6dJm56iIs2eS5WA0JGULSi0GX
cqUX3kdQZ+mr1jz2F+iO8J3ldwD3qk6GrLwMTGmq4TRL8QLejk9askLmNv1jj1Mh
Jtf8paU2YbMQZuC5dtL8cU+b2iENPgDxns7DVJLioaYKHIRd6k0f7O0xQz1UyIYs
0+KQmQkmfHo6umF47zsYjkWyqoyzHGbRQEdQ32fk/rp++AnFzRlcpykyioa75Msi
DgZfZMrXdxNYlyPJUVhX5HXq/uAKeU0R/uCOrSOBqt0mwFi+AA+MLJ7KIuxNYSez
KYbmafnZCfEqoUdaUar8nSXE0Klv3otapO7zfld3YbACmrLnG60vQNxkeZTzn2Xv
E12bCmLHuF41rOr/S3if7g28U5KDb4fP6PG4AGW80unxdqOdhg2nzZJb3NTKuedY
Yfg5Or/83+7i3GKfiGjiikXeNwLEVt5IBwuTF500ZPCoopPRCiIYOGTtFMvTb4Q+
at950u8Xzi9ehpgvD2VgPo3oPvduCAbvhBz6fzS9n/Ydb2vbng31zc4pvdTJcV60
swVNpLlOEyK0GG3JnUNq3rTWQ/AnptNnqJVa4K/Qbh4bBsiPAXRwfkmtKvzgY9ZF
z2AzpLNzdWuLq9J/g9hPPakLE3LZ+p9Ay3rhYTjWCw2AtiguCKfeg30L5GRbhlHA
6HQWr5YjhV9dGxge6q8bXknocd/9zn6KpMJd4jO+TNf1VRWsEyM/4Fx7A7qeeiZX
onh97xmKEj+/hoUMpZqrcpoLve4Fc57XWES+V3XlAuYEEPt786oBz/JouKNRa/U3
4pBzGTFrkAX0z2bfRvQNSWvyNwr3dPeBdfxYAINfokSqbbeV5T/AQDT3dGuWvIYt
rqhgM7sWD1jEEzdEo4K9HzaVds8/jHKvygEQ+5PW1FQQrJBoxG3lYIbGqy1AaPPD
sWpjAQG9j/qMti0f1tOxxGMmFR4lPeNNHv+RTX6pm+397q+lhOnom6jVOeikAAbD
KaGJ7ZzSNmp5FgMrXG0ygCjV/9wUjwIO0vOdCUWmKrNUgJNaEo3VLRYG6PvbTdFs
/mXBhislp0iTuvFBdmgCjZXJphmpxh1Rji3WIXziE4UZgFrfw2JBL8rndLZ7XvZw
8kB3rKqCIKwe1fUGUKCHgt1iJM+AF8FfeQiCv2m4txgYpQHJEDay2u66+gUzxgR9
uZCQLjo6VMLUf77HPOQyLsBjb0a86IJoyeKSwN3Xgq4ztvgV/E/jnea/UrL4oIlp
htWs7uoWVYZPGpABdqsWV1a/ryvSHCrU9//wZ2cN4/bxQoYsbzGnkSbpkQjpeVkl
UsdM/YN3Eem5NQ6fgzbwUp2Tz2Pm8VPY/Wiwfz6HSbFv7V9Wci2WZa4nbbP1cKnu
I0Aw6MkeZ/146Ojx7ff5g4pZO5SZQqM6AIAvkaFpcg4LnQ481xRzMI9yyV9lNbpQ
UwId/YDUyFylqH258uGGCPsAq+IVfFbTfwgp4d4YUZZ/1IdlUZiFyo0e+XSu3yER
vwV8aDSfy9oBJjTQV3Qec3OqzcC/vSjWf9hyMiETqnqmTrp8vJgXBgeWXFmTz/He
VJMivlU6fLOTfxf7AyjXvEQV+rFInZ05UJvQdv24ce7d9aQDH2E4WXAZh+aeTDW9
XTd0tHIHlP626/MHAoJCxwJ3LXtESIvPkfYeCIpFUyh0Oce0+3pf1riqg94U+MKD
iEVeVyoX8z9OSbEDBvSJBNf6kgzOn3RhPLtknSXQCMQz5pKKflAcMNLNlQZ9GrdK
vbfCN2CbCAEqgx80KGUMYfehd1kshGMPbFLoo1ME1LfTRlIT/Y4ShhVbXtk3o3Ln
j9g2foxRXMOO5eOwJ/HUTzm0U4veCko7JfiM5NP4nP6WgKCeaTULOHWI+lDtnJU8
8L24ZI4pPcr5LOhdGP/f36W/Q/vsb9oFYI3fg9Fe3Y6SGmUQuMWRmHDNrjbvI6Ta
prtp0iW+XFZJbHo37R3hOOps10ZYOhgZur30gX3hbiIIebjTJ1aTt6B9QcPs5CoD
qqFBVR6YjpMJQiCmpcygLDh3Rgs84up8PSogXtqB7kmRpouAGaVoJeYthfytqrqL
hsr3oPw3Uz5K3j2NW8tutmmgw6eVPfLW1yLQVpSUtkJkBJzET4uNXusVYqZDSYDp
9aT0bEAHG82x9pdXKzpAE8HuHsssd4vpQ8/vM3U/XFQymYgiUlWdyKKtf8AXgCqN
8apP1RSWyJ/gJ/5v9VMS06P+qn8Mo8JH75XURDLYbwOe3wcL5WyZ3+To24BVXB7H
vmZeVkThlPjWvwRi44/V1/Ed0nsTPxRyZ1/M56NLQ88GKFSZ5+N1pydKIteeobZg
ZUTq162px9gGUjef6nAOy2c2GrG7LAqFasThC4zYx+AtSbH+bdjgXFhCunub+n0i
mkfgiU4J8RvL00FI1W8JnVuWVRdxzBNztb7q6baYeMFLLHosExrr3n8nnxeERgFX
dA04PtE+JpDlNUEnJ6gh3vgVThPXM2GSrVabS9kv9JrW+VIJp6omiIN0+qsac5im
gYmLgMOl8weU7jVkPZOmLrE+hjh3V4lIgE2KErXPz6eeypilIS93evittQd3sE84
69VCk5LJeivTuxbtvjjGYFxPAdrl2dA7c/JVJ68aWQQvTWm0fQ7zQAtmEUIN1LHP
y94reKEUWWXi4kwYEz39rwIroN0IlFsyR0ArrLPXChnrKIBSkaJsvNOtW3wCyww2
k3xY3xbwvpAOXy5kOzanFHgXRaE5fv/ZtESSi5Ko+jzt/k8HcLEoD6auDlFoirjf
c1wjUNexrj1mowtNmMB5nCRbpur5nFTbMP7UVwx/bgLGu81gTIW/qFt/Bk0GoiHh
vCRCAA+EdZBk6z1MEmjHrs42lDv/Wglnfw4dLHSduA12B55a4+uiQd13o/G3Qelo
M0FQ8QV3tngRT+Tzh8O85IgphdRHlUBKDue1tij6V4d4O+ZSQ2WhghmIWkQ3wX6C
iO/2dPLaXy5PMI7WzgQ9fQX/18BFRxbF6z2mxOVfimaeVY8+j4BtmafsEA5wAX3H
6587vjKwP+7BD3Zb4zwhWRf3VjiN+YF+4lefdzOyv694kTW2cufrwJ5qQSV+BfxZ
OQzbrspzeUEB34E0GSwjNRRKRA3kGEft9LafGVPQWPZStVejE9uaxgGp+80es128
H0Taghi/5/bg5lV25od85q7T15Acqno6YCKv9KLi70rURuPaT+1Resmq/b9L83wR
dsA6tYtGMCYwmxjlkDPjHKPf/EKN5zGmfQ0gb/lYWd2q3R5KzhWQUe0Pe0qquOx9
IqJg3RRZH+0opn0vhYEm5bM8IRiIjq0McefNQTs2+XgxglaetFUv/KTQFTBaf6CI
Mwr4ooVkkOwP9psxqCPHrlLA5dVr+NG8SXdn2X25IAUR51oXdWWwWynV4NSqdyOJ
CGG7Wbk0YHInfjqCOX+mFd3tc3oTEuiNUN1J9TxthRQBGKFtkNaVQXCXG7mlxoBX
YOtfQv9QVlDU0r9id68AvypV/BU6hhVaK3sBfRzdn7VAjqQVAocrAiinQzftQkY7
PQiQqVu/IhU8N4Nouk1jmQvBdgnNpCreCLtHEAkKtbDBDmQ1mxZFivE6+H4xL47V
LbDARslafyRz6B+WO2+PuxKp6lEr6bo3XQbhkY62KEiDFKRFD+D4Dqr5pQAcvKaX
fd45LRyDX/r0OnhPFaFLZhOn0EltOdPjZ4tnSAQNh/hLO36LTSIrl629yDFH6NYi
q+JPM8ZeSx+FxQ66J2P3gZbLy1rCKQ06WCG2ZnJ05kWLyWcB+p4jgprFt3Rkk4XT
kz+e4gzsKfbhifpW81AsSSGzQarQOzodvEjyYkmBQIQLiOujLdaZKp8t5+yRq7DM
GQwfvWrPkzX1WnOTw93Bs45wfpLSFKWXuqZ3ckLjBuSi7HeinMc9Y21aCzPuqzwh
Wk6cWQe23rpPTg5wjaxon4fjPykXkGOYbg7itYjjyPMWlrSK11cj8hR8eXs2H1+b
SJvBuX3PYBuDYINYmgAqTUEs8ZJkR1XjKX+60wY7bS+sWaBtBEWi5rd6/Lm2fJw/
RvMTtoC7E3yZX8s07cfGp+WLX+3rwKUHx4MozcqSiuQW2ntApaNiKzASD3Ag3h+r
6j+SVjaz1TE98Q9+LKh8asorM7Oi+zrHvDd+/A3swrAtKSYqukgHcxX/5N3cpmZS
txsTlrqaj9v7C0KJDg6h1HzzNZJrtVcYTwry1CCZJQI408QNm1w3CWsWCiNFgpT9
S/24U/eKnbpFzGMKJ2i+WKbeHU50mFCZ53g+77MB7cduFD7MIDuTe+Xe0RtUh4v5
XS/31XnOzSAyC2h6xuNHMvaAdeaqRIOCowgE4kXhGszFiuCOvW/kX3PSwiQPTPUa
yjSVU2A7iAhzO9CYRqNcqz//E+3vB8miYZ91C53M9zxsocrCsVANywLcsohZfiM7
/E7zxgtLBr3BD9PxH2tP2lu9cbh20qdpB3McBR7hBn2XNGhG1C9xYQIjnarqJmjz
Zq4vKi1EHg//asP7DUaY3sLK+Y+SlPJf6VGhLTjmOYybA+bKImHl9qao/mmdILXi
YpZCSqdQB3L39cjcPBULG6D5NOotQypYI7PPBEfL1BK56UbqrjT6/JZBJ0BHnBzG
1JmKMexYZJ7zKCM3PrAxgLdu0Weob1ezFRDhy9UJiPuqBUaan6nCG/hUan2dG5Je
yjQy1/M/X35FbBYQ9dS5VaAF9Mb4s8az5w/4Y5JhxKANBGrJFHx8pb37w4OAQvCd
obrFrwxyP0ds/GV8RkucGPKOcZnuwRB4Pm63mCOLgXgX+Gq1egrsmWvxaFjmXuGR
wFM+ZTaU/hD4hBkBEI+kKOwyeNC+0eyvq9mIghPOur/Jmq7U5KTl1qwTjzMVKaD2
kXbv7DEhPx8TaFzCD2stXdm/epJiwdbIsIbCKyjxPoLvaGFfzi/o2MirbiilBke5
Ps/hrKd5BeP0JDxbDZ7B7D0XLuRoCSR0SFIzdsCDHw/HvUiGPeWk4HnJmdkYeiFD
myh16WybO1goMzinyq5hK1i3nRo88EhSi22ipd+vNIK1J4mC3C6LpSt4slZpM15t
i2lrVSiA+0jNgj504/mk0NhYfxIEMXUZSNrXGycP9MXv6DCcxQvBgG2Ed4sgMV69
SCESWJ6eIKesDgmB69mwa/jgQP5gQb/W2am2jAIuCrOp8cm0uFnsOl+CAZkUROeA
2iJqTJCWD7M5/l3XhhC//BnY0PIqwomkkeHHfc/B7PlOLBv1ogVQddAftdOjcvEl
oz2fE8lxOBTA9Hw5fPYfmLlRa9Ciecb4WwZfoX7ZrAOZq2U7zOzQdex7ucyZ9BuR
ZckiSw7NvdfOrLUJ263nQ1nSu0ZHnmPZv/2kBo8guCzcqZg6R7EikZB6YlDOKDLf
M5PzZgCfV9htnxK5dy6nOABQqnKj86EoxugS+AKv/SyQTTn6f9lAQLRjBweVBbFq
WSHLPaB8ryN5A925X4Oc+qsnPdQqQG1S01AYHWvgiRM22ixkOeBPd4n+KYAlonCn
l4cN9ecVk20XAT2dfHp3aAKYNXaHLBbc5wG+hC+dIOUs1s1nDEbbDUMeUxsFZFvV
OAThtdq+ap/MuDTtfbCes5d/K0MJ2/2Sew17KKl7VkIe+BjTfWESzG62rrkOChC0
uAUOqz2em6TrGsfZu4JnW3EYCVA+1/sZP2b7yyrEpBK0jixceWYj5yCJgsPjXMdV
tYD94FN//S+XtmN34kepub8DHSTqwoSTkvp5W4qAno379VnWlgOFcQ8WPqRAqP3S
KF0edcCh+pZTM5LrZ0h58mGN1JIyTZsOSnNwV91b1KH0JOua6Ljsb4ecP3B8GPCD
KPoWWijz3udBZWcmxiyJl2htp3IEx1eHoXnpfkGyxaxLt88Q62zrB6HNWfrJ2o0c
lo+wGxzIb2TuT0dFjWc07XJA82B3HQwIVi6Vkx77ueeqvZGm3M2mK1DzUufVY0+T
AtO4Cs8V1E+zpIQurfmYP6wK6jTSuioZdzq5grdVF44ORFbAaVCm5q/wtsiTuzjB
2W0UOHuvgiHZHEmVp99xsLoEo3I7gcN+CJXoV2HIcalk2PHu41DPcMure45X/ya9
h1unNhvPsg47Q7bXpsx0wv01MrjO+yQ4l4YUXglBZcqqqiK+3Anw+3AfenPNwwq4
bafZhznrJ81oo2c3mSevmFMZl5/vH4jU+1iPxR0GSWrr53oJigGQedh9ESPLQqgE
tIJezVdwMybUXZM4EcWwLnjqjifELLGY4mYgtytMrb4MP2Lo+M69qjO5vzyFguX7
l2LBtI41VisfAWBa+I0zboKEu/C9lF50+jbQhVc87/81CmzGklSr5WgRLnCb32KL
JtUM4KmHea1qXXIl9vS4W+HLaSsphGOW53rLLafpeCy8NMlTz1UaYceH+1ghRETD
TcQg2FPwKSLnkQ4CAWZ/5cS1cgpmFjoYHjBK0DCiPsHmR4tFm3jXTSFyI/tUaZT7
9pDKpjbRsma58AtnTGS7nbo7EYLC2xDf73REwceIQ17jkq0Fq/iVHNb4kE3bxzot
6UFGRsdfXL6EuY+iV+zxWZIu7V4DuBfFO+oBXMgQCdyJIemm5boEsgbCGiPaqUKK
vBzIl+lyJTxfyGL7x/CnhvPgU4Rk0PS2IT8n2wX/44YryBx35vlVEO0R7WE3LPpm
+co5n2gBQ94MF50WMAG3yACDM18ogxkOZdSKjaoIfbhVjaeFFIo9GSMbA4vkEaTF
1IvAyBBXAY9Bhwbt/6V2LBWmtMV/7uWvnAeK8inUN+nOUrd7SogSkydJH/NYiWZ/
i2itWyXWYbuqSURTNCDnKGzYQbz2C4NTatOO3g3EWr7aVA9ofd97wJkJ85Mve3xO
qmTZQMwi/ueH7GpWnCPfgx/LJyglB6IEUsAJjbo0Zz7xd2d+MWelfWV4NRn6xyoj
NDI5JBR1F9+1CCON10TpxWrEf4drzMZE1WKaBZjCDsQcynFgR9resTWN5ZQDjHJB
x+IE8YXITym+GSICDmAF5PCQiyWmRPuVsdnXUrpMUBlW8iJcPTLUu3VluXjX7XEm
c8z7rWE53SZ8/0tCwp0ZLpjktUSod9fwObMdxv1hvugj491G1jD9PLyqtMvg5BKO
bNzaJDphC9li6tGGT2pp1wSNPJPEkr5L25h8hDoGtHAlCvMJaUGnwRxqnrXCe1Op
SEd51ep/D2HAqGhscgbZyUUdXKfhOOge+lLvSirSqwnSkW5mFlyk/0xT1ASrpjIk
jiyk7XjWWYUS1YcgbZnjZwAtRc2suzhKgrFyzoAAgYAoMBj3u/C9rKCbABXQRNSp
yfoTWohYnyZpTuyE/kGMeOLVGrMckBPwddddPXfvWKCbPLyW/mQPmgf/8qKGC1on
/Oc6Qjzjw9WZE4DgKMsMA01tmoVu2bih8IuBv1b2A+96iW/yeIXoCU3cpqMWvDKf
fxq06iED4qOi4KB5RQsS5aBV/LK5t0diwEWmkmLHHk1tkd1bKJw+w2pVrdNuiQ3K
OjC2S9m7H0bKmdiowXqzfrq3jjY3/W182nMDE0qJ2L10VZTU2neEP+mDb3cc4F2p
G3MqbpFN8R1PkC1s5j8dNlyQ04OtNNGRktdaXAsZqrbty1eSccD8IwDuouzlccCr
QC0SgPykI21xNpH2sezJEGw6ISYl2p/uztu/mm2fzUb5qRfLGTtdX5D5P7j5Z39X
iLn7EQORATDwbQZxhezU8EtVbqJpVDU9/uCgZQIutaKl99EqezbxcZX72EeUQQa8
+R/GJQTj/wWPpefZNDE0k/L08z4XLnPYeWiERdztaR69B+aDqZYhsJoHOKTxDsAx
KWxzio94wVGw+HE3PJSB4kd+Y70OGttrfU15JQQt9cLt1GlWhgFc6psCM2FN0+E6
Zart0imIylq9g8/Nc1p6KgAuv9tEKT0qB2sWBzoFi8cMHOKfqrBFbNJK8IIAWPNR
0Y6xuMEynKKzsy6TJyzKJpmCJOL8PMQIFbZn6/KLCXy0dpiEPN7pD1PYZYcp/Cty
Zyh+5G4k5pHO+zFut+xAFinhjkJA/4W8aDYOHW2Q1bYSqPN0sFG9dxGUMF9FogTg
W/Qh7vYlWf6UvtIUbc+4BTjnUJrC2p5EQYlsx3Doc1tArDzmkeZo9/IY3dyBOiS6
Xy+s7N/MLcULR6YYUxQdtTfzD7OVYf9U5cOeOH+iwkbH6ssXyOACDhK/uiiP9SZK
asQKfAQ8FiOPMx00x02XncDHhiAQ+6TLTVSkQR94oTqhgZJnq1pdYzV1cK49r3Z3
/Gele23XHcpRjL3M2QQCsA0z0YSwQaCb7ujVih0Yt/NIESrXym4qNDs5R73p1g2n
wjvpdrhLR2vMDGFxdJ7tJDHk9SmcDXR15TRpC+p00prqcr2obu7TEWMEhtkcFPgl
GjCbTInaALb+IDxejw7NpGG3Hby4Xec1RFzYfqazBVE2sKLC9jrGlgXnvEA8E8X7
D6KdBchKPOG03XcdUr1O6sgETT72TFyRGT8bpALNubDFLlRKPnJQPKh2ShW3J4kU
unTs5CbXcGtEcdQDyXWZEEy4e+0tcwsbKE9sUaFBqdsVzZSeXAWB6/Y1GqlIGHIo
kgFJkE1AG72RM0yAvU6Lz1yhYEMopi33utza60AVwo3UvCjM07ypHEJx8hBeHRD6
lg+z7ayir0pFNOlJQTHCMRQ7e77LxIn24bqL5KkESzchxqmLxe0SQfhY0cr4J6BL
dVBFFP9thqLnJePgHsHIBUdBi4eXSADT4Wwwr9gMQN20LZbkAdGtQIYzITNn6rDy
ftq8+7GoGLA80V5d/z0biUDYKs0RGcYIF6Zqoy0NgdSmW8ar2zbxn2Y6gLv2y4cL
/GuZ/VkTqEiSxpz8/Bj7Ld12fhu6oEUIAcFF3k3auuT853k5Ufg1evP+U8NTZWuL
/E5aIiVX8Wlovu1EUjCF1YGfhP1vGbySXgiqCGArDVOD1lHaPQjboc0aCwK8ZeuE
Z0bYuFqy2zfPZ0SBPsklLSXDZBv2k86ATOVlTgBVGx3IJsEeZuPP9NxpnLG2jg/9
WUMvF6vx01Hw2bN5RYhaztg8XuaA4g91KDfsaq1lnlBmDgYhW9kXP8H5sZ9vVC5a
fY7DindIoLpRPx0Ij+J/woBbQ+ecRgAbCEBnAq47UxirqnLYbp6lpPVTwrIOQVep
TAA8BvXkw1XnVxepSqxm48jBZrOZTmQztE2O/CF9zrOnbSZcaG552sDbLpnFV96i
2MjVryBX0hJ3XSAr/e7JJdpL7vzSolKLH8eyD1Pt4Y0pI6ny/tAAGbjOQojl/ifk
dX8bLz86wZuFr77rx9o0fvNS3UF2M2BExSVwujajkhjLW0yPdlPkY0my2OmgbCsl
eBTQWkVGmvO6NG2tXwilCeIJ0dGd++oGAJrsl+Q99qCwM2T8n6q+UZTg5v/8O/6r
VwzrbsKnP/jwxVDf9QJgm4w6dcRlDq2VxBvVK4fa0kvqCvCZXKePi9DX5M1yWH7N
h3ty3m15FwO/AKystnnd/CtRrILaAJdX535NZLaZ43euzkQDxNAGDG78zS0c0jqZ
PNwRUpCfrPwuHfnj5I0U6kKlk6MX6s6nss0B8CFPCXyTqRU0mN4igb7mvAiTXR3k
ufUdhQRuSc0tu51vfdiDc1QjM8/nB33t8xU6y8XyXjsAeJ68R5BnYRE/EFEA37IP
gKoYi4YNWwQLZ4jOWmUhbV2+Jwhuo6HiLWFSAYoDvlwuqyh4daHKIrR18rLa6ojb
Aa+m5qXEqK1vqzCfK27DWL5QauDuvHNDXuk0CJjeD1R8VcUExbvU4PF47cgMbrI4
fIjAPuFf+tmL3UTglDsFSW4GCSWLPuJrEBaP3jt8l2TejEBnsFeR74GKIwRa2BaC
NivezikUyI0oqQ6PlgYX28/C3J2mG2czEX41y4SP1ecD0B2T2lxJnaE61IcDqQC6
8rKcJlsje7Cc+j7Y/xB6lHRm78dRbefMFJJgJdDEj7WfR2E0DMEnIz+XL2dlp59f
9XIVbrS1b2TJKCprX0lrthyxKPy4XX4n+1hEzrslJAI8c5StKylb+FT0qOAqSZo3
JrxzxbsfadY2BaS9K3i8WfLTtZ4jUYJA4K7NuWqEUNWgSnRbhftOog80JU6xD1D7
0vU/KD0ff5+zUKbsF+MH0lgkNsdPr1Qmk3StGz9Gqs+kUWazT3sAfC4NUJCm0IyW
HBClgS8trLfzNi2qpX5yZj8T+5YJZ/D6mNdDu9Q7jaeMDv2zW/HUuUqRQeh1+asA
ohFxoQZngPs9r+YCt83kS7hFQujuZAvUWsw/bGfTZvNPj0FLZLtHl1Ms10M4icVl
NOWOW9lX+Th0wbPgd+JOGDhbnSh0f190g74xuTjDYXChxLHBD6yJpzVeJ+0XJz8h
8h237+8FWtseNoqkZ3NEXlwt3w9VWjw6Fr0xH3TfCObuQVRBQbex/OgrgG3nqRoh
nm9uoSw4GKIkxW1xhouymShXRo/Ci3GNlRCerSXq8pKlcEeGRTO+MW3JZWPVQ6Sq
UoD/GZ0+dRUI9zxQO7+Uyi42qQ+mXuxptes6v69AE30PMbk5ov18NlKyfOHMM/wf
jXf4KPm0YOZC+00Kk3KWjMMiI/o5626XjbLEixFAKKWm9CiFg6qbwjxLfq8VwoES
siu50P86vYbMjjGpOHmktabv79/x7J71OU/hnpHbAlAQnDEhoBNAyax6JoQ7pTB7
zxk4PnVMYKfC3Mvf3OnHZuPDVUgT48JMCE21BdQHQq2DnGfPA+D6xEZoAHDoTIW/
ueR/dt2NwAsisgEj1h6hEDJWZ8ygqg1OLlFTwdkpQKY8F5zgGfBFpqK5lNrUTOmk
IVyQDUq6+ztJyuQs4ZYlJtGjdk/ZKnsKim5OsrsUakFGoQ8HJEhqqy7nBYJIte79
4tSw33oCjvUql+AXFe7UnOF8Aor/kUm1p80AMKsqM4tYZGgaG6TQ+nhfzHhKWqeh
/XZJKh4aWJUT4RYFlxyJPRqLIcozKdPLXlpwGuZr4VUxZU6YudPzG/bJETv1qQyq
/eZkaJ750E2FyEEnnD4NFoWpbUZQkR1j8Y17tYUNFBRifRQzX0zCBVoMuK0mv7Fj
RXXJZxfAGrNJJ5x4uOk24uB132xX/+gN7pJoQ7v/Al9cf4Gr9imkNL/ljTDHtf/u
KKiHzNuo/Mc29smK9OVEeKuwOc12aJCN7xSYUCCToZiPWMhM3x2iY7nMMyW5RJ07
TcKqwzmG7ruCPshuPA7uJIqR/cfnPXlvZwOnptEA4NRiwhPskjfK44bjsYRHmG3A
K0N5m2KVGX2DWTHkrfO2JY6kDAP5SsQFtRFO9d4D/GhnJxK0z5hM4BikUYMevSjz
B/euv6tDr0rg067j0KsxgV2CbUdsmMDEFcdolcUtfR7rNdcwUgGYNmOIisE9wl//
J9rhsSUaPaZ9LCOLmY5ZB61xgC4td3nXOAR/T/Xw45954cwBV/eN2Yr4KD2x4IE1
qZTovOZF0D62XZh58S5zSSO4nZs+H0poYhTvNpRLIbQOINVQlLlbjmCyvVJJS0ld
xBtmx3M4AyjJ4MOU9yRZX1SWWEuVhWznyhknGHUVcOIAi9hvd9njsqdXC8EKEGs0
K55zKUrNlJP2n5t1EL559WQjJuBBnMp+35UGov7WGjuIZwKElL36RhxffRz2QPJW
rP6QFlXBKsGGayCQeUXJrMjblaVsyOJGl1XK6xM5XkAneImkjrG4WNrCV+bJ7VAm
EyxZzUYfc53MzUiYoHK+G4Z0F593JpBGo+OpfmeMll/13Jv6YiSbeiiHee9MZz2Q
8+sLWf9ZYmnqi5OXvyBqSXVWnQMvNBR4AQxtfueH46jFyDITbZywkCERognRdzMk
3z9fNXpaIm6Y3XeLajdI62ODCONUvdEQBSew1hwbwJefPElLhJBoZbmvIGo2KT3O
GbrGN/qaqLCYQJQwqOtaXyyPq67FLW34nR4/qVI0FftJCEWqmqbn8yZP/4jIiEUa
yT7KZCxyn/cWaAaAMgHVjn3jx2IxmPMl6d3Z1936Sa4vmzKbuaK0uWckJAGfy7Fi
nlwiuRnFfp8MNXS7ukZGqw3SHNvEgF+UvqyXzTcsBObQkp+/dnuV+lQsjRBoOU0f
Zjz5xsQg1a2jUQEgNimp8Y+9+pBWI7qF+mDFY5NZkRXWsS4g9QyYukVRHVVSYrUR
qQctqj0c+vdb0zXvMFedORS4pLfUojvTzb3j1TDwehnpB1eOYN4Fn4yXqvm2UJSX
Ik+NpTIfX00V2DKVRwr8xS++eEXprNVGhRbvwdgKLFiXiPfUK7xyrSwp3MfgPgiD
BJpRQTJR2RRbX9hL+gyFWBACBDv1rm4iGskvAR3AmsNIWI9UoK5kF4uKet/7bt7e
aMHK7wxq9OVqvM96vFONdlsRU3yBbdZWdd1C1t53jMeO9iokmWkM+cwZTW+xu5om
TdW4RX2vryv6tRB3BJNygt/TYizgY+oM+6J8Xs3eCcPC8k+FFmu+pSJqcQ0MBUN3
ncfFoCV6WT1I6Ch07cQJlj6hPj1tR394nWHXhu3TJF/7JZPfJQS0u71V2DFYCH0z
ypC97mFCi7mA6o6JwTTEerGrKg87ZWYdHubqk/PsRpZ6mYh4qVQ8tOWAkX1Xyv6n
DYI+34t1ElK1SD9SOQc/H3wNrO/ZIsZSlbxuZ3ctwIp7lUDA+2O0Vre5vBDBkIcA
ETBzKX6U9q+Y8z31kfrsKgs7rInHsa7+4ma3ZewrGDc2+dR68DTQK+X/7ogOBE/3
ps0JJLY3rwT2UZ+Pt1Jl7cT9oKqjbJfphY5U1sQx4dD5FDbPh0FYdl7mN5Iaor7W
PIRl27CgNvsp8zkqNE+fpE0uaHQ8VLZhi78xUu4/Xx0SLgXn1+6B1xMjUNN2HI+C
+a28mah3p9BL0zc/QW7fgPuah+HSi7HqXzk/vVo2r0pkA59x3217l/7MgWBsw+Bj
DE59dURI77lW8yOuv0wBhCWY6naPAClsQBw1AdlrmonvkiKKtbk602rCZVaWCjl5
3ihuYpmQa2xuSQtERiprsFJXQhTlMAZ+2MTWLsIq9Mgvns93P1UWpnD8Oj2kN8bf
pRvU7qmOxcdrug0oowtKlhZnpirGW4IGeBLtuJ+isCuHUpiq1rFVOEE/b933or2D
j5pMG9zK4LA2VTCyFGc/MrFWcBJU7/tIJWMIQCxfnjFPY9aKQA8nzpPc+6g4UXZZ
iNU7kICWncAt9PDgwaV5xg5x/W2ZxwbFuInJFNnz4HAfJB/VMC2Gnk3wqmdnLu3N
YcpWohWZQCSU9vWNDg/zwEeeGNsDTbpvVCnnBrue//UxqAmoeq992nyl3xjEE/8u
li6bpT9ZIBiyEVv4HmCcm9XWEz6qoMGO2jyk2OnRQHPZg0hBy35Mjr5yH8W6A0Gt
1D2wp+Ku7Xh/QV6yPfFFWxYo8J+qiWipssOP22O/QUu0YAWW0UhqmnmUSinUoOdt
anghbmXdFwvYT8R+4lA1IFplEzGF/CNlp9IcoMf61stT9Kqy3VWc4SSVEr710l59
0O2NJzHX7d0Adx2CVXkrWwX+v+RAiU6F8w+hndM7SqbfIvJRL/iB5M+2Y9Kv2eAj
jFpdrvOOiOhAUJWh3TF7ZQRKixHA2o0F0nf4AsANsO+u5iJ80uPT+aOirUPZlVsO
VklM+M4YyIHfSSbGdeGXXHFX+gLbn4z8ad3w+9bP64IqfLidXvpA+wI2UJNHccyr
eiyEgotcdvP53ioE4EHR+XBz2GogEBkNxTA2mcRu6SA/uvKajSG1GrBil8HN0JGx
O7EcZ54Fa55xxprB2038d4NG2dckPY2ZfzPNXfplcwYKZYxhgtC/NMAZ6lJR2Eok
SAdMIpkPw/luQBCirTLMS1CYpXuWH4XPx0qe9+YYE656Bj5jlS/70Txy97y89SXy
hlkeG+y3J2Uerco+GuiQKyHHwSzVX2115veDND/0Eo49Xo31hkTkLE0o2aM2M85/
m29A15V8gfvaErzoaaaHweN1ALqAeSQ862JtMLXb7Exb9vKhcWGHIZsix39DO+kA
Mm460kFyCg4hzgCogGxtqPM/owbIJZHeGIPLwFovtSIWl+BuIlqPE4I2LnbkMexw
qga7QeASm4YmHhqo1ULjgsVRAilyqn3O8wJz94WECMZDB6lNgQCO1mu82WxDP7aM
JOc1cqnQcj+7OELpbc9Ezpd8ZBPziBj5/X4QWG7ujD5I4Srh713dT4SFu/3lXK/K
Ja7wDypfE/FrxF9C3vvAjMkt4sUjhhDDIOhcAkxX2dUcyExFqo5Zm61GkF58fyfs
ZZ5KXJMpjU8a7VVNYUJ28HnDKgyKMJGlYBy4Th/Ii64rHkKI2DBKSZAcJucdnx7n
3qUpENqIdufhLhjUcjntPsDbN65OTxlw6cdz1HiEaT2tmdGWZv87zWF6QL9HH814
zrNyMaXTj976MS+A0tHPQ5ajOXlcy7UrtRAd2ESOz4r7+o1d02uco4YhTsfL/Zmx
QDub8TPEvbvULMCQPcUeyZ1DcUEEkWPDMKCNJ378dV68TlnAIfDr6rXWIgo5vx4N
sJjD1fvw6RyRjp1lmDpBr/GkpLXYe0OmXhcwyPL39mKpE/G1a9GHKfIAhYZRmgg8
gUEWgjRBGgWaZh3G13wN4woPfQNxwtLd0ivQEXkO8wSVes1gpDDHsMfk/ttbyn05
Y3WwDsmgHvzHeWXnjhKpvH3Hjhm9E48QGn/eALbWC5ZT7Ppf+Tt2N8F35k9+DYtV
pxJTGcn8zURgeBslnJLBYHgqFGibJ4kRp6G2OxP/Otb2kKnOnix3VTnz1cBeE+Rr
jt+8ZBrzIIOiIAGk8b3HngBa7FqrgHKNvo71zhZWAdlz7jUA6/JB0x5NzInZd9tz
pkDBLXa6wtZlIyOnoKPpL+cMG6++dVxXwrSuM4j9Wap8ZdWNusQlq7nht9mQZ+gu
vERHGk1mUTJj+zBcajF5FRM0MEGg+guAN4w/Xaob5aMj7yNJC7gTneLVRsdyM6IO
gHY/awTUoI5AvWgkHEGwhDnNzQ2CDm/wPw1gBfPL1IUKYyUcgq67LcZSzUA4Jy26
limNXBXVEWZjyJCwf1embn9hHBVfNUn7Qq3eCe213V7ZQh/TMfoShBPP0HK3FqM/
vQRzwwxxEHSBv5Su7n4yZ0wTUtNkkSEBWV4Sl6wowcZYI+iLfrakcH4GI/2ZoES8
NWCm4cRCJiJWKa9ZujanKLou0CCgZF67E9INVJznfCbXLI1UvIqo+ReCucmw0Hlr
ndWZ7VckAvIL8Mo+4X8l3NEUvFBTFacAg5ryUoXjYgoFXjTYFFU3ozWeXitDgQq/
35XUkocaZwUmUP5H33UeLOHjgNdJ3u2qOsuHKd3YqeVqmoiwKcYb1CjGu7xrXYfd
G13MR/PFTxjGUPgor8tbmNgZwPSnD17wK6LxfFVlKZI+F1iIlx2seukHRXBmVvFz
MgIHc3JHW6UYJAt0bhJhC9GrNZVcHLIDgwmUsjUw/3FR31tfFpCd7wVCLrsDsHYY
5bL4cXNAOU5JA2RQk5fyRdnzAF0C7vUFszwexGVPJ7uJBSMXcmuU3zh5pft/EjLr
XTrOMaj+veBbKnqPatc3NjKGt9MAYBj9xRb1UoRzgEnvtvpU0q7G2WZ5aaiUMb2G
EnnvcrhlXacH9cgmF5YsQYKK2vVFG9pRNlNZRL19lA7hA4ykQ1c/hgEk9WddYZHb
ayJWim81gaqlF+mQ5Hgmxt5lzqbe5KI36UM4tLK7s4GmuBNxlU7nNMRAz4GdpXmx
WlFMn0JqOR3JxFPYS06aIO8NK3ia+lUCtcLfNeSpBGlxQJiUFVmTvWmMOBKken7H
AaGwVbA90Dmfy0lGJR3RmLw6dVFtIjxCmEEYON5NZwB0vXpPTAc3f+MQwOtoJnDI
la2ReoBhvuCN5R/4NHiTjvp0zizQPDZayZgAr62u1lKtTIm60FAMWRXnXor+N92M
hEldBoNrKvJ5iPr5PUgQU81gbte/OIS9yvpIygyZ+dTgtCOAYsTl3QQfYCGn7gWf
uEC/Zl/Vps4Im+JUswrWmbc0qm6QRmtt22gZZ7ipYJ+JQT7tcesKd9N47dpTn5sA
WruGtVI6NJcPzduP568oEWBRHWHtuWJhaIFrQA5Fflvum7J5GXtIgKbcGNWGJnTO
7HevYNpi5JCaCaqd+eqYkQOWxbbJGtxEgTbVkytKxhlf0uOlZUQuI8ypPT2faZl5
UhdG/gGgRUmbBq99TA1GP21qE7oLCkkmU53s5vvt/voDj/cTBL1Lng8FwHb+4kPd
RSMIH56Ylqm41Hy7iIJQFMAp9b0CZZLLMPPA9N+ZDVGOLyi4IxpnTrl0gsZbMAeM
iu4uoBmRde8vnW3QMsFz0xhd2lym3BKyH29y0AMpUpfebKWzc5Tef+ZFRV7Ezwk7
2LPsSmAN3+ylKzkuef6cLBgxZYXvoGAz0aJ0UUVWps9lBdj9zQtChTj2ImrjiIGL
yK9GTkQwUNLDb/0TUfZc/rtvq3UzHVhCCX7W+DLka01kLvP6mV+HBxF8jNSCTeGf
6nzcIz/N4pTxHEs5JUhz6/zzXoPJkB20oxiV+I8mcpKO26LRpbd0njy3iIlWcdj5
uZldJDqQV1hW8ogat+uKwuuJYekOt+RZe3e+9CBh/R+9n2IHUnUzfrAa4X25Tgav
kqdCTg/uR+SpvpbUI1Zwa7jwwHSeZSyF9TtY273VmS+wi8Ko6i2pUcG+9MhmpoWG
oK5AUZB+xOj8Pa8FLF3vWAc94d9TrQotpUX48imCYnmXL4nRKXMWU/DnbvIOgknn
Lzl9RtQiDqaYXLCQkrD02u85/G9H+QVHdgx4lngmrAH6WBVEasGCBu0rI6eKtovh
wduU4SmpjpNz4Jl1TZ8BbXY6/cNTzQ+e8Hgcro7SAjxIavUVhnTQVnQHPaIgabEF
bQjwlsJD73xvI9sPKuJK2ISgv/Rc3mF0dI7l+yWRRbibGkjoexd90CdZPgzNxpIx
rIc2jmbk2khmcBM+h5ryZlc9WhPyjb1ObxOdHSXTPRHgwei/XVI9T0yBoJs/0JFS
plsEWGlmNHa7OhSSIWhzGZOn1QEMbTyBL2xPrVHty8BC3RYd9FrSWv2mylscGPvm
8vQq/J88mxBip83qrtQvNUZNalgprFMWV7otbpWBvMVPnqyaaDRZjUy7iLkjxpA8
Zx/2fhGuz/ZAPO4kLCY3ONA8nw/F51aEcc+yfE9FqWaYK99KYFcCu57vdyt4E0cy
XQwp+hymLC6lap/iGxuFljfeTtRN5wpSTbChLWUbSlRUHpo4KTqJRaTTvjse28YA
xcbgmRUZxW/jAZPVt/xFYYUnyqAOnVsr27gE/BZoRZM4qx+ifbL+R51jQv70i6By
jvePfrPhhCvxcGr8swaKnUsT0Dw3VMx8G9ef8PEK2V+yetnBsql7kO+rFxeUVcNT
gG+MuGFgOqMSeyCPgEyw/mLLfpUYdR6eT+hADJ0W242MPxjCdwkAuFCvfzWMqMOs
lFD2zwGL2VO5HGNW3zcMxcD4jWAxWImsIJk3Ol5Bl8cZa1mlv+JtTNHBHJ8b2akv
i+qVs1BmFWjLhZfqcsKC0iENkOoCDuNoBxM3RjZ21rKVC/zxBURwXi7uX7jDV9Gq
A4S1n6kOdldgPsxYQcrwk9w8Ivl/NF9LAAUVqC/bryfoqo4xDHSd++Vzte7Iptuz
ITaGrPZPiQnvfHUJXkI7QIHECz2haIBXzzm1YoncuwPmWm01Wtf35ka7MQHYsBZb
m09gPUIFexCXx6VNag6z5pWWRiD4S002MzUXn6Adrx3jsYpZxOuVpwU1W0NfXZ+Z
o3XLarYTqS4Q52rXpK8hnxSGr5sNq37IxCmhigZn2m8KZ1kBNRAbSDEqxAoxKD7w
0/PWIwMbCuz8MXenIVcuvsUz0sKKC8SImwzz+2U+qG8DW77o7XFKcYyRTSj2KbkL
fFvQtyT2qP3ZlRTzu352v54SGnxco2bpkB74vusElpU4KPM9PpjFLTEZEu4VMf2D
IgbuoUCYbLf4sX1WCBcmhAI4kSt92K7QEPZ9fFwQME9tjambJlE4RVw8JZcujdLE
ZkLdoOtll9M0CaRxuTEq12t2H3m6elaKDE+N1gQEuVb9+QNPOdUzsqT3OIa0Thkj
7e9EYCfcVEHIUvQyj7m5fS0foZ2THJ2BV9v0VHZ4OMpBYE6etOU+rlBJQnmywpkp
BNXCsFvtKnMXiz3H0zPOJsp73KPWnTRPwsL5sZhDGAShOpi9HxG7MRcXvtLRLFU9
HX9/gbsn2Xne5IAC/U8UQNbGIg0BTBAXkqYOE5nBAoNKQKieCMN1m7+z5iHrMZ+G
tVRIhTbZ5mjNf/wMVbAHWnpfDJXkCR+2L9nyjf5WGNLQR+UEV7N/ssRiqMkr9P9S
4+cnKjUYsUXF2B52RYJlceWmTsNkv+ZposH1KYiyXBgpAnhzwjPoegHeYNiKdCpC
cNdcLohbMVvVYlt4AZjHUZWfr6CtBfzwksBMHkgyxvCCOklqLqU71y7CCkvAA0WK
dZz7Qot7D361FLJe/QXDJe732Dnpby4FecV2xco+Xcex9HIyqdI69XyUurz1uEFY
fUb0zH2RUGWY1CXTNWGFfv64YjAIs1q/gXgoSY7li9cuV/7Ef1AhflX2Ex3znLTx
szc0iunhPOor04AioODdYZN/X1g1pKSqoDxg5/RefAyqLv7TjREaByC76XtaNRFI
5szlxdlUb7g25hM8cIHRy4mDMPZjjvVqFPmyAkhfA6mXSazQq7As/xJua3TR5iYD
vOEX6I1Dm+ie9SbzDP+IthnVAll6Bl9LX4Fz7TtQ/0snoxaintfuCFEwLG1Xi/L1
esjbzEOVdeKuI/qgCof+Jwdf25dNZ0lvQUNIPqbm3kGrhmyhaW+3+7qjpCl07RZH
JUoiY5dHaHz8Q5KF4KzAlv0jncNk/zr7XS+1hVEsBsc+fJPqSZGQDnlNb3TiVLu+
86dZE5S8YGqc8Du+eyLLyA8zka1nabYbCq0g0dHpc09ahOgmVRyTIarrUC7UexNl
hADcKAKrdGYQow86nv+uk7iwm4ur+Zp0+IUV/4HL2K8x4JEDtQdcy0VUGiSeQRGt
3WaX4kndcx6yn91wnf06YKM420wYUUc4kxx5i6AsKpIdjF44o2hRRm9A3e+8k/3e
lAINLIrFoNAKksgyBr9HlAowDkTG3lsmRsvE62myy5DGjPsVBB13sFQPJe8/sarh
YhFjjW+D3akDh+QcA2+MWiKPzj5vIVKpNzXnq40aSfVxIV5KBuvXFg/JIU2hPSOl
BCaAhVoNYa8r/rE8LbVlsj/K0hVEUt3RMJF4sEUweBmO5cpYpCrGwsgGqJ4k1+Q+
N1NP39x6NUnJJkFsX2FDwKMmDMKhTlYO6vTtug6LiTcLLvw1A8NpWqOc6Z5iDBQp
lpNOQqlBWJ4TZqBKttqrqCHOL+NXjQ++NRlQ57mJD+fKA7L5DUyR6NDLa7Mys9+H
ljUdx5NVhcZnTXx9/kqULWdiwVrky/moyTGV3RXnXjQKR8uX1XOCWotCX2u58l6X
zCZ8zhV7qcAxzwYViQ2mUkFnyR94aPHVeyfYFZl7aJuWsXxNwhsnDGcqEeF/AGXX
uFYI9iILamDWaHaQTE/1SyclcJbAd8p2e9swZbfz1oj0k0S5t2ar+UruK4uQvQh5
wio7WhojoB1cEC3bdydOVsUg7VVuEky4wp1hBGnLMIxg7CZy5PLhzr5GC295b9qq
zcdc/CI7J0jCthoAhJGfcWn7RFBMIrh9plrymflEzdfAMj6j6oMxjbIOKwR7/V+Y
4Jc6sPEcEv/rYUxtVYNneNUij0Kulva09DFATNmNXp+ENwOTF0AtlsCEDwmrtQfV
IbXDBTBPMKIF/pMVCoxuHgSZ1CgfA7saOCUntzAt3RxJ5Sa+JBlabJhqsyTYNU9g
WBhDpjXeFiN40Fwj5i/x0EojgAiLArgrsC6MzRuxik8xVr8jXHWZCYcv6poZ4Udw
7jCJ7L+bHDrTjPhLEL+B5b6bDH1FOr6AgxY81ASaYjemkonKNjF41vle72leepRl
8MnjUjjorCfuvfRThaefLo0m/Bx+x3etrwpk9zYAWq9dRYxHjGRG8dbIyx6Rj8UQ
5nmSQijfTuuG69lFOxiwMD5yYfMZbWqy6Di53uiSjh7cp6ZdOXU01V4A8SsPOV7l
3zgHD8qhECIPguUXlr1ragr2/YkxEATfxmIoGZeNDbdnH2jLfnPy8IjutGD2dYzk
eVxoXSwaU/hssxaTB0g6TquchlNGKinZWyQr6MO2mOQCtkLjf81R7HNBUvlrnwu2
y6cw9huk9LYWZpOIsYosFem9Fs/RzcocoCoNI4ya0BtVBKVoUjwqDnLB87I/xFyU
inTsf5gnbbCcYFl7gP+vOQXzZ4N4HXMm3H0wnT4xBsaJBziX4RB9Bb3b/OrBDkLt
v7yGsuE1hKaCoxhFFObYjBdmNvb/9px/KV0jQjSaw4ryLQXJZc+cvgsJBYpII4eN
CIa+1EfX35TGpPqddUPfxzYH1D+J4nhhzQ7LU/3ZO5jvqT1/lc9tOKi01Y9hSUCE
3/GdCft9FFpfjWgf9trYtkZx7PjeKRWD3y+f1LkEyUg96DgjU48KVJHPZD49ufyh
pA9FwlufJOkgbbujuldLn7qJndTNnsy7Xb9HJVtlBHh+SbQJ2AhuJuEkp99u+0BC
Xl/rUgBq/JsdX70SaOzQcdtcZrMqXROwRy4BxpDgx8RZN6Y0+64nta78ywbmpUqw
xJhKgnfhwbciqKHDufbiORGN/nxBA9oM76TZ9Xf4ZoInpjkB19sUirNsjex4VziB
6BnkBNhSJ742Sj5K1m0RclVD8ZC8QwrgbWtii4d7D9ye12si9nlKLabj3/RMlYQ9
tFpolBNpDucFUSBGpfrYApA7iJUyqwYPR//y4/5N5eFcrDp+FEzIZRvAlKIW9IbJ
tUY5FZ32pttsdbia/rNi8WLyXUyZxMi627t8BW2O0QUMcesD2jSXQsWuukUK0/0z
9Gq45HlYWKu9ffwnHPjuRooCLYuFXAPWZWCqyuyyLoZhd54i9rEPcl6NW9O47o5T
qwijZ9ZVTyLERKLdljPfbr41scyavWd7InVTvellIiaOlebcs97SK5S9/nFmDe0N
EJukoHV+b2QPv//zstmmEbnLpVExot2peqAISx4wb70IhajMzOVm0drmCTDCZdi0
Zz90qdt6DkQtXFn2pYve289vGzZbLkUUhaz71ZKJj5nIHSQz6+n1GlAs+/Ban9kF
L54mSXAfwLWLnGNgbehY3f1FiehwTLrH5ajxGSLFWK/0+qC3fhHIkf9hbq9/+x8q
FSA2xfN+0u90juocwwf14DvP1IA9ZkuphsDPIU03W8weV4iHL/EQwKyK8iU11tG3
89eKa5etABVq16RKRwnz/RbSceRtzV3WFRFDrTbufzQ/nfjcTHOn7sU+51RWPQEr
ZfoFIXWk1KBsan9/uqP3S4QqQNHv+jIOZO4aECLEMABqRu+/RoGWo3q+mIHQadzc
a6wLMMLKxRNfOlMccbko2gMY56Vdo2U2hfjXbdkqn3p81dy3uLpwzAbOro511y0J
dWV/1P5hwFtysQ8NugHJjC4dlhpCfkhkGHnfML64lnfLVsPpYunMO8sqVvh2kGJU
2YB6+dHnbBh6f4b2J+AykXU7BHPUrKXadjr/Tyn7XDS1Y0ZIk/7Dmx60X4UWEaJX
woGnRVLyfmo4mT6ORfsZXrl/T1ietR2zbVxsTrzzrH4n4UWOY3sTA4Bp0ZQkQMwj
eC3fb/EqeXBOCi0+G8VFUvw5euTaOkX12yPyzFbiiZkaqrZOSCRbwVVFzrHgvikk
osTAKpdYUbmPGj4BtXi5oJhTJj9spOEruczS8wEUzcsmswedjtc16NX876IjIgCQ
bT6JvEN63HV1rYd2cLPIMoXw04BNlRmH1BnEXpdR3xj3CqKO4/rLwQ0I3NSeejjY
1nRT0qE5OQRl9H5E2w1msvYTlXvxCCSKi736gAvN2+vdBGCsC89+6fCqzVdiQar6
ii/XJjc4IYuyj8u9fk5lPmZj4NasDX3hvy9UkvF2t9wBh/GJkDipqfAZ7qlHK/4v
ZgmVpoYh44YSdfH5dfaI14ULi+pwVMgmuPB+VR7ZiCpEVhU/3kOBJ+T+hKHCCNkQ
yCzP7UrTJdjrC0BByouvDf1rPLvTeZ/jX4R4xo4ec2AO6F1tTkuECGC84rOVrC9W
JqByGJAQI1lTG0YWpx2ef/sagHZuaHrwpaO8m7YaEbQXo+arntYpGnYZejiskiAk
/rZsRmGhz1RFny81CICrZii0AzMcAjGpe/b76HOYYkumAP2eUrP1bmSaGseLHh6P
dmXhBDwqu/dneXWZbIuVkkku4gP0g8W78iuA4yhukfviF9o4zqIg1r1/XM7yLuZL
0eJpCgC6v/N1UXH1idzZOiWkdI40TyZ/P1WCFMSei1GNVyQV5Zzrdi6VFfP6+yie
SPdbIdWw6yydTQ0817aXYZLtjq1eQ4sN+aGqjMkGnC4v94Qz1VZ5keC2LUJMAHie
HUdBFRCe7Wg8rwJFmEmp/kIuK1N8Snri01e/8YRlL1bi54exHC16UmW0bs1RfTIW
kupRQMuWZ8r5Kf7tyVBrVSeg9V0jXnyNVNGepKeA2j2+8Wy8wvIgxL3khazk9RCL
NPBb8FUHLnEpWSHtDOCbM/hlBZVkFExi7rop9RHj1woMgPEV1djsmvcPCR+q2fXA
p+h040IxcJLIPtITqlnEjMXyZTOoJGA+fHj5a2N4I1W+NYOBKYQHdxuwOI5HrJ/q
PzgPHbbzZhgogjsN+UgY09yg+bpV2AYTJSbpg5dyuEj2MAtNHQxNNbUYQtPguCn+
i0Uh4N4L5+Psh/BHnmoUY9WivEpJ9OJQD9EIAjcvNP5DQNdJfJ3dhnNvpFaL+QWt
hQdv0uWUSUqUwJ4aeZ5ZtODvatep4RUMf7ic2nSGPyy9Ub/zEeOT7QSgXcwb/Ifn
/dIFlJe12PKginLCMyc9biJk+MeEIB5LzmXihkIpcDWvdJ3OH3mG4TPXUQgBBr1R
I+V2Xg3V6poZP1cYpLtuTgw0yanJEnrwM+KX9WOLf4VXwKpPuu1iQeK06iUu5o8J
rQp//eOYwX+fZUJ141OPOMKPlYz7di/BTm76GX2MJ/uUNdIt11GvRTmxZpq7pFM8
UM9OiDnrOFuRWJA5HsKnPXXeaZjtgRkBLpoCeV6LUGJjxaxWaYqU+zqJwnY/5MPr
r/W0EKR9ZAexUUJF6fg4vix57mWSRnYvEpM32pNp7161YXD2zh3H8lpJt8mrMZTf
mLwzZqDY0D0XHzLYfxfl/A4FSXxC4n4NKPJgSXwicsgEDPBxyyAJI8oQ8Zu04lOu
UofDuc+M3BUPuA2b4Ara3U9X5rE+pPVl5w/FvPH+5kJ4X7YfXNS6NrRdf2/NplvR
9h/nm//w3tlBPrZUPWBp71U40rUUy74UHMUA4AxYKMALHlyvAUWZds43bwkTOxJj
JDRNanvPGlCcrxUQ4lS6HHM5NW64+++bmIWgAJBoOBZe5r7ZQkz5AYF7lOGljS5G
5ruoIYA5VRhGRFnN6NSAP+eUFC8QOK9ao3oYyRPpOM+aCnzRDUVhsu7AvIJVKBD6
ZEg9G26jEWRJrr99uUroxMy28XNHnZjI1tUzLD/9hcL6St5A9czn5BAigmKjrz2U
E76jZiEtxd3fjkZqSz39IVxWKabLOldL4gTEPQ8OmGOdHxtJgVESerf1eFnyfqam
vXBmWfduxbiXos+i/dd08I06QjlbNsMTZ8Enc6iqejcQPCq2XaJyz7bRZpjz06Al
HjE/E/PQPS1a8403pYyYtQ4lfWYZd9SCsyaLMpW32IqFga5S2vQrcLKEXh61QZjb
KLKkMZu1JXI0xefqH3RttBk7gmTolpXH7PFsRJBvISCvOkIohl9vQKnyK32NbWOV
Rec+LgvY4h9JfpELSCcHo8p6l52K0cH3l+Ea90VkJ+lcC1+SQHYeK6UTR8LIeKFX
mO+sJ3CiEnXGyZV77IMOI2/Np92oe49jvBK97evR0PdEbIgPrKCx9GaZ8NICgYyr
tu7LF5cgrNktQwta3gsliweHj4WJO+n+0GlybQYF7fupfJdvGFJCxU4vQIVt0Trt
qqPaM3CLdEO8FHi209ZM0RX0diuqyQTg9AqNwWIqehpSS0PK4uMI7hHnq3v8ppnz
oPIuLO2EmLcLrEfE7r8+Vd2hrocUXsEXmPJToI/O1Yh5dUKpEkUFOaU0lMuPeGHb
/Xa08maAtBVCrtv4M5/eFLBZQKxr2Q+qWtMxxL/aruRInY8aF8iMKrzsBS+/vQsj
GpsoFy580/mXcZ+GD00nVJDBlMjWky3L4URsBrWwdm/eJidBDkYh1IxqwwSQZfpE
QvEPsMsl2Br5Zqlo8lnTl8PIbYcOO+Guz/FBKxXpCRCPlXf3NW7ltzv5puc+1Wvb
rA/SSOaiQ4sfQeoypXWX6z7Knjm5bRQ4EZpr2hYhzBLnLU3Z6E2qxJi24NQHyxE8
CNGocruf63c+jkgMydyrCAxQ3mUruee3W2XhkUHiByviZxNmdR57X3rPxw8ocwZ1
V3dfzjRg1o/v0abwuvmbADdHH/zBjNF0AVEMj8aSgQBsz74n4vfTFHY5CTjClnik
Kb4hE4HEiBW/toIhO8nynUw/NaU9rljkIO3yrlcjaPBiwDRmQsNbIEq/CLAWGMAq
rrmGXK29Y5T53BezakCdW4moHB/EnFLc0a42yvtyupVfTDQnPjKwQn3JZoHEHnfW
NjFrRCnGImLRysLep/Yu4sroV4OPMMQx8xY7tJFjcT58gJDVaC1Q6ovbEQwO8aF/
BAZZ7Jw3KzFSXY7YSg02lr4f4OyZlppynTgQjlIdK89PGUSu0fkyEMRGtrcRRYZz
Kx5RUs2tsD4ar0s0tATkGxSQt1uU/FVrQLQMZaZ6s7uumiF1Qt2bww0dyzsA2Ri5
DwMgX6Q6+48NMHPPWyXwTOjDCiQSJgYh2iuu/uzZM2zNx//Ctgxg9tW8VT/eIL/1
wvrmnRLg4SfGmDZjWeEGjI3P/1v7Rhg9hyODezuHU/HcTMBc+/Mf/SUW+lEgMOl6
E89W0hhqTU/Ay+Xgzwyig/hUj+WY4ncKasHonsghB7TGsgntrte51t7/EYd+bCd2
PJZDjP6lbZuUYbXpRf1nvVUZj2venkG5FOIbSZPMyPH6wqIKpMCQl6avf1CPBsvJ
nD+k2N6mbx6U6m9TNkwAsyvPBJ42jOJXQ34KwJ81Kskdm3lWWUX3/zHYaL087fo1
a5MGJlN/4Rov9I2kMQO8iTqXxnP5lGBzhRE1VdnY2AuM1fCNm2+O3LgBhsXa0b9R
/t7IvnwShH9OWpxRmFTRX/eXazrh3CsbRiwR08XyxhmpQuA3Wl/Z9V3R+DuPpBOL
SdQTe+O9p3NZfJqnuaJa3FTdFyaTk+RCnDX221/Zs635ZU0RxQJ4o9R/fG8tY6sj
xXJdBrslJgKIk3IHqH6K6Q2fFUW6NifbL4bn5oETGhZRbP0/77T3dk2jmUQHVi5Z
Ba9uYmLd6TFnUZ/4tDRWNECa99CZOIQSLffGYovCCU+mBwTNPxQ3cPyCVkYw/oHp
vLHwhGe5DMujoQFUMgB5Ob7PSfXQCV9rik7ou3lsLBtMGMCwI4vBAfsL8ysDopvM
FFxn9P+LEP5OSLgJ9oTNOU6teHzfMHo/4j4QxaMz3eM8Jdy+65p0kMbrXq2ojVTd
Ow4D2OALISg6ubrJTWY0eZrDXg3TmdmiKDzXa7H84L/UVVjkgwfR2KyGaDRBjcmv
3HGCEcvAZs61g2pN1soGZ7tFX/mA15kjzJL0ploNwlOeYc6FHM3DLxrJmVBESsYW
IAt1BFuMVWMTqutmI5/6faYPtqHq/n1j995mar9Q90TnM4H1GhiJ9BpGR3ShToyz
CeVC34sw8lKgM+vTbPGaAIeM8BPZ3j3r5F8/2UaT708foy/bSPdwOPb6hO0s7kbw
qtRHIkF8pOqnNyEmucZnJudhgyagC0xnGPP63eMdxcWqNuIJrqUZLy/Bc3h7yQnm
3yMVjqU/UPBvXbaqe9yXCA5yfp2neQLmigvfZ4iPY7XhKlnbNM4+f3K2kirDPuqR
APR2kSWhWYvchKxjehNwF3jS8/gpWS7DOYPrhOZWbsjN8FNb1PC78sdLLy/svetk
KdA/+QIp0D8XHq98RmgKfcARUU31K/lwgLrW4nFsnT/S/PmCcDI9R0HXz2s60wPe
ZOn1fXgLX57twzWvfadZmT11uYmnpf9mHawpunwmS0FLr6gsl5KvLWkWmOfpH1kf
edCRlwvyJm7NjRzhrYzHqclcuDe61BzfFr3KWOG3RKvbksNrQBNFv6itA6AkYnGV
aP0LYQbqPLjO6AupmaJ7jfz5OCo38fdTzsIVmiikR0RFcIp2ZlcabqqCT6SSMci1
LNYvNM3uNUyYV1XGP3FOy+0xD+c7Fp33ABU21P/qltirzvntyCw+bFwexEOLtBki
PTBcTat4zn96fgCKY/knci+LJuqjSC1XcsOhzOoItOBZIt/Dy3m0iqpLLGCwATta
wGZCTspKh3agm1Nn3tGE38rXkEcTVCha72aubHnwGvoZIOZfWyztr2w5UNDrBcTA
lP6/tUD2y8bAPTCF0R+xz/vRgYe6aBuq1Do6xW6n/FIxluhOQ6iMsDd7xzVdKA6O
C8GXzA4xFrTsIdgNUkN1m0+LstJf+ARqEzw4AeWeteSvEoZqIMCh2l+th80LpeJU
hDi3jujVnD4C1q3f9zAQRjL76kBQUHaMta3jHs07Lvyupg1xOeMZuEJhye4K5eR1
7/N5RXvZ0oEvB7Ti0uaN1267BZUBc676zbrfznSNUru41MiS0CFgX8j9mAQI1Upf
dnbAFCESrWxKvSpb4szurKFDtv/tSXMElJSst02UX5/nI49TmJvv67X7RmBbAMiC
6moTdJFTYb7DLRGfBwpyM07qT1n/UdkIWlviNsi0ZSNyHsqtcdWUaIZHcGB0/cbP
njV4k89L+aTQnljhJCoWICqvNRDpAO9TxD3vvgx0AUSJCPIrZMRJZb4H2NkpPjiD
PcFwSeNJQ74YnGXBUEGU5g6rGh1SQNCJ5V4uD8URDNluP4C7J7MxZcOds1tJjw/Q
I1poufvPTI8iBgqwTaGUgGF+3HLi5+HQecn1VpfMF+FN0bEwuXYCV7woSpVPNZxy
5+daWpNFQHyK1giPCFtZ8f8gN0in/hDWznQ6fKnFX0YHL7wkSUEek/UB3g/WPSGC
iIpjBfWRjEIqHAS5DBU0rdeUJJ4WtTb4A/MbJuUflFVlsOJG7CbHCdRwIODy1tTS
MK0XcUUeZKmy1QNAkAETF29jfWzlGvX3+W7cNFFQCxV4w4GhIwMIY2hHRhnbmcPz
z1EYnGm7QGPR+03qvofgv9/0eKKEwwPIjVxy5KKCrCs4B4FZjl297bpw2BIm5L9h
PYyKuq8w5pSCSqotrReKkedv6+oHRG89R95v7D2T/1sq1h0fKZIXSb1t8adW99Zl
dOwMLD97jVQAsiOC7Ic3RmvqM+iJpxy19On+Y5TeZ5Xx7/SNaJ+auhUDTMf5hlpR
LXVZu030qK3JLk0w6AA1GqlzRN6/DTI6HNhXWB3TbCpsllNXe9xAnHZ3pRLqOBH4
zNPpqbqrjTcCSbeU29vqduD0XOVBSZw0d873jDG5ugrviw5v1uPR/8goIm0c5Kgd
+Kxgh3a+Zgxs2rqqDRfgAlcv1A5YmRKOovQX3x/KGnjIfjG5GjsTaAT7Lyu2NprM
u4EC8ov4V+K1ewN7mt4lTy5+nL5G14duy9nFgYAUBoMFE4z1Vi0GkDb1XQ1nLxdf
8ePRAEuX3uX4MUW9QOss/8FtrIQ3DrbFwKyuk/48rKAXc51aec1DmgXDf1vfHBS6
OaB+ljuBJ4hq/5RIYVNdOVlw3b0JJo2Capk4S+zUF3gg8ef2cF6KfIrQHwGwUSQ6
koLOi1uuYvGiYknOHdjr6K4UrUz6vfAbESedHWNCHJoG/tee3t9Use5YxYvwJ7JD
I2MW9/7VwcEG7uE3YqQTFdVwcCSOAFcxi2kQS3AvudcQ/wujBnX3ns6fBzl2HyS7
1DDp7BTL+769wcfCnGHu5Ex0Dg3pq0QSW22t/ox/bKfzJ4HAjJGYUGOwogEeCLc1
yKEpvEyV4HKj+rVNorZ3C7kI+8fK7G2+TvRKn326nZqYDmjp2R+v3sX1lSOlvtg0
NS8D32vjGCxVX5FwxG/yCaPRrrZtGs6qGAhUosbWdtktCFfLHd0NtwuORhovt5zz
uEy94SSrvErrcRwGXz9fTqPp6F7uaPnaOhS5C8PgrkN2/tt+E/wrjTlOESSRb56G
JySZmBJ+DrfcxXAe2H/p4cl0wbzSINlUVEFooDwxiSppD0FwqtriENIA1dKVq0tR
6yl0BtY9jXP/8nXi6L/+ue6Y835nmhkNsD6cP+9ySlPZIRPTcrwD3pL+yVjPR8A7
pZ0CQsSmIjGIYEnz4PoS5WsCecXr2t6MTjJV8X5Wnpw9zD3Nb0D6y1PPct9UH622
0uFVzv22za7n/1866imOKweKEwgINqRuI9QgKyYSXzdby5DKyIYg5Wwtm0sfUsAu
qt5I0pjL9i6o1ft/QvzJgWucbm41JS3n4fp9l29BN0F1SUCA1gd4KuLdLbdxte8B
56bRaYRevZJ0ApuQDPIVmaKXs8BCuzLeaJSEaiXI284DOjFSbAVrCaToH4PSjLwY
46E4hh9rYPdVbqfCg9+qL9bZm+lWS0We831fLtioVqm5In2iSg3UEnJKDRWTSdkq
l6g9+wCOxG9TI6w199yTr8Zf41pcruvavLkTimH02zhRJsMqInxLgddoyBk35ULA
mL+UYTJS2u5mpcCL1IciJHGEqnKzhaPuCHYqe+6vT14B5GCGOZ66x2uCo9oQDZD2
p8UAwJLAwJba2IeG9XapZlKz19Tjbrj3PDP2+uq6s18tuxvXqgZOpWclDCnuvgTh
Ih9afj+zw98c0P+tcfpAi4y+A/l9Hy5kkr/r+JITPlAjNgnh6vkm+P9YKjuPg62Z
fw87UCrp6VrpKW+c7Z90NTZiNHw1aEeP+3K7Gbq9UQD2QDSR9AbwttAESk2QdW8S
YdKqDOA7W83Vdy0lwaeFiG7sBgBYiLbWu03s7jLqgbjvxYkZ6aDwTgST9OM7IEkN
XT9kTkkipEHs2r1brmhsa4qFQy4zcx49zfaF0QbVCLU4MZ5e2JSDQGJ+koy135yE
fjsn5es6meJRJjByt6PM25baqmrSNrkttWLiDVmygMwx/q2u2wa0VP/MdWKa8W+D
UdvGdMZswEcrUWoKGfV/v5tEu1hR+iCXLWqDYHMxYWDS4MPrM8E7FJVu9GPSZo1r
4pqI+dvA1mjyN0qZjMFBDKjn83ZtVzWbxk+4uPSqxXuWWfLsP/oPB5TWWiBHaG1v
LF+vWGLppyurQcy99lj0FgP/OhIkaAycr2lynXqTFpsOBE3iRUnY8Euaqt4Ai165
ZgAv4cNlhqykyLtAJlGjW/TQJDrJ3OMJ9yWE4y29qrF1pH7oeE/Rn2qk95QexSQc
XfKRXiBCaFWQh0uurzwqL4ng5l0TP6VjlTdiakyAmIcTXiPTy6uZiz+cuvv1Mmip
H2T/6YgQtonUra43NHtevp3pYwrJc4+2GM7GDRwT1mcrhSFTaA8aOov5yNQfbrOI
4ohOx705kf0h2lXq9txpfKwD/VLiulmvUVdCfjhDdKg0cHUfqXwIVKIfgKccD6Uf
oVuHvfs6hKk38a9xE+a8YPAeunnGa1fTmM7iWjkgRsmH8ym6qTkVgT09VguPFN61
c6SuO7qa3c3OUockhaeV9Zxsf7xVmVwbFZunDv7y1iHvK2p/pHej9DkF+Q5JwSd8
j18OUR0MN9WhdnO+E+1myMhAdlt7pH64cksP7UHYmwESXodVqhhNdonrD4SEu9Kr
/0iVnKA/VO9Myh4SxxPpEKYgcw5AgxKvw5KdSSt8RA+tghsctGbCsQwqDLXafx5z
lrX74ql5i41SSC/lhihLe2tLe4wNDmsdJp23ItgXLl7UTd+1XGcD0mrkSgtXMb7p
ARqrO3ZHOlTLZ+QrFPtEZQMx4hIyCpp5v3Ci+GpnqUQRl2l+cisI2WOn6Ltp7jsX
hBN84EguAR9dGi0V6qw6hoxlUK8h6UN9G1IlYqo7Rk1BXRWqgXi4NcSPfsGOzO6i
movI4al/9FKD3OlKGIJ8Jb3+W5Zl/Pa0A0+/FmYsTeljNUWEkbHxMyhfS6I6mAFo
GycxAF/lyeqHTjT6VfeA97Z4GPvj79j6Loj4/xgTnmyy5ulgFt6q/nXDTBv9u6v9
rdYiMrCnj3DQ8SRD+CQE4aTu7m0CtxdNfbB7nZ3sQhpvSu5yzSw/qlN5nu10FXku
B8OFJHMNJY946bPeu3e+9+LRMe0+855Y+bZ1gAqWcKfXVT7+GXuYGpQO9aUXpIE+
6h3yIm+qL/r1XF8DBjmHu6B4t5kjYf+GdF+tkCOfj5DSnkk0PesD8Wop5i5SMbzM
2wyrnvvZMuaxXZb+vD3+tb4hZVvKHg0Rvun1bBOE2tcoug228zwEZ/Cez0h/B5Of
BLVka0jRuJ5/rR0HCLz55qyqARIXKkUTqJFbupwUxFpclAvj/fHvYxQMud2ywlPW
sRtZy517xGSY3RDQiINE7e0xV157zaxweqgBX7lxr/7JtbxC01Ri/SVKN0VTFjHB
2upf6MNEQK1DAi+OSUVthhvv9NrERaynaTKXQKl0yMtDjvr871HPNalJUAeOXPaA
mQTu6n8PgmxSfS9uNpJkA1hdEEV0zDWFGDrcUN2Kxgo/vDeVIhzSeel6wWAa6CqK
CrGWa6ZdNQwXmPkVB/nb5fUqm3RzqORszOD/300cuOaQOGSG+mfsGmMjrGSPyX7a
yQujazx6kjghfTVQYxAW3flZ0A2FubyvYO7fG/+Mk7ouo+ul08sdkxXp2/tTmv1R
kjJC9mFSlcbJvBIbxGX4tjUpRG9Qb5iRAAi3hMzmcBeQPHeGeRgNcM4insDfmBxd
F8U2LTBzy7F5Nm4xS77sFN2A4AZL/XAZ1wB4HO439WcFXv/gAS+ot62VNXW0hcHz
4/nyWfF/2zRd5G4OW/GN/ZIR+tevo3S03LRdgEfJcLsltH1Is57FJmIP8XZX3xmW
cr3zTalNAXdoPUAjOnNGV3eI2QPxBLl5DS2ITxMkASFXcSj+x+s/IkLMXP3+yuZ7
GFBRnGhd7AfAKYMUwEofkSXJunLemGeU3tA7NI7TBsn9qXS4hw4v3ruf9haQQucx
eRHovXO4Rl2HG9Qb+CI6uZRc7sFLGbil5v3YmkH9hKMpCbP4K1Pm6m9uDZYI9Xrx
6XLxVu0Uq0rR/013ULlOPl3Edha3+a6OStBEgVDM7lrhBmc6T8E1ux/Zdu5uGQ3n
3RtpSiE3TJiCNA+AqCMlcOZV6h0u0JhJwt6bJprm6Pr/xPwNl600Z9QMY6jBAVa7
zAGbskeEHHZEFxf4a82HqN/KpfTS6z7a6AChhLpl5V1nQ7UvSC/5Wz1eMGZNoAq2
ncfh63NHDmazR5bpj6L+PzPYhXra/KjwD05E6lMxGX6FxSisbV2EE89pdOTfRPVP
gVv+jjbIrrwRKAL1DmAd8vJHOGgX9How7fz1KZ2LeNuwAQ2TqiWFw0DIKhvY3Lu8
n3b8aiLpkCcEZw724WZhRyHzVIC4I3+10ytvJOqRRe1dA7+XDU2iRSkzywy/4Ata
NPPAzhM9RCwcOsi+mhBuIVUnPAqrgiZnJpp78lUcbH+ExQ5WtFMHfCuSiPLmUSfi
IDz4RZFnJ5IOpTMybuvjB6vnhnsHHzF8skbxNjlizDrKPYWkyU9bMc01G/834ycC
xhqQbuEvGxAquDZMMWnGWM/RMHhJCgw1D/oyfoT9jY1z/YUpsJPuDWK3Da7i+I95
OUYotPCt+Gcbcc3W9pDHmH4yn8HnGQApHa/fWsuOOwSAmSvdAMSOIXCNnDux2qBp
3gnvPUmn4BasCtSrbRZXAjORHRlLz/0K/ZrmpbgNePbZZgwxL2gYk9E+dnnMu2vq
YNq/Ivxu/Bmz1X1YdPakFhKdv/nX6BakQE1fQ4W82fofGo2XHn2VGeunRh3tBSVb
cDbNTIDDdyBRphQz255eulAF05gdH80LUfamBqi4IdeWUVZD/PIh4QEHuKRE8NNq
oG/+4v/wG89z8hd6Qw6Xdx7t/CvuF/FLRngjo7D4SJGIsrdkAwc+1zOCK3fFPqi5
bAsrYVOCa2Nkzr8iOFlB3mXqxFR65pyP4MCcppezegchTBwwTXbqU2Zf58Wx909R
1cEZEhhi+WAdtDtMPd2bsUKWwLs0aiPppBcv7PjqUDJSF+2edWVoMSyKoUWqt+qD
epwzqJUkjqd/ervo/kWEA1VoahZN9p26adUyGz6hNLHzUhWH3kGlxD7e58/6UJO5
LS1O1yZBHBHiGvdcpcvOXIgJLDtPaSs2E992BU75ZSO46FaIMk76+EVxgoHDxLKn
QeZE6lnRcyP6w6gpaLG5KdKc9H2s02V2HVHS1ZveZBV+90q5f2e6d20fFuyeAOpc
gPuLP3UhNe+gcTKvvwBmo1yQ5LYF7f9B9Ny91GGnGPqRAp1HL3bydzfiYp6t5nyk
6JCY1JzrtcpJoJyUtEH2FYNGnJp5HT0JU3DGR/dl8p8u11pfowEOUgbB2f5HTveu
Edu0bj2eL7jutFEM+h6ldTMQr69fCGGsT1PNCK1RTtCp895uUVpMeu6z3UChGWbN
qwKgCh2N/YSYkdQgy8xGWkP3+KCeyJ5C3mof7AoqbEADbKGePhxvdXw8UCB/sWFv
jeMGRuFKSEle8Kv24ubnBByzU5pgD5aO11pRAyHwLYlFmd1SjfycbVk+pSaPD/FO
3nLInrP+EyfjUKc0PwAJe1dWqMGi42lyVNJ/unn9tZIh3/SB+yD001bh4tha2SXD
/xbVuNV2lEEArEx30kslSZefvaoZr9NnoqNICKoVfMy+zJC3eLjSXrQZvI8kXfvF
XAOUk7oS8qB+8SSI8+UBwjlEAE/qEMDcqmmZI0oSl+0oPnzQ9tTT7oV4T6TIZBcZ
/IwdiqclRF2kS5c9lhsBp4QxkzrcA+Y0J8JfwylSzSW5brt0nUcNR3b4eNBeWMRg
KVshzK4rdcYWndPZWXm6OF2hspkOzIGp0phD3EMW/d9YwVDtF5t/7W3jj425IXJc
XT1OtAIHdVnwNgRv5OwKZiskPsBR+fJZ/DR3O3IlHgfKZA0rOcsDWxNzKL/tuwZA
zDNoDM72YWDruGlEXUSpPelnbAHsaL8NqRP/16kgrAK+nMMZGJmu2/EJ+owkO5ZD
oHDuWNrIpqJ/9Zjn1Z+aGk16BnPfnm+1xg8E8yy7Hs4iPV4hsoCluqVvex6yoxCt
gUQtT2bSkeoMqxhLScPS0vKKKca8lIt7a21IJbZ7hZOhse8TRIwccxJygxvr14cz
6A3Cfxs4j8b6qEx3MuvVC+OkUSHVonfUo5scypijDfZwti5oP2Lr15UA+86gW1DP
zt5MwtcuurR7ofYzud3q7Z0Kx0wxvMUISMpwLNNlEuzTqwAjDugLRLveCjtiWjUK
D5KKX60RryHPXLcO7st9rTY6hRNL+Se79nBUvMjZ0iplN+R81O96hIpTGKrP1VzI
kb3rj58a5gaY7VREpGOl67SwySTIg7EzeQMis/18wgOnt43X9ECOAsHXANMoIobK
7mhTT4nHUScRZLHlpKuN1/WT6fxEb/YM+nKUP0XEwaiwnPxiuGbF+PLRlnFhO3X1
vPbZTx0CP37DJgUZFQqPqxOAIGMS3nnekaq6hH1RNdktgCIaN657cpG3EwUEpe2v
RoAgX1WTYl4DOhF4IIy1Gyvy5mrQG93EfKJBNeLiikCuziFPGZwurfhawFGUa+Ti
7LZlrAOKTlvqHlZhMu2UZWsFMxs/J5nkCT0ONZb0HQRbdzqWt8ITp44n146LKYHe
V6uC1wKvmh70+UdPc2sltbPQKZVp50YGUFhu0e+dONHwVn0suYdrUz8d/2SJZJOd
y9aDhM9j8T2GtLCLFkWtce2DXaYtrozqyvFWPNQS1Pr9Ui+YwLPogC5j0LNTuBeC
3Ijrjd6ezIcubY8/8fDKt1MD0iz1kPlBqvshnVk2fMxLjTTRS5qHiAIhsNBcPU3i
3/kEdLEoqlqJ7J5N8meSCNOQFeUFkcs/SEMrVtF4QHXamX2LEjCun3XHPxvaymos
gdVVOOfVfL3zLAFILpUj/nTcFtPAbV7PO6ez7jRI9Rn6EvkWSbMD9WmGbi3HXXvO
vpVlLSe91c3dccisUtYl5rd3EYORGA8jFnlylJKCP871qFswzCmCkbBeKNZghA12
X/gl2rURZoAsuBn8kZlzcHVtR5+20ga0+sdwPsOea7IjxOd/UCXXERndqUQ8/Rm4
DJ7sfybok+dl/JgHmMWAaK1LSRo5Uk386IetViKLh8MgSMDTV23YCjU8F0xWC5Nf
lvhZBQwr5ZZdCHAo1r8W/5cTAiGXIaRtrVH4iHOR0Wiwi8LSXLLv/aeHUZ568Sop
vAU+cblQcdzrRoZDSFAXAGkwfqcIIiivc53cNuR3V4Cs96YK8nUQW/d43s0R9M3d
P7SOycfjfgMxs5IhK0RscvwOU6Myv7lkKTJzyalJj5DRJcZeF59lwu241yqnHBKi
MtkSlssNJCetoks8FC7q0U1IpJfTpvLwPQhRB7O6RIEzsZlzqy/oyra6+t0Myfrh
LwJ+GzwJzVsF4ZpZWfxcIDPt1O9I1Vuya5xfRGtrUSIjhaLwR/KTSNodX5OJVvF0
/AR6E70MgR7HcLLyvG/taFgxUYPqhOL0NnKzRfY8O8Bn38AThRP2mz3nDwBYFdLg
5lnQYPaSZxyugWj7rTS4uqPSh/ILSfpdgFAWusz7zkw6mloWAn/75wRDuWOXIpai
gyf1TwAx8azOFTowmOC+ytGSOUQUyYQU2hQJnHCtjErYhtEOWPxso9DJyl3YwGWW
6Y1pA3N6L4cli7hV2OKivKbj+4X1iHnLrdDk+0aK2nbqk+AoqYPISgeZ+e38kcwE
RckklXZ324zr9OfHu9nnbS3Ok5rvwnvz2Wwr0t9RWFjGaC6RPhGAyEC32mz0ZiZC
Mv9c34wU38+InGwv5l2qkQCscnuQ0LUEC/51+JinYlqbeWYTH6LwwcjZW+krkPwb
gbeHpn24HjkflQGfKYXekUmNiBbbo/+bv5qwaskeDSnDqxXOhALvrakwIA0C5W6A
paCC8p7J0LrO8Q+VglVKKugYIBNBHLUU3WkggM3xWj4MY72Wv7gDzcfNZzgs+G4+
Udl+4c/0PA6zkkkgcTpDumEF7fmOWxjVEvuCt0hXdsNlZb0gYU/C6kMqRzScG7Hd
uaKqT7X/UFQAzmjpVmBp25tvla7Yuyb8XpHao0ZM0JwQfC6V1eUleUWxcXlfNpVC
SlOW4u8A2hmrsH82UOTRzRqGVtIXIHlx/FOOpe2NgjgDHOjyU8ePAVo8hlITNnue
bezyKqcba7v/pj1Loq3vIs+eIYT5QYePxHOL8rJV07n1M9sgCh7TketZMkb1QMbO
EVa0GuO2fIBW8TArVY+QbEqdIhq+QqGMRqFYZ2Pk9lUSI7Pa3teMxmi4q4Pyszxd
ZlyBV8GYEupygK2eYFmSVklXc8BjlwfgFdNo4Ge68E+nOi/SGhxa4IBOoIVsn34D
WcHXPZDSnkRcFIczqKospC/wfja8Pt4ddOy4q/D/Vtsg2dHmXl5qx/5oiqVTFEm5
zROTlQj3qt3qCLO5zhvDh21EXYiP7SgCzQ9Iudt+xbB/OT//Xf5umbu5r7Eh5mEY
saBgK+DCEabJen4YQAMNtf1ROfWpG8uv9+EFxt9laV5+G2v4wjgXXVDbgSmzwZSV
FgDCjwFIosjR9ouVfaBzW93kQH8vq5QJdxEDN74CrsRHQZNfPysuawgOJQi5JDZU
cS0zeTWYL7LPQWe5OeRvwtl3IGfRa0HI5sqTSi96C+W6rOzrFeBGv+LU0/YQYzTX
oDvWqdimTS8MIh9h2BDR6DcStuCapT8Mb3AWgoksGEM3tLwbvjMNDcu10c/0DoCq
hFmpHdNU9n3GRZYa24j5ot/+RBroSuTNvT2DtDPz6wSlkHrB+J+LLHARMhDAqq5+
OuDio/m8xRtlQbDbRxBNowSQLoM+rjTWQSsVlNWB+7gTnToc9dVCQJAEfL+Pg3HG
zhXqO1pOieAiHT46ueqv9tZqfGBg0HZND+QwvuA+RT6zGa3t+EZ6eK+9X6RxBibA
XY+quPJtx6vEv7LBIm2r0DFqsupZ7Lo7FcPmxni4+nD5tdK4r7mackZzDgCwy+nc
N6vfyXqG1U7lV/5wOQoqP5Ze3HkMgWrAB3y+L3aZCZMxabmG8f7mvneZy8ZsMfKY
h7QuP/wTNRXqyAOrWlU9qr37+YUuz+MJrZ0lCH2iN1hRP9Pv7cdGe9lEInj5EYmw
O2Q8CU4zidoxC8u7LBgqBpYI3+xdaXfa/6mPnVPk3cqKvxi+aXk6vaFTML1njJj4
PDZLNO1WKlpoJE8QVQajLn1uC1eiHgIlPo+WIvPvhNtCFRXK7QRYRof6bkEhgF4y
cGNewmZA6k0pTwHzvUShzvkWoRW3tx6lCEymO3yl8mRRoA/StL4Dh5QmBEn2OwMz
nHsBEvPjOUm9hB/MQvezrm6+RihS4DLB6Baktfnuru8tY+9MSsxsahdlCNKkZyp7
/isBvnqbHV+ZKHVXi7U0QS2rOAXQdQHh17DahPIUsWzgvm6Rm+eSG++qPYpvFjtL
U+1nHPqFVseA5UPo2CpAlzKpF8dTHu/cb4Fe/uUXuEHIsY73UG5zimfeMDsXsTow
SxhQaMP9VSthhTof0mCLN0+XcnPJ3kTD94GZH5RixEAUJ9s92sbGaA7cGF9RlIKs
NnoZ+diorvzSI3/SWHWxDf2GRzU2sy395YUTp9jhwBmb6etz2hOQsH3A31GvjLnd
l5ABSpe38LKWCbGxQeQlfNQbiBCey9V5e/iEwGVD3WvUot7jFmcGKz2MYxXcDZYp
YBev6aa7NHFYwyxnlTrudK4iN3ypPVcrUi28ZFkaeOWsltaABgZukFO1qvIlbnmS
g9VF9/nAQH/RiVqrpjE2YM7UEbI5NaxIVUvvcQjIZOulvJ9FOl8GrrnH+ZoMi5VI
GhbNSnglHhzGrWe8/TXuVM1IYYQKmgE6eNjU1n/LEv72uTo3aI1Eck4QEou/M0wY
T3FhEQq/EoS/GMEjGJPDwmJ8A/KE/sjJ7gI06U/BxKZs1Pid1hSIPnICLxgXYQQv
JeH5XhSeW98smxjm0R9nbvlg6lDKFej/Zgt+bGJGX7EbbQVH8YFB8MbXhUQJ+Zb0
3gpHkA4VY40jCYXtYQ3gm9P8aJK91p2hDmyT2ykI1AWp4pTTBmtrjk4IsRNiedxe
w6uTraNbcDFXI5cJZhX8GRrUXGzWt8Pk5H0eOno+nNu9vquj/fltlNrW7vf0+9Nn
Xt+aR6ysfgz80KNx4M+w0QqrR0vu/DFJA06bPczeU5ZwMFDGnXtPu3r0nry9pBgq
RAFe9AyVZA8Tr6VbuuMGaIL29hoccRhv9bAxu4rJY7iiXLsF+dyEMwubvQJbskj0
f9lNJ3wd6XOtUk0BAEUSjOxt0sgBqxg7UZg9Y5z9Ve9alS3mK9CQ30+AyLSMD6ly
0bTSjNii//EZ49Nxpz/c5/vP1M1dWYcRKKTUYBWcBtUmIOvOLUs8LhpBl9LdY/Bz
1v5YqzMT6NeHCl7ewZUOd9Oupry7DQf+nkGLkxsbLCrczGzeUsCqxp6yVdKEYT2a
194bnAEfOAvIE/fyns/T+jp8haV4x/4EYKAnzu+VlZzaqh1ejkw3zygMNNRvEEiE
Rt56ER3KCHCrVTCuANCzxvrGS6Es5m5UyOUxlGN6j4Xb3Jjfir/RH2AAnAXDshQB
42lb29IBbAlXCmWV+DanAkRh6Gtn6FJx3Oe80yE9N5TkGWFEoJhcePCrrDT+OgLN
VdRwq4ttmpgwyhiEbQ7idf26AxpaGiUMJvAOFDotzNcBWOTOnD2z7czi+TjAtKMj
nt+tcPJ+BAM8u+/7Jp6x+cRRCdirX31UH6dSUPoBWl2rsxsb/0L1h9CN8AFhYXsL
P9qGfbSML0tlT3WUnIVoIKLkOReP8z8SYaunVBl6MJ4gAxlJsxyS5uPB2fOXxYDX
jgRw/k5RkTd/m4Qm9yYzcoz3B+rOzOUHmTVmPsw4dR63A4aICLf4eM5fIViAAiGX
TGSqBgj6AT4cAwFBmnmRuEMEemdIfFcjaJtZzdU6Ai7F+RnSESpF+G1sQZ4+KNUX
DagP6EzNt23SodWpJvSTT+gLUdtQF5TASqvUCev5U7XWTnH7mc3Q0Ewcd1zEB/eX
siSFV+qc/7IaiD5fyAqNtWHo/m2tRO2OFAixVfLVRyI7y+gAu79HG1u+NBwvzTZc
cBXgBcjyVKPs5TAWKXiFMxXJto8NBZvK12dctZJGgQ6EZ9aC3huG5WK7yIq2iu+f
UOos7pJPFmLESJ/ob93pnR7XtICLzJAA8n6NvhLU5DweuzVmH4yD7vrpj121Fvxy
2FsywilD7SKICbyqz+gVyiYA+YADWkIiGUwdtgwxW9NtK+oupKR9QLRJ7BkdfrqM
RwJk9pN2Tr4L5p/RwAfkktC9OnJLmngLRKi1T79Tz4+ig6ofbCDt0uJQKRFPQ/aZ
aYk9wmh1W99PG2Dlzc1IIUHB/nw94UlqS1zEQanLzIZrOHT8zKJ738iWH5PAN/9f
QHliVfwiUDKdAZcu5C8YSbbLZc24bc/J3RcXgFZMCBoMCKKX4XGis2mZ2gFdAePU
C0pfIKDbtSunk5hGmLIJ37Ab7GcUeNUlyFXmYPGAtEbnfV7Oc8P1Abq+rbe4yXzl
chFvL9ASimKU1dm+bna9YvdiTH/zIpsqn/YMvWGm3KIAHYqLEyA6sNTRvip1M9jA
70Bia1MFikdSnOgkGp1kTwx5+tmUZ2qanqfuAI1yROf3fg+r5uJbSdZKf/kPBO0n
NkMatyHJzPID/Fbr+zYIHRnXsW0GmcKh8NgDIPZtf/lqormRPLbMVSEZzFO9hhk+
/7Ei9IwTeSnjaDYVoQBfpqOU5Jw5as8oEhIXwpCeJ9WQUlhc+2VjAwKFtiycW5G9
r/ljobkWiaGw0Wx/qFwK2X4siauo1KH7o66EamOGeQ7olVyRRisJCrs9mM5qu2qV
+RDG89L9Zbh10i0++PwntZJWBRMbvIStIzToE1VWEgYY5uXOnwTlyiVXV/FabDU0
WwT0hZ2BylqruYxkFX73z3mhUDu3d6KW2W5hALX2L5jTsekqjr+CBoVCvQT79Yvr
3Oo2f2NzLcudntrVBX2Col4iib2IN4DUduhuGQY9B8auK+0EknDxbs+H1Gbz7eIM
mJSa2cP25KhcY7grWiK5FG1pO6wMvdyXnHF+AILQrpNiZrWZZxcCQqQmn9uWhoEh
M0Mz+DFZ8Vtq11W0jZMKWiiwOcIJz5Dbie2EsOxvANwEU3F/Iw+cuQjcaFb+/wWt
bnTvyhTClh+zPGBsyHpXLUJLU9wmTnJf1xtIdZfgpp2uwfoMef5ehzKQKZJbnWlF
EYhJMmyV96ZYM+A01pyIiGjo5gP3tOkV+i9wPwMBS3dSwjoulOcl+akTyyIBgEwG
R+jtPGPAXA5v0lqHIvM8zaGgzoj7+JdrWv7CTygDBjNiXKEtY6FKl2ZuzOiilWDk
lStt7mszVpbM2sBjHuX3Sc652Qprf5rtvbsNXreEOjk3FLXju5koPrARONoGOTQK
tyatm58TOKT5Zko6IU2lN8fiX/R6aQBk6RheEeD9fo+jg7BtpzCMcxOFDLHcM6tJ
FMzIj3tN1vevJN/aOnrGS8DFfx9qPEZ2o8YXeaZVoByKWHL5FeVUjoBejJ80LiRG
MFD85G/DFGSVYhtypW3xEwaPOuZEnEPQi6kpNRV/qAmNSkXPZoIRACjSSc/kPeAh
PrScrYeKwYuAMhDmLk4uxm+WmgYI6sPCAH36j5CciDHhGLmZD8lf/rhxQZERCh1A
gpNE+oy4ysn1xGKqxK9sq6W83s4+ELEMB6xGpd+oQEnoJ81m+XlYMi8ZsFPo+oZk
BPipEVj0SNLpw2LMjGF2sB8Dr+KzpKFdPxF6UOBB9Nuqop7cMY+EzNZiwhywufF/
8dqu+dSXi1DinXC1LGV+WL4+VZDyTwfkwQ+Hezz8UAjCuTEqGsY39ExP9hcMsvs+
38bHXm+qMieK5ibIWvWaBGffMgAJUeVE6inXwRJxhQhXx08y/ImEiuVbpFcghY8B
jWjulZSqbJncVC29uCMVuqqBUoKimU2okBHdAU5b5R4Nr/iLaOtz/afUVvrZ0GMD
Nx0RwR5aeEaCfpngtUmyR/wyrLEagQw360bsCI+Fi3CnsKUespYpP9WJw/ei2foT
uiwMpQewEGskke8b7b4ly/i+X03yaP1+Sl6qZdh6/bCtRDM/X8jPdzlDt3A/9Uhb
WSvecU9DihFyWNvtKbw2dPZ3M7NfBTSl8UXixvdBK0sqcNF7nzWcl45ggdWMzFwM
/RMqcIQQs0kl1muLOXl6E42i6CkSvfj5DwONc56sWCj6/VUqXafl6/7YEqrGWMwC
pDnPhrv1zZCeynE+0X9PnV40eCvrQkEtQhtBKQov2dBBBvnY1qqWpLonRhnOEynH
8vindpgp8pAljyBOBljPQAD/CJSo16QP9eF/u+KxP4Ua1sw4F9BDX3YDieyPgy9D
H1G87si7hEBm6G3FqSIijkiG95NFSeo7ApiaI7OVGiVT+tt1opPe6h80eW3KQkh6
VrQU6N4P9vDlSUbtNG+L+jvADsDcCV0c3E7lrr00ZjNOrFxdYRMImhBlLPxvp633
N3Wqs1lOzyI/D7LUkUpaimizrrCPxpsUJ3Zzjx1g5+nYMswMHepgu9rr2KOK2Hey
47CFnaP/qTDeQCvanHe0GrXfZaE3iOjl2w3EQt8iZTLZPmwLd8cBz3BN4i733e+E
HBB0MzCDt58wSTGa4IG3Mfe38eCVBElMCJqOZQlwfEa+UUhS0QRZXb9cf5sJZWwX
F6rcsmXPfuFOCDhCH+UD+LL8poZvmbjYxHbqS150g0UCCKNYugGY5uvv2+lywyYZ
FVowGZF9iqJ2JUWYjWLCVdWfHieeda7AbZ+641SY/gKaDKzwGcxxHhRgIBaPziCG
o/Xjy0i3AFZCSMOPhNqR1cNyXtEnmNE0fp8UjcrcITg4qkLlbbGsdRRXdxilmMtS
ItIK+1uIYPdEAKMz3Yr7UBIwyjnO9I6J1eo6KBpuozBgrInZ5fDMjQXZZcOAaJOa
nEcNUeDYRQxevx1LIMBwbW88Fcj9y4kBdIiULX/dMba2vHlvz9RGIJwTiD1Snh8q
hp87p7Zif2aElBLUZBZ4PvsS5Nd+eDrThpV/tqwAwJmTi0LwCb7w4ZBRRXm789iA
dudiAXCle4NcqLI+1Aneuc1RawwWSxRr1GTL1Ns8JQu+Mq8CdKyHuEA7NhZzEyNz
+0VAq0Ug/TrRRbwVJkDSZjvxPHS7gun0RRpUs8QQwj/JspSnjjk2EIoeEZ8ZUjsp
lSghnGpXE153hMafxJ3XnFCw8UMfzWiZuMdcauqDtxblzJh7TSNISeJlOYZpYNV1
tLdUsA0JEkqfBB32y6lgi6KD7wknBudvdEGAZE+zmrpq/+JttnquIqQsun2yXFep
pcMwI3+8KJ0TAlf22tFpFqtJlEpRVjZvk7qpSexfScPTbNI2zylfCimXfMdd/TS4
3wBcNV1gshILo2WOyk/SgYjubgSFYRL48wfHe0CQGs+Gp5jy9sVbFocg9OkZgM+a
MFBTVmqJB1RvePEfByr2JLsgdNFdiDi3ityfrtrBM5g52q5A3KIfXTm1GxVbBE/N
W3Xq7W1IH9YmAmvc0EyAvIPnXhHexACXzRWPq00fsOtenEkgyMoDRK4zc82bS/Pp
1SI9MXuKJN1BBmYBJH53vcXBeK4o5eHJ+pO023cjfcCiVQ095inVDotuByT1AtlV
wOgxBZBg5O8WZ0IybREMyIoEW82P4AdTX4/F/6OaNhBZFfAppysd28DHdRpLxk6E
RyUucG+MK6ZT6xBo+fP4Ltdsmk1/D+12XPrF3Bl5sfDlHiyPHpuQS3ol4REwz/Bz
BUY6GbTUW2kkSMyMQ/qoH59A0NeoU1OseSyi/Xe7iQLmoTtMUj3TX+BHtqRenM5S
GUyzQTD29nuDTAuC9maIWcku1NCEoUX/1Ic2JqVQpnDs/TnVFgM70u84tSuOet1j
uu5Jb4/z7n8wDtLdWsjFIvjYazYYqGUycY5xLg0msEcLySRn0JZEhNTvaIPr81V0
ajy7S9M3BJbQ/ta8L+irgDwqXzIMrq2vczA4trVA2w3z9CFr036+y75/ltr3OLvn
rheWFyMWTqsFeHzYXXxMMGCrGoI1TRwEhe87J+HypZr7pHWt/ZVLTj6RNhEasQv9
qPdLgDijjnoMjxFKNXCEKQ/fz397IM895O5Mrj1PpXPibhElY4VTHR9YQTp2uX8S
rciq9louJLTRHTv5jy3xYT6+fYYROBGPXt5qvq+NLtmhaYtKAGnfuwVKVl41E0oW
NV5YOY30q6FqwA9MhemNh4G+i+TYOMNS33klNlvtMJEFWaZsmTwKJU5WH4yC9EUm
3/nl894vySkwItBEZsP6g9Esc3PvNB8Gab71xWzma2oh4DoUDDTRZoJAx8izCiov
rPLz6tC6T0z9Y0u8/DQTYG/zkOMCggBCEIK8rrg0O0UhlHRQiHKAsyfwrezuHsAi
4Z/EbeJYrDd6d7/o+yFDMrT5/AjRriYQK6WZbnzZLlwCLobS+8uW7JSKAxur3fzd
dnzi/175t82dZXt4LgorH6PxwV7TVuqZMAprbmi1J/0mN2+WTerzedx0t4w9QbZr
V77FLkE5710chEbeddMwPwrtwS+NRBswUnUZe/BzphP9q3z1B9q6L6z+chbZkdPi
p63p+GJaHdGmRKamZrcyLT1FcEDtAlVXahCguxd8GPhYX8iLlDxRVXchja7vSIuF
fQtKgskjnF8qlF+tVktYZyYQjisz/DHWD/rv/QdXCAQDcMkjmMfOi3u/OyvYrnHs
s1MoVU90sJhe2Tb6uM1Rl0yunxxG6KBLasbcHpPJGk+88eTt/SCNZ6G1UklzGUWO
7ZNYBpoSCPTThR5lxdGXkRU+I/9y5CKZHQduBxCiO8nmB5ySggI5V8lPm6t/WSVf
mj4WywL43Axpc0yylFnBirae7JMIDRRWWFqK70k+a0Jn7PMj4FY4YuENj76HHorN
/ajGKiI7r081BDl3XskqHtC7YUdJpUMBp2kXSrHdHQ+uwObUdLcNA5Vi8CMnC/uw
6Af693rPt+5UXHueD8RYs7IAV2Vt6Xgar7+1r+mGtMqxY3Y/oQD8RHDFe9TDVqK4
xfMV9A1Nl/bFv9BiTlEkqPqVlvIIWJI+t4T6elkVNrJAiVV31tVS6hT6c6Zmtuar
1ggKz1EQL/gU67VJgkqC9xW7qWqgGFWfzfLnUPVEYS0uzB6pIw40zbOQDUZGMkQg
RavbEG92FmL3H1xrlRju7IOcpClsKMhsQPtnB2dcNDMhpAYDBeLwnal0IRGrXT6m
+uW0Dscvwc1J6UjRaoo4HtbUNEWlTpmQC5SGE+oQbtQCpevYkBkFwm2NfjPCfVIq
JgGlOSaiiPenkJAt7yGDZOaoTUCu2t5n3qXvmj8nVVLdHRsm3KNsKQ67Ri/yIfTG
kHqDryiGpPYZFma7n5umGVRpCAj38r/JLhHUHdm9T83J3rkpDuwzdFpXDQHw/FLS
WihEJVbvYn1ioEyE6CQjadj2QzM/PJ5/EFKFzAYYIw8tMsEyrSba4kyZiNbMuY0B
gZuupX7RwJDzTJ+jx0DH+w67uAGugAALK1ANt6rOu1keZk8dt/v8sM1vo1Gl9ONw
OIdMJTcfAIVdZEJhO+BfODfm7I/2PAJY2DBchzt3qoRjBclB1tzwqgxGhd0SgcNN
XBek6LIo4AuISsNBhgkhIr+e+0VIvM0L50gFTyZm0UynzgwuvYQ+UfdrbGOHX5BV
r+dTZ80buJgBthA5yFngk3PwPXvfQZtenWhDJoEfnFYU+Xjrl4Y1QIzGhdYlAnLb
TwycU3WsoRarWZdGD/itB+bfrglYRymeJs47QNawQQCsJ3F2r7bxYSSFWoaKpBcM
DYDkSQQdhqetXPIwkiAe/PYiKRD9d1bvXfuBhU4wRCo+fYEomys4lhPH6XRZ0vET
5LwvdXVfzJgFjGxuG+winGMzyXdPm6XBlsUfeNTpm2AvLIz6e5dd0l7KKtZLB/KH
KALDX8O22zGbkk45xt20h7Co31GHVsTRcqMewM/QaVcdnaV2kfWtwbbLBkM65oK7
Hn4S3nVuYcapkmDU4QLGqXwh+YJL2NRRyVMXUjvx1MqvcIsarBith3IksSv4Uy7Q
0jEzNmyZtlAePFyxy7wxBcILeSfsMKDFFFNBO46TUDPkvDvfMKKgOCctSrEd14Rl
Z/aSKg59HFqi0aAtNyOj7g1FHAQGKl9O6aU+9bFiWc8goCNbXddEKAd7yJbpqXfI
XhuLAYQ/7omCFYr3KdE6F64Wnghc7d+k5A5qBoA+GA3ozVq/ImKgHGHGiROZ669Z
k2/5j85PcBsoBlgzY/vppcV07kHTbySmaNJoO9aUYkV15rMy6awMKElZCfnroKcm
tKCunRZrzTQskNcY7uIvknu115HQg8dPzSSg3qrjjdEBmispPeTfvmpEsElUmHkm
/fMvc5KxqQd8LTLQXgSD0D5hURW5OyL1T+eGjdnSZiuiA/qjrWSnL63kk3cpDxTU
mzksO10seqULUj6krZh71hg5nIP4jaYkCYMdlhxJkVr+l1F8fkacD+i4NlE/wP1h
8tKm/d8ADp15sOzTBeu8L/9nYg/Y7+U69Oa3iUR/tCNFPkWZ/lCn8TyomHd8GTgQ
vMxaVvuXSGWOk+5ZZUATNOFe9rOJjz5UrgkcbEVr0UlKH/5j9q6mbOj5annbVaTb
/FspTwVA0UhEqkPYQ6pFf3ylxB84xGh+VYVUCtdeL12zexlq7tXYbH6DFEA4/Z0A
ViXSC5AKIGknXMK6tT8PnI3UavHtznSKBee9/8yShfWwula+3jWRKXr40X3RlJef
V/qgtslbTcMmnSVouGb/jwCQ9m3OAVccNudEHhC0BFce3cX4f2A9MM9Vjrodl0dk
rU1ooyJYv1QnHZitOUvyPRNLl22U+iX0xB8Injogfk5W9G71wwHgI/yD0ECv80e6
gpc0MAQyYdjdzJuSF1flntGfsCq++yOuC7lslhMjBMSaUvLXXU7FzLy5A9DbKnfT
5DT6/JTVPlmok5xJQtCnNUlen053PeMVgG3yazLT7wckLgRHqr3Po0Fp1eG9WfSy
tb/GSapaKH3xv1/Ow/q2hL/iPPZ61q8dI0iDRqbfyrk3zljVSRSwY0XRlfCE9S7t
Bh6zIEKCkQZAanNBao8k3qKsA1wYWs4DDkhc9jwSRKLi8vHMm0Vv+Jv4TnPPpjNd
osKwmIWd5U+BUJ11aH0TFfVdhcN7+tHMx1zY1e4BChvwduAE9o4osAis5XakC2iU
/G1gKzhNIMBcmsuN9NIPm4aPcbkfMMo6GISPJaEEIp8F5IwYAKMDfO703UsvGmiX
PhfpIw+6ZwRjEYD0bAGuBiqkV7dDY1PBV/Lglw1PYll1Tcplg8TtEsZUrPhemlDa
6HRiFvhYV881O0s+9u8pMPyS+IJgBOAYAPHWm/F8ntMp1JjSlGSOaIjUpWFhF0NG
hZH/WkzRyU7Jzt5MuC6WGFSMQAXylsDPDEoEdv8+H/+VnqgT6OO0kMm5fKghnDWb
QGLfQzPqZMt/7El98znQHHPHBx9iI8ChScnBH9oaOcXIOkD9UkmoT5Xgo0OfR8XH
w8aNGfSRwEUVk4880GClr3I9h7ORHC7mubya5wNtV9Y16ax9RjcvM5KdjxUPnK9D
+NBtQdvuGJUvDPGlKRKubXRh3PUgOd5B5hlQDei+olohodmRxFytN13iaHvNc/tW
V5m90L+09qqdBOPqCbzYPjx7EspJuJuGGmUHGmmn/dJGPwNnK4CX/kBiE8Ji2AI8
UlwmhVrQr/kLGWJWXH1OctGD803fhKzIuGhVNBSMGQpxWFyxpwqEF7V0zfHuTcX1
TPvrnaVJw+a7o/Zx0RzB7M1oWB6Is7gZlRJx5Eoa3AFB/jW+vFpbKjsAxna/C0XE
m4L12o79nrw0oeJbaceWu8nUIQbs2jBp4u3wXDRLBDD1S40cxKlxBl1iNcCtEyv6
TzDs9snS1hnt8uEfd9Z/q55gmzQDHuFV8GJaZw3tYgfkBO3Zv5QwWfyPd7A53GDx
7ntZ4a30BGNGORVQ+1cu2czlXVDazrtZUJYhEKnwF527NoszWTcaUVEpvSg6T1hq
O3Q0XeQRqHYuTywWBalazNzgjGoiNvbKYFyFy3NiKQEftFQAXdSNoSsGmBy/YI4R
kMbnnXbNexl+FXvYIDD0pYUacANeUYBJo6Hfyf8DPonkytdXfsc7b9FgHSXeNjth
SlSsqQtYF41JVj2hSVh5H2qWzscOXPDpEuBDi9GaSUZg1kNfsecgpNuxKT6DyNlk
AoIxKXUFgFVEh1bPtSbX3UwXeHd2cUzQBR9SbL2JR7LPmf84TY/m7V/5JkxIZwj4
Kr7HbcAk538XDdD4uhd9KgMyzctJKBxiD4pQ7tgee5vpuUFDed4OfZkfauckEa2n
mDXWbKCq0yFp2baF7TQdkALuqJ73VfGqXif0yvwRYtT+LDD0Uoa4UiKJmeFbyEDV
mwuIqU32+FXIv2xA4MmbUoBrfV6YgHawaY9ntWQjRNnMPo8q3nhPjFNW0qyDalvm
dWvZYCYU5cdKoLZhnsGezEGNYxncijudJFnN/FxAc+lJr79KrunrLDCSx2zYomYk
jYGXEa/0IoWzNsSbHUrloicbQvcGCYr6wghDS/xpWJSQJJn3yvqkw8EA0hghYCuW
bpMtgKEgfEoeo6Nqj5MjjKbI/WshXk3aaaBMLW7hka41M5oqJ4tIMCUbcrKjB5+1
uQTzFPlf4s9A8Z10zy6z/tpEmcuCcRljaHwvb1Fg5shRKr5j+8+cuDVCexNTclrF
cXyK/p4Y2dXK/8U5wmUQa0oyfXTAHRpQTQo6o8cAIFQPmN7W/iaYzmo0cYzqE75a
y1wvViGBj7gCd8i04rwCNdDFmzVjaIALM+0zD7KjeYSPVkx0Khihl49+hTjC/jEW
VVvA8bLK2kOGC2Qp3Uwqg9i2PQbJylNK9yZ6k8OZtdG9TJrP+hX9ax5+7lZw3T/L
CU+QVHZmweqBvihym8mKWQIpwGSG9RxAxMagdNVa7YwIjOK2Mpz/WSY5/GnNrJxZ
8ULD6Q91Cun4I+Y717mGu5LSHu3qh1BVOIp8LdLXCU6r8q4jJr+CJ5QB/wruQSjp
Jw2stwSvyMPphf/+Eryg2uL3e+wteP2c2H9d/vDZTzJUjBb2HJDTpe664mbpn0K+
2OVfdLwBtqYyWml5lJ9nn0Cf5DX49/h1D9ucrPNb2y6iaQ2IM9SaV7oF/QSevkLJ
ndnWw0SQp5iM27wV+F2Kpmrfcs8NOpkjrgdSeZ5vY3M91M1aRax/RWFxiT0r9Qta
AXgo3avy31y/13RLyTTi/mErel/vM5OxyosGc0G2iwG2UFevpS+0fuLbtv/r+Pyk
nT5F2/dGOzo8/d2XHCA0T21c1Viseabg99y5IGiuLd11mAgq2kn0deb7UcAbSGeK
yL2DF1KKadwbpkLk0WNBJjcD46ypT4Y9FcY+BVCvSM3zTFYVUUka4t9fwr9S0uKY
5gd0R1diLSzYssRTl+Cze4+fAjGI6zVvZMP1jde1BuEdhoFPdUhkr4BUnvsfKTt8
eSDT6AnfIxZzLSU2tW5kd8d0Xqeoa56UrTtqHC5ef9MI9vyQZo+XH2x3sPJwg8cE
Yp4DVqlRpi3BZjqwCwIIzLnDiHSYZHpmLVBu759r+fZkJb0OmCRu/CLVwKizNIPC
+6Aiel2mWsYeO6ato4uzYd/M8seGNJvLSY665HJqGq625UqhDQY4a6padiYvHqeL
yAo1IT2CSvC9+ABx2gwNasIaF7Kzi97tdXlFCFbVj/puEnlTSWrNvXMb/PjbjMt9
SRYLV/3nzJdUUMYT7uYOTm3ysLjnYVJJFCAY8bzprfqCnLXqT+0rA4H7nFENoEZi
fA/65HJ2Aih/3vNFrRB6mfxjRHVNqo75ESowbRDhiHIzY0DdsbOLW58uDnGpbld/
PIq7F1QKdmZbPQAXnJOIC6ob/HxfnO5SOZK8qqZ+Ao/irzi4R9kOne0GLOtJlUgv
c9FI0a28fFQRfO1gvkbGDp2i4TUyZxEy0QpxDS8vNFIyvyuKcO0yMhNPJUhI1NaC
dgLJUNir0K9Tj7PSRKzIRw49tPl5/FBE65rrKWhMqZAaH+deQuK4Towa8JiFDPAY
kxILl2gy0RLbGNGnh4zOgnib+O+zyC+zJnmBo+/rssbSJlLMz88O+TrdtTMiFa5F
IWRKrRIuWRjfUKJaBUmOFgLbLs9o7ugCh8nza24yLGi7jxeU30KQ3pQq1PaXYVFB
zUxsZtcT7+YFTKqCicaym9o7067QZSws1vhXsWS5Y7HxRF0wPruWDGtvoWs4iZud
NqLHdAHuCBsbpzHXQPGY/IbmqcOyR5cC6d0wVLD67aPBJQtddSrjDQogHD40GmTP
Ju1BbN2T8SOi+PWPj7XUez7Wj4aVnWPNaH4Jp+NLDxIPuiQZs/tJ/7kZy3J9y/1H
kURACiUT+9rksuUfKTtgt3kZLuhZjAXvUhTNXCR2Gx9bqMLnBuuXWOzkOrMUfMiL
l+7EI0puiLDM2N857RWLRLbc6xS7te5wIFDE4S2RZ+ERREPX4x/jrMSYhWyGvOR8
pAD8ge3OBma/D69h96MPW9k18J5oWvOtQD2BSu14yMZJwrDi0AnTLviFZ/yHWP4H
Mxl5iHGvGXpGz2uDeakTRt/VN96GrrMMzrWvBVbJ76Rlw42+Rh00hXjWDQIBILy3
jxjd0Y+qIvBlpCWEIRIkE4pPpNVWXnM3Id41dE6i4CWhndo11HqyBGczvYl2fcZU
v35JlT0K2dqrQmEiwV9krJN4rxXC9+innxUZIh9B1EWUbK8hz7OMZwnk7c7twiXX
Tjq1FIyJmocg+NaQrrRWjQik0NXn1iwbu7XKWApLFXu5lD9rACL1DeZNTlDNQIGD
9U4EI/tQtUw8dt6yELtUFAP1da2n41mviE9vEa3IbVFn7XpCepaQKnLgW1ZFD37y
9XELUdJaoNU3/Ka1fqrPrkD1YotmdX5c8/4tNAEHmj7R/oweAeDLfw7kQUkqzW0S
EaFfGhhcU6uO0rw7gFJ2c9dZEzVevIED91Wx3a3oE9AZJ/N0WhSNt8lYBDod0YdO
vpm511tASR779pB73jvfYErYIQiw9Jfc6gLTGKhS2ye4+D/mUy47yO5cm+JgGvbv
OB5F9DKvaj+CMV3ZvxfPhamW4mtBkbJPeSS21d4VRv/nrgXwjs+3sPEfnKVEDajh
vHlUItsbPySymc/Ufkv6jkXENrxEPAV5U8AYYaCj7YkbgIokYo5/TvxaRsh5k+D7
3zFcM3L/f+Wa4kO6XWuVJ/TrRU4wDEuvhhAESnsiW6EnGljL8p2x2+NSw6U89yiy
AMu1tvGA+e2iXMsuxqe7I7SW38bzJ5kpAndpF5pysvgTVEGg6G6Q/P9sutdCi+zJ
9wFoil4iPcO4xxODoXx1yHQC76SElfZ9ol46xv6XnzD182Y/uBh8sqaLvvttbnsj
nV5dS1Cv/h+rZy6omwqK+AOMf4bfrQVL13zWkX5yODljbRiWZR9U72DhnGjD/fo4
fr8pX3Jk8UPkjnyyZmmkrCRnDIqRNmTo9Z3s/qgTMxXpFcL36JFlCOOJzUXCcF6j
usPyGap9hpEloYB583crGEm0caOX4rMxtwNLH/qndc52tRXa1hRDSSntftKBz8M4
JEfMr1NHsgDzhZjLCTCVCOkWdN04aOTaMc/2+HCvmo4gqROgUsau4EKDMauJm3tb
0Qss4GCfp0F2SouQBvtGZqPXNEoyyl/hBEJdb+n87JSk4u5I4bt+R2Wa/lRbnzPz
UDqsY9mniXPZJ5gXUh1A6acT5lpWVCVnpcZO5Fkm5NLdVH0yX9w1uFnArvflLXNa
kazv8UWhNtlBczHaxWUPTlrnspBI0cJD7UZpwpm+/3eAOwt5oVLpjtqMqavFEtrI
tgzqsPBfAcRdR3XZ/RfQE9mzgU3HHPwqSoc5PkUnmGQYI5Ae5x88fOlDcrUEqOmu
o6hv1l7MyVSK7rsvIr8IKU1ahqJ/xuFL+jlqLCviMNSOmoSVt6GLKjcLzK/2thqZ
yRYdPBokDcM6Rbr16EROyg7/TJxql5+Dr30lT24JOeBzD0jww5G5adRJwAlGruk1
xDguLUUNlUBWWsDC8CCuVwu2TcZrb0VLhUFl0CfjrIp6UVjRPi43ltOPNB3euIan
pRBd9ckeCuLsXdL4/joBuw3WdgdjhpR9am2haEK5WSuSWHFaAQKHz7PGPkMIk+iq
hZAjBIs3huF5T6kOSKX2kquhBrf/CBICDgRgE6UDF4EEVJQdoMTFBqyFK4CFJtlM
uAxAVmITwZYjm+Oi3F3zQFI+JDxXWNjbmSK+A1FpyHqQgRhKOPBDQ8gOfYwRysfV
Ip317onzDkoplo02cFdtoed6HNOo2JEqYFKAPUYVv/sUFzAUiXbaTCUhHb7ky0v7
P6BkABC5v7rRVNWxOSdpE0g0uSyGhN6xPLVgAgMC9VBVVdKt9uQHwrvHI5j+MtfB
sMTLMKMf6tgI7sEeRndCqw/O17kPCrZsOq9cz9hwQTxSUMHyU3LI+VvCz2qaVFbS
PdsDNJ31Pym58KTflmCQMYA6YgHfgwB7fc2TkCoQo0F7+uc4avX1DRCxfiTR8/vJ
M4LvpTH4M7iDhYuI8YVHiFyLREeUvjYhdFKDVQ/UEk1mSzslhdXk0r/eFZaoM1WD
eyddshm70WOpaX4Tps9yDVSeKyPTMJu3Y+eqg6yXth+Tc7RcmCpdKfx5C04BsEqU
fqgaz7e1mKtrYxotFFfh/77h8pIfNf5JIyK8++03Jq+2/fxLGd4cyTInzETgbL2I
GybDL6ZdcxBNiINpdahybrH5m2cuHgZZgXbEG5U+gQ6DIRCb+qAgY8ku7uA0kKtW
xlLwH7GMihXQVCZVkwDlNAkuk/YCDH4vvUiQH4S+Ed+m1T4lBnxlHiUtvkNxVhEb
IR1hTRAIkLxv7vdyzmOnmg/wCAiVtL0mQhHDQ/cKbU3OW3DXEOykhn3pROdKglsf
TUsuFct/3WQpBEXUdUUoiU/KWCJCqhI4hDAh3mME6F5BLcguejjw5FC3XJASP8tn
R0K3KACW6LumnoLm5+lxAxT047NH/zHXxtIfFDMuXshlrh2sPTvY14dDG/4ltWMY
Eqn0EuwuF9BRTwVPWxRIQudHS1mD5kHn9ucirc0agu+fDa4oc4CdFza0+o4I4Y0R
rqEQszBUnHyJnwGoJnm5SvbJKUy7NqY+Qri2syMnSTd88qrrD2UuW7Ipu1/ukL2f
5wOHeW0l2eE08oV7nBNA5CGIYNK66lx4mLOdgzsuZcc+G32Wk1aG6y89jcNFy01A
07oM29HtrRjbpIBBZ1EWQcLxacX2Gg7Wq+2acAMFyOvyCCzIg6XGB37dPyLZVv2+
m06xSQA3WQ7B2BZJ8+faQ69dEb+/DEABhABRPu0wiAbxtTHJdbQkH7YvWusn97/M
Z6d+zOrdevlZUFNo1GPkrwG/b582FPAoyB3WJbxz/FKgl2AHoSP62lm5NgJXQkkJ
qJISNi7EoGmQXsArEwnFJdwzpvx+jHlAjH9F5gUrfcrOMrtfPgD24/z5DuOC7hTM
r7ityyx27Iy1HDa26hYuk2heS5rtTjLRy9VQZSpUrU/uqSVJVrWfKv1DFOk+q3a3
rMBzDh4Ze4lNgRkihvfjj7a6O6ivUr3yIgBdd1WJkkWi/UquP5syC9s/efppu+rq
ZQHpaXIAHeKolhTvXgzVATHyfGj+YY5j0AjzQNjYxW3mRxi2RZei6C9aq9hxSXH2
0mOcX+uc+qk4n30apJkppOrnZfyLiDS5SHP9da/bFIert2h7mswupdWDnCak0qiz
sAgpVCkZuo+tAcsHLDHSOwSzqIJiIHsNWdb7wIhlglUABUUl94ZpZKMJH9FUWsrl
raDqwiGNyd1oNZMnbGcdHDo5BqS+mdVNRKmdkXDgrW+9PEEpW+YkjmS2LNPedRxb
/Z+MFvf/zfzOcO5x9pP7aeitPJtu3fg/6KPUM6V9Zhk/8nVLg2JbN+PkHPSTA357
HfzugCyibqeeTQMSq9ZFDL6BmVpWTzrsUlJjn4Dy/vw8aoDL4o6ysV5i9GNQjAdg
Frvmm66yT7YAZ7QMaQhZwieXQN/bAKSWeaQSM7+UIgNEFAObvxkrPka3fTbNNI3h
sMFL89oYI0G2DggrNPEVRzICXErnEvFUWBSocuEtyII0aERVkPkEeAUIROpTXkSY
ZfPIGHGSDAVPbczMe3YKpIpMUVBltyr38WPb1G7CvxpbtmGNmCryAR/r+evjgMma
2PXeRNJf3lqZmLLlZBaGNNcC/h9JvgtQCIKCrNVTNK68z6UfMxMBrdDFxPZgR/BM
0UxKTCRUNxRVpiA2QmCpxgV2lp+bdT6tc98Y06KKb7i8odE/YPuhYIvdSX/gS/6q
HXbU76QrY/t0WEmLxnMCn7gW0rPvGl+bWP8ukhXnYQSYowGTZF6RufQ8HsGb1JV/
/vef9l5YMLNhAmvXzuoH5HygW1w6Wfq0xwqjVOxTsHEBZDDEY77TDfjUs+ZlCQOO
oHedbhN8fFfL/WIU2+6RLI741tmVR+ty+vDvar1s8UkWZaOqfHO0/OiEu8k2rQw4
mFz5gx4SkNTCEnn3kZr91L6i26pFQjOoyoQi1qlUjIWmkGEVOrqnCvVy777phwXL
rRl1V22BKvz9Avccpl6G+DvkHxGnNyA0G81ar3xC33oBNRVeenBeCyKwzOieUg/0
847Fx9fOxIiPC7OnvjqJgDmaIjPqvIM0C6aOnoJFlL8PHDDnLdOvM3SfwHVkDnDU
EQC5VDeRvPceX6zDx4jmFm1LMfIe7Nf411AH/1qSr5QDVGZgaOq4QE9UWVJdS2lu
POAsVSA1Cqfuai0FVUTvYs3jbv+30N2YBHx+SXhcx4gRz2I63tisMtdt7EdkBNV+
zfJAsQbf6amILTPyOjI0ktdMjUt9edkbE+T2peVdYSm101wtMfpRrfQ92jZRrDlI
msW076u59wRgY7oyYGfAOZxVtICh1cv+6Etj+Yl8b2bY00kAzgZZ/7JSrp1lgUk3
EdOjmGrgK/E09tjFDWOjxVNfLMCQpdYgG74/mFzprIZPX1LRB5YzeAPUMKPrnJ/C
FbDCMDWq86Sp7yVXgrD402VJFXUxFTX/hT3q/9S7YDh062wAYaBnVPVX3/HIX1ij
1HadjJ1vu19jklxm01V5XtX2zgWqeeGTOmHpDaLTKCU1UPPzTecZuWwQ2lRdXnYO
jcotMJXNwMBB0CYT4fe29V1d5rylhITpB+O2tX0l8Pt1vmUrNyzHhieVeEKGiJMo
4vdis5POGYUIeOiOeCnPxWY8nlcJhKfA9rFYBBA7ClU28TUtCnD6tuNhV0FzFMtr
DLSQcavluEQyh/oLEevxidHcEoHLd7QIJqdou56hn0Ic8kBUivogGIZU4syGArYL
Ov71nqhFmagZJM5Llq+ObmWvuNg3P0/Aeb8hZzJr5jqUJpDM9tf7DTrFlQx8V/Yk
OrbQbpAFpIdCIEvEpmsEAqjoBmLHk4eKBv0wCHtwWb3oc8gXYEdfFRgcPmm1b1L2
6lNjNqw2eUC8pf1Kijv3E3hxaTi5BDKbBCD075A5vQh6V/YdvkaHNqoIMlfVl+iQ
NhrjpDeOa8XrALhHcCesDCfL/HrKj8zy5xdLAxFQYpTtp2HsBljTL8x6yZm6LZ2I
ix0LOj6N6tRkUafomUgbOkI2L9vwDdE465pHhcZrsqAR2TkoQXRr4RLw93WBMV1p
LDQNkRQq2Ljdty3zxQ2BwEgAUtxmnaY0Il6l60T03Aqkm0mdTGzMN1V2ITgMSYhO
GDY9ZYQj4v+Z+LjvXVPdRpuNi2pwb7RAKIIY+ld7qn9hLQHp220j6VvU3EZmb18W
KYvfte9rD8MRQm2oZtTt98mcyapfGp8czjSiHOUkfT/Q1JxopTKDfrL3Sroh2iUv
YZTqDm3nnyT2utod13oMh9TXoIRaAk81+OlArUu+tBRcfiS7jVCcU1HNS6YwV2c/
w8kTRuLRyQ71TrI63nkwbi8gXvhiAA9W5AhKjakwt54nQiKxMJ2yZ8DjJ6DqSG3v
8GEWSNqu+U5QhybdYr7+RQnsYKZ/idweCHEe31pbc2+t6xnd1aCHr9u2cE84N0k7
/rr0fx+FtgimGvG8+m1eNWDblJsVc0LAxU8XM/u3c38dzkIhYWgqX5mrcF9Qe9/B
R0pDyPYiZByD9uqopnwj2G1M2WfKhFQX051wJkwRfDBsXPz8sta/JIQH0QlGBAY+
3uSbt5PuOC2Vlyv1Os2L91/DPUJA4w8A6qGy8xbqi/4/FFl4lxedXg5B3cvxFJsT
B8eoGitEGWPQT51Bzh4LUFbkg3mlHrqlZVEwBH1/RdJSIP66rHNNYwoJ+6QJtQT1
JLLqv8gNWOhxZXhiSAZM+t10ZQaX/h4GfUsZ7xBOzLIK74J/+NutJLW8irlibXT/
SvwCoLwKMpdl6jqiquTm7qBhcqb2YUNfQLJLSB2iYVMQhaxrG1FNrXbsTpmxSELl
p2IpasibwT3BX8BkXY3unw94rZBo7XOjER00ph+OsnID8C2z7hqt4CoN5AaE4ipG
hxF8vdWBj2Ucay+asYSUbrQzezTj8evV4iSJN6VFO8cWXJlIBrBdDBCFx01bC3bO
wfR/lnKkoyCq0ytKF2RP1ysfbDl6ULRvp9qkkGiPbHKMttTQcHGnpv++eLIWqcRw
SlpwcLBsJ7PkZ37ulr3q/3GK/9xvcQBsrkv5WM1UO3ectofdlQFIBa3UMo/HXE/O
W6k98lQ7qvTYXvnHikJH2qtkNZdXLQ4Ru/zICMR7rfaTt0XuXhZU5epiG5MznedQ
AqitiTImeFjJkx37VaT9k6bfpFcWZaZjoLpV4+bW7C5t1A9P4b324f5maYWr4Zfq
eEr2RvGHYpj5Uqy9lALMkBcb0U3m0MBrGXMJ2EHneHJWTDr03CVw/hpDPupSyh27
WhqeM4tG1jut+f56Fk32+6/HAesUcb8k/W9VYWKNbqBBvD5VJ/oPflkQNmlr+U3t
fBF01Yt29Sdiqdit3irpcjMEO+vqB/WAgXI8f9oJmiUhwa9ugPR13Rm9d4sqRrkH
pSsh5pcUMv+7Vgl77S/j3MJ/8CiOmwNx9jqNPFNCrJ3TOq9aTl4q08wkJ3t4bKAl
mRlMsTCpgx8AObZVPj0pY6lVx2hljTOLLnbrrgGaVzFFsDCVNSFLlyzvUzsYxHw9
owlzlkAz84ovSc6tCiB5ppXYYRD6C//qLxow9HBz1BpQzdIwRjPsbeSMs156PHYv
OkS8SxACZCy9axODuUU27Gqk5OUqlBfp0IzSDdpkvXC1YJmG7R4Y7Z0WMWmpyDKW
VlONOH13pMdvUrC/1Oo24y7H863qIPmYh9xbGFNtTB4LXoP3pBQ9rnIxBqf2n8+s
8BaBKUGRlQxaFsWiBisjlPAu4TB1tqkPlOGKnAuAt4W/9pGAbn/gEv7rx+6+lu4R
Mj1zk9pbIDbCIukc/uUAykS4ax1ClXLqOSgU1jfxirdiPvN2Iykd3CXkNoUZwZmi
e2ggUMbt6q0jjavUBle7zn/GRIqQVVhAj9zFP+Fhz3zS+/4QGDDRjtLZjO0yUO47
bpUsYsKhRc5RZUcj0kbjr/D4vAfqWrZqPmI+5LWJpEHLyGVekAWQ7rlRcdtZJ2Sq
c63ZM3qqyOkZWw7bjCoLsd1vDBgg/j5kLEBsMV78r1s4uHvtTYX23hcIz97V8/KY
Qs/ZjEIt8o0qiD36zpaxNnuLix3b3ei0dJTIsXBFA4p0fKYH4wshJpJzexj6hiSp
S/ODI519R5MeoN/avxeO1KepgCoJKsXK6ekVpIRpe6TIK/RBAIA8uTkrwC5Oc8G6
TvpzbezLPo/VFNh16lMO1Q9l+7BibZNQzt583OZrxkXKoQkA4mKM5UJwgZFNj2t9
zu3To2O/9QfDWHX5TjDpMwGK73m5bYlhaZ6SNcBI2flFSiseGQ7ahc39czUle39r
s0p9r5T2I25WBL/7LE6dgSCrBhKRLg9iR+/nA1xFvReudKU0UsYJW1aav+xCApYt
a9hIz2BmWdHxZkq0sn92gnw/MpHd9yE7AkXXDDLJtRcmSacc619/zTsIq7u5c9Qu
JwMc4BMU8LMyvHomxtJQg7mC6ZWByG/LY9cnDWVz9kqdOfmrCPENq9oXRsrdwEYS
4iniiIdn9esZgpmfYZ50D8HmhSkaSPCI6jGymU0mQQkt0EGoYIsOkgZQQDEmOfhv
2eZsxAydU4v5C8jr1acEC6XTsCxtClU2sBNM0X0FRzwsAjgzAxTE56iHDf5JqmhU
+zpQoF82qoYNCXVx36T7GtcQo7r2NypAfJKlVvnzT8TCbMJkwR03UJI7L+TQFWlp
+yiM8ubS8ibwtLiPQzIwg1UDSQzbIQ/WaSduZhrWQeLHy3k/Q2VTghw3g7cYKmGM
YlAau601JVTlGAiIJAeWugwQC4wPBM0z5WfllpKv+OCPMt6uv4Jl7CAYOGasWrr/
FDu8mJPqSTflUpTGQ5hAD3FyXfbKnR8KOlV9EHo20DvQFudocliEfJ1yjh6lT9fc
68S7570sjM4ABJSsnkHtaZv4gkFxrtHb8FCHNAANCEflteBF43xrdTqbq+wFGs60
2/Wsz2txHk/T8wn43Rl0zLhtoE347Dd/EGws9S3/gyqb3rAzU6eaMeiBvSLUAcjx
DshvbXa7pEYLajUHtQzz3o1NFSpJDGIxd1nemij+I5gSKKRVa8uNm9fIvRjESsUi
H4R9mD9PU+lscKLbHUtWeZJeIidDJ53M7cOQ2bk0fIFxMgU4t0Z8FjV4YIzarrs/
O/MW8eYfgcFFq2wEUWvq8Any9Ak9PkvpotjDeLRnAFP4ZSS+SGt/QdJCp7BNkkLY
0VWZzfdGCnWVgIHzGC3DNfSa6RMp6m2w/nE4VBDuaZuNK1IchhFKnqKWV349U8em
o50eog+ti7pNYKwFyipTS6bmXyAUdq5Cc+MoBlNrJzFAoQDEZqsmJ8OOusRVjXYM
OHOFjQRAkjBdDC5S9Jea5ZFUolq+iFxuOCDrMJ8UzZ7BMsjDf7netx3Qe9UkHbrA
1pyw+YY3LaAMiHvMZzf2OQyvNs04TySIxQjdBe6+MGm9JjEE1+fhSlBydLZFKqLd
fjkI9MRG7klwKVG9y0TfqfvnIS/I4GIMr0txDOO8knkJ0iIDyhcQ2fVbw5W+nMMK
Onan4ii80yqxAfHjlGOOQdwWV600z66XxMKBo3uaxOyBFBSqhEX883fXC0VTQ5Ac
fZp9xk6yRv3i5LL8+EJw6+IDF9BUaHy9tlFtp+fQpZhhSAqoBtaksNx+zed7tRrW
pa3TY1eW54xKe5HkexVaPB7TRArzC4HgNA+tjSoIBEgc2TTtTpRp1TroOVqYSLzK
mQr1Yu6y9DL5qOCVV09AWnHoM8N5tKWoKSzlSsmB1qDuIeCV1j309E09MpHJxOIJ
0L1k+YK0DCM3o7hXPTKJDTzGKNn5xUE4qvlRcftw9z4mYQ6p5k7wo8QEE80nYdW2
Y0CERz3UAStLt4VG/oRL/uSg2KWBgaxVyW5esFStYtBszDBVjta3o89YXcmuQjes
/Vpz+tgYdA7o62I70WiTdjR0fru+se3IWuaHAYqtB0MEkcX8fdvhYXcC7r4re63v
dQ1XOwkTFyz/pJkUZ+IoTVxcuV+iUZR991CzvHBeRwP+i+textjaPAf85/kGt3AB
qUSHSa4Ti33FyQq22Y7IRkDOqdczFCUtKoQm9OAwmII2AIejwaeEAe5bbW1c1egR
NnhnoUZgymGtYvr/YfLtkI2bPgRpitG8dLZ3zOV6Rg+jSvUB/pMyG7ktYLQLZnDj
2hXUW87uf6AQ8kfkK/rs8aSCSsAH3sBIMGn32WmH911eMYLZE0HiK3LQHRhQRESL
X1ehXFGiy9J2gUMeZ/5qavcHG3DAcR2GjlZHCPVQQhU5hzPReBskbDeKh4rZi6VR
7khk25M3bWMMxNustYOcxQN96+78UQJ/DRAXi4wYTCFiKjWdM0+4qM571BStJkel
VJrOUByzW9+7uXnERJn98vnw2vhnPKngBxx8syA6kZdVz1MQeBc1xC7dLEZHlIRy
w6FpI33qNJMokhcLSI+1H0u42Bc3+pa8z8D5Lqi45Hw/3EIOVxOkmnJUHI9Byx28
vy6v2+CFdZwEVcSnM7k5HstJfQ2Y1lCmha2JbB233shsCb4frOU46RRlOW249KR6
QhaH1KzZD6lp5U+zw1hdiqdanSaKDR98mBf38gIMBYOSnJYv2F757/jasDl0l0hV
62Plg5+qsdbdP/SIWGaqWTAc/pSXXvgd5gBP3ygagNzPRa4k7Z3MMOMsh6amXIqf
HkwpuZA/w6jhBD0onwEWsAk7R1GKIJQ5SQ523E3etuBRJgg0gEOMgZADMshuZmUI
TCLoKxc5QelS/xvJvirHx6t9VW/k/R/oCKb2m0GWLKHWsq+ryybIVejV6RfbT+5e
qPOtSZayMr6t48DVSUl6v1xdksxPK7erlVejwm4Q8orU8eXSHcGYKp+EUDHJ3Dfj
j1+TLzISkRV6OlBKoenuczX4h4WSL8s/CQpxMBhOpeKDxHICYkC2sbiaFFLSYhbk
LT1nxONEfqlEsAVzIuObrMz67OrNWmqqH74vV+cl2Y5b6zr01J8dkDf0e81Z+Tqx
cGOl1iu0Cgfw4wumtljJX+kuVGrzhPWnsYadSQB+wlP246y0BxV8tMGPJ8/PtHT8
1TgvDYaKxkV5OHxultMUvfHHbmKN4Izopi0eAVxOEfL7tuQMrkhTqleGX9C3MHcz
mRgnwYTh4pmNT6KtUq9R6zId3fXmqWoe4/2D4T/Gps1ZI17552peJ/iaUprvc2kd
NyiGs1jSemSYMFI4p/sw34V7TVH0W/CFdb2p8PzmzxhRC/9IwdPvo67NE5Ofnz9P
yrlNkw67JA5RW8CZNytPmQ8emsHbeeU/wO+4VoDHTqbUdKKxuHoump6+5O63AV5Z
GfEOIq4fmwhKdYZltCHZ14o7G5fI7mzYOMm32MKfXXUxHgfkjiFcUhFwT0nDEB8f
GYUDqLuCjgM21SPqvlWbqTfMDBmcRL6x0qrturgMFJPLjhCJpJOyMQJh1ks1R57W
p2zcByrlt6XO2jdRSzeGbT++0ckxGQtED2gmJPeoMEc76DO8pDvn/U++HJlJYZA6
+wGPMVghDoQ0aAPf/XVw8HvNOOdC7m05AnnMnIxcVPENoNIue2YPQtsdRi4S8ElN
TVmLmToRxDaus+laq2TuK8oU8Vcn9aO3sOhDY81BaXVciajDAMJhmXzyeiWSoNPO
XygFa86B5YJOUAGNjyPEaBMbaE7nBg3a8/xOCyZPyPFeuTmiWKjEAraduBiMLKrY
N7rjRaZ2Dm3Yr+2dnh5L6gsOJ4rgMoXDboNgKFITBw7WVJvS0KjQmsxdmpwctp7I
hRFfJ3HJG5oFeIwi/kVRDHDcaVw08hLiQg7O8hSWkLjkabzYD/FhR8s59SQm3XN+
qHv4XsZkOmuRFVqC+eo1r1kySWntUfwX40gMsYlv1vPTb80JLnVbOJb/dsEY+DXQ
9ispXZB12Wo9alr8qAnITS5ofZ1+OT0rF8xyCU9syxJddsvvr/0PTwmUeoWGqyHP
KCQJ/yqpIeqYwgDu8jtvGoVso0lvc5zCWLEWmzYUVLxjwQN6NyNTRjFQOyWyEm+v
wl1qPNsk88XyvdDh+CCJFFWYB9JKRc5gSunjYwEwnDzuEwLtBcGOC7RGHQ/vyaPS
Oon/SuvfjslfdpZ/OZXPQMF2AoZWVvO6CuHUBvS0dxoFr4cJCVDfly9lB+v75HAn
4pxeTXl8hNE3sTpySYzr8wIxoFaHD7nDxMJsW0KYsrtk3nw2+8qIHc3NML0mTNPm
ELJEfGIIpWkt9uzYktcNTeYWyp7zkaSizPLZt+D5gtHO9M7XZQFUeBMfJk4NjpVR
JwL+41hCh98BcaHYxCfpgsu6ZVBTK8SnexvIzK4AgEzHC05D1Uw833wj5fmkXZFT
xiz1UuV8x4IJ5cCJmVPh6BiExmer8U9wWhqg9KTL/3I0Uaoocvdf6E5TIiuZuMbk
4H4BYY9drfOseSmZqUNG9+okHydpIA1XmxrnYAKELWaMizctie1jTygjhnXnQMGY
hs4SHwC+lWQljuXx0FbsaHYPVEcaoPKEyLa5ChZW0/3YwB2HTLTmAjvx7LyyidiY
Z67oSqyqqtsEUIbyT7E/OS0uCJIFmpc3lt+OGzyWdLom5DJVXgVgEX9iOmS3vn9W
NRfsjoNbYN6vK1crqViof3PhlWWs4Ujo01zcCxhHXlNgqoarciIZDGmB5XB/HaoO
ZCafdYTa8Ed6+mS6BRHCiEoEGsTbtxZpdyt4LnhSGb/MN9Bh36rj9MZ4tnHxocF1
3MRs+vFEX+Eo0TQe6dfss7waiOcz51Q6NuUPofK/14eNg6FMaIsbnKbefCv2bD1P
Qyl6PBYn48QKre3mYRgMoBl3rsmyJcUdILW+Thpl+NuuAfsp77jVKVHTf3JPMu/+
V1UNlJoZCVeTWrdJvlR7G4V5C4bUOx8psJYwysswlKYUZf0mjMHZKKlCRbbairQ0
q7eCdPHjEoem04QlpRh88Q52iG8dIH1O8EdFX/7tRUX+4xum2L+Xw5DP4Urvf/N1
jxTeKrZr9akejtkd+9JsQ9mAJQEANFsIdwiFX4CIYoTraLuKHQ0vcRW8SNzGY60f
BBxfEnFozqoA9XU1v/DKlrKvwkLqkd1sXCg0wPO0t7SrvB+2XJ2mnS0io4wFOpBj
JyLiJgYqtjyeB1FSAnQ/QEuBcwFQSxj2Mp9068XF7OsTx74+i0GkLz5RCBQygmbi
hec6Z0K4Mj9VZCAshCBPXk0XuOq1Ys2mm309o0X/Y71zZ9fBJgIrMRAyHqGimCKS
j5BjXy4c54Q6Zy9ENjmOEU6OAeCPJ93Grwu30DJgH3Ly76WQoLLVjWPVoTnEKqQc
gYC6w2oVgiebH4Y0NFFKjVwVrJS8TbKZAs4/zKbJ4grF8HysUewoMAVQiJnu2OIw
Ow+RCQAV1E480D3Cgn/HNhp477+qQBZT2LFwjWcT27cq5Ilvwq9Tk5aF9PXd0V/K
a5AXQh751ODJW3gGWy0KjdwEcfdfhpRYhFPlJSdPQOzZqpIEewuBWoa7IRwsECG6
lmXqHScjL7H/oxtMSvb/zyHEKwk8565kKXZ0Tp7zQ8yRL0wutIhwAjC9zJ9HyLrV
YJNxJUrD0Ozw7DSBqKLcQ9RQP4gswtduEzT4Ri9L+1oc0u0S73Iy9zPJQ1qctl0Z
KNlayWJ/TgS3C65Dl+iZ38NacAqrLleXdYYoAYhc5Ly5JgQbgdfVYsUFsG+IWfMs
GnME8wQokdD3+SeLF+ZTXY5L4XzWs4dGTAyPvhYCMU9+J7XMpgVWs+U61N7UtasS
Y2qSq13C3MBsB5fuSPvOuYdCw2Gxw2R+eeHg/YPRyuHb7f5JikBvXQs/s4FA8x3+
z4+BaVxG806hVtFJkGeCakWAsZe+kigU/AyCHnKIDpTJZRjVC5mrruJv6Q6U4LrR
6ZVGIfk2OWst+/Ww423f7M0zao2AzjQdKQMCFKQHj7Y/8A4JKCP8J4Yt3yK8cTdJ
TFSP4p0RwA71JiVYaa7gZHJ3NSIxaR4ZfXhU91VIO2JZcEmb2xBlu7NUx3ZmUqkQ
0NlTAX2+qHZURrszIv0KoD0kaOmutn/uaC3aDNyfe75+A7aFCpWOg5QMLZ5mtcwj
r7NieE5cMspxXzG911WXrLPikz/LlLgQ2mqeb6IRD+5fRN7J3fSEofqTDL/EMZv/
Y58Nwx81C0sNzOTB8NJkiuxurf0P4+cAKvaB/Xr6mC0E20AjIPqlAySABFr/V8QC
rTQBKv4jC4jJaFLI44qelWgrMY+WqcBOIiOvpILnWn7eIZrF/FGXzjAg3xN8uVpU
6ZQqQLlg60YqyTiXdLa+im7FCJpVfUBIWjxEUo5rHB+SsAL6EJlXoua3ZK3GtJHo
iX9cg9sR+sS60/FdaQepAPR0j/EUU7w9i7SJz+8ntHJa+a1C7NrLp3g2MukQVBmY
Zr71jAgI+iNnpZFDAjR6Ie6DMIbj8HQfH1iUuTqukHndUx8Ms+VLyoheq/QEiP56
3+rfSeYd124cqMpIiH6v9/YLujukQkKTOsKYHSfCEVQeWbmieh33idC5aonxcMiG
Jke2r8x6cszivhzkWf3MVJu8rXrPeDk7KzOj9IqTS/dubflk0CqoRv0fcxgjyFs/
5laCdQcl0wG3k0f1072m18ieQPX0GIAbRe1i6IlOyEUXOMqY7UYaipZqfvDpSgpx
8cFGAuXT8/ENgXLpxbu7fP7W3jdVkRz9CKMve3YaIWLjJa1Unli3xCzWjgnQ2mBU
ej/OfUbmGeXLcEduSAiJVEiWfKt93qDDYBEPck4k46MiFYNH2U+yEyGFZYSKzff2
viS9aTl+PWiTcBpOGjOpZ26MhNUOkR9Rz3LIAGGG+eu2pOVnGDHw3ygFu+R+2J5N
8uE8nbeR5qqvDkm1W4OY7zREyfTmQoH5w1wy/TeAS8RwmG8exxRhuFcBUNVCgTz1
ttd2RQo1YMSpVem2Plb+1Nhykp5ji2M/EXqupkremB6I2b331sgkFB592bgOvIPo
nt6ntql1r+Plr1xi8OmdZjILwC6fvsVTMw7Waf6q5PyH/R/lEq9dDAwgNwAUJS6f
2k8w9nfUMWmz93W2VvRiwzuoIs70YZECKq4PFtAc1dDO9O8l+601M/irR56mt9B/
CN7divnMvgAk5Yb0RPIgleJwABENDGjBM+0XvFQCmbgt3y07OFURqmEg5A9oKf8R
7N/Ak6fl91cc5OIorcwnBbkh9OwDzlWWYfk7Q7G1BpYuzELI7R/PnRzdNLzJmunE
r9pbmsXAkb6xUghkzdXoJRcfBqUZABAkMUN7/bH1WIYWXywYFWPevfi3E58bqiqM
Vvm0bsNTpLv+Yxz6qXGG8/QcaAkpvlS7tyeq6ld6dQQUbb9Xn8K1kBE+0HOWE0iU
0t4cUAvxVmepmBlE3ok30tcjf3FhZ5JcJXZLFP9NuyKXzUHlKNM8Ob39YDiv8gS/
cAdGmyUSU0umbmPAGvuhiigR0EFEgDnLwVrr4NsvCeQwLXRfAmCVAaC5VrfwLRfa
/uboxoepSSFd8REgHQoa80kqpGAZpwcBnDC/TVDMLbK+q67F+Su2/WhInt2eq33X
L9rZp5IwYA/1jAUkqHHOoQn1xXE30IEqFOpcuZbRyk47vGk8wwxb8UE/TNqtuilv
vEhchLH5zv5yQD/9L75yfW6yUw9wHDUxiBZNk8dIAabzI4JAggONOu3L1lmniz0V
0B8VPHyxQWxBgmtAQwsm8VXy9UPs/WOKpAgw5HWXHYuQWWJ3ZISPqOhgI90uPqOa
TuwsI49RnqpHbO3AO07FtMUK2WpIkN2AhIZ+xsUpTei6PyqvgXB/FgMXLuv0IWtM
GLsb1mkx5vuirKZBi/WYd93J/+RLuB4lNh+TLxp1zwP3sl6rFeWnIF5slCn8UBFf
GckZME16NCt6v2Sry8VeGDJCpEvb0ctblJ/P73+j3CLiIyaIU21IF+2GgxVuAFSe
KAMAzzci3byYs627ROK1Pkm/y1m6bewZrOEof5BvQZCEZksjilDJb/FdBiGs9IWs
aiHi5Vbco+lyspM0Dr89oYsHwZhLmZxXixv0IaLTK+5caAmmj0qUeLZ8rbm/5mlW
nJ4N6IRefUe8KhkFIIKhhm97MpCAJIPbsSPyPI+2RCQHwMLF7sYko6ZO551zOZta
ckQyhPtb32INkrS2YFAjjQoY9PLwzWcCG6DYba0k9yxWlcZIHidzvoV8HtpPCLg6
7D2z2qJDiTVnoDoidJx9bSq9AVXsrnkJPkQRQaCOeJmbUPdlXi470CV5KbPpkZqO
4+utdonRhnuJMUpnJTOxziwTDlZaGOSVSw0QYhbn3gCHRMBYX4CQaD1U4ZI7m46F
kFRuDIRu5zuHRZj71nEbD5UzLxH7Iq69ALJ9++nONY3mPgc3PVG3WBHuzsRVktHN
TWPVY8HHCKLQI/0261wH2AFvmO/hFZaGVRRDF/XNhP/xEz4xfJZnevh/A1YFouXA
R/So2eq7CIRsUUZSWhB3GFZyIONx/G5ncr51s92N0836K/N9h52TLrstzxAobrQO
R5bhROoc8anTRzFWmmSb5O7r/8BPfznnvMkFXqPkJ0KphywcdZXdyLY6oi1ipQ7X
0U0oo8vHJrT5CiRwvTNpPDd6icqIlfBiWHdEpkEIxi20a5BA1fPWeR1p3neqTUzD
BplMf65w9n71uzC0m/kMgqBgUeA90iJN0cKenBXEzPtSM1FYyeVz9JCrAnZSIr6H
flp6JePVtbfIHNg2NhCyldhrzJEMUiI/PFOHvqDg//3ipZPqLDKhzaRVWdCKkNTO
BFbHoCpxHJOft42bijNFbKZlP8q4bLDWGVsPqf/kYEahyCNSHnNhxezplBkwnJmi
DDKOfwVTBuRYQMQQeyGTx41mHUxZ3juYb+bglxLaUFTLYdZ226qVHQFv6u7YE4Dm
3KCnJ1EOr/j2agNSpfxaUGGSBSRQX5gf2lHaUNpUePQb+hysMqV7q93UDCJhGxNZ
IcxHfqLxdPruK2o2O49GEeGUYVJjnr7HCJndYGiNaiVwr9ZYuhUujueblPoQVjPR
16hWxftpPweH3ioGPCS8UTunHzzNUqdjEwsfUkaaoQ/WhbT6+eKYo7Nqm+/5xAKI
kLFXmMGrVM8WlgMkdMLdTdMmIcvy4SDOjinPODd9NIawhFEYlX8p9qdDdI87WCRn
GKKvxnlW1XChd/YlLnaSm00rPdoY60j+9VHnzVCpxJ9DhFIUHfN3gdjcervJIW0F
p8iY6vq0GhPp8tlCtHJMpCGTMIO6pPEtbz4Yt2XNd8uSgmnBsklXHs90XqTwrzjH
kW+hPoLl9XB70U5vB9cjiJtwJsDk3GeDfIo2wr6XB1Pubenvatk8jNjWYSUg1c/1
pmin9sJN91Rm+T2i7Cu81yGY/RM2mA9cSdo3qYtuXJzxOMkUx2Ic8VPgT4CbPkHG
EbmJGtrP7tyCCUDgIY7Tr/HaiiAn9TnBJAyjw+WzhePA2MGTQoQYYejb5aw9tK+Z
68aRsIwsZxw0GtInHPz/j+JdqX0tym3KPe5v9mjBoEPtIzdQ3tMa8PUlQRBfahZy
5IWi8mCRBpmLmVtxvfNgQYt2GxA6AsG0Ui/YaNxTBydWsqUBpcSrQLfYz5cPwjLi
0Oj5LVmhA7hRTMy9wyCvDNBuGX4HY/shbhfU8tIJNu1NRuf+uo0bAB7FqxM3wN7n
0DAnsfEfoWZlG5CvFlsR9zLvsX33Bz1TyQUuTC8EiOYO/ZJojwO34jpEIagJ2G9C
rkGTg5IB1VzAc+9/UY3KWHAvjQ8hT2iwKH0XF8Pt6f7P6uVY7UDfcOUffTRJwNdx
M4JL7NY5GUrwKZUBwJzDJUUNBJ3EZbn5Fjutr7uECVwOTeOYle+qZu0sNPxRUiKa
i94JK2/1kLwdYePR8SH2SBFSXjFSEU/6UPazHI2SzEmohXrkmeMVfccd7aH1fTRe
MC2yCtbxAs1rIFZNJJ76/SDkBw5akgObJi62knu63fqkb/rarX12/AJ+VDCzIhDn
ExvWPEFnwLM9bY3p6dvZeiIOnTxC0LAeC+2yRJ6nqr46RiLK8rfQcanEeqPFbb8t
qwFu9UTSh1zPxiqUTZ4NcKC9blud8CY1XHNBOR3wPCelwtp9PbBh+BkGWYA6XLY8
8NMk6NWD3SRK2wpfPaBlayV7V064aDc/gU6iLdgzCFsPph2T9pJ4KKUMB4PbCdIB
z8i9qYl/ULUXtIDPDiNd5C2eHbrNo9RCPews2ipaz6AqBkmxBKFqcPkczsMhu0Dx
8cnbBr1Fq6eVCAqf8Xo2hXn8cFCcNkdhOeRyG1xVx4oXkHbQCoAMcPjAJZmhNUQJ
8Nc5EDRZDF5H4Po9sdl+Lg3Ot2YZ59023Ob1mNiz5YFEFieqwgTTY947Yj3GpWbC
28fcwWAQE4OUQF5mR2olQTFxHYtoo06GJxWwTz72DVZbq9uGY83aUjB7T+yETcB/
EHTQO5haA1tWmGdJthNA8Dxi3Lr3iD7NxCJEOQmbIVUSbAcnmsgx9u4iMFDqSDsl
vVOfjs4qK8SV1BmrzyiLo0BIk+O1u+8pPxzELXkeyOCZz245Pu1Wf8neI/j8h+Fs
vzIg3M1gNnpSZxazYAzgcQr1s4M4plBHBcQAt5ioWyIVqvNo6AgFzp+aTdy5WCe8
Y5b9x32QV4Po5bUykix/yuXAvRhdGqdnmbsHZtka2F6THCXhFJPDDHHADBqBU3xl
0913U/s1nYi/lsDFr9vYUaeirhlq9W4ebAZOaZPlbwZ9QF+y2U0EJPq1hrKCUpfq
TV7xUMLRS7RGD8dLvykQ5hRilgC3bG+lgG73qc58MwySdMK4BK+bE3O4s70HodJI
tJpsRE2tiXZVUOzfL5LzfrMpPuUBZyxryHl2nwq4q4I3jo57YI3lKC8gGQ2XSyUV
vvDEHddlLCKOzDI4euU900HCu8+SHJmgtIG3W+OiM9pC72AMQ+G2m9KLtmJsv0qp
JChXTuu33HQWXLaGQfwQwHlC/yZC5qi52Y0uZbTZDss4dkpBn84SH1GJXj1xoj3W
eKuQdzZj/iyA0xySwo2FZGoZUVilh1/DCFD++UUI8XVJxS5C/NzsJ1jMYT15LitD
ZMj6P6G5mBvrC4MwK+lW2L4bbYRrXEcTwpm1udCqrwFURFINeh0a9OQGHFhFakpe
IT654kTTjas8O8Zmz0/D/XgKY+t8K7eXl0TENtQKTYcnQiI8GW+SDlD1O4XX+SmQ
6R+Zq4cnOQ67VNHzlyLezpSITPkDBl4cDD4p4WJszYLLSuYq1ou1NnRhIYV9qUDV
L/cMIshknRrOPuoO5Z5UdQggF7tBQImG/eVaFr0eoFd3+J+Q7Fb3eaZS2nsaNDlx
Fj+/SLgBV3WU55L4LCAWv5b7lAA5YlZT9uLsb0Y5v7WhcO9eA72bhN0S/BJhvfUm
K2jDEEeFFnzrhCO+HD1He9VJ4brwL60WcfJY9rnO6tUNFvoKBi8YYTXMaOIdQDFd
vjddkJ2/CI62YMeSAoUH32Jka7PeX03CAOu5wOb42WdwTh1/CVAHTLjTJC6DeXml
QWUYoqctW2Ci/rptU5mqs/VZe8hJ6A3x9YH0HvWWu+oK/Y0cmzmKwTqEFPhmFE2d
mdG4hSG/rn0ity/+sco5x8wfLr7xIvOJTHhvHmltsbl2Jk020CTBAWwiARUKXmTz
xGtZTGJzQ9UGCZ4MaU9UnfBzRQuGXEfJPObocWu3/j2anGhfA/P0CEBfXd83a3iE
Itm2rlg9B6G8pucRP93tx1+h9tSwPEJU56rrOvU07CdQ0hdVl5YxMrentKf5E4XW
3Mbv30B8yflKBTL842W0RM06RMJH1g5xWYtlDM6N71hxTW1xQ+HRD5uQ4VF1Yh0u
VegFl8Urg+MiMqsZzCwc0yJQtDUjnEBEeaOcbDpVCIAVOIxxthtvoGYSkrrMcW3Q
qBVUxfHmdpXsHTBEKesfKJT6kwf8qHPlfY7TbqDWSe7fObQdac7I380nIgWMcmQR
M7nu5z9pxvisShQW6LLMSyu5UnoYYdAYNaEBoEExwZY7jw9Ew0Lutln0iBHrmzah
4M4JwYKixmA64lXvKVz9/VFZHFLxff13bFUpFcgLvBnr2KIkSx4dKlwyNz81FJ0q
1w7Cf3PRMGdw24jJNpHjI21WdnIsNQotD8mLihThcPuPanlnij7ielGT8i4nYOag
VKtnAJqSNH5NfezRGAbwGdbIRFkzWaVzdv6rlgoTmDUWSmduu8NetjnsA92ENm4h
8dBzazDdHYE9COhrPr4hx4fQnosODR2UGJaLhY2d6MBkjk55XnDkBsZyemqu/Jky
5xGVs7gsF312ubnF4V1LYit9/Sy/khQvHCwjpGt9LzTGvbJS7d5ufFFkzdoEZIOo
Vt3Yef3EAoYxwZgrE+UXKdoAgu+XlwsZioc8XRCJF8meaN7x5h048pqJJFcP6uQH
HP1pQ7Z5xx4gwhERsiL2iuotfBOCQSlOhHyo9IBr4ca/jOHE7mj5DTFCcEuNKG3m
cibaTblCyTxi049VC1HiBr6YRgNn6kWHQEf/LPj4gYmV+1YOiPxRHKdQ+Poqlysh
eMKJ2Vi3T7LM4XhV5AovEjuCIfPQ12Z+z3cK00FVflNAqFD8a8Fw+crbFYtzj9o2
e8pIGEpJlfBblEHQlP2Lxqv6el2IqZGqYJFxCiDCkHOjNMGp7mOw2JjgPm7OjXqt
85GepnDGqqslD+ftdh4zTeUmgJ3gJuQz4+HJv6Gp/eu6dJ57zr/++ZKgVvgB3lIJ
TOFZvjIhQOdQDTOrU9aTzNPh/OjOgfZQEg+LUTrQSknyNZp6LlIREuPA3Li1Lbw5
OrngfWGdeUAqMY7msQRxEJHVpnUnmAlhMGL2EazG5PEn8FSbFYNajDaBXkRfAMI8
PWwxTKQEWzEONdmpQLoOR0ehTR06VlqCPWF+DLXvAteNCfrUzfi2NUIzV8G1x+bu
GGjTfB3fJwfBRadYP4az7pvEoQ8ULtYXaPeM4VHtYzD/KuoHNj/ym0SUmwOl5sKj
UKcRNbg6YeJiETAKwFIIHhIP8qqgV/mBfywUcVf1/CCJVJEKuj+WdtI2b+MY8G+l
ggEuS0sjCTCkXZVlw+s0Ry3oj/A2bcvylja6r5kNCtcVd6CmGg6YI97Ge02ggM2w
xCrKCKJq5DZGoYVy058qadPN2cmWEz7VeMglOmW1aKag3+khDR9LuDr8ceIQ7FWX
KtA/5DDmeHdFcHS8/mpnyzo1WFJSi2HP4flunoUZA43Nh7FZ31fpzmIt/OX2zPjy
lR7VJbxzZyZugkKo9pa39BMjb1jOoK4fgBSxYXJrtkoJa+g2DkaaeBvlFYV0W504
UDoc1xHjpi5nWYHFb9QlCPjrSFLdbU6eyOT/FdqRG8cmrI/rq22Q/QzFaoEV6oEs
yoBmxxzQ5l8ju5uZTLyR6t+ngbP5xkbyhaKQNSA3RW2+7mLMvuKLQ1kDlhc1AvNf
5RVxC/i9DW/6Jrcgswfe+NjS2yl9VNmxqdaOaO9XP4kAbdxI36cEh4UFzcZ0XPra
ua/ZOtxoAgZan2mWc6bxoW6g5Ix0E1U6rMe529OGJqkyptU96X4FO1ZpUkXt6EBZ
bcghIffi5uZyxx1evBNqcN4heaxOXSnrkzI2cVFaZUuMl3GJmW0tD3UmjjxCOpK4
UBLUNYjRIO/yPkbTcX+J5o4jbGuskqX48b7s1ZQMXD7GGWqYUVI0pv4cvIg9fqRO
ltg6SKz0gchZYjN9tF5aDAFBLS+iSC0DLivjd516O/bDAlcGaED3kf880C5+ueFP
Ey7p9UA9dyDckpkQrWi4sb8H7yNrSzhGHzWiv2HX8BwxlMLqMhQxpoe9kP1+77VR
ElbM1D4EP8RNQ0NRaGF4lK+1pRr5x8HsLQdsF3zOjPixbixObC0Cl6rhOjuDiAhk
30WXr+//7b4du9Z5aO1/kwg1zim0k68BYPPjV0Yt2ic3UbZKifRCmcE0ptM0VsZZ
cb+HsI5o8d+yBbwU7fKe9xf/8oLN/TTddlcPDr7RwFDdEcXqI7FUDN3+ocj8yDhh
uBY4Zqp9GYu9ZkrlYGsgL97s5igZDzxn+XcwYhHgXYAx+zAtOdoqBMFPEtWlzqkD
tiitn+azd/4V3/vVmEmBisMYd3I6I5spDo41simWl5uNHN6fvxfXkvzzjR35Znlh
wqcTtdfHyzNNW7Wlwovsd4aNrT2kvPKfXD3U4IdlK/l2s645Ux89s3IgYJQwXaHI
UjnjZoy9tIClhIRO4eEAfTBMb85cx+uKOwcVXj/FWs2y74u3w8XmHLoCQrzQdSaX
txBpweG/uxL9DN8SSlvw8kfWGbt58KLF9BxtZEykIUHVppIm/znyKFpUZdacA4cC
gg9/5Ww22GSTI3GWu64b8VDHxGuUYMXrR/IA2tJDcbRb0IM2blYBCjXhCQa7qh6j
PJE4BrCWUufV0wCiXwMXWZzd+1HuIqvBowy3ixInoaMAkPcoEWnjEXgNdKGYBlOQ
rMhjca4ExgKXx7Am2b/NbZovmpwDiYUFLxdcxvlsglOZQr89JENPQb2G+HW0LHe6
Gq5CC4nlA+Uqmnj3veU+o1xC1OkjeXHXdIG7C5prDggkjJNsa5CEwUF1zZdNayQ3
pWrAsgJ8mBOa0FpsN4PhABgT8EGj8JF/xsnBHjRlhQNYk9ysn0/GQNp0EYhEHH6s
R2NGTilrIEPD3u9F/M2qMsKzDrFJliOGWTJW3BLdr+ZjSE61BtOITgWzSTzCrif3
AufkCQlfqT6aKyi4g4PWNxCQeMcOWWUmPGdipmv+Fs8Sc6Rsx2QWRNqje3J7J392
vO126QhLcgbUSlyg0qkEqcM3znTOIxwQpoqbKQKwNEYtfBjt8E4CU7FKc40IYsXp
fYYKxot+nm530eJOIUITjeb+NW1R++zJQpZpphsCK7yQ0HakKUgmQm6Jm7TmYVrW
6+LO9It1+1tAas17TwerGhtOy68tS6GVTejEWkLPxZmpSaWz3WI2AiLYMia28I3f
pRFZpjzbDtx2sLz9bsuw9IWc6uxyb0zGM+XY/8On2dkUgaDLOzbFscK+cNp4hHAs
uSOlZfAGwDgNeX3S/PdySSqzOeZhl9VssWiB7RA18XhmrU5wGzGeOtWwG2FD6XoX
OIpQ2RppEx0h7Ol0/bVPwiP4Je04/6AFuvofFFGlbRIgTybOFQ4sW4u/o+r9WGbS
mwjmeVWmplh7hd9+8WRZfIweWUBXeXL9wqpEEWUmKs5gbXffX3EC6HHL1NJr0hm2
eU6nFCxpyHN3QQp7SgvXo8CfFIUYB8IOouAHO+J0YeE25R26K/9BBKgOiWPfpCgF
OOsB84TjlmRBw2p1e0KfbD4J6rawk5ZaqpKi8EWP4dYleklr/DGyUSxN6dyM4Zf2
EHzL6fYF8G+pSjSu+i/dkZZTZoEl39qShOnGXL0KUj2GfjsO6A4acv2WZpKY9ZTu
m/5qU/+gm/baF8gGr7MnDjps2s1F1qNtgC2wSrGa9E77DvlJNkazQjxBPzSjynXh
7ik0dsEBOFJFbM3axlpKgqkjC8+1Q9muIPppYaUkGwV9/6PMlgfQRDXWyI6JH1hI
T2dST/GRedbE8ydEjR8Bh4HOnsczRVKwfEFyWs83i3sUH9SlnPvYc/kkxCyAnHZh
2HesLdU40hoQy42HjKL1lFNZ2Tb5AXH1NMis9xzN8UpnWCs3NKPYMs0YR3nFnq04
5ecdApW17+aUcjsmF5pWhOg5yUWwCRSM+Irjl46LeXwdzuWUAoxPfdwDCRaA3xoP
hUq1nKs/xxjMPHWwmzRg+uZw3kuPdG/0on9N5/T1gCCrMXIuU7qKNAur0AgVmmWO
zhKdAviUa23OR5v19DMnaSHXzc0UJnUvwWrmI2XQDiMJFilUNnJTkFCwDZJq3wLN
7KuNT+ZUnJBU0g5O1iPoyW5LNvRqGfJG1RGleJwB4rJP/Sr3lDbkwQyebnepYUky
6LV3ERNiBCedzHLRM/n7vRFa2rbAQhQmgXwCujCYbCDLDUzCqNWXW7469QFArJ0u
0K2NCGCJ2LigD1f2ff+ZVFOgauVVv+/am1kSQ8R/6DN1wBJsB7YyTjgz/0HbVpWJ
Ym8Sy1TsEzKKIDWFCX07eG2H6bp+ujv+DSSZMHse3vtOJF1E5lstqJ6ym4kFGwkW
tV45+vtDN9xdp+u1Z6h07Sud4q3jFj8iTFmbqNHMmNWJdrtdKMdllXB4voyrfkTr
CftWkqQqA5qFJHWrgz5au7Xb8IihvjZB9hCjz50rNKcIxjFnj/VUz2CFfC06pUGE
9gX1rVoYZqeIHb9JjWgC8FEDeDjSDse4fV5vsfUkqzfPfQ3g0WcurcoLg1/iQ8bm
AjSk3E4Vt2HBpvEpqCOkJ5k5QbUh7wsu4FY+7VnGK1qt9y2rgC2i56gDi17lbBCC
bSmXCmaa6m9RPCDRgd4VZVxbe7aou1i6QRyqhmI1YgG7PFZL0OZy31FyLyERcJyt
5tXUPzBI0fwiTtW7S/vIQxPYSVMdg5P0Jy9PRDV6/mxEgMCXx/a91G7Q+Z0fBPWI
dAlTY733nuwKRyFK0zVoyksCAjQ9Zj6va0D0bsYEFcgC7QY/8tOLKHyBLOV5E05I
LoCt2+t91wy7TtuX751sKthImWr335TEEGkyGdXXUa4jkRQ74m00Xlibsz6GE+u8
jgJ8vZ0/LCX7nqTVGMW713O3ijgcmFctUxi2wIxIUiryaJPWxfbFPU8sMSM+FBqz
sN0/dRGwxLEdVDzLqJnRyart0XbL7Qmk0mojN4RZ8yI9rZLSlXYXjtQ+8/2nyt6s
/tugNwZS7EORFUj56FrZ4L4rD6PDA1pzvXWV0ZTmDvoMV1iWbmL/CnkhWRlzHn1Z
/71+dm4mua1XlOSznebMYQmT3s1gQlTvO5/KBFSa9ERf123LQtdRYYFWPBL3rXR+
4uB+suSW/9iufYYxl4YH0IS075FMNsfXkF5/2SHKGcioKSXEiqUFGYXbXC7N+jYJ
A7IFMNT+p/IgeBKhX3y0bWXlRY5TlrTB07Jpy5DwVKnz4zUT5PLbxNYzaYaqNav1
JJYbjputTxevmgNkFE0Q5MJ3F1ymKCVu2O+QEBSkB1/eXscWw6n/aldvCRQtTq+H
yDkPpZFvZRcsADO7jviHH2ovi7kSoa/beJIXfHUBPmJJtk3IzdzfONGg5fW+q/xt
m3wgopGP3NpfBdVqEj/W1IO8k/Y8BKoP6LFgKA1hyz8Yl6jh3kwYmvcdFbq92AZ/
BH7TTzkS0jvOJq7yNmcYoe1Bh420pHk5ob+jLa8fX/6gafTT3PSwLXtAkDOUqavn
F8Ww0i1JX3lc64rCKzgtLQInD4AGbQZRvSS1FJumntp5UDi1TYWQWoJLkt6L0nsA
8Ro7Q/3ireKEgxLMgl3gFfCsWsGb1HoozQyIxzGrjdszvuEXcUzabXRphLh+D140
O+TlylDi9eZ0EykvbD2m6HVtAnagOAoQX+mUilaEJkwP85fqWVtzwj0Zz+5Zm9cO
aJoeTFu2TV/nV5GPQW0fXZ6DodBhtNN5Q6twHhu+SNBfYnrKQwVJYYw8nS/ywQoB
oN1E7ZDsVSgXIf+CrcrIxZIIEArPcb2vkGdo39qZuASCvVdcDI1ELUzDWZbDlTC8
LWIlZDtajvmUIpTZud0MdlWPlC1KQzjS5/DioHTdgSqWLHCxlw6AzTRXpID2/ru1
yI8kHmtXQQhYFAL4ZLWJIX8qlH/3sjv17Qr2KzS0302hm8KntaxVjBcjvaLEU8Hq
7bSoDivETYV4HlIi83BImkz1b/tZmSVTdrFIt6D9iO74IcniCJ5ajtXDhzTQ96gH
XlIGZlxTEJElfueJx5+DR87+Y/Hpx11+iUDWYIvwx9jgAf9K77rBmMZerHft3jD7
LwbVkezP+KC/e+K8ZpqjyWVNWenNIsyT3x8J/tg8x5tF+DGISykrplmebwXxH10k
WOFwYOkJOQWGRX/HNw4AlVH6gMHBXILf6KymjUL6Gexf9qNvDUyLvLAxxa6ZwGHj
ww59PhI2tdA0CqRLS7LDUW6N97SNlUraDBXDPgFEl0B+4lRpHvNU1yLSz4HmPK7i
bhJd80c5DnUWnBZ7L1njHYhUp2e0fznUydpWbODzZeDA9y9gvXQPROnDZuENC670
bt1bgAvhsDsOHl9nhbkCKJ96HyXzgMc84XHary0/HhBPYyg6srpCqu3Ixedm+Mao
28fVxOUBg/55IPJaCxSw2yEnMSGcBRXlTBbq41EGPI+fPT/pualJRSv6FS8juqIi
dNno0SCL/ZLtv0TiWv4ae4EJP6rxqjriUZ1dpSyydopHu4rkoFWkChBAd5SWUV74
tpOUYDdAIpEOZx3R4BFYePE+uABXtSvCnaOrHbedG01V+P2TFuZ359EJni+z2Mp4
022nyGc+IjQ38xmk43bgO5VQABYUAoOyMEj+Q0S0OaTpm4DgzptPwMs83E62jEsb
8Y0zjaax/KU9bw7UJLUbZMeAEUL5aLkt401fnZj46DP60eJDetR7SpIsiKzLrz2X
KIk1Ae2cz/d7fiYlB/4i8t0dHDxDmy4btOCdbFAhJmcscKH1jNe/1DcAMpIMypI5
wbMVYWwry5+ZcjXZ/1NB4VZFV/77nw7ZWij6Z4IhHjlwhhQ+ZyKBm+ifZkFAJoYX
rlwkpaz/VIrj07nAHK1WVrDNTR6QJvP7bzIlNuRSnlbyo3AVGfuS85DfGL9Ge48i
9TXELRS1T6U1oXvOxRbGI+7sT7XQu41OOWicyJoEvgWby7XeoR+830+wPRDMgOel
qyd23wuY+XYUO+Ki0IgaxTx2j7oFbVc1fIs3hXP1ErVk9eVIxmYAaEv4PLwJ+K85
fS/l1tzQ1cs4UbrA9XZU/xPhFBE4ctGQJDxYt/w8Irt53ZAa4NKyiVuQAuB/9zL/
Hc5jxnLnI6Ey0Ts22eM/l3bvjTz7llSDbQuW8k1yAD1zTB+VMEimouh9L3BzhXzp
27rSgpg30AzdTJvKhtC9J/532OzjS0zkXbbIfcd9YIlREMN20XikIdko99tAes5m
X6M4VdhrQ+yySAC1phHuF45WXhp3IVCeysrXS64HPlXDfGzHoSwi0/0RtHXHoy7H
/bqSp89cBz5Hk41XJFgW9En0LeahOGwcGgHLAXeZZPP3v45HQKgZJhiIUtbTcJS/
Fx6g9TdyLZlE6QGQ+r96N0nE8OLOQ5g8oItYG5wlW/vDZ2WX6Xj+tWuv3+YBrJRK
VeubCGXkimTv3NK0okoJyhom+J0Z8FLY3Wlnj8yDDO5EAEyUFUQyYlCGQ2dfmXYw
pBEVn09hNL++FvUVUkSixoLCAruy1z3TpE1ktxeYPtIm7jXEMwYEo2E8BvfCBP1k
uNMAFWewX4FDH2Y3Ftm7RZRYzBuErY3jpwMLYg1vBi4oIhp5NVK/5G4BBr8fReJJ
Hm0VGV23Od3s8WLir9Q6NCYcdMy03cJdpnqqvYDTzzsqo9wJuYrBKAj80mIO+1lE
yXSs9IP0uiR7hWy/pnfTl2/IvmNvS/L0wWhz5je3hXdF8IglWpt1j7CLuh4rLFLj
nhXWda+ZjfUn45hdaoJR/gjEKSykD3hjrNIkRmwxmqdPQt1tbdeCtEG52XlkCG3T
eMmB0VDel40fl6rlC+XWv5FgnGSVMegr5hxu4ySEugpdXFX4uM/ByJVGO368jBYF
gSTtyZ3azrBkWw9VtJHJWx2iC5HNIfCVAILp2Qeygaw1n+466X7h4+DZ/6hSvjs2
eLocOYgyR2/R8IN43SG8MFLKuJOKQoKkhcTPyXpnSxVdFjyMlbbixqPMjxK5v094
SKEgQewlglMCMeXiIgxQw4FTKaLZfzAvJN8AQjhmao3WF4LIEhC9O5Ll7ReuLeZ2
16ATAhppMnRW8mRCOJ34mFmoMPGhgwRiMxNpBFhDnhVWHM/d0HpEpxfeWLC9/PTs
LD/vFlErvtzNcBE5q0+1yGxB56mxnqSti2RU+aOKfPbg3J2382qodgsVVsl4YDk+
qbWHT960YizBh5jbAFU8vvTswaMg+p9Ao764h9ETpqhnvcDbuHR9u8pq9D1Sdcl2
cnh+0OcUye6CHRMKKeT9wLab12ZQysnfeB2C/AVZROU+7xji7DaCZaEZEPpL/6al
G+pvl9Owk3ZxJyDpMOW4HtlpQMJ+KoWAVOaJjBqzQX0u9wjksNJk6eD1ioA5cFI+
tn1tum8dkWWdLwf9v76g3lkKdACHM/E88C7oyIOwzH4tPuzo8zYK7OwDRvykz+O/
9TP+BO4v/TeIoiFI0FvwLDnGHwq203TTfhgQq5snbLUBr3jgV1b4AhbOwH8Ekjgs
c1jjvD1xi4tIlyJ7a3C511s1i0t4uF3hMPuK8It3nLSyjK7XbBiBjfqDQdWd5y4+
Q+zrTAjsGfeq9ipRapFzCA/6FPfBCX+yQCD+GSilZWyRSGpI7qRXgKZXfqQ4xkww
ZDf2cJQmjxHww/KILhESJKxZyugdNAKBRe3hDd3KrmLfjeHBoTteO3XsWOvioC8Y
lEAEtD1mf2s9b922MU8qXr/Ep2lC91mk2IZqZKkZ1S0PmN4yoQeZxXBXbQ6xLK39
Nxi8XdzJ6mIxC4t98puiQYVsmctDzJc5I5THQqrwFPLIRZhX2cREBiSWFJqgLLPK
ya7tPBFBZOxJp6ivX1Kh9Wf+fDc0D6WyiCr4U5wPFwSoIg6etS8FQ5FDGoZ8Oqdp
oGe0uvW+5S5kjU5yQESnOjKsoHMPbAhWsW+VTHvgPzi2AAdXkTg1wYYVgXpRr+iZ
ursq+KfEAPViGV5I90KaeFRwms6Rx72IuzNMvEPagEzS2tKEZMK9oe3EzfSlN9NW
nQuYCQaQj/Bsqf8sD5fR0nnCkumdcTJ0bhkXMZW6wLRdiAeSv8Vgg2ApXS+PT0FU
ZGHMHRgBxpzwKIn78lMAFQpYVgmfzwMfOhKqiquJ77Psfsl4kApo+/slzS70wF1F
ITd4/jIdmpeI9OMjyqAF3G+TGBJJXAxa20HucM4dZuqcymlrwZTvauaa1VIW1G71
YsgjuFoKBJw4kyXRE7LklXmkW6BziimO+O7u5DooLP4BkxKcicuRPQ9q8LJpEf1m
r6brCTWDPx3HD/+s54XnED4rSKqyPGjqoWIq0arZnFFd9Hx56x6+HdFdD4lO7C+K
BgIf5zTy4ur+ubItFi6dK3y40lLx1hFjCqFJ7WcqNQSHFSo5YznzB3yO3m1ku1NB
nZ2CRADaw2xR68ILGwTmLX+bnqkQkNk4EJfzCoQ8TIk8E8t0Sfu7mjtj65TOESd2
FNOx5t0O2IL9r8p9mimSTk6htWQSZTXYcMJ3RPrYJpWVCTgmo6WukR8kMhT8l3c+
0SpQ8ZPnQu1+6byfbYyvMOFeFEda8Qn0Uw9E4ZHtUGawI6Kf1wSPQVmZl7Iypbgc
rUdr/ge+jYr/DFKbylnIXrB74VcTWKcoSfAvPu/83p/62MrlJv74jFTYPldsc7Bw
Tf2Mh3J96cR4rHQeUwmZd5Kh8EBFwxcUU61wPQ4gDhr5txpmhXBTS12u/oXpjF5l
ra2AGiPz8vP3MD26B/IrYNNwd9vqJ/VywnJrbd4q2YcF+mLc/jAfysZQvAfJuf7d
jYPAlRgseYg+wueuYPh4sXqFIr996IQOCotA0hc7SQur8Gcnz42craRyMwj+2XXT
n0UvbNhFmvWWl9rC2brsXIyM8k98XWuAKIvrSC/FzokAXXCuRmCcytAgC2QAI6J1
9l6iYsx2Ep+DyuMZzzqe98t4aph6KE6u/77zsUlNBQzUlEIgeLzd+LIFUV+kMlv1
tmqw/CBtPKZEtUybitWozcZZ/q1yVv2/2pMWIOKXH33iwNCngSWTfLE/LqvTQViD
YAAReUhWweS1hPXpWCuPBTzyYXYjaHTEXU1XGX3GtN106RruAuTFQfs9JfI0j/6S
OdvV2b+sY00J4rTvpA8fFPRIK3K3BGOWFInDocAeaGGTtCG2UhhZSpL1fo5cqS/7
SKAsdLMvRr0DbGiucbgq1XlpBZlhkwjLsD+w4ox4JqO/LU4AdRxh91B9++pR1ZcB
v4BYnGAJip/NRSeVUwiDW8JpMqQANtJdUaJjXCwcGQA5Dyiaaqoj5HnJKwByMMjq
6ueW8r9Q4dLbMJEXp4gUcy7G+v1C539taeVSSSF/38x0XpygORnwHVhxF4KcKcBa
9QZAELSdfGVPBvaRP9vY/8+xjAMKmbhgRXKLBRTPP8Z2REYEB5UglVWoGZEa/uBF
ySyvffk2bvUcpnBU4tHyQLgXxL/bHC9MZcT+sfC1L6R2bqUDdvIFJVPkzgp/FcVA
jLiLpdZzFd2+NC7uojbVwB0TNaOphi1dGotipLZVOLBeCJjfNiW/q09KlpXAVf+F
0h/jPlBsxyuNOomrX9qOlYBxQn2kyvnZdXeYcefUaR92ACVn7GgfGJ6BaZqrMUyq
JgMOGRa5+L2eR56c0KmYOh/ubXi32dOUb41IwUFGfNj8n0ZG741JG3Exyf6TmTNA
dHdNemIQTd9kW+iYPPKCQGXlpc7E1t7jHT0PZnqUn8OnIxWghehKZvg375cZGfWj
8JcOC4MbM94BR36G9APz2dfrijwaD/t+sED+fupOF8FBy97APtU4KcY0f0d2M1oA
yqnKTDIrZC4FZ9rWKysMQ+Jp/pFEv17aqWYyGOJf1mr5Ng8+aCkjeXktnEArjqGg
nJvmb/ksc0q5SH2Yc3GYdv8oZL/FyZTOL4wc4zvQher715V3u/UGw0J0exNvEy8b
0cojKpYD9MHeUZmpfCQ1w1igQAPHi+7ca4dmt0gxhDlfRJSBfQTadHr5MyBaTgc3
q89Z5Dchq8Rzj5bfGpepjW0eqXQpaTTXI2Y8wYCpQcxcGVl1wBjua4ZhCfr5amB8
WZWoNwheQXsyySpm4pwO9kINr5qsW01JYNcinmJdFUzDc/qScwUgrBWM0Ckvm5u3
x6q4QkGPXoqTAnMOTNHm3oI5TEbmTofnJO5/w9no7GI+D8kiCyRba0+v3iiGMaOP
g20FcWVMwmIi8i6j/yirv6r1eaUEXpfmJyhwso/cggzKeliIdhH8Il7+pKZV0s3L
C1eYtyObE6sdhlUDDevSLS3mqetf4DyGRD0b5D8wHVvkDdC8sTr/zfe0Ug/+hEe6
Voj5g9XJw2dCBqb1UHGdNPWUgBpkuFfi9yt5gU+QD/IatVYnivc1k2XfoxsgEz02
pXAs6gR0HBBQ+mXSYbceR4CV0RIu4dkkRvqdyDKKueLlMuBlQPaEoET5f7FgmqGm
iM+MU/VeHRuOYypD9cPrpNIxzzw+BW0K+b3NdFY4/0+WNFTfW3VwxOronfFycu6G
YqXz0K7ZQwK5uAw/dT7tGio3LNjF4EhymzIHupq/rMjFt0b3f4zxB2jx3G+81cFE
lwDaKS7XHqa6vjqZVzCtMJZIQd9x4WxlCY/l42PyQbN4X4qGdA9HEXq7nxSf/H0j
BGnxAItqJ9ueHefzdqCPqvrcgib/KUhhxDVbHlWs37y7/gUBtLNLc5/EIqkyio9D
xfdmXS9OPxptkIl9IQ8JyD3YKU2of3H6ah46ZTeqeIBPlt+KXhg4/FV/6ogdGhsc
vkz1ezcMRvfwXW59hKwm50AyqCUw1TU3wzh0izcWpdC0KFYs+sRpEhclnVYHJeq5
dkzXfjmAZZwCX5aN3JSFOb0draxd1JtWFEpiGDFbaGLh16v2YKdZy/1AY2KGc/jI
VNS0D/QMZXfaUO26Vl5l7+RVn3l3SyIY98fQoCztvQtT2EQYgKxTiAHYUZmg/avF
a2CN/qRR3ni3eMdC9VwYkwNEaoVQc075//P9H0hhpTrY8BBb3tdm3D4OLZpzM01q
qoL2T4Ckm15sQ0dqkZsdyLMlth4TgIS8i9+xPvSswrMsVb/htSDBqd5w1hG6kqKf
dKRWqzeEQB1yaR1x14/p81eIteM7D2/38zoJxZXQb0Et/aeunzjkqDiP4hSyDfrg
4KodeXhvqw8oHg4FZvNBI3ADEG6LwVipkcsCvckfXfSreJ/T7DAgy1G1Qg2Dzj1H
e4VTSSW9Aq8G02a52yfn0cEM5xqqRtsoiaTgF+lh4rxBAZ/Q8U9JceYidSanAuYr
b3f/SaF7rGXeuZuYY8u9s2rFN6VbOC6AdAFHzbmB+KTPO2W7iQKnBK6g5al+G+UV
vtoN7v+c41jEaQMMNxD4Dddp+1hsQOiHthUPOwTwcH5YpD+bQC/WWhrYuSejQ8T/
mZks2I8fjB/g9DBGrJM7WgujOlO4ZHZCkuhJEmrNvRAbqkOO5h6v195E6J04XVu4
nESoTb/JaGz+Bxiqj92YiNxCHsV4EPrhIoaBJ+PQFtXsLSuzdCC/JVYL9lpog+3m
UDLf3nAzexRHD8UpfpTSl5vssR+QQkVx+f7o5rjt54PuCU/+TJ8lRSnSFrEc2uPF
8C5nWFqycS5BI7MaofOTsqcFfXwu5ibPTV1kUVsEnHgOVbUqn8pHscnPq9v8saKB
XJplS28ZhfdD2MaR6QtmdlcG5IO70mtbhOWu4xpGQIaSFyeR6QYSQYvRKll+Z+QN
wB7CvRmHTf7FE+237rvYWWVbcv3LjQ7BvPDx2JpljeOfGDxmJYhJl9SG91In/ymG
mqRHsfK/8COjbzFFCqc2J2K90fcB+fTFhMg6kIAWK+kAxy65g9H5gh2Tw8pzqLiU
PE15kISrK4GzcogWUtl/3sWu1rkDGGeigXKZWGLG5muImQBCD8FofF0NB5XHgrgR
Uz4sGg/YODvazX0GI8HwA/K2amqdPY54gw6aBI+f0Do6ayrnqPfIwJWzZ5n8FyxQ
ugSBDjaaOpI/ry7dTnOUkC4qR38bdAi1Ur4YERbB58fMP/yVmvhXL84xR7vBYlwU
RpB29bImTWKDoyzAicpCZB2KNUGh4eLzIHymfvL7MMbWfcQFINQOXDVBlafiiHHB
nqtWR0MGSHBFHbtErgnX0mlVf/cJXqgi7IzoNzDjTQYRTbXoHVcdUZI5FBZoCqbV
+odBRFshyBwJy5NM73MG7tExxuhK+oXWtDhrVpMtydqj9uzEttY/2w7qQHqrqB0K
lZQD8ecJNYa04iQU3KkSglvtlIMYw9mX7KRRgb2rRNiTKXYKHG3vxLxidPH61fWh
H9/DCnSmt36MeR6A5BwE+dn5cE2lsac53GPE6gDKCqMAiqDYdfn2qH6B4BlQCwQa
reKjbgfIEHarHIeohvVMqQ9GTmI5NGhXYrVp1LNg39j1I3cqACAAJp1gJFgzc9Lo
oXmrl6kqvL5VMHeI41z9TrpRuF+QuGgKCb1NIlbCw34G1AErloIAtWeVCk/2Tusk
yAALK8TzgYqjE3J7hNv0vEfY2qUx87XvwZur1hLleZny9AlJY+l2IpqyHkqKngWZ
MuEn/bYpqWwarc92HUAO2lW7Oj1wfFZeI23VFsY44lRknwTpRB48Tj3lk8v/Vmpx
bN0z1Q7WDRfBNgWO/A8ONIWWfR7XSXr/zSWv/pE0URxsM+u4LNPka78RK8vO7T8Z
EJ8p25loyCufMJ/dBWux0WzaEaThGT3c7rwYYWJgYPCXlDYGe0DUY/B8YpN9pIQ8
NMA/uN5nTbMMcbxyKcIOJmZ2vYDZlgQP4OA/A2lTObs/ZdCBWd3zPXloIuTd1a5g
hDqBEhP0cLoM2eMsHpLxdJg76PtDtYUGxXjbvaqGG/qHfl3nrjqnCec4lhs7pUuO
8FR1efrvuRwUWqXOK9cYSsYrHppgc2b704I1FRmF4JPtSy0jVHD3gNzAZoHmYXwN
NexfJPxW+64qeu4gPylZvvbFF5tBf1Nx4K6Y9tB2eu8R+yd9CzrPLy10smEtwTRa
qmo3zlkbUib0MPBmdFlTtBJyox48kw6f0UqtHVFigLVf98OkpYUtd09q9ng5zyY7
AvelJC22+nLyAmKfrGgaCrceTfA841jgtsoQTAYci1KotkkZSi5O+su/LFAtQ+Il
P9I4ff/2yFhaoQTIHfcNnvgzntO36vJMVT5N8fJnNLyIYt294CDph/N94Cmqb5+W
myy+61ZWCMMAGx5UMEL5oji4BYKBVA5oiTQc6OeW0ISs7e61WdJHitmWFuALN5TI
CFIQNgwxgWch0GgVMTpc81/XxaHa5gqPy+Jt+ebAIOhTDvJ9/DD/v3ExEG7gEkHb
q95V6E3zK+vo43kpNKNa8EWx/MSi4nuDB4AjXrjjsNOZv80KLQbUDHfF+pCQaC88
tLxJzr7rUep4SDm23MxznfP1Ub8S0phsBKaIFKencUk/lffnulqENbNpv1d4GZvU
+hWLAAIxL7cOXfSp/57Mt0+2HvJ0zmTbrdY/LJbtm31B+l/S7rVrZbl9NbOC1hRP
Mbqa7P8rUSwLfrxgbPiqZIrI2jUjmCOIFWIf+ruHkpkzTYgH1/c53wrX/QRGnDQH
FKmuQll1q1/spH94Gv4k3dhlXAgmroo74MUcOaUkhpX0pUzhtxVKVq7tYjLaeOT/
r/X3w/noUaiJZ5zQI6ctck2a5ZQoEt2PhgXjAKpkivsO6yeON5n7C7VD9rcGgER9
UUEAMAduMiFlY1rcrXlkhKQUwkWuLNQh9KmTlBRiVe591avo2fhCPxlSKasGZWku
0Y+YYau13iXRkTLqXyWRn3u6gwOuz7g5291LwddJAHLr4i2i8NSRVbzyq9O2QE1X
RQ/S3ySB8MXXA64n7JdiyxKBH6Uhwt+b6+ZH/Nj/UvyVaFI0MNISVYi+MZLsEcJX
GWi11jnRoC2hXrrbD0hWVT7NGfNMjvPDUTr+P8SYBL06vF4lgxaO6BZqtVPC2xkd
QZrmLYlq5bF0IFXAWAXHKMKzR2n1veVS8S1XDIo056H30YBfxHSfZMQWQ9h1b7wi
F0eCwwDpgUa+CiM/+XfGsuMbxfCpgX0VtKqpMmaoSTy6XJX0ohuNihtVaoHnCgKF
2Wdd40AWdpil2AYSG/h2ToqACTGC/WeyS/F0cNhsYJBLxfAvyu44DsNnBg4rGXTv
yI2ZOF8P/8Yy6349asU8YFfBIwguNhWl9gGafIJwaYE73y97JSb7yw/i4ZVcShBM
aQc2jfx+09EiEqJNlJz4dhnP6x59YMjCSRea7+afAmUCjz+LYmzg9lbIQfmmfSyS
/9z0URy0U6yY397Ld1F7ashGx8yeKsU+cm80O1tI5mlL4Gu3OkI6u89LgpohaIkn
mcu31QXTTvsufuf139La77xbalBf/Ndf3fPHGguDG3p9QrYEkXAb4mTa376Q1SnD
Mo/OdqPIS8omwc7nol7Cf5QRPHH4RxRSA0miPj0Z5Fhd9Hmxw7yo/VJ7laKn/9Pz
NbHUqJ91kLl1G3UvZ0rzrSnywKZtLWy2vqo77tJTEpKW46PI2JPB7Qyaowqbon7N
fkTE+dnHwrtT5FTrIS35swQjG/MiJvnkxce+RJVqZE0lU4ReymggQ8GLwr77WGEB
gB6S9JFlQSy7J/Sz59gMkME4AboMZBRhk1QQVBcIgGsTdsSTXddfC7NfLGDl4l/U
ybGeA9Oc+vXF9vfTUz/7kVljmqsaLPQ4NUdsbglGJStrnaB5c8EHVQ9vK1LsUwla
s0yjQl6jPNEF1Gai0IHZpXxLxVV6pZzz6PIAFa1KpXGIfsFzb8tnytArjFAjlr9e
FU6HYkdFiYohARv0L8Ae0NNen000TZ6ksHgou5YZn2fgf6IWdhCjhsOgTgD+pfdY
fhkH7zH5rI2r3ccCq7PcSztiS3ZqC7JMischOpQcvvHMtlC9v4o9+U6OBEivTV1o
qY6UqE/qyu2PsLATuZ6rvdIMSUt+bx8tSmRrhj4A7agcFOAAGoVtsw0zf5+J/dMD
YjbkLdI3vAk1cxrXdynDhifdrv8jfYOgd0vzzYutr+hJIen8tq8gWbQucsbC6FcS
Je6Lw46jSjRJshfW7c/qifsK0/II+5eBaeoQjn7RV0Qnlhjb70jQdzM+VcDsPU5/
/4CvkdQWEOwkd2rBZ4/K8W5Ie6i3NnJTeHc2HcHzftz3TqFfgo4c7dKZAA5cDKwL
RJIkF0fMo9McVQKNCUPdPfFFM5F7ECXsjjCxusfXt4pTTkDzf/d9s4EkL51Ii/ar
j2rfZxpONooT0n6NvV3lwlQ7wbk/4ukxJ/T2fLPo8pCq1AZ5cCnpEUoyPAQl7udC
4eANaEwTVdqN+jYga5OFtWo+9ZiZNbGUK1ArixTRMzgFBtQrkCTsecb7cFHelnoj
QWARW5Xe/D8MiZYut05gpSUlnQbkefZqOSDYbrhaWuAT4h/roB6PHyy1y6IWJdQQ
Fgv1PgM2i4jXc3oQrCPpbNeWTZzbEuxuVtHb9yzhXAB2hbsyhIHPOdTFIgM+k7Ei
29QtxxmFM1I4j5nrMokp2JdeAhq4U+ebmGFhWfJ2Eet5fQXecVEipMhYpkCbi4ZI
65saBcYmjf1oS3z8lLKZCqJbiavGdlyAVb2l4kTHjrZZewFzVQcdgh7NmHpIUQBs
edHzxLpXXR+WCUO96i7YBGCrJXbIEWpxMwRAYyKz+a3apn7jBvI3cw3mSam0FMB+
ZTFZzS3Z2A+pEytgQOfI1rzSUrO9x2M4NsUW+PwuFDsIOytccoDepfDiq0qMdG8L
/VlaXX6p5ZLVfAEZuSZ80MXD6mY8KpkYl196JeZOKEnP8wg/dDy2RSo7Rg6OdM/2
sZHON3rx1S4lNfYXQSjVs9bWiMpTrTzBP+56HPfVa5ye9T8peMT+Qp9o65mcf4aR
aIrUSMjRPtwuloI9ZdSRKYyYvqf2i/dldrfEpf/zL5q3icl3kIMo3++a1x+NErHW
98xzFnzvtRN2Ty1i0nnxRnMBGTk/J+uOXHYDG4OFW4D3kJ8oBRJck8JvmOYzyazg
6zb9Q0L1l3k2d/XwUkDkQ0OR/3HB+mTR76GRGjCRnuJMz9XeelWvrTAVX2s76Ota
OmhkTa4W9gBD7RGi1OQhlnmPravUQOMP+Lz+jkPN1UKxS0uUS0GEQn6Y+6AEcXci
JXI4p/Z7ivhm5nzx0zAeGPhfdJtC9liR0zoL3CqhvkOMHJNT/hyW1Kmm9AeKZ5ZE
UWUoH4coCclPxITjfKRei6YRBxBPkUvM1eB7XctCvB2ltoKQWAyo7lDCyRRstwNU
TGAV/yOWBpJ6DCztTzXQsIPdo3VBIpxobUx5mRx8xAJtDBlFZ+kB9juTEQuuu2qr
OqG0K6VLcoAb0+ToTYeEymto4/Kv+GJNIJYkt/BPtBxNiXXnEFKu4zb58OKhRn3C
A/vpyeFjr15WwzsAW01BBrlwaGzjWhbDZA1BjgXVOUj17W37uzPIYxq2fyzDykGo
aOVUNFBIevx8962/gczDkDu6/1ppGpdZvtoziE0EVQgB70yaTR6g+dMuYc1Gqj++
K3ZbN0b2iC4KERqT8LNWoOadzziI6hxCMMWF8bwGvPrCIGBlTKOoBoRS4qeGPCID
XAY8LT9mdzzEoT1SAzNCBXBWiF9YaLht0myisr5pY63EgBwZJEirx1F7W4Ni2YAS
Y13q3wpCJVE58lswFy0ir3VzKQcusUHnNFcwLLBn4dSgzqTOngm+2fzjF67V179H
9TxLo8JF0tw9U89w3qi8ZsJX3jR3tZRxFFMmAYcefR+dMyQK1PQ6jDNskdEdv00A
v0vWk1B/kz5dWBUFJ39NKf/L1R4btyJmUhZFUjMPNH5mRMwv6HxcKlnGfyqbCISD
PTCpT1S61o/B/hcvYaTbXghVSdgM4DtXs4KkDT9qCvHcqZur0i3Ln0y4i/2rkoc1
0s8jfe3zhNXWf75a03GnxY4kPgFB7qDTq66CLVUvhm7bUfu47LqIE36w2Q7cxxVx
/+c6PTNI64d8HeAJGVDr/+Ukp+xQWjAVHPYIml9gYUtuUdHNVr9/FXqZ440hzDMn
D0b9hIz2OoecC8TDEcs7n4luM6DjeoG4jWTiOdhAzUd2Tkzk0kEPvySbCElHltqw
LtLfs6nU3YmTGVX6LApEVpBysw3hEWou5rdO6JGJscY7NqJhNM/TvHc6Tnw/sIRS
Y+umYgdYElPoVgT7sjvlc42/eG3RTt8p0tt/KAvEp65hC1svJeONzFt1NwgBJ7DZ
RhQDoimQoMOakCQ+ugff2qBMyIY9w5VUGj+IJJItDXRzl3RjfQq4tqyfr68se7ID
6cssPDLbUoq5sg07RLlgn3Pf6BZtmqSCkmsMBAB7UyWe6xsljiU5dl9gP2YCr+iy
D8jkmEkfoQartOUAOlek518Nn4+7SKw7e2hM/ovadDKs+NwwAAUNDaV4YM638P7k
ZoFDcTY0vuRSAigzDb/XrvjSrF9zsG5PoxEDiyI2oPYmBym5A5d0m/dBLom+UzFu
LgA7oWuJ8gaJsSzwO9vkM9i8PSaim4DcudBZ+sIvEF1zAOvoWi4MKFONNK0lhRfs
j3p4HvKuQXEemlnfmGT0nsFo2dXIqBijoRLu0E587V62b4bJDcYUfWfgNakFQwur
fH+gC4DcdqL/SxFt2T6g38SwLQMmhr0fQAzGG4F+VuHR7iRBrec0wAc0J6EpdIx0
1C1j/dbArF+JL0l4yHvRXv+aqbCoaU+rhs1kXmSNQquM6Q60BkvOqTpBQmrPjAAW
qKV0v+xX9YdpW1xleHVc0bYEFN0+C+KNH96iZn6F/F1v8nXOBpNGVvIzKR4PPzQk
LiAsr93BIUrnVY9L1zrpDVGfu0/EirbcAiFUkNhi2s2vOw5fxLdCtreVbQ9gKP33
hccWDa4mINVMRUHqSlujbQR52EMyl73yd5Yd7tpYfo4M/yysDjeDOLTLJdAyB/FR
Eb2VDDcYh2pS/Ia5B20enZu1haqjcrVHLQM/OFl6XOmuBup0uGjez/qySyEw9MwH
8vHH1lqa8qbIeRmWDWtOv6SbUKHf2A3YzDr4tho9bpx5ybt3hdfzpQAhc3KMUHlq
BHlhug3Zk85u1Yo6ALxxR7yO9vJPScIxAfyKuzNhvE/OagM2w7OnF8l5Hw71MlO0
AV1EcQ9jwQMWxw9UpnzjUVyGbm2IQzUQOuW3ImSGqD3Hdu/zlFwVgQKSQKAG4ESx
8GBgCtVSnnVIzh3aOgP56F66/IfRpoquD3gEafIRtlxRq/WbADVzOqXl9DXVA84A
PMXKBMZSYpLBCnADcSzkAWHoSJh3Jx+ApFGZ+Mj/Mp2Uo9H4nonGXJ0rU9tax8+N
ULT1vmcf5GjQ+hfdmClleUaqvSzJCv6k2WVWGj5GODRw+2UxK7z4SmjRSugCjiOo
kHxng18oeGQVyq+JuDIBKI2IHFFlTJ6Pf7lQTMV+1dJ3EPvE6EyWM60l7vPG3OU8
bgIKCq4dRnAndYaJqMG+96mPRRFp52qPxXCJOerMy1BTiHG/WjSZSphuDs3bTRvK
AVXqKLtXuwD55Mr5WF78aCAv0Tjcq2k+CnzxT7JjsJIw1fQxqt/qyW0Ws3yQcYK6
mIKs31jvAprqJQpY0olSAkzGPA3Izi/2I6+BTZKcTKnS48pjUIIa6FOtWdyzfIwF
vSN+Ub9UX2rskdOmcopUqbtHuGDcpw4DnkFGLNhuoDqR1V9Ef26WUJ0+4Ee2w3HT
bip3vJCqou5NcsB1eP9QL4CDe3VRWysc3hQLdoaGU37G/adL3eAUZC2tKbEOy24g
6XXRsTuumuBtv0SxFuMisk2+GqpIQFzdRkiP90NqyLGnpSCDBWTltX1z44y463Pm
vIemjxpVcNCm8ttFylwuzvPMbCA2pGJds9AMuuj80vRnvum/wdJy+ax10yR5wtdP
UMUWIrEvE3q6AtbnuZ4Ty/mDNkKU/E9Qwb4NWVhdFpOqT+fM/2e8yNwE66tKUJ5m
6zqZtPZXgGFUH5yJhmQawNA5tQ7hmwY/CyLqBraUaAIGwBopsLqoPbw08UxQWCz3
rckAz4OzfiAI4ycpYJtLUIHJfT4aj3G9705zNQUecBpADU98X3ijHgMjph9jE2HN
9yVMcM3GrCTb5HfVl942RsJom2bMeO492CZNPqLiVQcYMpvpF7rpL5c9lPPkA995
/N0IHlvvSQa7RjZoEL1uc3qPhqduYLa9IECIm8fXqlI9HTjk0iPEC5R1gbNYpCnV
pVjru/GiYMSguG3/1rlPQUKlsfUZjTbH+fYzABj/gkDBkDkWyV/1ySb6Yc67RxBp
3ijojA1EzTVYA3CCiyZhxjyIZi/j4OO836WwgiEXz7Pz6+x2BGQbWXtNTBnm3j8S
H/ysiZ27fe8giTTYnVxhQc1GLP3NWWViQ4a/U+IgJEG74J9P2hv9ADrJgEPEPFPI
CWc9J1ljGnb9YDgfyI9dEnJJIkVp9P1uHwE6VQHhh4etWU5MT2+ulJIqG6OhS9hW
5Ogj47Cp//sHrwljW2iAsISaP4GRWTaEQHddjFz4vL0psEKFJsM+sq0+i8Toamp+
yvfnME0QDpjCPmqAhY+b8Enf5+1lUJFBf5TQ2mRbqf1Z07rILP5A2Mc1VcA1IKTW
JY/d7pUyqUFetufX2NAjp9pCjZFqUcoaqKMOmzfFhskXVrOqGTtpzP/A0+nJvmLv
cUlKPvN9HEg94JQxboGBWN5Xamo7MdfiaztL72zQx+qx5qwFmE3gXozFyRt2SXdd
fAVwxaGYqMhFbFmZX2BSGCqUPL636xArGHUXHxIqEfrPCcft7wNqqegc9jhfpy67
9BNd6xkjvDrtLbINbpG3lBEVO3IQIrRFIf7lcZvTXT9QoEE3H6c4JaibA8V8YRcA
EeD9jTV2XSU8wRIZsgX174ocPod6LNEWdwrqbol8omoZ5VU8ttaNBRLzgnvNc/aN
BxuEpvSiV9k2OXSHfSOv18qd6kaHorbb3L4PhS7I1KeyEUQArChUdhYbRd0Ycfsa
9WcXUkBcF9vO0AYptJXSngYn6a58tiiMFjNNiaHAKdSOczSjwtiCa8dPxUaVAki2
w7SC+GHrHaIJi9Z/TlNgqeNIPi3TCP5hvrmDK4KxniMAbQGOyIT1ae2K8JiRyvIb
ACnzOv1AJ0AUk1uHkvhyQQrHRgO4OSbJ4IccH+4X+YU+XNWwy1oEaWo3IeX7//gV
0wlEQbClkzmVBoXhBDtMC0cX3t/iz6dNMaWF/jInnurW43Vm3u/mxulZidyrTQHP
OLcWHOE3WGwomim7RC0OBGpSDYuyJWgdT+m0oEj1ZFDWB/GS5Sl2pXh8viuckMc9
0ZveHvz+3kwJNo87udzEv59knMr5n05UEr/LhjzXpD4ddzg3kU+YztVQHopEVkeH
hWqYkhTymoafRQMpCAmoSirMBqvPPFukPWelmZ8+Dve5aAvWTNxCs9x9PViuqJoQ
5E+8CmOSD5gTrl32pNzLxSby8pAagMNUGDHj2p3wCIV2jlAPDHW4Wz4MvvnyjB1u
gJttSiSKb0HCPAxdfi4oPLtTVMe19OVPXGh8yUnM2Wz5qsClOTkx7sXGrmp8K7wH
hZjd3N9WXS9FzROJaO7xGosbrt3QLIDNF3BObhdsFkVzFm0QDURP30c8L/lcWyHI
66DVm8kLiLS7xWXQV6NvYo9Em7JBbuJOR+D1yQzQxl9WjgsaQEcikiodnK3EKG9o
GSO3gdIqaC3uGV1nxZJG0cLCf1TNftSw83wfFJz04rGCOMPIL6wiKGJA/aHLFYIJ
Xj5Vq3l63FoiJK06DEsknRePZ6I28LNhdSQYgoUlmUEsr9E2DdSW2/ZOd4rzl45h
KIEIUuM71aiklhd9B6fgkhLHmjVa40TtQrFeIn9KHjJ42307dMMM4MGOISuAzEsA
hEJJOziGxrnHeltGzLWv5J7tIdOwpMOGseheWblX5+w313pI4K76Vcj7S/32YRmq
OO2G/n6tVIcEr4vnrY6TeQOVl6Zj1iXjqML2NqVeEX/vPMmudH5idCzCyNS98XeJ
fyQO90QMltEHej2DlwIh7C1ZFcO8PLGvRrlwERH7Y39HZGquvknl6SvTe4jbJUxx
3Yp8wJInVVa0QuXVxjO6/keZLg8GSqmeq3bjoYwioKefwHKBHxwegsySdpATWAZS
S7vGLUqEDAJ2TjPAVOACg5QEZ1o5bEVeT4xiq6nG2qHOov2ZYlo8AT5OG2PDpJI1
Ay2TEcdIlq8ZlhvDmHebXRs7SthpxHgeyttz7zFdHZcio4biNYWFHz0gKUkXtOnF
nEbaTNjfzgvDWXmGC2dILDAOcxuMqQsBDheIBJPkn8FNZ4s3i2Cc4VcsXmq0OtFV
EhQe5QO6+gDrdZWMU4MdZJfRYpNl4xR2p5qSRce3W8nR+IqCE9DGONlc9EOZhHDN
PTQmAKWB0pAqxFZoZZEgRWPseCLsqyys4nqlpR6LVziFCH+UeU1l3VQCS9TDFw6m
BPvvnFA4WwG8p0pAGuaBAVFNTc972suHFlfJmdbV/JvtUmUWudVzp4xDit+xvgai
oAomrBaPlEEYnapLxY85Zu68+sCghtOqsdeP1AENcn19jWaG0jt2j1MRZP2Aijri
iwNiMaAU8mllYF7UY+iQSl5wfohKdB1v8JzAwFitRIonn3eY1aUozEUf3WN/wNJq
HlOVTATS0XInDL5TnNjt3V1kwt9UaSRdPzJKVq3LRJk7+YIDmsK2oUI4dkF1HykS
zMADEmwKm6NpkDuVl53VdB4B1pTO1ZpJ7smv7bpz/ahlOyRxbktZovAmQa2pnBQ0
TYnY7NV3ARcqwxuAVwNsLjjXTqHq4BQB2uRAwzjNmmKSlNIcuImydzk2qM2egWRh
5rLihk2I8aDEzg6eDrKWFZIODYM0Nsjuuf2LHGOABOTOUDgRBjiq2Qw4o/zf9HZ9
GED2P2rnbALsm8ir9NHs+Fk685hJhH2mvZYD6AZHGuays6ipqOC7LpP+DnO8gu/0
DwdkaUO9nhIdTuzb8D1SnoLkfmZHZwmzntLjNWKk9G4wBUBSdD6Q+K3KDbQ8K4PQ
C7Ggt7/bytPTaT97RZHc5OEo6iTau7XDuvcDSucotBDr4qPQzpF8rHWfk14ikeiU
5nF6p1vL9Z78NwQFaMe03g/7VdMal/PyrDcCe+7VcI6bznNm+fIzEBVTNVHev3Pi
dkDkFdqnPkIp6BFURpl/cBzUWCQpoZu31Sbq7Rkja1bkYOuvx8sBn9F+7F9sTPti
zEMxUf84UaibleqFEieu+4ryWJwW6/JL492q6xl67xA+Af0pS10m/REy5VdqCm+O
tK7c1mnG6yv5KtFntAPHM50ubI2zumZeOi1tQCN3ylVPMajDk2ep7gvAjWztRo3k
c5XeMmgp+o8XocvhVhJ4k3OkobSfw9DDOT7uMGfGHChCRtafDK3x4AZOKygJOcDE
5aKygkTWhAwpYyEoPSQ9CdCEJRPWwPg1Yti88AIaRF9l6Pgs2MCEqWrsXs2pldb+
c5ovie1iWMItZ7VOBUDowLSAxKqEn+qkAhMPWp0FIoBKOjcOrehEFN6g90Ta4qod
gbi7dIpTBrFg94yrthEW+0ZS1qf7ugaxnj3pgH/v08IUbtG1b9Q4BSXfJqPG9U1T
O9+1ZT8dz1Ki0Swiq+YtSmfv+tOE0G1InhpcLiTh40WIXihdU2FvXD+ylJj58uQk
LjmuqQWseWTm24CCizQ8kNUVKalu+sYV8eR9G2vvBeb4TN2XQl2Rxn+LUmfL3yC1
Brg+AC5k/up7zHPhvjmQ1RwHasTrYvmAPaqnvxeSjGkmWWwpXrPxdmANh5djqReW
yf4ENroV+NyMqnGeAOubrWjgSrP8kfv1/LmqLloCker3y9JQ1Vws6551s12HRIKB
nzATuJuj5CvVjYu/+C4FZNOnu/2NNOSECyZlxBryH/HCEQm3c+Ul+c+HOFQf1Yb1
Sdwx1ExuOCBt/CETm+715/9+DgwDDBn4Dhh/o/lyiWbjBMxEaMFsgCHgNWRt01w2
QvlUUJvIUL4+X+OzferiHpNSikX10uiLfJhraK4mMmhNzyja8Bpa40hcVGwikCIm
gua0aq2Xohre0XKUgDZA40SI94Y/+UHDodO4Pqg36y9rhOJLMLzxKmt//QCL6TZs
iJO/h6lBykAUO9996BDqPRGeDJpbfZSldpO0KZduZsZ2K4P7XCS33JWYzQA4A8HF
aDOT0o5gk0CnBIG+S9i8WA/rSNtReY6Pf5GeM2jYkjXgcqtiIsxL2Rgq04BWfw5q
y+T8y0/76KZjIeSNSmHv9vlTTO3unPDjMuP7Rs6LkJ1gzcP6VID0CvXsUABlVaY9
Dc4CQutN/ERC1QO/9em4x5xto2/08mvTnuXO7yBarbFXbRE11ps3HvwH6mfSdNVy
2/+bT2CAIAPDBuC9QsLhr/zdTSqpK22llQo5IP8lcWV7WEV0WjRvfTOkOEFQnK2e
V0NtCo4+Weun42bWVWcUK45wXxgqaOK+LdNBRgN5pPslUQIE6KCW4LYmu6XYrGjv
aOEQ0781yYDlOfTr1s1kLoaFPsWoh9vAwtoj2GSjsm03r7jc5v9fI5i8wu81Yjba
pU01yv5lSIi0fckFGtrtnyN8jlWIrRo9dosC62kwfQ+Te5PgVlHib64xg1AT9h0O
XiypnYOOXnrJGj28A3vgOaCf1n5Its/ujioTFLHmLp1DZoWLF37/6wtM7nQRjnPw
OxqVQ/v/tgjDC9hQU8RMKRH4YE1sKFSbc56OT/+rPWmqG8M9T3zV3PmWppnchM7h
a9FungVqgx5pcYmJ8BvVwxFYvzgG9GX6hbPUOQfAPli89vnOe0pfKvQmGEAeD7Ze
5qEM5bti7T0yl/ukyoU9oSIenFBviDi/zGWIEAP2FgeYLFake5h/sxir2EH1fkE6
iM9ZHKODo5So7faBz2DsW8eOTd4bMv3w6VCUw2GLx/S7XPvQBOiTLY/JaN1fZboe
XM+T74oOtAjuEmcfo1FAftskqKeww6ZEgjaj4HtQPuFxI1ApgD8W91oHwz+Ua6fM
yG4AzCDcEL96MBd7mVD4Dk70B/eEc5yOSapZ36469+MXB56VINTFbTuelzcr0HFo
YBrllW1kGjWY0czDO1EVqOVqjrjObf8eGeH5dGg2WzsolKqsD/XrJnpKSbQb3GWV
WNlHxkqG1f7PQtuawMfG+hzbSnmFlZW7gJaOCqx20bXNcHwPKJIrRHRYUtSsP+un
5RUA9RsWfTlv2FhzYcGFuftHfuhu0ykW95xmlmoHgjEVbqkSREx3mmyzv43KSwAQ
6FSRhMTSsDA7DshneA2L7ZpUdl1Wej5u6YKRIsiHTZ1UdjTadloB3Tfiuuwx82sg
ZEKtlFjoIpNxajNGZHx7hE2BZcloTY78RHrPyXfqXAXS5sWu8uHIf7T2HXcW/yG6
rw1zyQ6beTVjm0FBTQhqPivAz8FxseUvgBRFF0TNOub2fxGjfCLcJ+TQ3VMpcCLt
CwkDt/PJmXOpCg/RbdeF6bYNc6FrHZSDiKynvkGqNtvOAnsHHvXs6X79hTYkmAvS
Sn1aj4lqCpOnHS4IdVtMyNchhbKeFh7HyPxaRvKz4X4BI8rLLSyW6JQV+16J8GtS
HjxBE5ou7wp53gMhej4l1VHeYr++2oI/tZTzjxn7LSc+yXQQyI5Ozs+bU/66JvhC
amTo57Z7LundEI/U4H+m+68LNaZImBwEmYx4yGDWcteQMq05/DpiuYyCgVxFRKgW
HfdVlUvfWG5eeByv08ZWuue5A3wcfAv309uEhgi0Tx/Z8yi6x+PPqNLm+WIzClhw
F2Szjal4wTdHIs+l8OtXInkaYYH0zxYLKO7KwlhKclYlQMOjBt6lYo1h8JTXDzQ1
TLjbR7OXR35hM5E6TVurz6DGN27ch//m4WgxLyGgt9q5EIy5QbmBCeq3STEvfmjs
lSiW55E1Ou4wywrw3JdlXmdnGXjaJVgxpjlJNKhPzc2Y/q2DuN4sb+Uv80uKdV85
JA3v7K0YR7Ecp5eKRJBpnoeojlSArnIp4wvUnaFDpkbxlZfM8SHB/CkY2vXHnIVA
D+qrH7yCuBwztvsIPyJC2TxU52sjl2FxfWGMbZ5nwN9i+v33dpu9bQoEtxpK18V+
YL6k+aTPWuJeBYYEcaD5Xq1yYB4hFPvK0GO0O7rT8m1DC4hWJjY313xWkz6zdvkL
mVsAyEZU/ZdJhm8BYVGlCP7dyEhpRL79W1JXinViL3NK4TK8DpBfv347yYvivcVr
t4uOLiC72gPvWJvtsnveJiewJ5wsQLmYumRTcmbpywOicObsubhNL+pWsYFLmtAj
ENw3hE1BOitFNDOYwPOO5Tje0cy6WxwIyqBOB/AdWKhr/8lvjiCgqVnzihBaR1qN
/ZcmUzilNrTOs+NvXIeJX7+UgVV0LwYUVYVWnmo/GTzAQENx0YwrsXz4wmn5M12t
rAzriYRXTWICXD7PdqmS224ynXhsoLqu+c8BsHn7lF4lI/4mKmEIr7eYojvV2Zlk
OGIghP6P0CLoF4hi4P4jIuYX7gZ5GNVHJxSkryrWvcKO/2f9kBG+1PFffLdiWB6n
DvGeHo3Zg1Oq17vvKe2T+Hmq+lSB235Q+ATSxdb7Fl5CW/9DrTyoerf2Rt7LboM3
q81DnQOj/1z4ehhb75xi9frwNT3IYxGhu0wkxENzg6wqDlOqjsT7LWj75FPlSTq2
x/UUxx8nJe6H+2l93m8DYCwXMnyJ/jtLi3LgnMoVm251avebUaNJg7f8+WGwnQ3j
Y74tpLwFR/KZFoIZX4KdVVit3jw6r6OynGo1pSwMRCXKzr6hIVpU/hewUy9Apwi8
lkx8TJkPNdGlydNOHqcDTof3kRN2vMPt8Mn9LV5+OmaQnPzT0HbqnA/2bh5Q1+7Q
rHjU26errnyxhq44mJkqHQd8dvi1TTSUzRsOnk99W/jj+uJU5npOOMqIwH+Wp5UU
L5DcKcsTaGMbteb5PwTPPj3cPtteXByePWKU01Nu+wDF6LHD1lfCxZbfCbbk3bm+
Od9ZdcgKsnyKwCVq/7+rn5uzcsaMIc3SWzXS+R1DJXYSEW2Og3JcG4gaRZZM/Tm8
D8b2sp1MIDIJGY69X6lr/Xgyot+OuGOrNaX0Ytpl0394pfR689eb7/lVO9YQi5A8
uV1/gqvMp7U/nSD6lOI384jIlev9XjKU7BV4itt0VY/BszHHLWLSCPQpjapFegy6
jjWWS3R6Zd25PvgI5JEjlLN7/4KGIv1x8Je4ZLUqlqXYkYtomP8OiQf+/xGTcmLJ
ieLQSuluT89C08i7Ushvt1ukdCm5l6cERNE1cTl/e0vTfMQ5Wn9m/XuPtP6+IrbE
JDTRT4rB3UO2L+BYVqaPv9pXhDJajxjeuVoK5V8f7fFMWwyei9kIIAIbOgFS9Zsg
y8t6dYJbezktNPF0ImTVVzlOoG/4jK7Nr31Iu39vXmmDnly8rBJVLgLeUuy+Jv3c
ihNcvhoAsrtJX/ovPFIR2i7VfYYpDndg4GNzCdbUdZs68lKXebxtewK1RNauFofj
tR+VXYI5wgQuZbepUggT+9uix4HAK0l3MNODZbZWHDs/9sI4nDuDdu2SwnUHGTgi
K2U5hQcayjfZSWF2BteespV7X/GoGkcsyv962ovDDYbjelJQPoJJgSVPdjEjjP/D
WNtg2sYbycXf/PsFToPzovE/gVXwXXBBHilYZusqctH7xqhew3jG2TzTRBti1EGB
bP1nBhpL9Ae296vpFaa7sdydj/KzHjVm6xNtY1NTijpguMSRa5cYdsbH2/AmGpfr
y0FkhKKewzdRaY9yLXp/EqWCOWkdj/U5QbisWBLIVxJh1AetHxWbszEIEdRRiflZ
QqlwbkPYsRIAxmiyDdSsvTbfkwl2eE6/jEnUNSheZ7x9/MlRdWuKxU0wB3IB71wF
/CJISwe3T0Q3GzzwPx2RErvAEQIniUfP85Vt9CxtEGAp1TXAhRG0uHKl0E9j523x
FaOdbkA7DZXVPOw3Tov3S0ILVCKWG3YvcqQLWh5ImUX01EJcTORBw7jimYt7pRhm
ptlY98beLsXPuIdxPEQU760fWTypz5RoF0Er8/Se9Xg4vLSAOkmGGRNwvAZ0YL0S
Km1jh26z948NRLltfbWTvv8HjoLMCUXzSGeZv8vBuLVO3T3yUHoCLMU/WWjkV/qV
Uxg8qUzP+hIliOyvpnjs3XnQFNnMJ1357A1yGK3FaHWMyVW3W2uLKX4uQY9P/0f4
o/K1B7JkD+GX/UXd+cSc3WLC0hpLkHwf4C/0RyhCru/OVcKHUoseENrrIMUAbL1i
0Es1w5L3/KgSyqq2oa3cfqxycZXRm0Xj2Z63Lqz5x7wm5H6KLPpVChg5NHrgBRA/
EY1YxKTOqJoaiSYd9nFxqEJJx0L+jFc7i8d66ScO2eit7bS7VC5h7uYId60qAvmU
0Ji+1MLGlC7CKxaXnjbNa/WZt7mM53MDqm1KlUUDMrhmD6V8COgEoYlhWjPvkC2O
fLWiwq8frMrMhWGvDRlgGboI1S2/DyBv0Yg09eNcKbgmpbji0SWG/7/pAylSiwwr
faP6Kf07X5J5i1alwyQeUBm/TyrhvLrWup2sd5Z+V/ZZpnt6fTGzIu+7cvBanAWH
7os6fkIOHL2D5F347M/yD7NE60o05fFG8Dbf7HrHlqEAWQ5BEOPzzBoHqDau2Jzu
PIEjSM39svAratOyrPKsrb23v+4Yf+qdkqOowLf78iZsrB5eemfAHg6bNem+GZqb
72frOe7Z40Ujt0cCV8WGgCPv/7C7xl6+kF8Su3vW+rLAebS93OWXwt17RFerwtJB
e+3uJR9G9cIAXi13M+3fvI4wLXXtMYEPXsqrhDpSr7dLXxUUPpeURGC00D9F+C1B
gAWKxRJ0879Rn34EMTaT07Q6GAT3y3uOetpcgBLEmF3wlwkRQQLYF9PYzve80Ksj
SeRNXeo/PntE8gF3cTQUccWQbBMLCvLoZqT9f+rTij+OB7GQKCvkbvso9L9j0bJ+
tEHAZS70LBLgv/XGeByeozzwMaVB8+LFmeZ0pT883T4tmEnCogWxtfovjDzm6cRf
mhLPUUWvE1n2x1gpdxXD4L6Sow7sgHvg/nqBP9O+RiWpbTb5jdeRcUYb9I9hm7lx
YFQhp4EvW6F54dTRe85p3zPt/gfwkInN6m/i5Sj+tEjGYE/ZSQmFn3LyG/tDTmCd
/rd250rGpmcWauMJ2tGP32TIjn8Jdx2P7I4ZJ9HxO6Xo2qCh79l+0DmNgJIa9QQf
OdXv3Yu8XclNufXiqZtOgPkKVlS/XcXPYCqJP70BCqoHkVRO49Q/8mly9giMHXxg
1Di6nsD3tLaDHyjIROdC1TxIbISTmPkqgnPj3+9tonj9CRZKqoJy0iJs00vzFUsr
XZbb9ll0MnA5zux0B9YCk2iWioTioZHPHDpiUwp7dtanFkaMBEMlx7Ua/yT2ZqWG
3h+M1fq1tWbP8T0Cl23PT+21LfkI+qXwFUgNnGve0qYnDKWJOpGW3DX3nUJf0PRt
VAbby3hSNDWhp+rUtgUsx0z8CMQQ0HkTrdOn3RpGstff00JEF03zUra5EygHoLcH
nKYX1UMrb712Q6U/rK/2SvY7sgydJXqynxg8T2JmaLXzR3ZcXM5zEJPLjGa/TFWH
DGPUpa2QeydZoppiIEcC3bW7MjoYXKNTjaU4w/ZCN63Irz70ebw3b52Hdebq8m4P
IaB9U6FXe8lEG9IkjUYtgIY0K8Om7wEOr0sWblLS0HmKpdl7iOY6iHcV3MSPu5TL
kQvGQEJxDS8VEEOnpIRG8bUuqMemLuJ8Gt8qF99QUatUbLotm4xKnRs0gnUCOtvN
l5tw2Wfz+2j36ax1SgtGJUYLZNc427S7mkJpR9CWRDkl/UU6bsOR1RE1dXTEje06
/VggdnssMjwXg0tvIJxpipuH8i7bwohhJgRWFirQtxTCHlqxNR4iUnkBwbpGFbwB
2idW67rWi7661kLboj8khx+31puM8I13fz4zfA432EThR3H1u6Wl+gy0M8g+wG0y
u1w3+G41mQPkRchrO/kIHDuQI4k6Y6P2Wm4VWxgeV++3KjAWuyR19bUmp9z+2vVX
aW5y9qwhABji/Eflz/y//LpJTttu6kdnGEjdy3AnoGZiAoM01LOq3caXtjXrqFjn
SStyk8IGj5YK4icvbSBQXnmdxuNicRNFWXQY4Mi61zht4AP0Xu+XUvNvQs3Ko/GP
yV7JKMuWcsaU3y/eGSipNUjslGaMkwigPn5WSoBHchM9GpOXpGVY+tzFOwqJAuty
ewmxHUVyeK/lkld3OjuVgYVvEc+2O1kbgKjJo1RmfRWRYT1wj+ZpHABizyewAQAp
+RdSDdkFFNbzih3Id5v4dGGtRLzz87LQSlUs55oPcHGQuUqqBymrfq8ty3ZVRb5N
G0RzHWaj2lIDtDvzEJge933YEut/piJcknazpbtfV+3hBwCHC8mx6JDxm7FoSYpm
xCcIHaDeCDbvLIjy1ozX74VVszv+aWC37U/NZsSLogNfDQ9ICl6TW+O7rBtVovU+
/JoOTjcD1ecJ+cio6mlUgkI0P046laYwbrzmEyK8U+s/R/gRZ4dFOVMoKgG/PL/u
/Qouv0nTQBLwOfzbny1Q3mYJViZu36Qi6Dbhd1FGCqelzdxg6BMXynt6I4OEt0ey
PQA1qsAfa74Q43pbkMifu8o2JhfXl+myfijnkAybY9Wvonpgg9qNQ0ugAcWDZzN6
CNJNBk+JVVSkU0HosGGgSQsKN8psqBHQWp0Yw+sSh9iBe0YwqTg2I2vvrNmNhuQN
999c+ebZv3YUgKYUNh8fIFikc2j03pa0EqIz8ZjjNDJbTk+l0cW0SvbPvIKyvGtW
1OkWD4wSfqBFY/UVbwY5eA8u/f9z4dQdaRXQbgRu6AGm/Ksf4lHS8ck+mkl2IW75
OiiLG9/OXcSpOo7VOeupfs6M+WKcXw2KvrhaEohgznIgZMzMsqS0cJQVL1cbBEb9
wIpLpSoYSXIwz3Ju54nmozmaK2jeOtFnmLpBZYdNOA5Kc+j89ARe2uJbsmQI5HhJ
BlIAnImGhEecPG8SVlOKfMbFePcl4EPD53DrEAXlhZVssfadoClycVViaAQBS2cD
QFDhk7GP1seC5tHgBCQEQR6ySnEMP0hd5E3MEL6+LFLssOxmWVQtIfs4Per1/I8B
6QuPe+jzDDI4xqMNHzhF8LLY+90lm9XxV5XCh4YYkzR2+hHakMDMR5irLgnIDYwD
KWw2Y0pmBL59e+zgKlsYQWykBgjspfEQwa0ifp2goQMcZowAdToG05eDZAy52vjh
ObOVHI8IfOHKiDYjzSuHzhmIfj50NDDNsPMX0+UGQzuKc3OwHg7fINk3TEM50ygX
gucxauWtFRhd+hH4p7+Sz68c07EQ+N1nlgAZ/wVpwbwZTrrjNsVDzT0Tcak87Z3Y
YCk7YM8r5K4O5PATeVlzCal0BL8lC9PhLbyWONj4URn/Tg/iSmnR6+h9+2jHX2S6
cAD6BQ7QOT6p4exhB8Ddsg44vHdjnqgUAHXo/8OG92h5emQg6KG/fBCXdfDf+18/
7pzVq4tOVAM6US9+b2u6bAguoy6e69eeBVFBnjRSHqtoy+sY4wGsC5d2Vw1Sd2uK
UXNS0lmSETqpUXsSag6KrJNGCeuNviFFwmzOkI2x/4FPmpiMHi8KkXyGgTlEdSMn
2DKE3gWUwReqNBxL4kvaxe0pBkQSWKaKot8oosjFZmSyo5MDR9ZIN+KfxGQWDUcI
wFot49CpgB5t/QWVFnKXXtA0ZAdlAfa6pl7EtSiKrfmZwQuW4r6h5J/qjex5hbRe
FgAW2E3Pfl9ZZ4vHoH//1d0XRt4MqcCxS2LuHnBcxMztBrkwhicUMIJimGHwSj4d
1oPvYK7SWtfLv31HKyTeZHC8dcdKE/5JLXFyFMonlgkmR5AoTS7Q37ZUXbA1ueaC
/je5FwuThjBXnrK6yThRkTQA3eWeOFs4VQ8N6wmDThiq8abuSdnejTzWf8++MiA/
rjn9VEpguNJBUrM2XxrkiCmv/gMxe1drPqfm2949fOtvc2pwEJhUVF3DikTJtobA
JyjlQkCX6qb1GNsgcdnieUobaNNvrRCJIfEebsmgbRC7W9ZDoxHJ9EYPkc7ToAj2
iG1naYT7KBo5vSLASyZXjtPIqdToiCl+fUl4nPZ01+Chds8ATzdvtwcPsuWd3rlW
1tbkg/DggXT1yMkoUpHF1eFOupboJ0pi85TeyFsEgurIqBIaNCLh82KaVL+oiG5q
YLz9+/ie7L+J45s82uJhMn+o/xUkun8qJCSlPdoa0qK1g9RTn0TAvXR5TcUE9goO
LoerQgh+nK74UYEuhzfEv627ZC6rNr+3Q0+3uF9GIc763zttO90r/3A643IBM6gu
Ez+3+0wCcgTU7rgBSU1IKOdeqLvl5EyPYVpGbCHxwXStrPhrHMSQq3kqFr+EIOwa
jayeM+E2VLsaA3sdjorcYfNlsR7C4CA0BPCEciZDRA8zX8fdOEK4G18lar6wK2/8
D8AJSUWbczEcy6Mfr1kfd7aIMXSa+hBKK8xEBl1Tnh9F8q6J8ED+QbaQf+oBKbsz
pCZFXsuOS/chlS1YWpos3+kCgtpxMxtA2rumLF6De1hwzh3Hn+Lya64UVwtlSCyy
iXXPEIDhXPWZHWEyAFMSChsg1iA6fdPZrZ4xIz+sHtmXhpx2DJ0I3jTQONWG0j2P
Y6LROAYvEIaPpsJJUhaAXs6lx5kuoq7L0pvE9G2dgy9vg2sXbf8zrnkNwbqCe0k0
YjHPQns1wZxrJGtilteSvJXK06vBMSQLkOWy3wjcU9VwguCEQ18+31gPJVBbZPsb
WgZ/3B3QTMwO/LkDyyCVbgqjexNAfa+aXLJ14//UKdepUcjjjBxdocUb3cRsIjZg
4MvGhi+yEBbfVUpgPEwQiNOkmtrdNmBcwZpB+PYamiRwRK9o4HZcS1FI4IqBYDIO
ZVn9aEUa1aBy9KTzMXnPrcwfDXSQw+BtQW6mazgG8hSExvhbBUEVGD7LQ6AlQKEl
ujfwDUSjbM9Y3aY7xT+3uvSUMXwpJntlCW2sJKbmWv8vrTLQBLl2SRXZZkXsQH/Y
rDkdOYeIwumNVzBzY12VrKT+n7gPuZ9d07N7Svpf5qHBh83jh7cSfE8xKWILWdVY
Rz+10vWHKUB+ccVnyLIVLloS4AiMF6PeljdQosWaCc06UCSNSESshWZmSPxGWS5D
4yeECT1tXUgb0QJbv/5DuDBImWqta+f3RV7G7rqScOrBqHwTMxmeotdqXpjGpH5h
TfDE5G4vJHCk9kYwQcm1aGtNuacIyjjjd+OL1jmvsaQQVQDDmvDNqAGuC1l4Wdga
p20YKt1ZQDmuRNsR7UI708yrXm6ixEWo7TWgpXQzFuNCZ0hyACIok0rTWqr+qBxT
ytvORvDnKhryhe41UxVvan1MUN3D8nsw11+sVGlWCpc8fi5AvExv1UpHZpLmebXt
dExlXaSwHNHEr9mpCb34RMst4zq3/0Mxta50Uu5ZLEEZc004mDjj1n0N+gzKyfob
nhqipjQig5tcyq+VicNIi+FzSZqWrKP5GQ9tQrc+FrNg2bBoGj0ZhWYGDgVc++DB
8K/IfssydTabZT8F4wpCGpC38LTFGpxLcRyIfDEAVbuTdeOJDsE4igoq1zvtSwiP
yXtQGwKv15BqMwIuWlofa2JefyEg+OaB1Xunk9s7NtDFcKikf8c1BqvcizOkyazA
TgesQTDUoeThX5Js1ByAo6+SZSyfuFPxxLcT4UJ2PYSuaym9hmq2QAXYVU6eRjVV
VjM3AVFKoGwYrwrq8ZijB4pO4TL4itC5yvOw/651r/gEmQpajX9FH5I59kL7rRCQ
RE73PHstTe8NsJGsd9eW/11dm93UID+2dzBAt5aIFu5GkqvraV71FplFUp7hxVRP
El59+puNhASA0+FOE8GNZRr1a+nvh04jXc7u+l1PX3Jz1ywwrVLZpOmbd3o2Pt/6
uY1iKJk+/OggQeKSDdBkB6zetpt7ucRokt9okhhNqjAwIlWdjpZnv5ZZo+3EyjI6
W2gHEZPYV8gLUnt8u9dT084/u4cX4rSpIGs3KVs1+QRUUXAX+T1GUpmQJewmSOvU
uL4PM9UNqsRSp9715UFccKMS1lJXQO1ZZakw5AkgnDeeBf2sdIm3tF1UGM/trZtV
w/cDA1hoHOfY4RYx9DFLB/dyaP/YJFSH5I02qv8Ib1yeUT0e9SgTkQ6UsAepEjdL
6m8nYDvDjnFyhvOdFPusx//nxOymUM+E2KrOl/WrlRr4q/rKmqoatiqIwuptdHaB
APSizL4dCwtwgy3yKDK8P6fRU5cCQsYqMO/cyhdLHDSFUOC+86xDHK69xmUeqSLe
rod8FKsifM2O0lDpUvX+Or4RMwPJkP/cQBsv1FKGVBeEaiRMrehWrhx8IdCXj0Wz
6TdUa+kIlB+x7K991BKqrXRFzM8wclS+gs/cNjcXVoIGMCPJyKAod0YYd9WR+kzj
dbb5trhg8b+or1wVqZte7ocP4aYxXwFfzwEpNy12CgqvQ/mP4TpEnnaq13L1iopG
4ssBR8xouhvVDXhFI1fHMTsVBoQa0zhao5vSm567YD2VurGjkraEJGDfSJG1XZQ0
FnG7n/bo1yIoA1cxIv8BlBACP9uFVoZVgPX1lQWVJJi5nBCr2+DkSsUkb6wEuALX
5psdgN3u26cWfMbMjQH1FuMYhQ6KiXIn0RBymB53IqDpdZ3GcNQGgAS7BiC1e6LC
0zDSVMB2KWHihC4UWBW29rKrJk2aUCcDjm9VUzvwcFvvdqGpOxSRWPnYHux4zhUW
zGBrPKKC1oXcRfidTW+ZDxpO0NXQ660KufK8F/7XLunSwC5JEw2YlffFO7glmuYT
1n5Pa/8Gto35yiTftnVgWkjKky3DWZp2JTVIXXfnSlEqTQjXj9IEsGgbzPGPFwP7
cLXsdV7zUiSZl+udOPV2piXpJNx0NuPbCwGafkuvHtVu8UAv57rof0ygcNRIDG55
x3pduE1ZFHbsfoCWFsEaMVnf0vv+SbpS5/7IBQzntpeAk42Wo2LWkhK1yzYnAmEt
wcGnkd+CO2uHfR/D0aNzymM8fS6Bk69Ancxiz+yL7+DHDAEUb+bpDdQ2wkJkDo5N
iQcVADY3A/1k8HqvtTtW1QdAIZFjiCjMAN7FBidAvb7yNQ+AXyarM5RcgOJzRy0/
kZUwa1sNWRc2nxGO0IrV69uM0ujRRhLfrVaN5EVm4MuJQpUwOinwZhR33NBWuwIm
c3PcXhtzHaCDq5JxXL8EX0wvQCZI6GvEn7qBZrs2ibltmSs/sn83Ir2A/GN0gPlH
svzyIxaDAVzLa5M9LE8uwEDd+DOVR3c9ohHQPPFtH+zuUAfMF1yToKfQfulaxrj3
r7nQcNdbIKi2jPfpnHEFmQKC8TO7qWTT2ggfMcXGhlgjwH8sbtKzIUfVjy6klLNT
WevVAj7thvfUlM9FtARwqo+sRqWw0lZzEWfmFbhXpZBcHWsBWBNMjojKHDJ88OmK
eB1Sa64SQg+oyry8H0Tydwhy7KPXXKrlr0XMYC9DE8w82jBc5hKKInJHmDbd2R5j
juBhkH6CgKLmBpNOYT1A04LCGHQiRzzVgN3wqMTaB7+jDe0PIpaAm2+OCc9MMson
xIHjdtFjgfIThBrzZYCfJpOf/In8cP0cH8RxOgj9yMl2lpg6lmNtlHbDqfLTpE2+
V3OUnlfebpVnoSzE3jZw9LoOvaujTqz6Ou1uxni6KakR2gK/ZIa+u50pQ2es1Us6
bv7CNPIEqtO/P6pVnhVBwjTsaouCvna3Ct72c0J/s7L4UttkjwmFNfikadFBz7Kl
mLsq5/ZVn3zkXYbI11ZwYpzwJA3/4N26KeQFbTne6v0HwOQxUDnGm8P/44CbjwAh
MCyYxZ26QL3IIQ0YeyJQeAt5FTw6Ao0TQu4Obbilt8mNQh4MQI6vAyqvLsMTSPoG
vqrihAp7c8CqgY4SFqgjhOrFSFKdFdrvSUhvp/PLLKthrKNeHOH5q3r69O2ToBkV
jLRsSkPB6k4NMQvBJNVh+OrkZKQSNYfVXdC+sM7Dodv53eg8+i4xWc+N4ke0yo5O
W0Q6t6hxzMvbTMG+yBH4cP6Tae5WQHRZ74tzvbY4zOkQiCM1QWzFYxvV4ekEteGf
jt1rsnsQ9Zdml4+cghDES72v+z/ln/CHJ0o0OtLwed4BMUUM/zoeb1FQQCHmxBoJ
P0H7Geokt+UKyMFDlMlGQkyQLZMT24oocjI8bHzHo/SQ6/oxo5OfaEMflLC2U5TT
U0DUJTcqm9+PZfo6fzsXNc3ip0/6W1ykKhBLjs9xpNi9RRy7RkyZE8/mpr009jKr
qaAu/BW1lD1DPAuAn0TMgSdOXezvdS+0ziFxibw8z+GMwOm3UHh+UHvNzfhgdl4B
ab/XYHngVT3VNH1e7bYxjy4duHTD17bQc4fcQbukaCzI1OYu2qu6tdC0sNw5M7N7
69zaIm/CC6lVfO+WytYNnxH5yOqP47Dm3NVRACfDdezz4wEtpWo42FbuQ8x+al2N
XDxUZsg6oyOaASbIVutVmtGfxxkDyK3CEn8oaUPH/kZcoDrSeHCWxjgYJ7qkQcr1
xtbzsNT0rRXG23D2/9G7yju+6et+H26Tviqeo/IRHUBPWwaJC8vqC3YoXcQ9LF4X
Ct8ZJuiZ6gwwvmiYKbo5kPcFY+Jfet1pc1ScjNAAbiuuO3ixHG2G8xx+rvi5hgHs
D/35ObSLuDLWa+WrmD4RMD9j3jQ3tLyMjbGtIJDaAT7N0aACEttQs10rjgvM0djf
AToFM9muE8n5sZMLzuh3UGppMEqKefieSLuzBssiz+sNpY7I6h2k4PJR5fHrsu8a
7EFWrGh0JHI4rmRxs1Jowp+ZRwDVF3sxdPTqg0jR5J4fFiJdihDZkRtQs8vBYRuD
MoJdvYc8Y9EwjVlf1ooTE/IA8DODLQVttqvWDKa6GRcw/seHBLWqFJOZAk1GJwc/
I2JVTllbp3Ui7eWPZTvyFe9A5XpiJdVBAfaYiDsLEeNFq/CRtTzOS4+gvCnObpZw
sSQ1R/B1bMVyuhMfQbZAPsVsX1+jlmNMRRWTIrcfsyQMPaoBy1kWTOmZNSNs5mdC
JISBaazbtLaITWShx6+wW1i/RqoRYWAPAJgWR6i97vtraUHNgnOdrYkE6TPJiQX1
D7GMyXa1x5FD5oR1kbrH88Bj01UJgL+Hl2TXnkl882BapElgyqX2caCq2YGw2dQH
18G/LWc2/hEJUsBZVmiI2ePG0FwpYoPqiTG6py36y/WSw2+jfParpFGP7UJx1Cui
IOr+mOIGzmAIVuYi2WJwLVNZiaofjqSe6HGFx5UTQZPjJ4XxaVcGgWaWwqxS14SL
dxKZiQ2DlsAkVCh200i61b1fHPacaGu/+5kFD/8NmGk7hMOZkXzp77xqjlJFuOKF
YnpRCM+gr6bwwldG8IQdfvEQPtO9Y2eyNbbh/ZYr4WU54VaKa0unYLPgUZh46GiX
OUbGtDnHTlyL5zMC6jx+poPgCBF1fsp9hrMg79qEgcRhPk03Xlljkvo7AlrgwhLh
tjHVI4/TM1gWqwcCgAnQNQRd8RZKnUcbKu5wYfbnEnn41N+JzdBnn2ed96skp/UT
s+A1su7RSO/D44/53FzMJBEiL9saiblh7LIoT+evw68HRD9xU0fQdmHvre48gXew
/XbdTx1xCktWjOOwqgYeBwb+4iGZCz9UTytP1YLtnO9ilv8c7x7SAxEwROovVZMg
aWQ/NseWhhg8FviytCGMZtJDy84scnwrufvv5p8ISekQQzT3nXdjmKeeCOa2QIZw
47PLNN7JjyfsclafzwRZbz9yCVyD6u/Rx/KmEyRWVrOyDy6+Vay2QQWlYcE48j7J
gGZSp82phlHvq7zImir1Kqw2gFohH0ujGzvI+lNVzk0IMJrPgiKYPFbdHg7wZh8T
AKNJrD8CW4FFzxKvj4c/kYIjEM0FRIcbbPM6kRVM0WmRRCb+MeaKE6bn3b3nD4rW
U4kg1Gd4NorgDvdHpE6clX7ZOX6xR3zmTDzxhh/xuv+5K+o8X04aNrEfoGqfJBKg
4gsjSff+RlSXjDvfouawaoWzc4hAPkUg9ZpG1xlzE5AD+ZYWYaDD8WmilJDDCXAk
9XBF6YCDX0qlFDUkrVWGNW9lr0mgHQKGqcBkEeIFOUQYqRk1hrIuZKC1MvbADUt3
MiaPmZ5NYhJoTI2YZEmMjp/iFsI39U8kYfGBDzqMo+9hYuq9XByIQgGzCj2yjkg6
rl2lWvd4gq8vl4GkiczSeRPmDRpFBOlPCVOKmnBiLvkv4Kmd1/3GSMLB+9xxLVP3
NLIqE2Vs91bZSVeyEMmiDvAWUMyToIkm8rP6IgOdK6o1wC0zR1kGgi3hDuJm4VGs
gDKJIpBBEXYTlLT+tQ6GjGKRjU7ZijEZkFj+yPcehuS83sQYq+d0ktPBN+rfxVXM
nQqIpbFqho13QlKw5VO0pxsnLlSzTXQVOZgaAk68dBz3tQYoZQGVEt5hnWJnUj/I
oKsPITHcq4jjwMrCgkMk2keu1By3RuFGHSxBDw3zx2PTsF6KEr8nKZPXb6ZtJ91y
YG/Huj6VIpvbfCeJpIbNA5OdanJm+Jl+BwHjwZ7fVY/gzdD+wM/6KsEpvZashK6E
ASyE/E2Z2+Lczf2L5Z9LTPK+V8EqYi3ViU4zfTi3iagnb74utdJqHSV0JLDuKEQ0
FkLAF0z1sxMyH/hJRFp8nCQUySq5Z9AHB5+Lq1ddeSGv1c3WugWGOUCXR9w/Oy12
hok8pcXWoCrBMCS2nloPE5rT0nNji+EmvK3W07Q07LbsiPNBVokpIzMG/0UnAR86
+T87/8nEQtQQsNFXNVjMmR0ggEIzWZ5U8wBHz0ZnSSLatbDi+0+HRj6xt3agB1oL
3iymIhXusD4Q593aBo26Oca1ErUyTemtXgJ225wOnIVzyBvpjDeLyyE0HGj+s5XN
9599LvlXwxpiz5NWTLqOVibVvxTF3Bd50UQ3mxKNOr81nmiIKLzgggf1hcStAyTF
3vrlEUNoylk2StcyUmQWJMTvzYogdWwAglwftSxxsg3USeMwqTfSRqYdMKQR0Nc5
yp64IrJRwud5FWQgT9iTOVnK9s+FmA6yFbs6vVsQAMIo85R5zvP+XDPPVWnE1lbf
LzrIGBLvH+MIGh7LsTVbe2SYLUvJYJaiAz/TKP1tJiOzAyCkv1T/hapLRAifBjWc
W9ow6n5/gRNjxwaIZUhMaMwrvaDq3C7uVKZCycFb5sy81SIA/gxz2v9p2NVCuU2d
PzuRf0PyYoJ61+36mnv3iUtwt0H5poTmJY7rr4gqzlwEfi+mVcSd/2fu+c2eNLbL
Z+SK+Df+70pPouCFs69CIF5SLIhQt0tU0wE/eV4K3g/N4mNlWQz9W6ftjjBJh1dH
CHrkSCoxde/aUOYnOX/TnpUy5i4WC/yCCCl9nGNYifQDWowrH+iRDQs+WE93buLz
+40VYs5SJZ6OpeTJZdP2uV/ybVJCjipVjecJyG17aNx1mZ4PYQ7MwnY64QOXeqe9
7182GVKGJRpnpmf8z4SdNVoOEBieOKjUhHJuIQKSP3i+zsyoI3oroBNJDPwqrLyW
5CAsONv8gp+XEIbi3xCQU1bUMthcCPRergVhvOpZviBhm4mIAsTHuKKEObqgn6z2
ZYQsjsNNgB1YpHcov49hSH5cpITh6E4PiXicS9YsS1GGjLgr3wL/BRx6AGs5C76r
7WvZ/T/p948fGovUwLj1VUzmoZw/GapiySC5MYTv3Gwf+vy/tjMf86ZCHQp7zIpj
EVB04puL1vBN9JopHIcF9JiQ3QtpvrqjmqrY5xBCwf9ExGbzxwv/0F25+/yYxy22
q/A6BWPuICghwkVsg1bXtjGUMXUsDNoWwm3zk0LfV+oTi9KPnXF+ZfsGYGZlBE3O
aRkb1wCkQsIcwsZfiD0lOX4JCWSqNJQgaM7b8PLPxuFCpKXMFkNnjw+Urh/z8K8k
wMKPhSs7/1CgK8v5YON5v1D63Jp7Hx+VIPyGWgz/Co5/8wmpotY/MZwo01qrKieO
syq7v9Bhs5FJWfuJKQGP6IM7CR28VTgNsdXpsR+gmiJ0EbwQagaTS8Yn4gHg1mcg
BHbHqhpiiyaQRSOJm2MNMU2tyX9uxjwiXXE6hy3jXnI3IorhKOWQPHn2bRFY2ako
btxZXQcd2bXl8MoCzf6fx6x4zoyFDUGGiCpJQfmNSd0KNNTn0+bmp/nqZ2lcdf+G
YAgMumoMeqMJqiceWjH4EwyALookUZlcuxjHj0zDiDhT62MEH1bxSzEEPjtJj0bf
KwCnmTmAYLCMbWXUI30e4Gku49cvD9FvB/UHndZlCl2FB/aUB2V06uw590llvpbU
6OxP+DENGtYnXkPGWAvSudmp3pdJcy+0K6NPsMiaO0eEoPdhdRdXk5NNPMgzRHMi
jkUtgIT2bZiP8cUR4IlR1LX2l+UMSelqKUHYinEwP8oYNpCekIN1/OdArexSRHME
BXGNc4FaKE3B4CcF8izgUfZwHxlZzbz0RQIrwAkSK1mQSRGrP5DqDIHbPE8CVAtM
DVE/YThaoytlh2AdGHwqJsYqjMbWfvFa9NuY1yebVb4/3ogZ75rSwhhcD+OBwwjK
atvK6ebzxfy7dD4Yu62wNX7iJdcJHBQpS4aUronk02Y19BDxwNSQgS7JdfBuXLFF
kdE5IbUBfo2uQZ43B/+GPmmONfm9684WbtmfhJ+ems+01wscsjXeQ5N8n60A7En4
vg6VFApiiZkFUW5T25cDQIOL3tq5mEHlrHaIVOBwun2cQxrow2Hva7/0D0XdDz4Y
7jiWmRpxD7J5Ef1esa6tjTMbxQ38KlD9EkRXNvJaoHzzC4aqsI4AlrTuMKBP+rCx
GKo5qFm9KEz8Vy7gBnf4/iu+F3R+SgFF1xyJTJaAx/oXAgg+ehM1FJLlCeNVXNDd
8u5tkhmbeOQtfPZehZCbiYnK9AbQQ1sqk43CEwBmseT4KevlzZWJantTyX1D4cj4
6whXPwRiOywAsUw+fgZfIFD21aV/sqtE2X/PdRjppikP5uJc5FrNj9e8Sd4JTnF0
y2c2Tiyq7rR/yuB82fEf6hVDRntWw4EeQ+j3y6/XnIFRIyNb+6zl1025+dAvKWBR
XlIAprGs1BzwGHJXimnXkRlg5uGiJEvu8WWI3jH1X8vbhF2dsOhcjLazzDfCGkWd
nehtwONPIvOwNWcH3xPKZJOxUn8j+NoysmSxqb99XQ5s6Lmoam4QJHfprHOn5JY2
HvLSTXiHtInLOik7Ahf3T0J//Xk7i+U+AJ89s2fEpCKhZcx6QbM0AZtFN7Par7bP
doCwMXVALDn2djSvW/YauB0hBqL6tJl4ReGSdryrR5dwzhshsoeGcHI02VQng7+5
kUgNpmhhDWwAcSvO6+2O8OM0mYdA7OddHb4KSip6/2lL0C4+7yK+FhBX4rwC0Wcj
KQGsbC4IFZYWpR145P7SWyLq4rxWStPrmz0ml7ba9Q57PcjPllMBW96M386/IFRz
VVOgd/hZ3SXPglhiqQkW7WelL0jjWcSGDkCkcwWAiywLbnsXM+7WPo5cY/t9mx/h
tg/aM/MVdgebQC6MuxQHxmUheFdi14iy35fVOXq8Fno9E0xl1kF9j1qm6m4oweo/
1xKp2w6fNx+eOHqmxaO2cgx4cz13dp/DMcHZnOi/YFYNiN4zApfQX0fQY8oca/bS
YDbMv7mEV2tZjKM44519dj5Yg6J0lz7ZidFVbRR7r1ELGzylKgSuKMefnlNvdS5r
T/PgZPhacaLwlZZW0+7vbsJomZiI3cJPjkeX3frLxr085yEVO/mtHwgGFTY847ZQ
8vGL69peLcnp2QrIQpG024h78RrqtWmYWc7rS3K6DHhSCCmMNLzqx81Vivc4rN3w
DNKtOxmpUFC1Xf8SV3D9MaQiVprlfI9Gwe3lhsdeLweC7hVXnen0ru8phmq1zhQp
p5WLq/gKGomlndzqprjxCv+qx+fghCQRDZgIxWU788Yw62KJHCqyd8fztvJt/WrF
iNPzRsWWrnhReosAfmYPso+oBsYRINyA09EhRigBrw/cz78+ioLQtNBNCz698J4H
sAkCig6ILY14n1+Sw1efUyVV3DrnAUl+jPv0rp80/FksXp2q0Z8C/aDVMGZ2jIaW
UB+bhzT74SZzV2Gx0XaWt6KvSgSDtc2YD4/6tucudny1BvE5Vp5KrbwpeHxQCoC+
rlRsK6iNBTVL3imqB1ZGfBewUWe6c8O0mL9aKFuVfVl7IBWP9v+KJpJVk491HEj/
de9j/VPjuJ3Jj60QVXjTdqziK7OtSbh8wsVctnthbNwA3u1tAy5eNGmZPO+C9Txx
THSo5x6SDpz358aWkfWVItNeTCPlQX0X0CoMtLXKck8j+JcPHUGjTNqIX7ITBzcN
eCcaD1lDReH3V5ijFqvaOPBflHVgF9yRithcyTwrgv19OeHPUp3ADFnw6CWOJs2r
QbodsZlf0CbkDD+f6EwqVAMlC2uumqih1bqMZNVY+9hY+RXWrSVLntOypLByfFo4
uVoN/5yir7LLVbgK17nHEIi2gLRwGjgEJMo9Wyh6Jk+lKdbduhHgoXk+QTkCd+uS
4ywUp2+D/FeLPj03CwmEglfIMdfZUX8+0bAJwZHgkG5+zgsyOANP4nMRtJq5MZyf
0ynXTyC93mRSeOFW1rfj9N6mwUSjek0010ojWKFoe5A5S8TMd3etfI46KhyExBe8
cmrI0KRAgs5QzlrDLr58VQC3aDyXjYZN8Bv+f8Zfv9QDD4+sQifLAM/PPKL/CnH0
ppQSAjt6e17A8S6F6s+6gQ14QdtendpGLsJAEB2T7D3aGEi8s/Ut13cnprszJP6D
ew22g23lNS6gjDgyUv0GolCTs8rZWmxFzkIRBRpO8QRIKwJLp51dyBf7lDV/eRZj
F3TwTQCFTNwkFGHk2NmHo+8MWkiKM9sEeb7RDJ5Iq56jRKqUAeHRldZuKE/yGyoa
hB+VipI7sQsXYpwQBFEbNWbip49aqAa6bcIBvqWg27WuX5ZKREeVAoipKDVO7drV
/kfja2NV8AeF15ZUQX6jV9ghvL9IKuGwpJdV75RyZj47oQrO3cUhlruCBilwzx5l
ZXWJQJ7rqcDFRUNt3RNk661YBaxKlcpC9Tnfnies5jt101+Sr4src1uOjKt0xzEK
dkN5K3YReqDFq82JM7n5v63NdaSUd76nUZGV2jgVrvWqZ1v+rWJ/PtLapMldy5GL
3ebW/HziugnMLIyMTr4T/8wkTjtuUk1R3zwZavXJxat3082eSq/kyglmdv3WhNxa
753bvIWJcjiu00KrLHgUnn1l/2wZcKMEYKg4qdMDKgtN7MeMMucDoNwEI0T+ZIRb
v2/nqrTFQ9e4puelgyrCP7iIktEr/nD2u19OfxoCu9H6uYVa9+CbFpri/AA+3Ujj
mS/+OOoHS4bhF0RdlPDE/9EYg4ZAxO2PSDoA96eaO6RtXf/5vYwJ2O4V53NER3ye
nFGlxNZONoykvsBJU9SUVGkQJPKEedY5nndwe3oIGXVhEix7HTX8ZYD2xpmxsi2n
z2MooeNCtux4YdZa2KGXPFEmCGq8j7FwLBTBWhoPKWCYUoHNuheI2b8dWl8LKnYJ
Ht5JgCW1liC3x0nbkLo4D+3IqUBZlnUAnkQHzFNGSy3cvUiIfYV9CxoKoOe+SA8x
fxmcgv09NQvZWFu3YfQnKZCOlqfvkO/rfsR9iluWG/GBdWuBCcCCKYFvvBpeoLPL
2jH1Pwb5wR8CJhbXRQjD3K2HO5irwll6HWk1NgUUh0mheZpDuzFoHjsFHE1NV0cH
z2O0PXkDxdwoDfs7eBTrBEVnNO9Z3VBLLC/nQm7x/scM4u/LjRJmZL6WIWjZiUIY
eUH09aod7IdTd3Xd2AaMyuCyL9ONVm6W57zD3M/oMRpFERkB3UJKs31cEM55G5kK
WGn1LJy345Mcuf7HVzWhe0lOpQyUJ+O+szPEnFE2zKiYA+N0rJygbJNu3Xyn2dUg
BL9kn2xQo82Gl1VjW9UsqkDTEYzNevmOVebFi0bWASoGQLSOwMQt7/bd/bzX78gW
eK077NCKJS2e1gPC3h2ZREqNTiTjdRuRG0XoiD3LBwZ137wBGY7jK4JELzOLTaNX
SuITH9m2nEBumYzOtKbC3p5F4CJ2WAZ1YjO3eDJn5VypMy9yOJav+zG9o5pfvdvc
bH5ep+MzqflMyaBEwzS1W5AGj0GBeTjyFd0AJcvfF1kJpGJ549QyreKJ5XlEPKvs
qr8igGxSZB8PB1AmAA0AhvwZ7TX57CQ+LR+wSgwuKJA7e7jgLTYbjBlpPNsi5X0W
ZgH58I9qu+7rqdUKEp0ypcOjWc2zCCXV7cQwouC3RbBF/8lLuK0UUlhObC2IY2q9
pXU8WPnNczrNG2Bu83v8j+hbL60uiv5Z7oM8a8QrjOYBTUAiInPFvvTi147x5vqQ
pznHN/XJZQVmi/8pfXA7ZJr+OfHZjWixTyXHjJO7oJclu3dPHNskUR06e6PCM/1X
5CHZKBmtN3T1dSNeiT545c4TOiCyOKB4fmM+favop1HGAyiO/GYKin3xEyO+beH2
Gc5/sSPM/FtagqpsmiGorDIuU1D+L5QApFNs4Qql0erWVrqlnQCAzRCa4oyhJnyw
A1oVgx6UiAV/Km60xlixtk0Y/Eb1SxczmxepUFW1vyHSMHviP8dyGOwOXbPM+iZb
sBdGf9uxtgeWM2ydO1arpEbCghXCuGUtp2O1tAAB0sGChRdLlHJYhu9RJ0HDAirK
Tx6tzxz4kDFNbH3RIhzFiv8Qb8UxYWtiZaPTSIge78GAgUDHpS4H8I2shIsX6D+v
wqSbgyua333Sc4H0R1m3XX0zJTBVkiQVAkZ70/3s3OXTZ/x8HbBs/iQ0F1RDWj/f
ktQdLge4hYw0Vvu20GeAQdduGWR9VzPoOJg2be9zeX1Ct4xCKzWgn5F2TLsDPerw
EyTh+35p2fk9drJLvIrDZIfQH/otiyB9Vb8CwErG6u78QgOWwbtU3Ca48ZUaIw5s
L830pYBB00Uu8hQEXTaz51e0hrABXQiX0q2bvhpLhY8krRK8lYYJ7kmP16Zcv+Nb
5g9SsOTR6ysZy8cNop7rB/+XayX2CiuTtrXwQJPqvYYkI0BaM2z3cK8UaYA1UAhX
lKW8jPQwhPXI3wQ9Cw8sTuGqBaZuNNC+knII6L6UeaufDmPEVNM/+LrxGAWx5xIZ
MLyHqDZpplAKhiLOSWJpyQndgGHWfPROABKSpg9QM8hj6UOor9YvLis+N73qU/58
lsFqVAAm/qdBxBInhWeLsALaPkySmvPgAuoqU7VO7sBlDCTVlH1RRb2RA9nD8ZVl
Wa1jWaHuza5YvOY+GgE+MxaFcN8jajrO/ZIwGXLVeJ/3xLDZH4yO553TroATTfDz
m4IoK7+QP3+33vKdOk0Jaq5TQ1YLH6ZM8y/+95cYU6okJfENVVIK94fc0qjhvY4/
vMO2qOjMkf31JkCaDej142e0nifoH279BtU3UEXtK4eKWKeo8BNCkBuU661qav+j
rQCjPUxaB0JYb1n2XDFqkLeI1m1pYgNNjIw4Nl0/2dTWdWzqgD0xzha+Du/j/R53
aeT12WFxAyrcgBSgvhhuHrsPEpZRQw6FQcPcEC5APyL7uCcCLmc5bpzRdfuaafx8
RwHwoUc+78EaR7WhudxUg0rN4aC3T3KIFIiXEjH8uDT4OJjhtSORoRUeDt1gQdWW
a6TslCKUbjUDVnntzKytUvjjnlSkjVWLyO7wwdgm83TeatSntoByCEc/WbpaGzQU
hUQQ+5DuEqnJumZU8mjxObzgaHq8MyF79aWKeUM7kO3oI6rLvQ1vJqP1L+uCf3nm
fFsuS6Py+B0t6Pa24gvFjD5A7WJmOeKkYq//XRfA+0QvUYZLY0Gf7zLMuHJC0m9j
F9ziIZqovaE8m+2agrlg40vcRHchF/PZdXO3pk/5PVnOd04HlE6yZZKMiT+sT8lb
olXR9Qv2BZ2LhOL/4v3HE6VcF/hofgTSW4rvbVcVKZc7XjH4esCF7n3oCIqhc5H2
kQdehRadOmqjXT8MeNw6ZLcJbm8eMpg1TiK9mrCLN88r2EHzR1nWih/RryDDE1RF
IF7fDlA/WOBP8c/StbLalwDlsqlj+E85eaHbklf8N0iVdzy9uXP94TfSE35y3kew
VPwkHoXQlupAWgAk3g8KwYfDJl1tvK7BXAaCsZIWEDbt0oZliv0ph5Qkoh97HEr9
w4wlroH+Q6DxtsevLpQYR8puv7wm4lezCd3YcMZWkdEWO1P9AXbdJqV9Zyl7h8Y2
js9+xBvUH+QqHnBYTaSeBWELKPx92pq0hnpxgnalxVuZS6X/NqSqPEP8AehrBRGu
DLleLSXQ7STOo772ml1I/vGsUTrdubs9Z5xbGBWCmAo+rBBqE16FkDXeAF8wRHJe
rRMKqlqigI8VYICto34KNRH7UvK1LoGhQVmwJStgycK7XyF+4isOdizugQ2BHGP3
NdKuWqeX08IQRXCu7c/8kneOkbZp+CIlXi00Z3Q+ngBoC6xn4PVSoMYIXnrbalNF
ky1a/E+sEukKEHbtiQCncfHgzMXvspeQMR5GtxO2jC01+usuCtBCfGyynkwnL8Lk
TUYzuOCthP0qsiHEkevB51bzawaab5VH7qUyP3jHD7FTWvGlIlwDSZ0GYxy6/u1M
bPJXZRqPau+Qso51XJQY199KaQ621lu3APY9X7DOfXGu3CE5rEdaf7nlmqfjRVco
RGRwQOzfKWfwT6iTwm1RlMbTUEvBQtUYRqg4osx3TJ/t42jCC4GG1Og0t1+a1eeu
D0NxIKqBbF4Q1Be7yh18LPkQqcWtf4O/5fEYpp4mJSfS5EEmFpiABoquQY4Bn1jc
JcD/3OOgodcnUHpaFzZ3NOchYBM3XPktlBb9lJLqnDtwbKcMumalEAebjhKRUlDC
gQXxcRSiQNHfj+UOem3zAHgR6VoVj+5AFJd4LJbxZ5kymF0KdcOun2vc0kU9RdWY
YpAmekyDO+zPlw3Xo9yfAaBkoNXmtek62Wrfo9eEy48AH/igBD3nhoNJo0pw1HCs
GvB+jy84yw29GjWBFb3ogOxDYO7XfqLRrzdaE+DRhBin6BlB7k+/kJFjm/J/kUd6
dszl2FGKyZJ+Lggy/vqKH+NaWlOn2DYQaSe/rDFgB2Z51ZSu6FFe3Dh0qfNYqoej
4wuHkyYcfcxGB/ctff01I7M6RbHoU2Vqv7XVGmgvI/VERovOlG+pIrhjuAn0U69n
dQg4cFUmki1YZpw58eFF7BTUZuSi1tfwy+o7d7ImLc8N53yxc3dK/axRkXiUjj2g
4BYL9FcQf7uUP8BuvbQdIBLIHKg/SH+8N6lHIS8fS2OwdSsYSit0qX3v89DDvQJT
yO0FCt9C0KXNDBrksVL45vSSY4g1hPdUMvpvPXSm+oEI72InsR9SEjZulFnYykyO
M9pR7wj/5GMmoevyp0ZkqunSHeRr+cY8U/53Xd8gaQ9GXzHoL2jxZG8W7y0CEi3u
MNxoZ3Fg2/pZn0iHApiTFxzWIphn5V3swbw3h0Mn/FPT8/KItbHM5k/J0b6aZjxQ
8YXlXFqilQ8a8D/apmD25UYCVKyvKLRl3AhJV1bmmBA/V4ZFpkKPjOmoT2KUTTAT
X8UnH0g+q2VBoS+sFX2RUM86cVbUzKSVQczvCSY9QtwIts2sctwXf7IUC+ztmnLn
u30CpG0jpqqQWGFrYcAZ312v061ElaEIh3F/L1w78Rvazy2iN08DHU+lUvfzGiUO
UnHnKDkbznMPOU5AkYbe5h641pJwITHeKhP7hgtFULxRmdk0pSYpZMgbZHR1IOGs
+y1DDWTWkeWU+yypjNEwkExtsWaWnTAxDagnGUAoCW50B9rfUNSETV5x6+bZ4fyj
uvXcSG1mr8Nt8pbXSJXWuTMGuR1Z23srGf9+aYZ563fmWdLedfD0lfDhDp2T56Bt
Red8dRnYvUaGHz8NQ7TYyTlsPqYNVoCdWNXite2Q/CRKl27ot9PHySUiRn8yd/ly
/uXojYN3Wa/HKRGgtuwnGraokMUXNhQWQ4m90QF/Oai5o0lCyEdrEKEob1HHxOFo
Zx1zMtB/RM3wM9qSmc6nIL9XtUulx9YUHjO7U7Z3StH9DCLfRtT+hwjCZk3/NYT5
nLUSBOkwJvg2LsOhe+P60H/7BoOgAW6P/0PYvSIY3NjBnW2KrWSjHxGBE7gTdeiw
mLNB8TCLpAXd6/Z6FIC3Q0/9w3YQBeND4f5RcH0TJfFDD83ys7wVzo997BhNOehK
bzWRNgwJ0CftuT+6YWEd1JC9PEnOAOXfxj79AUj9X4kBs2pv81LWBxGsLHBByOL4
JKu1j0Bso0bCLgigP5sp5dvDR3ItCiOEv4Twca82fn1bzr8bM/KGela1odk3lz/T
1zVU0jPF4OWA+amD1wyZjLDmJMQP4DCQTci3kiyejd6GkMmcI4KQ5+x1IZirVr+5
68I2pLEyWUL1AwWP6P0G81uCl4hoMAE5WeRK/c07Q7I0uRUdncR9CnFKE6TqxUej
YEYNidYQ5GYRmEFEySbe56LgJRx8hdwaLaQxLmo8VzX+JpVxtjuDaF2uJPSabrQJ
eAIDnIIRaVe4Zcyju9I4hg6XE479V2xHC/mk61swE2EvgS++2sihRPaLVXccx/28
3UX1nA8310wvX0tjfCBWfNckH2vZ2cWoPCmhG7J5uPOPVBR8TDnAWJTa2tsNX8No
VK+Cy7xf6cPOcSDs0SPNbZHb/FMAd2VqaEbf6mxk0cwA556Q35ukpNIP+Kc0CI/c
V8KQC2RgGd20Z0O3y1frnQ/fkwXUw221fHvpIwTgCQNaFjWaypg8PhTQrzT9ZsN6
DOmcceYizMj82xvdt14Xqi0PbUEPYE10j1LCa3tkyTyB2BlcYnuyYQIOy0P+X/hx
zcw1o7CqaDUmY5hS8pGvdYOWo4gsRxN9PoPzid378vHWaCAk+c0oJGLJbrMYjHvN
633S3dEwotY3HLnRsEZd2vg0Zzka9DLouW5kXzVfs+cJw7wY5IBXL8faptYjz74e
F58cgnM4vMGdZ7JcuJPZ4ziA/Cxg6BLz80SjCmB62kEyKNLRKkVP50lNhVCUXhG6
JHz3JsCISQsGx4zjczfBGyaPi9M9RA1bjMCggUrFZpif4xqa8EWO5Cg82z04ZotM
5HXMO5rLTZqkLXPtqBYclyQt31U56fRDP8jiJ1g5EYEToGmEgDrb1vcHJSSp1rM0
w5xuUSYyyPBY2RGmhzw6YlPjkpOleYaXUUDaiUEift+X5C0F7in3UAiZEiJ5ZLD7
7KwYNL1mD2Y7uOuBXLLUwW3gHNvNPwBgdcnM+ej3T1W/re8ewS4CJnrKoRhJzESX
84V9lUmBfPyPvTlZeWiP93+7+ogZJIJS+MDVI6L8TfADaMPYzI7E8iP658BG3Lvd
JMc6FC/8l7P15PVhV7Qqla4evkYSGOwqkQgHtBkOncftDXsKUO2GpAMTxIfKCBJ9
SZuaOos5e19jYnlY5s8V9YK+Ehxz/R+8enZp9+CUr5/8WMP/fwK85gV9fyhewzs4
7MeO2ESzg319ZKKgkZazIpx60N6fPaV3XGM1ABjCOGjWGkHV31iiJRoXGKTz47zG
aBBbUVCSLFY5uMscOaItaNKt9NuRforzoNehWP2f0hTGkqbyjrHAVVklg/Q9RvW3
5qnaBbJE6PIzY9XWFdx+B7xdYdxnELbqGCQpfoYrehwErN13fzhanQqk4NQIC/T3
duZBjnKlJBlFGxkumYACo4BlqD57XWP7Fa1Gb6T3VZdxw/TaAN/GtffDsO6TCrKz
ap/KLZDrFMQX7uOi5OnAE7KPiD7KuMMrnhqTV6IUaNIUIRcdefMSm6qve5OYRhJ0
MY/5ZGGhwy80Pqdk7pcQ9I1dZ/68r+q4iUHOrqydKFQZsXaA1hCjWCLN1WBtu55a
eZT6W93Q2EWgA1s7bD87ekJSDs5gtzNpUvBWCv0LHcIZO7b3zWbZokPk07Kl6lKE
7rGgDLXd5qqy7ZKPISAT+Kdz6bjaKI0OBYIWu0C0LxKz51UUYIdSb4bpjuAiYs4/
+XwFJKMijbA8QLu8JC93rds26/P/3KIJ+EdxeoNwiOKLhje94U6qdtb+1I3qhOwz
HdH9M8vssWKozQo10PDj+XzNjtsV2DCvraaI7+bzSQvCBjMcoerbJQPUfKll3lgS
MQANCX+L6Fj7fF3lfQT6HnATO5E4Bjl/UNXGKkSJMfFfJBlLX49n4xUpYqoxC7r8
mvvmMlTXpkC7KLBK4PyBE/iN4eHazgn2XP2iHvMQ2wAD+ehuz/7L2NHh/Qxcw436
EXTwqAs8EE3gx85hEG4E2lQzx8X8+xF3kGvfWQKulYQ8DWD9qrY5mV14FMBbWPV9
FnV1/HHBicupZzSRSXcwh68m72Kg86dhN9y3tH7/AXTjJVh5w9P5fdbj4v8hT1iO
C+kxdBEjm0iyC+xa8i57jCig9dvT26h4AYBn4JB+RMNOwVp2DN0mdCNEAt4sL0+b
ng8vzdrIHsvVkjRidgdK4UYTwHMiXHZSNzUNiJoD5iLxWFFjY84abF/CLZ+VqWmB
GkJQ2DYIB6gRHcjsNBn/yie/5PFt4ZRh7fSQdwwE5u+4vWnNBdOyLt5tlJHh5BH8
k64s975VtoD1hFfGTqkE/+se0St3fS8tG8c6VhLF/1TcjK+7LKSFIGk9eiNTV/f+
LPU85FwwWw6hIdVPC0iE/GgfrRJD5+9kNeXfJknlBcJtG+YyI4vnEiZ+b8IVW+35
4GEXgQif99DDKWdo+12QjaZWJadUBWXzdsZt3C4jFA7CCFUzD5HMKZmLPJBzbL4Y
IG9J7lAUSdBdexLcVhYPK29CLcbRru4u0Gc3/PSk51XH8EUcqa9HytT+aOjnuZPc
WQBcg71uAYQML7xafejTkBjdQBPtfr3C79slYwiF3ktQMQo9UbIFPirg3OlFsYbH
XBs36h4GvAHTfeKxPLhSQwMkoF2qKSVhsC14vm99ECF30xDrN6BjdA3NDnwJp+VJ
dOaUodgFrN8QAlq/q1M+NJuUg9Mn7Rm6guOTp6aPdbgrBirOo1B6jTvtSrEXai58
B3GdchwtJ4rMOmqoNJyrKbbwUutCq3Au+fp8W0+RI+2g3JDPUxZ9139USkpOPdZO
31C8BDf7sJPXDuNxB4e/JNvtge/Xyz2SWl8pul9Wa6W7IzQamynf+DPdOcbUn9NN
T3eIazi+SOSAN2BD19dfS6c0dxtYB9YyPLA8mTNaf8mEismu0eiHQbL+dUBTy0Oi
s+Cw94fY1keBH/xcG6qrYPft3GMtXyTMWBiO+C0xe9LbLruw3y2ONFvF7gXRLcHB
Va5nQGmXFuCd8frWzLkSUe9tqjkj8OouEyTHaIBOs+9TyQ0fY+75j09DWxVZtS0Y
JGIfA64a9TVfPHOtwLF8p/UptgcshzfJOetvvzIwz0K1JapV2s/fWzsfPoqCXCdD
o6XIg2RxHGAdzJPQ0he21txC7uPfEaD25aoJzsiMun1C5JOi9/m59IZrKepOD94T
bxc1tYSH+FvnFc77Npkk8piY9xlZOHP9p5II/22IS/KSKr9JFt5qLKA6SaczSZu2
bnIMZZqBwdN1XrczMNI28W3yk6q94vFomHjzxM2w0uTjYAJ06B4bpyL+TUV8EfER
Vd2BJF2aZ6mpxtlHsSqWpPY7xums+Ouqcut0NyUmN3S1uTQWqR24Xk+shsWyxXY9
UQrQ3SoTmg/I7ULKgu94IZ8BqVaxtD8lr83PhpbAAvBQpmKJnIckzZqk4PoGERC/
NWewVztpaj4DGZonnDcoToBQAtcbBWpNDIqwtpK1D4WBL5whxHIuAU1QN80sCdsq
hq+Kw3GVX5i1/LZFYsdHwlHA/07ZAlp+dQ7OK1gjc+bcec1KObmftU5bKspVKaRA
OE6sj85JjHUPCiphTJugDA82EdtKhrILC9rHN3PsTpgEv7C8x+PHyGuOM2RZcb6S
UVR88cFgXwn5pTO0rgXcLQLD1TsKxelU6aZB0M9mL2v2d7BJwUl0Y7UIJeGon9jb
vB6uF1nRWIdDV21jKyj4SX9UTKst/oKglxL/AznwQgd+IDPtxBQvqUjqe5H8ZXlf
oEA9Cet9o4JZiNn9R2LEFfC6cRtiQF7YtP4GpY3mleEwzPf5A5vcPy9tMdC9LRGA
qyyu/zKkZeUfGPw+RtdNowm8Q4AlvUkFGlO/CojiDvCJUD5h1AavGVmUQf4JBpkV
Ofcpm7Up1787XqdtRvnaDovk6Z/QajTshi75ogF/U2Ue0xrH8Br15gKnkOTA1cNQ
hPDsdr5j5NgBK2c81MSKU72TzrMJLqOkZ46wxcY/6/V01QgGxNXxXbe+g9q4Aj7o
T/CbIWyZdCGMj/6y2kXHrg3JJSmAxR+YsugKkQnGyU0dj4R7GGrgCzoWtXTlXNHX
U3eHWxidhHJs13uDgaCE0KJvRXkULsLP4v73BurB61+mPooxhOdkNbQYvQbFwZoC
eK3W+12aG+lTHcql+yCmIa1tnN985R+WTsLvc1eP/YgDLViiXMYBFAvumSi9r9zE
dKv+gRjXsCGsCJr5JF0aNRpdSSYpappnAsXhvaPmQ9kDOQX+Hug+R2BL3j0ZiGlv
tT4atahgV/Y1LUeqJtLOxBH6NTtqFR6LIhmqa4kxGmNWM1gMcHlOiAPkaoW5x2nB
vrnCGh1+v4BBAHErfkXIgmb5umgor/qh+7JTb1Gflph3JAi9B0/SOBzz2XWcDL+T
dxvqKsEdWyVYNhx2pJNplR1KRWIuDNijZnaNODU5RcPU6FwYv0hJS2TvZ30qIJ6f
K8JvQQh7pFacck9qdk5PQ7z5sy6V9ClerVuZ2wDnylGI/++sFI5yWtEWv1BjWemI
D+cW5ZiedUVkZARfPlTkH6vnysdAKthQn6vxA0NOFv7sGdBxetvvue9xTKGFewg9
zG7iKuIZhiSDnzQ5vN6ScVtt/xfw6S8zKT7N6vaBn+akhvQ18ug6G8if4D3Dp+lr
6oMxsOgqtcW8VFHrVlpTKFMYhw9K6lEQy4NgOZLCz6O9y2e22ABBWDyBDlDw79IA
9XbL7Nofr42mP2Re/AMyUsRXn4fU+pnonr8r4qPOyOh/z/rEXDdXG6TSSJe75Hsh
EVMMEQUbAaixhMJnRfXAvsVnemXQV+1j2nMYv31ub8k/+CaIc039hEsEPWPlTjlr
qHZJRvIjNWUjx/BCYm07N4meBhcUMRGPXip0xehwQWz01NmCGBmEtjO5nigHeDGf
+dXC5lfiMgDnX7rGS1pvm17d/Q/XTEjmYo7ZJ3+STQ63ECHjnEiM1Z7Vnx++wTbK
9AdYdACUnHrM1G2tykJYshQtZ4zthkzMoE6/pBW3DKnig5TKj3v1isyOR0r/nKgy
fJUUe0imuo60oL5m7AmJRGcT9paCVZzpa3jDbQ1ozg2MVf9TVB0hiZSQlgT14YyG
Prx3YrQWhMhJouEr9yCdiPH2X4gtb2ZpmgLv+A7yjkssVpdZpSvpsan4Fn5X5H2/
I4JnonUy6nlcxo1pG6PnGWeUY1JewvhJ3cBsLZwidxly7/CNuYVdYGyahSjqrpbK
WcXQJQijHA7PMjXNxhvqY75zyWhR2ANMqX8C5+OQc8yS3x0FrZsKuPJsGza8yWW8
Sy7bD5BHZd7WqjKYL7sbFm0LnGDCGz3BO0nyfNBj4vI3K5+M7aQEkKyPgWcK1lXI
+ixqFVJGI+0ecbJKt2c+cIwekICgEmH0VqEC9wRBRFTjS5SnpZTlS989n4ju7zRd
kN72BkmpqF/+gzIZtX6Vl33gILy/PMgGbKxdgWvHdqBaP+9LXJ9CQWWZXYtjT+PD
3MIFmhMLg/aR/YBSErefq9dTr2+YJm+RMacUkWnYG/6DNV6nDExQqGo8sXb4fXWG
xNVD73r+4aFz73uQ4D+42gIqJ94llBdB9oHXIFnUk2eZskO4kvUUx3+C26es+7yd
zV9loxhl4DMpdcaH1ZOsnZbYIoqYnUGZR57pntyj9E+stj3qPE/nZTkHfnOku/fv
79uO3+sA/PuDTHF1FRt/QtTAxLxH7Vi+OXnM3eJXjs1IZIrPQL3o2BP0OkfbNrjo
x+9Dxlsk4hKlEoe6AtDuU1OL1+WncEg49pA2XrrlHrziDGiF2GOB3qe8IYnGOzj8
0+Ao49WaFycPAiovhmmhN3nwYtovfNTNmt94DBZU61QqR4QVWP7rL79GJ4luX33I
LoI2TV+UA1fqSbAn881OB/TPluejqrf0p9sZHM6b93IuRcOT5Uvx4RIf1wtkQH+e
DubPS282EPCpSUUGmPMcSIMlsZBh1QX48BhxHlcQrTSaE6j6hF1ggYLoNtyZGyXi
rRrLr7nz6xwqzGsgFC63SB4SK7g+jEyxjjyztwJnTzcb7PqdIKstKhn+JfDx/Uwf
Tj/jhZuWiSDFssnvBDryOTPb6HmpheQtMnEaLEH2ys82uiYpJ7qrdQRCy3SAFRLa
qBAEJlu/vpvF2HDO5Bnr2uCoWlCfLUgOmjYgdx7XSZdJLYHDaFd+RJvdya1joSVq
45o9c7C4iC38YMm9TBVBJW+mQA0wYv/q4cfuJT1FuwViPuYGrKdpvURCD+wfFIe1
vJCeB3yzpPp8DuJonL7hmMWUQuQ339YJbAmVHIdwMhbrAFYoUpDsI7mXt5KnIgUd
JXAs6Jrm9W+YBPnZiWt3tKs5yHRbkiWWCXEdRRyY0e6oXMvtd3ebkMdLeNwRoWTq
qnh3W9HgcWo0Pw0Is89ju498lLG5vBv4MVY9Ne8ob+gmNspLeMnyBX70/Do5NRPf
BT9yDutSDU85/tNY38fFc45i+wIpVr2Xp9XE7P4dvQHapk9fcWar2+CSIEc60YGt
CAjsesS/OVtPm9EVLz+IbSbzlld3/vleqi57oShHag82YbkQQDdcHr3kKWoUaNy0
RdBph4qx2jHaMKVXKM+M6eEXnSoDnTQ+z56w+7rJNYaDJ8oOr6avxbu+4mPtRBvM
Vq5eEFRG8Pf7JFUp+zWF5B3hytjOPnnLXk0EQpdeCgLeF1TWXklcjv8J1uGaJvqJ
TYcLkrG0IbQj7AaJxzz/CvEtTWmUeq7Al550Ax5s+s+WGpQNoCsSqYFf+MeGV6ab
byYebCCnzKa8Fzp8Cxqr2BZjDjgP63qXbGMoP41SkjPQfGMr0e8wAlRv8k5v4D8c
hEXv58frJcsrDRqpW6sFkCWXxYM770Fk4xPDcZU8x5EHtv+A38rKWotFJq9jKegC
Bztaf7ux+ShjOW60ShJpYYxaAsEmEmTRw3PcJ5uOHX+nxUs/OOaL9PBSBaeohHYs
eOd0pLCorbJz3X6GM7nlX+dlk0MhnGYhUFLSJOD5MBb7FsLyXgb5YQut+r4qd4HL
s3lBhb0oFy8CWaVf+u2VuA6ZwooAaF80egOyESxxC/zGp3UruDeHU7qDioXYWb1L
jqoizOyc6376Jcr2GJTdXLxMETnvQdsQEJ5ZPYCZc/BmS8iVK8H8FOYdwfkYLVZy
vfXN/6hozhE7rJ1xBP8PZaJZLsgH2/ZuhQTr1JexMdrhXqBduGXKhTObfcWIBY9U
rF7q/vAxFBKICiE0eNc2+kx46+yfumxjVBp9+P6VsgoQzNLpoTls6zbfGIC53w+z
39+Jhr0/OeWKO9UcubHsFLNtwHePzDDnw1S2ytigLI/6nxKymgHEkQOdD8pu0wvt
vmQsPXFg/RjBmK+E8qCEGt0fAWn47p4RlrYYqqvEr6HZyQmrk55POfNINPfnOFTi
d3Z1EjLfBvcoQnVSP8f6ctNiWsgwaGYQe0V20nTk/rtyjnwR3LxyU6JCEaYF2T7Z
wyW/ZfgU4LCKasZETsBO9IkklzCE5J4lQaYRz6p2hPZLMaHwaM+Y04a3q8v/76lC
x9EAA5u6F6K5jMOCrULrWy67PlZWg1zfUvYSZgElGW+/MB8C4hR1ecDbF3fhP6RE
cWxnVT7W+gK84WstrWMXmxSzChcmosVvMm+1n7+6W5hQj0+G8l4pUvrOhW9KpIES
as4J49pqeBOiV/8Ti3gvuUq9YIzno59l2+HvUJqCjfVQiuirBi6cKjACInmW6Jan
X0BaQ9Q1Yp5hMC9BjfBTJWRW9SY4IziHyugpzhd8HFi1/JdT4WrzKRf/Le40md9m
jaecqGQ8xNsDJf9NQsU8zz8manUqW0TasoTffJr4dctwx9nvUuNiwz2/sSCbTnIE
dup3NSHPqditQghsfhsHDmBKsCFdQ/1MY3H32tFQ0MvVGj9VDibPYW7bbkrCIAge
R1qOd2rMRrKhUgW1F3K6Vobb0KWjNQ5phk6WLMuFscMA9LDCeR3k3kjHbqlJxEO3
t2AyKnG9XvmODKiQHxCTP0PcN+iNH8ECNRFHC7qxspze4aEYbA2d1AmEWFJdhHYR
SVJfprOba11tx6UjRy1jSVa17dVH7vRmBkFeBEiaSocbTuWZVUBm8atGZjL1p6j9
paugQr1mBtjiICERe3WXeN2B4FYg3QL9DG4mh0Z7WtSLWGZHRkJRC/KE0EmHYc/r
+w3C8T03tnMyW2h2lMo3QhsFMxYHygocQJuMuILu3Mfsy/mYYK4esi5j5gM1yURA
zNyGqK6PvG+nsmOUHZiuy9Gzd8ZGUSmtx4zfBIY4iIL72UttumLPRaMSiTP+0hnL
YDzIkj5C9Z3X3hoDnhwFhx/W4dU+PNM/GVRwxUgqn12OH7rOOdz0dsbnp9tfdyGm
TJpa9brUpJieHTPzI8Bnq5xZk8fHxSEYOiMdVTieKUia+YyvPsACkKRVlmBoeEgC
sGsad62ClI4IEzKxBG8MPt2htN++gMKhGlRO9hSCW2miKOZSDaC0DsfdDDgvz846
J3QGBhxZhtw0Q/AtjTyiB4Pib57bjK3pd1yzvi2nNmZqai2K8I+gcoSMckovt66L
Be8eDb9RlUEhk2GN4PUBlhEbnaEwQYTuHpiOczVo7wtfGRWKBonYc18o9YqJanUi
S25EyFs9jGj6VXc+nS25FwAR39LRWuHxnNCfyCsYWL5yjkqRUHXlxog98tbe3Yj2
+WZtCcq5pegzZsJZdkQg+9BEMYvbYGWkDJ700MRIi4ZqoPudBc1KJiZ0s3LZm5dj
Szng6cDeBD5sO84gWLGgyhE5ABa33/TQo09H35UowehP7lpnjiIHNalZSykV56Sy
on0tgZ7mV9bpwhp5aVUCNLpU/a3BtUJJHXe2229ikkMKjnvfbwKkKf5LkCxTU2GK
RaWW4nwjI6ts8693qOLXxWRIFUHv4z8kuTxytdncAU2UW3C2cL3ptAx5CGHC1EdC
qfIxWssRl8RNA310OV0/FqjaovCnUF0Wwqm5J1O8TSoWKuMZMEW+NhwT1bvIIoap
klyzJlaL+a2OH1D1jhiRmrlB1ICtl54WsjFCtu4njoEPvbbsWtnktZfFJgVHJgnK
MyGwD1EUTfn6CRj86IV1A+adyiQoE73wJhuZQYtThEnSAQnmWhE51dq43N9XGIEI
jZGw+TWT/agEaFRDaVr/aXppv26fzaoB+cLSNfjbBOdZUDRNHsUirTztuf0HJYGp
7g4xc9XNqcXy0hde+ygLX/a+3GxJXWxGqEH6JUD18OCzFlZ9wnauK3pEyx8vUtJM
HOUkwYUIcTcGkHCBXuUFd+k/jxvjqGDeoXTWnXzvO90drkqM9EzFhdAVowzWmWJ6
23t2FT1wD+Fxw56xY1lYU0qwTJ7dh7FRDEd4NR3l2OyyeivcS0nWryX5F4gqL2l1
MUQyxTCMN2lBj+m107tG7Q8kL15pXHqpDBLD+zLCMjMZshwAN4vS2jbtMYh4qNxN
kkfql1Ean85wbOEfGPBnQnL6+uyb1PZXJ44H98boKC/T1QyPKzz6CQrkfJ4eNEIV
Jv+IE92XCznaIs+lkuMwLrNSKNGvOlSXikm8QhzzizzD4hcFswuI1yTI8u+2yXx8
Ns67TLbdBLoHG0Jvhnk0sC8nM2PHBpvIXBEOIEtw/KCEfktlwmghOr+r49dxJh4b
7fuJR8/xfXUTVPqyVJk1v27E42qFWb68erCzQ1AYLPa4IveuS7CawG4Qm9A30EaA
LHDffLnKtbTKYN8lsDsanIBFxsvrb/Y+HO7zNTGpcT1QbT+7XBU9KNoYL07Rayge
7Pt1Y4vMPI+yp0B4yBuOOJzlrbsqaeuUxmRL+n8apRiOwF1llThmEov1XLF3QMBC
vhAThjU14mYIDi4KlqdZJkzi19WoTDPDKk5IUoG2CyGLestVLJcUtKn/R2RPBA/h
x8J9J+1Ip1thnbgIfY3FakiMWBvO0NI7wQLyrUILZGZcl20NC9shKrlaY9ktKs9t
uaIRMOE6iymNItZd8xmbp0v9L9yj2ywZ9OwGnWxW3UZrLDDYiwwkhLKSZC+F8/Xb
HW9IgBrfGz0WUWbiPlWPIVFHKYWH4JDeFlljKrNHdaSzgLTijEXkL+Mt5uE61JY5
mXybexGcJv5I/QXgttU5J66E0zAVAaplcfWiyessBmxGA2r7pRbNfB6+dvlyaJWc
ScilOXv9UVAIjrYwvuXM4VCmKpRmOHM+7mfD4tx2N9I/4/f2/TXjyL5lhlfJ6GbV
GEY1de+f0hZHNlj0eOMB4ZoQhDBx02uCnuxwV8WSSdu26Y9GBZXKEBnDil+1j8RM
Lo5vLSTyrnzzFG2jj0AdZ7vvhlm+pvBKufPZbqnM7cryUwUX0fXHVVqNrRdBvc9k
JMecPR1bCvHoSgUlVhNMNmNKno4zzkde7TjjfyWDTnUvD+6mhD78IgKeJU10nEqc
Pg1vJBqegA90XijIs19DDWjosSQjc2PHOuhOE5byFBrniWiGCR3liEfXJnUcIVGq
XlUU+2FC0OtwpoSyBdtkL2NB8HEqAFjY81Ulxb1nsikdBd4aG25LlByn4z24ujSr
QTE+ZORGw9uAkY6yVmbyP6RsUNe4FtaOOGw7abXmFg0fsVaO1nCswiO/NNvIoPJD
YzVykzNrEWT3X5dA0fZ85wEdsZnKDYVs5Coukp50pJD9cOgYFZKmYrCgsTOznQxH
c+gsqh71DaRbVvvVK44QP8QzZnUDwxcLdyqf7fLttlBVOBqp4p6DyjH9D0prAil0
98di4O8Ac2duyB+PJ4BMiKpa5SBENsJdWEjuUXKo2TWL0bmYpBIJ79x1Sl4EbOgU
D6hYA0vlWxVZs4Z5DFeV2WYpH3pQJYUME3NRA4V3gZQgSuhjlaoYjK8pL8VZygp+
Bzds+gb4DtZFfp9XjFTzUJLS5+E9JXG+aZDsEV4sZi0E4gmZ1+oO8oT4M8OQo3wp
mr3cz7bvcpwJ8371dFeFslzuWlaXyMqCJXfA6k/ReSWOKRYOzcuujGEixo5dAkyM
VvqUP7ySImcBtO+7SyzBaBwyCEOwTKDrEdLOT+pyzB/aL9vIFTiuipKSdIg2Yrpa
/pZmXwM4nYZ8NvO/upeRt3Y6Q7gtdfteRmOr4jyh/zd+zFTd8+B5uqacuMVZQZIy
DtgXWsYpaEZhz5lwrUBTB+dEFxt5KORY3WYBml4g1+91Ic2ij0Gqn2ci2nXa5Guh
/jd//MYSxyUJ2KXdL6/n2LDNXlw+Z8drUBcghOEcgchL6cR4D/VgXvUVW8k2UJ9W
FjtyECeQ4gLJgmlJCwrZFBBTxjNIagSHacrDtIt4x/WhgYrVS2ZpPzn9LNzhKj5p
hS8dKxEY7TskWBVNTLP11HJYxiSBDmO+Q1UY3nY5Hipands7LdsNSxjEn1w+vpgM
jRxqmYUoKd5apBMidc2B4AN6D+fqcpxo7vTCxxxtfxRkreRw8X5OXQPhFgDRbiLz
yYJjZOqpasdjJo4EaDU+MB2s+ZPPLQTMKZSmyf4AjP+tKwOkFLn+S3WcS+8717U/
LolJGB/ykCGz7Xfb07QEaE3m/nnIOdzbB5Xl9NpialLYE/7vquDteOe33hrAJtvo
2AleqDwbAZ3BcfHWa1dprghcFm3RQ7ZpNTxKCnkKwXkuwQ3JFKDbMpbnbCeoSJ8M
JEjVu0nMd8HBW0aYUdJ8PN7aM0GHrGdEsy69scQ9hIN1jLkXGYX2xLjFP8zW4NMn
nsLRiT5YrF8Sc7MQPVXepFXV6DborRR6WAKmyepk0OD5SULl5pe0Nt2Q3ol7vQPx
0BEvS/wNjAHKY8TgLoXioP1wRMtFFE5YlGp9LjiYPaDkWG8ODAZZWCGdoCsT/9zh
E4LWTrZlD3Z4oDratBgJ4YlnNqcpJQEFIa4+pCGHwPzaSAEbrfpsJPoz4eT/Rdkh
EI+DBOSMuO/IhEjo+9YA80pWoOry1ccrY77D76Ua4z/tk2v1pb7LQgPZzRMMDrHh
2xz0r77azTBoQ78EhqvJJG7NwLQVhOgJIhYG1pvVDz411S/NDzRyFKqtwA4jjXgz
C/vOys0D98B82HwiHDTWIf+rsS4/DJ2Ib0hQa/vW3DF3J0j2kK8SPeheybPC7+Xu
q9HW1fP3Y1T39X86N1FYwsGOHLCcjAdw+FCbZuC3zJdAQFn0Cy91g1dOlxwCHajI
/pZLB7Ewkm0CdSdUMR0dFikK6+KHxtG5iVRnHpctBdOOpd/yNnzJk2pI6ade50wI
RW/3+AbySSzcjnIWPF0bMIDaSUz7ead9iUMBBbkGc2VA7psfRVogmQTIwkRzr//H
0eZHpv8+6hhFiDfOQTju/w0qocJMSUuZYUCy0wRVveQIyNp/KtR8wNGLQD1jQG8f
e9RGy5xTIYkw/b+EEBLFD+1EHb/K8p8SgZc/ToZZ06KH746qsOIcpNcntlPrCJmZ
RiP3iWpLjkGBowyIQ0W5pLsy00OiLLaLnXtNNhpxy31BiDYMavXEw9qEZudhFmJW
abInn9cE+bSeiQ42fRCTn+Oy6AJdwE6hcbyoxwtsUDd4VmkcfzgscMg1LSL2/4jh
eUHNP/Zm5d9MSkmgpQmhJANMCH9eQvoGM7hCIk8x81PVNOck8ThPGHI2wA1N0pY2
YK3TU1AQEDn8sr4Pu6MTMyIK12EeU56SM0vp0hsmWMgrBysR2ud2T2KvXdhLTHSp
TjMq2cxtGdam5dSrBmODcDtpaRf+kf6IN+JzbBLXlOWyxLKFvTZR5Xp6iL1QOY4J
mv+KWCh0bO+DQeJUtaN7qxfWO6W4qyOs8rU/DHycuOidV6sI8QgxJnxAbCDJnxRm
uYlHsPyfGgs19wO86/lrCpPNulfVwMznnetT6Dc1SBAlcOcZZdriwd9ZfhjugwOC
+wPSjxm5Zzy//5ou7zEzjgMK8/hc/W7AL6Pq3EyodJz4QT2tSjAfoZbRl+hinIf8
qzzldZRJR7moHNFeTZMVBcb2Vtov/Rez3KIveFNzKhD5tpdBabjAEOMFheHCvYwK
7Yr3sRrDV9mpGw0uUnhdMYGF50ed9lydzWI47Kus3G3A1SMzZ9ZC2klSb2FHUZKo
yw3YOIqHJhuKqk0MhzGIeRFATzZWDg0qNEVsNy0q9qP7du/0Z9VNFf0jS/t2kRKi
qxL7noh60Po+6OTpJqDp+DSZQfBg/jUwLd0vbEP3dXsNeoqT/9t8YMBYnRVu7gF9
1BMewn3IYE16FM3q1MAjLmjuiBiK+HXNFqbUZdl9mGpJ8AHrl525c+OMdOwrCD2s
aN+EiBU2CQLCl7pmDmwPN6QfMN6ahzxvQ4Ke5sS/f9B0jIpgo/1SMs5uh0s4dVZ9
nLA4HFDU3du5VqjRSOGVeWmAglgMTr1OloNhJjJaMgHTrJVM9mo6a5IkplCI2B2D
j86WmlWMAs4CGbQzxxYUaOgnm+nv2CP8ksb6+ac1p3C0pPq3lBxyfI8rtUfR6UYO
AOdIteJEQYRJbA71nAyOp2DFDHShZuSP9hw79RWY1kU3BSfhoFQWo5q5hEw1Jrcm
SfEV0MaFlz4eintiQFM20+dn5fpSa2yE2F0s5upMDOwhnAmg4F2LFy6G00W6UuHC
IwrPwI1HQA6dULWMwG9Ch5m4K/TP3UXWnDwQ7yKj7Yssdd3rEkW/gzX5cvvgBADt
WGLxbpKrO/F1mmeqf3vs6dnjYXVd1oC9GeL2q8NxkF98D902SnuGghuJ0zeQ+6vy
HIGrHXy5RtgWqZvoeyi/t7hzZAtqqX0kP5yLlzpkgDlgqNLpoN8eVarFKa2e6h94
AGnvtylO2+b5khraIyLdeSXUEwQ+ZFCF6Panw1P0Q+s/qaN1tkUY8QmTcxlXSSww
jZQw3ASjsW+DmyrxXk9GZgwDZg2DotsOF+GXIxIQo6OmD/3Ak9SbuA3CmE25xk6Y
3NioflmArdvgpjqb/FC/0dKvqUPsLoNs3Dau7CLa+Volr8RBZwID5kgJ3H9MOkfJ
CseHcQiPyCUNIdGzQnhSsZ0rLjIgM0475IRruo2PkHWkd0P1VGK2UwrCPzKNUwTv
YYdSeMnFLSgK4sT9pOpjCrYERe9rwCTk7LYUzim3W/wBDJC/+GaqvsIjBUARxKtA
SXYVhKYVF80UAXbimdn3JYYwDBhntGFuQ7teQqzAZYs0zI9T5VL+iimT6Wpxy664
ttvcIdOEPJVO4J2y/Ai8xoiFkNnjIKS6p+yDer6bS045gsdW9NJeJEUwcBoGbVCk
6yg7M8AG25GaaZnH+yxnZoFWKLm5jznVxaLWk67wgXDSzSKd1WlzpdBVKZ0VKRIh
fKUJC+WWhXfaaKPEZZVT0Qc93BEopvstlvinjm2t2CM/NNKXZGs3SSpKPaGJM/3b
4suJIGM5PLMuJIwk9+n/emFQHDxHmCNmw/1kSsNIWHScI2CWxMV0QunXO65CXmG+
SIShQBNSkB0oLddkEfxEPBAEHdFeczc+dbuDfOkBDMuZch427n8bawam8JBV2ga4
47EzX5tlGMj+6zmo3FktwcG8Y1L+043WrLB/I2UAuFznB+D5Kxr8epZd3cLtI1Sd
UzY8TYHTgQKD2CkxU/ubaM0qWSCj1NPyR4fIWI7I6VhKEVbTjZ39YNmxy4MILt/D
4kkto3ENFXrynyJ3N5JHZGxI52uquUWFkwSanRCF9ybh8h11clnKkaYN65AEVvLc
gf3Oc9KTqKtDzvCZukm8AqYl1Po9mFwo6jGgsZ43l7eTs6sa05kqPVcOWmnD0lk8
L+OBq4yy81vA7mQE7Ee4pQ8wpRg72kCUXdFka3J1E8dO2fLco3njy72RZaP0UO3e
U7pdzLYynJ0lco8Rzu52LOPUtvcK7H39SvjiTuvkv3yogfp0YIOvbgCfZNECI/Kx
B+ARm38qw5XG/Oehk/XWXdR4N0UUL+fZg7rB6vnRBWCBJSGNE8ZCEjyzomlKimtU
xFK5I/FhyuU5t/Y37pew9e5gu6fMRbPrX0OLiYynLmZOMyw58MseT73DMrh6lGwp
T9IO2XgY9nueuL5MtmjArxnlBFUXi3sUAX1hdSZGppJidQ4XTX8RQmLsqicI1lne
rE+wa58h9dQaXTlZ33Yaq5SBfZnx6BPktdy2HEa2W4LbX+P84UI2pVqdHsIQvzn1
iG98dxilGJcjlCYno0kMACVwpDw0o51X17aLjsWqtZqGauQsViCps9p4X4JkV4Ep
Fgv8Yut7OeWdV2xWzmJrSWexuOh4y1XvTYmJqljPLzD7aXMcERRRJ+XZlM8QI4qI
SfVQnmBtqnc0X8UZZOH9jDlDF++lnMdvcOEEcmIjhAT2urwa98BPbpVrl7i8YquL
tgq1kukZ54wf+Q4NggeoceNw845iv/ysO9TrNU3eKwcLQ2GBVXfYWTDOSzmWTTXY
nMqg8weHhLS579RwdD3pi4P+aGhfesesYipw7AHxsf+Gpb6tbsGBTp6pYt+SK2Ei
0qABeMsxK+EgrfekLWbwOXNoXEvsdSU7xAleNWZQdqhH07Ag2Q7H3vghGcLSpiN7
QKQ3hg0Szj7TkWHhXJ7ceoar2O0OxEL5iLFEVvqvmUdyIpdAklpL6+n92bjbrqUF
CT8PQRMkDMgyQ7RRaNtW4S3wHtPNqfUz5++O0oVycHVFQIn83yjqbyCWXfcB1Y3T
Qzs5ni82XkQx7WRYtl1y9GwfsN2/Z6LLP6pRygJBXgyPlOB8SWym4ddgQG3C0n4z
tXMcja5dTbMbM96nX4lAwXv36uCt9FGqKYCJKpV929IvEt+xeYOL/1ZCJjz2kA3b
zSvYYdei0YB6kM+WW7T7QbKaSYTymNl8EcIWK5kYKnNsbKt3PO/zzl8qkcTjpDvd
f4SQy40a/8/JEAIhPt4puL9TR65we+YQCKnavNhH6x32hKyNeXy+G+Cffp0gR2mV
bB249gmd+ig8LLitP4xFBqjMvTUpt9kDuo8z3qyn18//FdRjOk38u9ZpaLyguDdi
li8JW4dsXsaUk1dVUUlhbQI+JgdfX5LkOyxFcgQNxD4CHUNcQ59KZrRIffuurIig
2XpOURFxNUjW4GKCbwzlkbUyYZaXGlylWkDM9CbbjAHJLKaZ3XAWXAsXR5od9YLo
E6mH0DbI7G/KV1WNBhGggicNNVO7Xej66agDb7dB1HkilG561MSB8mfyu3baTnpq
4HohXRRvzzGMWiqO6+ih8w6o0GY5+tYSSdGEzZxr3bwj8bJwZpCqRUcS9datPrMc
icWI/CKxHhVk4wX5Zcqo2l9gaGzXZzkETcjO9fgFXeXmCXi1r7Ymdp0zv+yluxzb
U+qrf9GnWsz2hSrFG+lKGgDNBGaKM5JcQi3QJNSeS/ylOVTOQ4aaaIxkI1ErDxDr
MIgqkt2M1FdtGhXjh2qee07fsO2IE2LnLxwjrRed6xz8wM/TVRoGzdMivL2MmpEq
0PKZ1lYc+gBzFw8X0MRy4PivqhORQkUHiJczaFlbKrxqN2V5I9OTOfBJwi6XTtsS
cbXUblN19jotJTK9KMRTW48wmbOuJrCvzq4cS8eK/cXV7eqTBVg1KHD72FEwZmjT
9zfASQ264zDnDDa/W7Y4USXOjCWB/oi30QVKAElzu0nBr59u/EpYjFHgnh5WxDOC
tRvS/nYQEsa0brmhEXaXh/1py+XdZ2yVoI+Y9FJ+SCvaDrR5LtaHGRZeBuTC0VTM
6UHp9PPXIrF2RuJB8MH3Dl+GrZZGvUAosQEgPPfGEB+3S4ldS+UtWnuhVeGS7dwB
LEDG5ApZSvglzT7l/6Cki7kaG6kNZFOMmg0EhcEWDDZSUHIfk5D9WZR9VypSbtrf
QgF7LX3TgKXsOxrfT6e8fJvZg5Xy3nMQes5Aa3+7GZCKDEOOUJ7Eje1RgR9I/Eqa
hiqVSdukgBEvXVo0QhbUhWoWDIqXGv8kz1ld8rYWrfh2m2Uow0aVUcSuGtVRrc7w
Ak25numvSvedjIw/GHvyLyT++qC2ZEFrkKCAtn9/2nGDDcwBdnlHtwEcIijatJhV
/2Xb81FBJArse5i2hQI14IUupAw2kRmyKu72rN8jB9Q+nCkwEO/hR/jSJAuEF/7C
e7aRvDYOtSymq4WXRr/Kx+Wsbu7WkGu6QmLCdY79AiqtB8xz6NfYHrQuUm1z23Y7
1mzcafIJ38Hs1t5eo4NBaVn14318lUHkYU7FoaySUQs/M036vagQaX9Jn9QjTFm0
6XH3Hat8RHazUACS+TbyM4UZ/PnaLMhVMo4paeT8+3qBgW3vKMBI79gLjvmNqPye
5khxPeyuibjghYYMYQwQclE1PQROCHecf4w76JjxqFJr3EFE6+Gf5GKUUAFR8pty
XBb4JwuJaiqVgfz0ADZSxTm+zNBWx68nICHzRVeVEgnx2MWKyWsPH4y4qELBRhTA
QIwNjycahzoJGYsdylRgxkED2SkJzAJFeyhYgg/J8V2xQTYO+XT0q0BStsdpzPWw
JBVqRYo5cDQEl6xXrjF1UDtGb/s4QlniHnWBly4DKPjDMC5Yn2F0Y7eSn8ipHqPv
dvK+y7T9r2HdxgXf1sC52ePE09FP09dlvMl5qyaPAs3K8fQBjZkiLfFShVocC5n5
C7HP2pMBqxL2Y7SDx37FLdC9PzU8H/1SrgilusY2b2iWoZp0ZNhbt3upJeKT4Mh1
rAVMsTGJszt45nbO3H4VRMyz7l8CMHt0/L9rvmOlZ/46ZVnQRdlqAdnWGTYF4aZp
Dq110ptBzWfW3vi6XEmdEvrQmVELCuKEuIc0T/JyyJYLHsKhvkkeTqcgvx74f1ry
jw321hBbgEZ123dXPcCGolL4WE+zjh4l29GGzLNv/BOYW4t7rtjuKKrvTiYrUeqw
g4aRRQt+YGWCmeCzbXl5ULgQIgdRTg3oat91FGIYove2OjJWhbsBUHT7TaF1Aqes
x5v+auGTwILB0HQ1xHCxEcOMx2xKG/3Lrk6AWj6NRr9VDgV2PrhrdDLLodYSs/Da
wHhJJPLCkdEXQFm1OZ3AVz9M+XBG85KP+UuvXNyljomHHhWlr+5UoSihAwe5Tkgn
JlQSVaSOI0GA5LRQZfiSE1rDiMBbhyxzueOVF4kRznwUDwQVDpuhoLET/uqHtwqI
5cu53Xb+Q++EO64VVb6DrOLV9OQ1gxhuLgXjMcXg2tAYXHKLg0V9sUOg74r1Y08i
j4nRrOUz+YCLAMdWt0QWTe6HU3OJNwao+/I5++Z9NikSVURL2+BZLTXuucZ3eIyX
CShy/ne+O0rft8GLXnBY+g6gIX7sjdpaU8e6wyEGH3CZBxVWPVkP4XVavi2SA2QJ
QFtR1xLuS3gPnp3Ag6dMsLRoVgLNcfjffWh2Jibu/hRtw+AiTLNDtKAd+9Wx0w6H
vN6zhbvOnYS7xV0ZWT3+aykaULLmaG6z2k3A0j6dnD8xWH+aslkPP71jwkrbpUjh
K6fzObpw/gU7PdnPqFyi61TLWahzVSO38WvQtnotyxI64RrjUhyh/wjjQc56foH+
GlFa3gIHcFShfvBYtaJPd5GnZbG5QbpNTSNjc0EtikIiyJ7iZpPuo5w5gVvmd7Kx
jDCD6Vpbybq86O8Sm30598H8Mb+Rl+mY10NaNT18mjnp9QTQafAe+QPuNnD+zE5b
PffmUbpnUZejHIzMQ3XpXgNQ/9/sogFUfSAQoHNPYRvLydkfTc/WKWfjIGhgncyj
v1cUMnUgNhUvF9u4UBTkSSPtll+LCG88E5D/wPRac1ueNHqGZ0hF+BpZ1/A9DKuv
e3G86vlUHTqMwaY87ickMq7+rx/Hu/pwFfbtXzVyGEv7U6a1tEPEr1qXOsn7uyuB
0FEfL5LJ9kQ0+joZLgjFBPvA2vwJx8GmSGmbd/71l0wKTH5jEbhtpGYBYE1CXamd
FpEQej5qyurvtzbMte3LefLDD02YYvQAUi4ETFUcn5MfEJRGttYe7FGLX1QjwF3q
rswtrvmZt0/L1NLZqSaH/jjDHFKBzPPpybcLFbZapHmMVAFOPJSi9dIiGqj0PWAh
bsx35Pp3QcZ2LEG3Ng6+tw1kOiqYYPDr5YPI8jiK3r+tuyhh9jWmJbZ/9RUb1jH8
Z+LUTwA8ZAYfbCVQqRyzvWBVnFPMyRvotkI29d9eIl2BwH4gJ637Ld5LETCO9hvL
9UEYq3wXCFtEU/RL4A3hZC71uRFeR/MYkUwJZFmG29DUwY3tFXkWxvY3u5ujL179
oH3hRQ1xwPRMf7ZYIwV1egWOk8O0Auw/UAv7NHZJw7aHy0LVloms12ZhyPtOhyl/
LxDLCrUIBBBJ+4Ij8OqY6HSFV+wZ5OJSdTstcuUR9Q76UfTfhAiHsZbnpR9OAy1A
jsnI/uSvYDY3r0cUqKWj5cg2OkXt8TAQq0Tv4LEmp4e3GeEC6cpp/VDaqzimL8e9
7G3FhDN0XO7ztuowEpj7/xckogfELBNgqnnzs36w32fTf2gsHz36KSKuJYkIUS89
H2J2AduiKaN22bDeyEwSVrWbTrJhO6lcPO+5ansJrtb44eIsRC4YaF0cedSSrUyw
hU9nyA07Sgt0amlHYfPdpJe+zbgAYn9QWyFHf1DeHOr/o2WV3nusN1gOHVyxucRZ
zJPfd4adew5tyPSmgD7rMGK92Q8IB3pLbqFk9nyb8jS8MvfH8OpUjYJwcF1G5DOd
gLWw4EmEUfVbmhZxNoa7+denl9L+fFQ7QPCEAcWw0h4EhDamLNTa4Smq1iw2PdQM
WizeBBtQ6r3Cbpbk0ICubWnAwMQSg+kc+Gk5w9efPZdIE4SeOsGwT422Aou1bwlx
hf1FOuhpk52QMeOnb0ZGKOpUk/l2kfJH+fJryqaAAKjrOb6tYDfd0cnYgjrDlXpz
FS9HjCQ5L5dtOrBUcZoPdbx0LFkLvMo3DXDZJuXLMOfuyTvzdN9z5u2ldSytZVBN
hRaGStC872sn22keuQHOQfb7ApXGMSL+wPBaISXfI3bhLuiBO/n83WRBR6BLg+tr
Y/1pfaYGU19URWhGFTKQTUL4t+oKajMx6yrK6kKK/frAMpaNrSD3cd3ccTc6h7Te
WGeL0BgwIB8w6w9ohcbkrosXGVd33QO1NQxbdskPR7SPkDVzvmCV4fncBGCmokjv
ulL+yIV6rn6ut06+haL/Bju/ApX5MT0MekXZi7spTeACOPs+lwN5iRN3g92Ofvpk
opyWo5oXyB0IQSMV/nKBhfctwes+ytdGg9sqaXtiLRPxViSJ7WqZAPZYEI9c9gMO
mMaBjGQbbUKwRqj3Ux/bN5G+jCQwtH82ApkcbWlcD+h7cDlju+XHVIT/0e2zVroX
q+JAJrC/2yPlbAhyyQo4r90se6/bLFlLap1pz6+6oe0OlXLT2QcLcJRhCkzLIxEN
L/Nex0veqKpb//Ebc20kGN/Je7pBxk81Mryu/Gn6EPiupIw30xz214oeg38xiF3N
GR1Q3JqHzerXVldJkLO0K4GxxAHgdzbhweiv+XMW/PmMRrigeGhqp+w+Of1gAx+Q
ube4+fCORM4S3YohHqC09Ak3CTVQGMG6s0/H978+SWITWLENlRwYbL3nA7WnU2lf
rJyIYN93KvO7NmO0+K7GgEWO0JJQWmsu/K0HFoPxF5TigRAIsJEyaXQvJz9m0/ms
YTDflJf8Jz+n/2S34e3lh+1PR2UcUxoYtHyzUG9ch83xX9/NtbO6rv7IIdTgmRKN
b0o2tS8hzDoE7jTue9Tb0WEvD3COgX5JPNs2bMcKcg3pufWZfIBJKdyANXVVkWvr
0MbdNABJiT6x4UQvICes/mn+WYHPTXsA3abdHkKf7GiCNOjpdw6nHSZMVTzjvowp
mNolCoRoUixiHsVmwzGxnOC4VbcDUC6M0GkKKnlUSU7JlY+83tOvphNT/QyhZMWe
PihSmE/77F9QGX6Bio9yb1iYOCQ3SUJ3tWgCpefVM3jg4MrPekHMpyejHvPs++pl
H/TnxR/TlMgZISWQxJz6imHCGD3lrvQlkirCX8PRD8tjW7+Sq7k163x0J+rDZmKm
dczMP8LGD570e6aaxrTlnVC8QuuSO1Aj5jYim1hVvKAcJx1f6kTLfckP6Tl1jQuK
lU6CseIuloOCuVFJTweZ0bvBH3Rzb/YSGfVNH3ZZxpR6rVBV5212u7Pqu4fx8fQr
gB1J52HcTxEagvOb8pX7WqDDdQXb5eqvpKy05J5PImOtphs+zECatwzhsT7vweFa
a3Qu03TOjIGgQtQNF8f8T+LTpvw0Kx3bxGCmMs9QmhBA9MYOq0eDPzKJhts42Nnc
8/s7It19P/q2202IudZqNQIHBu61wdUgtdi0Ry9ccc272PDaD8AFcnjdZGrG3ACy
7jN9bJbynRPO5fW8DPIBfeYbl2+Ayk+NKvCiU+r7z5HmOLdAEqyHyWVCy85KUhjU
Vkt2KUxygRpxBRbVS/0P5Hw5gQahg/cYwvXMdic/v+TQKADt04dTXzn+EH/G2KdQ
GHIWc7X++KJVRuvBcAVPIGHHC9vd8t/0msT68LYHjfdfvYj/d3cu91azN28cuvIs
d3BGWhy83Ko4Z5RTW27NwVmz3ltteYF6+EYiBAg0esgCU6uL/XB90r4Kijs4ujeS
hUGU7DQ3wwfEa7txSr53wxfWFF3ak8vv47O8t8hc4YHfkbig4qy4gytuoMbBNCo4
drA27ARQxrYeVx7PvtToJgDSTt38oacsAgflAWzo1IZOjk66hMybcZBmGHrGNCMk
CEyOXsJ9HgOCM/QLp+g/160RmbwGrApsGdJXZlCj7d3LpTW9CO/5JLsyb7aSETgz
rGLgiEsTC2z1qPzi3E+4y/K7WsSSH6dkD46wF731XTkVPU2I2GoSHo4zRPSP5JOC
EBPRsnBkFoPh4btbROwP3dH6l4SYBC/6dtJGC1sZK0GC1L4FifKKIwBOEDKIHOgf
QWINzSccLhOoNVpfA327pGCEkQdvZ4EuvqvDhy3tco6XEMG+pLnATcLILtbEjGDa
7aEkQ7VWEwyxsujXBdqbonqm9yhrJO62t4YJcgmgwKzxpvaabLU8WGfSDCOZRd2J
cRRFTNkJ3II9g+9PaXB7MdZjuTrbEo4aSdq+rW48v7u7Jy2HH+vTMyaHqvo/KiYD
DVZRPumI2DcB0bsaAY/UzZIiWrxUfvUN6lIyzwEIi1gYeLTFOknkzBzpawwOcXKt
IAViQSyLMBNzcrudWAPvy7fZC1TOG9Cinib8WuSJpxWDl++QJ+B/hn8WWztY2ZHm
2qZDxZq9b7pySghv0Sb8lS2DNydV6r2/5mwwvs64hK4LbzA1NwTFlMEbgjagyyQP
34nKJXjlhgtUtNDmMxCdGd1Dl17CRl+rcCLaVeL2Dyl6vbTBfMQ5o51xa6nIMNBa
U/JotNQHed2s4trp8d9dNIbWMqn+m5d7/JipJZCsDMmmIJdFhBrtEbKLMYagJAYK
/E+U+Dza5EsvBsRyn6Vt3ei0DVZBjUhcwIW7WX4axKzhGH6NjMUDzPqWS91MXNk1
cmuqBl8q8f/LRIGapz2R9QVcnIFFiaOtG+VhfChS2+DQu+wW1Pwa9XFQVN/vMsBK
GRm5l6WOcY4tQG9tbmrXVrdh0QE9WN5jF9PdaFqTHsfNsVQzc+Fr6xNRVFGBByB3
r7MyUk4i6ntWIqAOa27Dey9gq61o5sfxnTCEctPGRTIkTh7is2OxA457J3vdXxLH
ZaoJAfZ2Ab3VgvLiyUSLC57Bb2dAdUGH020xvjP8fNLuJwxyjrYhidWoOP8pyt9U
jQ4Jdbcusqw86BuBXtbIBJLyTzc4PK9xfmiqiYudlXe8SbLNEumU/mA2r80tca6Z
vNh2DMwYFAVgBQ1t48BZufrB4izBdYJoV+vwuvbybkU7R6YjvU+Ow3+RuqPTdudT
k7bsBOYerzptwfLWkEjNmHyYguM4oX/GqorJ8laGdplrE1oyg75guP4T6NEAybsh
bmsIwfEgvATSF+wU+GBj0Bq9cYeVzZdnpK6aaoNVfyd1AtKUeU5AWkFF/Z1WYzan
UldnMmj58g+sJilAuuy1IIxJbn9E3An6YUDdz9SdJSkXlcZ9eOmzfxfMbxShYWqu
D8gXuqCn9j/8llAdzHeRTsAYw2KAQy60NVPkeJW2Mn+1TTm+Ha3PSoTohEC99i35
q6ZE+CN3HkWzBCJ70SLKQwT3hjun3NAYsQ/VIF6goLp7KEsT5zSRKDQT57pN856M
sSDof3RH6KHrD1FLf2zBxOEp6cOalvBVhtlv5nff0FrJHlYknI3sNipR8/Xql8ro
7NecJ5U0Zu1BAJxzTca+YOlzbQdGgowLcIKLHFbpOoygpoxPGlSrug4+NQbpRjJT
4AqGnMpGLsX2csv+2Zb6pzJMD2Wtv7KUvS1+WKzIO+lQBTnikZdzs9RU3J47JQzk
GbBqzpj6UMcOiSXB0nWJWq59tdpbAcpob2B5582KLORGhrcnZ1FIm2KYJFLSZ+69
X1A4KWc6RFQbiGrk6Ydbi8Bw6zMSCShNh5jTKDkw7iiXCooQa3mbLcfe2661gPuE
Mo+vusEM/mCU2DAsWuzbZ/7sIcWOrxETB5f3fJJBEZzFgbXzUObzfglSL4W+9zt1
YDosMsGFn4W50a8w3kPyqQ2pnGSNRNXnpkbi7+SValXb4EnceuTPzpLZ95JB5BVC
KGJ9Hni4BSuTzuBmc8BVGa6ydgZMcoxrbArln1g3V/4HQFosC1aoFR3w+3KeOQtZ
qWXQCqgaXF6nsq0S740eXZrQJ+WL5npdtzKI3T1v228UTxhJ2w2FTRHw4nzxgLCO
sjHFTGbOvUVNvQKZ4ag5gP1L3/p0IOFeVqGjUXrheSBosWodZbSBk3Js3Q1IosDW
kA9yytOImTm4AFLe13YG5M4yYVQLazHOvoogunZ7bhuf11EQNLH8ftzS5G0T+tsn
W37U7Vd5+zXJVm2ZFRgnsdXk+vnHdbf44gTwF7jMt9iGmjRrrpZRdKrN6eEd1fmg
VMb68QIeats23ZDbPDgqsvlFmKvwYy25FV8xoXs6lIuKcdEe4bTWpY/gLf36Nhcu
+kB2B1+mmadoSlnF8c25puMXPEj27ZMcELvh0QoQpLiIbsKZSjs1XxSVEtyaUbJE
KY/9feaSTzIO6rJETe2+pk0ok87y4IA2uLMja9rRwdIzzxqLi1XC0TngBOWuSR9J
cig1AMYJxqc0t85Hghwsuf4DI+t4rvsi6GCnIrI5g2g1NMR9ChPciWCYHapYwM+e
Sv2CxMjn5J7oYRCF/WBT1ntPCTS7xBFbTa3IH6TljhmTM+aoSsGq7y37eH18KrPe
F2Jsl4JSTIOYItc44JAD/M4o7gcLXWKyYbDplfE6UtJBzc5WEC9cPt8qbUvJsYYi
Vl5XF0ZL/qvMIjrpRWi8WX5asO8d7XjAtBK4nl1XEX7IeieX28cZ8VbZnc4JJAMz
cxj7eARLzcjHshPPuNmqY3aCXGCJsYzQGXXc2VDluX7fT3mCOOSUQaJfczlVFGSk
4qCSk3jSh+Iak4T72MLhHYiEeuTlg0QpdML5UiyCMQRwhxP8y0C+bd11iH+zBRz2
+SQnsWgcEgYp2WAVHWvEWaWfgeg7P3Yf+BvNTmsJnTCa6CILFn6VC6YZd4UavovD
FVY1oInUBfmLbhK/Q7JMLXHO48d01cbXWrQJMKduDE8g+90PGMfHtn27tJGsUYMC
+5N4c5Mal3wDm4ehH0wk3wZjnxWqeAbN/NaLXaUWqveJajWqz5blLpJGcbV1Ybwf
P53KaZ9aBNVCbI7hBPUCO6Fk/fJCf2fLdzI6pSAJKZj3Hzid3/grnahmowRL2lA8
7PGwCHxOw6aVapX1xKTIfyLHCc4WfHY02tztrWaTros5w8LwfrG3rY8UfBJgCT3t
H/h1INeEv3+HeCJrTCoxn4tFbQEXd3Ai+vNQXP5EM4RHVp21hxzH7RzTbS3J80qU
tAk0wqORzJhjaawTgXvPFjsVvDOUQ0pEiVMIhC0hGoiBGpdmEgU9cPs2WX+gCL1r
w6dL41ZyaTNSug0iC9h5/J2Aj6++O1GMZbn+9F2bSq+wE3WQwNMgZGVOOAb8J7k0
+uKwDqHtYEaIu/yVVfbHdSw7nNN1codpNyymkAbSWd2tmc7LStlUR71sZ6FQ48j9
4lpPTPeLr/aGLPPXmUp2uIygWdxcbsYig2jvrfZR1d4CvRCYUPHx94W+y4I1oj2n
Iw7Dp/9K9/nUc6/WftoNITSPyTbieJAfMc0ITPKq2ze3w1qcCxjBKBfFZjvo4cMg
HSPzWV20nhj6gWT3iEd5tBspwyXFS8KpUSdT5aolt7jJFKT2sBjWR94jQwEmbYGZ
+l4gCObpwmdYuy3B/Pdmaz+4pJWOBOnM/nJ2nRcdjERwLJm6m3/0lRRk2Bt/Qo2Y
BOmHrFBIQlEQa789ZLUT4OwKB4X6Dv1E60Li5XxZsGrreniZJwJST2j77NFAqC4A
chC9udgVisiwZ/Fi2Og66HbsfBOu6La+LzMKaQBIP4fwfYZttm4szDTITsxa/oEJ
mLAgRfi1d519gCQribUHMKU/uO8lbfQ1q7BTgLtnlIw7Fmfki+mIYRLGArZHDpnT
gY8wlXc91XXSdflVjrgkGS4r+hu7JGY0bp9qkgfeJvjuXjBXcWcPZ+qbOsfcA6eq
t/DUvpJmkXIE3iUpmb3d5hz9yKes/RsaT0neCUUAY4jtU0PFvALifsCwfKSHeGD/
clz6S7cZ1UzEpthp50sKtQUn1VNi7JAjL0J0bWrLMHWlcZST0Wlwy8QKg0vgtoti
vr+dfwQckSQUaO2pKE9QXj21OWvCdtqnGnz0idFR6+a+4C0Fbi0qOmaX2gHI3Zb1
o7ihij8EbcDVLygtmYZi0MOGgOIaUGCw8zOCvrQUUoe21AFwMGRnb2epvTfYyNnF
Ywei8T2+jLivZ4xKwW0GwzR8vJC9YYlfunhl47rwaq+fk3oSle0d93WkcVtNgCPE
PTo40My16zgY8YaHys2P4ydIQck84Pzv271ppTetVpkDaKIlbyjNr9oXH9Zn0spt
Nf1Hkkhotjunp6PEQ6KDqeZAU+OuYdxCwDyvIzUN8hokdKawd+2vo66YBKxH0TBR
GoTlJ3jddJy+dGtlF9h6mzO4LDupMpnvtv/zCyYCJ8sQgYDHEtCSFhSbho7/9ZC4
im1tdWV33O6Bh/dXxGDnWfpYVrgMRXiaGUA1pk4CCt6aItMca4NSICxJ3RzHPkkL
lSCo4AHe4g5y4QCbNtENTgJug5lsgH2N7npT3rKglbFCkeLzqUoBQtJicnOsTKUk
UtzrcTlOQEiJVLTkuhf6YSXTMuFioFnLZDTISSqLFBLwxu7qdlNHOmv5a6yOujsH
rA185oZiWGATAmwgPOJ8dYiqJD5tfCQuCFeg3aN8CN7p9HOCIFpvOmcYn2gcq+VR
z1ibakDUjaxckVFE61DPzYzqbXqTk4xQSbI7d5ovUS3zPWhBQF8e4FRao0Z9VnLd
dHBgv7Gd5Ju11lRAHGV6wyQNN+f8ytkX0beImGEvBM0KFJmkQPqCSDc+E3HSpk6H
S/favyibAtoJMrFAwaWTwWE9bXUm/LvBHhyzA7K/1DDd0jGPSSj8QnzXw2EFprSy
PgP+vY4c/m3eptdfzDrPkQcDuw2Ug4P8RshVid2piqhCeqfHinDEOpNSZRbIQ5TQ
2Q58SZDA7t3MCInGQtCWkMJTNKVBwE4+5r26cp4mmStnMJHaAlYJKE/3YhdEXoF6
GIjlc9+Ga7bdFyKIqrAC6TmO3Da97RO9TZTPgQen/amw4lhqmAgRQgH3Sd36KI8F
UhWU5NIy2jX4F3kHbJdk/uh2LfgwIpUpoq7L3atAYYWlxXhgqie0BY8zWx/4MyRY
1qwrNgN47lDmZODsTKa4biBKCzNct3fmKfT3cscj6Qge/oqyezQUBEzmmCNuaHnS
m2nT6SJ6i0cOSUpAj3Y5ymOWMFgkp5VMkYMDRKmhNa1O5kr4l3xUQT5QFj/60/RM
ekPIu00XtRkIF+xkUQ3ov+htyZvQV3UUHRDULlU48/4srUgME7Ir2me+SP6+nlxG
s1SdwgOTKDSl1c7tUnsEEA8tBnzgm6qjQG+x9HT83OTzXKLWemXjBMsCct8uCRfS
O6ph4NF56irINfjLfXsNxWcxxSAkmyO/G5Yk2Gbw8MGWxMm8eDKHQeKVOpQ1H3jf
qoy3mnJKsHHIXNmTRNjv/2LbmTLfknVzc2yxuJAvENtCZa4pXzq9Bq0VIlEgbuXy
yXbVffsNVUMLxgHTWZfnHtvXsFOdjs/lLfNubxyUhXQbbXzfEZWUdrRAxlUDag88
WmAPZi2Tif/C6enpSP166BZQua1uHSFV9+nOvASKyyM2vDcHQ486ZKJYHfcbtCkK
rRKq1LJQmUoobXUf49I+VBVoUAKqiBPhTOR1iLXsG5tkzVqV1Q0ShkOQmE2ctVCM
2bjn9P5pOOKYgTYHlxp5C2KpeWJsw/0iZ90ddud7sh3k/Kn7HAq8ZRIMPPn868eX
YTPV9i+tGFaoEEwEVgCTiQU88XMaIiujn40fJTHcjEwt2JpZp+ZHmT01w2w/7AkV
11rO1flID8wvNKycAIJ3OwgjVHQnzNNkdS1bf/O3FbR+lS+UHGd6hjY6+CG2jdgJ
S6UvXJeFXgkJkwFDgQTK5pjSqoN94qN3QaXspfX31cWegnYLDnJT5GqORuIfzDCX
6S2h60nypN/TqLe0n/9mpqJzik2P4vh+EVfXNuzIQFR4hoNv0HWBu+KAXXmzLj6j
86I4YUrKgFf2hVsxQbh3vDovYDe2IIrZGwQTWD9Fl2IlB7z57xCMpfsjQejyG0eH
6qmfYAaKoui2Id392apgNfjqE5hXKCgZ+dP4YFjJK9RF3c0ZOyBT/nwScbVBKw1K
2JESKC5GV+QKotf19XeHcEG2dBWitERHLvKP9PVblYZHwCTTSYwaSScY4HpJf/If
aGFnYVn+51nSX279HYZW5758idiSt99RWKcEhjdNldnlP8A35QjFglcWe31kzuYl
Rxa+Jj+bXMx6t3qYrpCVkjY4uAev2jdToIXo57qLqOtjhZPozhEv7dkTNIDerw+U
EwoRxfl3XxH0d/aAHWAyw+DroB9O8rzPzswktkGoWojqI8VmUpeNrny2bGI/mNPK
x7NHkB9ojHLQOIyc13tB3u9h45dL5lOTy/hP2JqufVxLFAz88Oh1M/4guxVx+KCU
R4DchTlYcKrzbvMjYu1fKqih+lVAnmZVhyX3o41YGD4RDuMevOkL05AcoquFKXnt
5iig3dlJTfpdY5SyAQ4Zuw/YPjd2QfYZpSay2zKyAzEe+Yb+2Gty/Yqc+7UrTXhM
ozxfNgKNsqC+cBSauRPQUEv/j72bribOwhJnzEM6mFhTgCwy9j36xBiG0g0dvfod
ush2zkzszdCQfymvul4lm6K/5+JgSB8Yy4MD68JmkqkpmCTjLIlQLkPh4XTeIW93
VzsPPVPOl7ltTU28Frtt+u5r9wMOkOnSuIJYDyX7HtY1ECdd5wkd32sFAj/Zc8GQ
I+4EshG59cGFLnpFbvCdzsYSlCvo7z7BLS3zDViQEgVLb2AlX2a/NLUFCD1MT63Z
CFMhlgoqUA02CTbyJe+8gaZKrdUiktfMmyuXuOIHvvTOLn9NAhb9Wd/3uuMmjfJV
up+XsUpjdrl2JjMouY5Frr+3qjFL9lBShZmfTZ4o7UoHDmdDVEm5Zs//pJTLX06+
9gUiyoX98Zx4lnK4sE7SzS/UbByGBMCa5xJAv/Okcu8/DF9OqUfIVx59Xon+Do5Y
ZcNvEPXIJ/sCdx/Kx1pFowdJvKcZMXspFFcRvTJlWr6jZeO3BOga6vDOLvotdzVU
AU0bqajbdZilGBLB7vEvQxzdBbym+jvBelRL4orWgHkgemV3PNN96YWPbZ3DYqV7
IHgpisbzKUXYQJBT4Vo1cJi4sgvySxTl9yb8rTZ0Q+IKuSOXF9pdb4RkMhkZPko+
SAh0hnFOuux6hIo6nvNpVI6wH4JWDYnWjFPl1GwlUfJ2WJmDQUkHUhogOINNg5+1
xa4siKKXV5BDopafE7GGiVT7F3YZE8jWSpbX9BsidRmQLab0K4nm8ycqvW5fFe+d
RhVmFRj7GzY5K2PBXPJ2W7XOeDjmbirZPgEvzKtB1pbFtOMntAwIWSQFQCw4C9bT
ZlXWiHbY13F/32kwoVwuQiIBtf/Q+vc9x3jcglr9AVCRdWMgUBbtYd4AdLU/nbUB
DzD6SlyN9Ml9A7BFFHGfMm0EM/aIqIi9jPpYkTRT2/NEnCotUrwlxV8Mx2CHXhIE
AJk1UgdvzsX7muy8qB3ihdhuAJDOpbbSOUdaHCBsuv1XyUB8VkqoAm0qMi53MXYm
v9TRnTsIDdeeIrEzkH4HUkKWdO5qUAxpRPrwhFQdQx9WoeaSEzTKoaeAojGiO+CO
CoOq3ulmRpI7Up8DnlHIEwJASIJVccxXx7h4Z1RFz5g4rbxwlZYGrX99rpSVhTBP
2FFBnHrg2awgJaRTDu1suP1JNWaFDtpcJSJyNkRlroecF6hLHntC5BpqbQHwzefs
Ry+xDLxRgaNQ6kXrzTLnZDpwWvAfduJbyoV7Qt518xq8SZJ8kMzMPEeIqD41LHbK
YGNbY0Vz7XogC4T7UMSKcKtrHU4KdwI1+SceyhYE+dWOiss6jDEwfLqy+4fGEWfM
Q+tAqtyZZEc8mTeG8WgjGpi+y4dd/YjoVrhyMm+ajznqyQEyDI8OHkFEqAHccD9W
cqsjdOn8baY0AQ6Qf06QnogHbM6MbXhR97DxV2FH1mV588WIMVqACzfVxCj7oxig
XhYFO4VAIYLPxmfRACy+pynmh0mz7K9WpvR73ZEy31XgNIiKOSGvH3f/Y/jEVHjQ
7c4S8lw13ASO0UCSn1n5wQTRgy9OilXXXen5OFRKaul1JsUw1UvYMnyNIwu27bVi
7E9C98xOa3TDIKsEE9P7l2SyNUbKRohOaiUjSYJWN19x3dXkITBDUBl7a0RtO+6L
lHjxXY0vADsXcZQN5489SCli4fRfQeV7TVG4W7zBxe3mHwdrn6tEpf2lZzBibsLn
gdo+72p7fn9MpkBNcjlwk4mGYhE7P/Qdoblo7YHTUWzEiD0pZwWN/l4Dci9p9sW7
dwqog2Cye3GRgAp2sKZeJbjuG1ItnEH/sILn0ri9GqRtXE/OZr+yBViO1XUDTfGL
yk8Rj1DHliFUPgajNbZj7i6OSD0YGJDp3TFw3IB8LazZEEYXEocLnzRBmME1ib8L
gIpP65898Uu+mIDV+rMCZAaxV23GFqDTsNiyKBe6Yrg7IDzzmTzNPdnUfVHU4nLB
6682zZMF3Tv/FlQ95XV0Jx40Ry2qPbuavNm+pMxJx6fIDY7GePlfMlR+3lVbuPpr
ax/rzrlaGN9xXpoTS7YN6VgbWjzQlk+z1WIJfA9s3h4XpHs/DN7gso6GDu9stbkA
jx2n9J+K9QKY7WkwM0nK+zXymCfsQNHqRCPV8eljuNqwhjgu/hi3GNw4chpmfoWc
gdt2b+G7dLa/dYMLMUsVa6qb+ukcRJSuAXU/Vh3InKISezvg6Squp/U9FbOh1fYh
P+qqKhyhclyG4lm31F3CEMZjmQBJ5EVVxSBrseprFWPciV8yMhdYvnkGPrhugTyX
bYbGboXM0+S31dvwjcSvZRvRiLVXZqvvw2+Z1/JQa+KdQ2goFahU+rwmUObFVPt1
EdFOeQ2VfVqDaa4b9lwNf5e8/0j0712XpPhN/j90+f3pGD+KvbYBHO6SELj2HmwB
erhd8z5UmAIqRn/O+19f0wnrrXxMSPeLOfxCY0oMiWUSfkPpOnwoFeDV1Gf+yAVw
1UGLZM5/ZURefjEcJsl10zk/aBEu/eRdUn70ZI6igI07CI/5LU1ppFXZVVDs6ULf
v2fyx3wjYbjZpjv6fZeBJxeRmjjwo1UOkLDW20OQTYY/FEvycFEmRB2u5JODyZEh
ICswagQAJ2t0MuvF89HeAHSYDoyrSOnSxyJXycjZaE0cufsKgUAIVg1LG6dFihdz
qx/EYSWaHDJCqrVK7N2czIA+uCEEgsLg9IA6MGVrZKQ1jsrl6LARU/PPXkSEYxmP
PZzhreGr99Tqt1bn181OVQyp4a6WHcFbaPJ8SfRqU6DnVPcxsJC1xTh5G+4b1G7t
Nzvput2a6ydCLyS7Xi7x/rAWUfNGu06xQB9715Ptk/6J6oW+g0unQ0S70xa/VCWC
HzgM7KbyOnW5JIQbuTvASYaO9NjnhEPT1eHMrKtYEUpXUXFzBKOplpihFKpHtHmJ
dUCYbQf3EW/M1/x1XQHP1M1DYkVprHE25QTsQkTgzSReldE+wVhfNgNTJbSYONcb
uM8lr9FbSOnlLh8o3MFHmmqKeXYjK/kR5Ualyds4nncwiseobZsA3LE8YMKz1CIw
wYHNyJxE+EP8v/6x8tH42NaRAjPLHy/OhWqdsgvlCK5xKf0SNf0JcEK7Bd9AdtuC
BomoJRLSxMg7vdR0FF6UC7h47+zlwWp0kTAdsMyJOtYApm6vOCkJgNhfbsXIqA2c
Wn6rvnzyQnngxFD74jvnUDEPqf/Mb92Td51cIRaTolxKUKjsmAIoZSZjzj9KKUcS
LN9Ynb2YOLb6nXYei/HF2pY8GAGBoW9e27XHKLNxnlsw8d8gxPNJ/eqxbIvTP01D
tc59YT4K64f6S4xPjf4qU3+KKf6BrDAgs5gN14UJe6+4JJwvSYhzGU5Kba3iYwOu
mIyUnzu5UDaRfZnQriIzrTwPgQZtCwoGGwVBAWlipaXEeGr564Gc+5gyJVJwcMqi
79xJ4TxqGjaWyIPmoDLX/QCUtOL+OGh0sX/DQEnReEkxmLlN4Pg88oFQq5jA0pzR
VgYJuT8uvm8k/lfsrjLGQvKFTKfivHFPHZtFH/8K0u3DX3FhBUlj19kwIxSP/YAr
V3J+tVY8fparp/dlTV/tYSDXjhlh5b2cz5AW0uFdRNuudkkbwjO0SJsAJsEAsmFr
kLCmZgdmLStPlkHeap0qzm8mMQcfeIP7fopSZUoxWlOaVD/+ycHI5ezIiumZGuhQ
Rblkv0UqZNNRZMt/MoYmg4nDQ8ZaPdeBUPaLILjxBCM8ElTkeTho0mogO+TMZMTj
z0ZMkbqTHdm4XORWD9vELJCXh6CKOILGp77Ba8pICx9Uz17spw1dB7iBHaY/r+iR
XdhN7sojctMbVLiUWYrE/9xO7c04WTbHZYswX6/c7QronX/splS07wuMltDIm+qo
1eK+fhg1AlphPVRCGkhFXzlCfRv41IgTboog4g07MZoXLD2fyk1VoGo2KdtalYiJ
MfLVSpniEl0uAwbSevyu5UB9h9uGlaoKx3PM8Z7FGpKFcI71k5QiV8po2QHogB9g
faOM1FSIDEmTOrqWpkEU7/Xrx0WOGKA54s4/7hjJXWvplBOFIo8pIpO+VJvXHPWG
KRoKTMHDecR/AAAJlcyerTKzibnaGt4dq+gLVISy1h5VXD/Fh+FelE/YiS5bCNtg
vSDHuMFrLapbQ7DAifA/vr/AYgsGZEY5d+RAnfGfGXDm7vroOKijVUqwTZcX9Ie1
maXbqYhjVZxwdD4P1CkqMu562oUP73sflk9jC0XLWpQnVGS/olgo3PVk9+oRydS6
e+3agmrwfCf7k4IOA0IiYBZq0qreZZ7tdF0oojKyjxEdMyqctuo2ny6Twu6AlSYp
mL5FdAycd3ZKjNwKkQgTFMv42S/s6nkCUkrSbnEhI2TaNcFTeks9frOmst20bHL4
w7S0UQf+88vMkCs+cAI51i6C7ioedcMJc9PjjK+A2OuUsfNNuTHIJmYWVboiZdQa
uqBRRXh6lllliBV+zEHgHODc0PXsSMdaYUK6Xw6JJhnqTcGttuzg/0XnemPPOgtM
6E8MA+K+kNOksfrOX2LYXFZp8CD4WYfV/+ViUDkVpC5x5/JhXPixb1ZmfkhVV8qN
7g4rvpw7xCrzAe3KxPqo3gpAjXhMwUhUjx1+l09Yrm8wXNyriW5j4KkBcNLHjiCI
62LvlIIcAXw1rMhsLzd6QrzqtOiqkslHBwek7ZX7z5OJqWzQ0lDtyxM2aWGmSAz9
l+0gZ6fbtWiZp4YM7ytZqkwcKSH58uYdoTALrAnR5t3/DwBOd9sQ7dwhXaB+tI8K
wp0bsb/QiheYNoqMIqSxLD7tyoB2mPEqHFpK4PsCiqqkkG6DJnCY2ooVa+sLNyGM
K2+rUuMeeOvyUslHxLWNcS1/KI1ukbeq8wFCQoiRmc+hXvy3fDoQhRcRnhvP3pgo
bTLZnLYY0GdQGLJHyINc/9ijmu98s0yXHBZcGArZ7xozj0s09F00aCHVqYbeobjb
IUH9t62QFqaK1WlblJGQXYQbm3rCRiNQpuYT0DVCrSrGehlnYigBCzxpzkBj9MVV
8wamQH2sYMkk8hJi4SZFCe6iIFLtNHJvGwdpKZQNQA7Cn/D+x8bk0eWV0nXRcjZ5
mBpXnILERuprHtF4yYluB6eNJ+Qle13gtxwSVdvbaqeMo6ZclNfyNV5ZPHhicEGj
rbnbbBi+j/CpCiDerjG7XPjdVw9t4J03vm2Jj9ibi0NQ2ENedmeruyn1Nu8aW891
nr47zo7hFA3yn+AZjIiMfdmT84gxlLptIIk4DbO9d3JSjq9XGsJgHSlZv08apQR1
T+uNifMbk334BddffGTyWwJChja1/s190Lh5lFIhy22oKGrupciUodW8rEnZZT0N
BpJS/H6/MiuO2FE+tC2cdr/YxcReEhn/5bR7avdqLlCN3+wjG1w3JQf6UQhYZGk4
2KCYWOecukt6h9N1qzO504kf3CV9FFYzeWUJrIPgKfDZ2VdE/O8uae6iCqM4JfX0
4WbXM9vyUaNRN9sKPLe4XTX4NCK5BLgXpk4fkgID+dzRAyAJspnrXrqXCULpNdN8
H8j/VtgwenNRQxohHmnmuusgHTUxx/yAnJcxgK+zpQ9Qbldoio3nVCImLnvOv3Sg
iRPgxlbxtAyQKPiOdydhypmQn79ZzrefJZOTqj6sHsp3SsStoAAo2bjZTis+lnx8
kI1HPb8vGBittMbqnRMO+BQavSDT6jSZjs7vtTpKLA+QctBjpQO463ZdYgGFYSZk
g4mC08l6G77ml3ZopgA54BqCeTbC0FM2X1w9duceruATbyq5B1VU1EoFcXVVf8l8
KCUastghI/fmAgZLQwovA9/bPAT6yhbmaYvni2w4a60zb46IB/b9QcmPt7WIWy0X
GzBFdt11uPgGZuZcZLxw3SqDZh8aFfV97oYrycXsB52x8Iv3w98lgohqklbiJNsv
jpkEQHr4xlX4xHa3XDhanQaZEzV1kfmPDyZ/bz47VrK3Y4nDaT1n+9Q6ZK2A6/Od
pU4RYuF3/SZ5Idl4AA3JpD+q00ZcjCTFq5ijhwiGqUy7CEnle/Aa6JVE+M8aMTeW
0omSHUzSMKHbi2zQgEM5zxS0WWupaKGGu8OoqNJkO2c/bfYHOe0UabTTbcRLvLya
8KvTJgVe4rV7oQe+YfQtXiYd7ENFREdiWrO/0V7F0GWhWJocGaJ62RebyiZMraIv
haqi2zGkPlM/LqNokP5rVtHyUOrvL5T2UAli685iTn/jWMb2zjMGOPlsT474IPJ5
ULrqetW7Pa0F54R/R3B63YBbyZwmoFmr1D495SbEB+XGlz8FQd2GrpFGswYIwyOd
7JWRYG9Wij/juUHUxWAVdLDT/3I/dI9qhLREwwt0yj0WYd/lH9pBKYtN5eqOv2cC
iTs0eRxDBACkETr0aYEbU3vQULsrkgplRB3p2E0IWLv4AsXsRxqzrbMsjA/yFZVI
/hc7hqes0TUBk2QoNEntwsp+OuaoQfgUnp51ulWGsyqjYtXI+YZczzz1p/QwpwAf
kpwpANw/6uR++TrAJV0LwOK0iLINCfdAcda9Di0A0NQFGYvjYfFP6WKyscfpYRrJ
38+CJrNbU4EZd0J3Rsa0TZbKqZ+A3GZsBviCCxxa7G6KUt3gZNHGulH1uZ7BKiZ8
mtUCxN0JTWeIu0E5V6Yw2ZRxuuEJALlJi8kLBghfkojkey80B/gzLqOXwfAXh0A+
pCIklmwKKX827DI0HOJhzRlz/Ylgu+96OZTkkR/RzKdC6pCucDUJMuAU2PvdaWRd
cyDQSn9MNXHuTpChAtjLebf7BeNqOQZOpEktbhaCLqAh29qm0n121/VVMjQ5U27T
Wc9JrxTAq0IUVOekF8UPLrU2SphoNmeDB0x0+IGxA+U+olri5Nbz8bYHCbSnIeJ0
B3Hes0cvcHP+Qu7/1ioT5VWiVvu+8+b+hZ2koFaHvL2AcWLToUhifjW1uw5SUk2Q
17cCwuvOwslh1oNq+rM59jNkOq1cDik1hNx4evZeTG3ypgDRGm02S5fG2EADdr/Y
7OOP45xTrYMZ8Hemjg/ynocwB9vbM7gjoHaJpPRT9O4btc5w7UrtfGMi0UPO8NvR
fPmhlLKcDlMYbXEpU1NVpjjW7AVk5NFq1FSHW183ujpW+st5dwxIBokWX7q/B1HV
zDhqpednI0nXAe/2IMaWEpcRh5z2aUvZd9kewG6COHXsPQqb0QpUaL2bEXTBPx9S
JcOYrvRtyr/9n/swXRQCOoFjnH13wKtjUDZYol6kC5BZ2lfoD5Ffqx8Mt1pNtuD7
CeIW3R5a0UK54hIwwGo+vZ7k9YPQxFgutI7sgvKZFBUin8Tesknh1L9SA6M/bror
o4HXnnP6y0JLxr4TKxSSJEXJzOrEIbVvMAaUjO77VzjLd7yTlY3107igpcrlpilv
1Rp0faBOb3CJE7g2pXj1JAa/U1pmgYcFUzla3jKCbrz/dwh7QL0Re6M6vD57PfuG
ssUeC6aXY0Wg/kx2m8MZgbfQOt6NDGMvMWyCszU2Lo38TVYkqL1cWa2rUWgNC+Ff
NLMvUKru2KVg0TZTqLClb//3RZESzMx5sqRcjFRRXlM7MmK9hCxF34fxpY52J/XI
Sf26Mx2ugSmxX3IV/KhF5dkUe8YbVHce3fp3tQHeIK0fVfM3GrCtrlNgYeMNpWUx
TL/E03Ry9JOZAfUqQSKqT0zMImFVwcQsi0uYaKLiaSkGoXp5Vu2pTzVd6oLiwuHu
xCZqm+HMvG2etIFhVuBBRr+QiEIaTgv2owMaruhbD5Gu3HJ9arMF6z5ulJ8hzl/0
TOTOSDrVYceLSL0yPhXy/+KLEeRo7/aCfn1g02hnAMwet7AabYsAjrEQa0Xfkjq/
EfDrMM8H2ctbiLpKY6Tfbt24IWi8xNyJHJlHo5CVcCrcvCorpM93xrC8Zl31Uk1t
V33GyQ6tb8ZrJ7IyMoKJFdWvK+y9q/pu2sZSaBDciHtoDuzXEAcCl1xv36H0yzpt
1dLFCizX0kSztfq5n2xu53UE5/hmr5Qgm+6dpsFBirr/zC+Bcudrp+tNIshX5K/v
XCiA1xYx870acoFT4raiPsAshToOTrx0Cxqu2gY0Ut2K8OLuMfgPNS+ee3o4caWd
nQ9D+HvHPSCKN6++0sucNOYi2cKMMGsV/jWK1gjcVag3b9MNsKoNyybd8kQYXBfT
S+GETQjHjkcD/aD9JGK1b700dEWdhjeIkaGh0Xwa4fRgMXWJ6mSCMqvqoEeg9+rp
kg1o8QnLphe9yA0Ja/BOB7SrjaVYoaQaiFQXSP3MleM7QJfLzc+ka9jL9QW1Ult0
FPVGRzcAYZeNm1OV1xkhffFS9nlsWsB6/RhSYpxqANzLG7kC1G5sC/8DvwvyfKgv
PXGwWehNDxMxj0uB7bu/0ZjuX5aAoDhMiKjernyUc0GyprgIQgevGoQC/+/tyW+4
h+NQ2jcFObl0zuidBQyvdxr0yQdjan1YEHDRAivR4V4DLAPWx1ej2lnhaTrsJsVg
X2Di3/AmMaukjQyILvIlEdbZ8WC+omKGSUCkEWkHZtnIV1iYNJe8EzOMyCH221l8
7+8LU/mScqxijdNXdTQrodK0UlTg/H309l9inAkeJjuE2ujl/iM9vId+zp1Hrb/I
IY/jUC82Dguxt1i4yCm7+3CXJQVzMKeaWNZHYXq6M+SJH1VPP9XgkEe2vQMj4zt/
cyWrBoWOar82CNvbQcDy2XqKVXQUbwsHn5SQCGaKTpY5iarZmVIlZJ2vmUJEMuFh
XZaLek9f9I3nD1Nand3KrV/5TS4fMb/VAA5n304F1kAFzmvHUbEI3DhKtBww0scj
zBElIMHBqrm44RteUeRhM8RSPwqMYkdUqEY80ZgeKBss6u2e/31HboNGpWWNntZL
FyRfTkWTYfjc63fg7Ap3H1ZRtPSNOi23sw3YlBv9u9cviQZJj+psJFbJPg1et6ZV
diPSfnqa9r2Duhvy2E2wtQP3Z+hTj0h8vjmFqSQPCamLbZB0ycnxWg3NEhpTBqH9
mdL5bhwsiHJYnip6DzbpY6LDoPvlbY5kAWLbYRaWYoouZ348q9T8yuuXCmyEA6c/
zY5r4f8vKwSrdTveehvJrtq1SpKGCamx3FLCql1PueZNEi8zWB1oIEq+S9zE1pDR
R6udn9FtmMvj/Qn94XiGYSpNz3eb8smfZi1JV/cgehVu00SNDHCCpR2UqstfwX/c
43HyQJc+8aipPpcK1vQTqNmTPX4oJfjJgGkDhSE/QM+WtL9dcrNC/yE7L4+p0hUc
BfVCufwMOsNeBVekKSvyR2JbZhGljgkcE34bJEu5NScnqKTvT/8Dit1BJnKp/O0I
6kjA3eZ80f1cQmBfvVEwKwMDeCwSP0cz4CUGuayWVFLsAaX9dFrCV+5B5clXu9ch
8fFB631DIlqpdmdQRdTOvC9dn12c9zyOJVFg7AxvbymmPk2/lmK/4sRffRUCm0It
d4MVQRm+TOjV0xjnjRcp+DQhHFTNJuI4fYg1f8+sGbObsh/1blELEn6xEgj/B1qR
Euun++ou0NSZb6ZYNMivkBct0IRgXGc2llfhQCPGonVMXzL4dGNIw8uP5H3zzfMp
vSdZWd0FYyrN+BTOOijpmvK6lE69/2y4qyGkcy2lRvkvulUb2i4IBqJiD/PK0uq6
rQsF//JvXkCVlUCYGQi0GoaIwgTIICAVx9abeIcqg9RvhtRGloRnzuLI/QHon9KU
x20IsCccWKeUO5o4KcnQuat1b5pM8DMIM+kFyGL3zF9xlglayTapsQ7fqqvROdly
NKF+yRIwqis52j16MMVpRMnAkeD43oeUdUjL8wen/4kAuwEmiXe0PRPCReZY743L
iwrMEj8Cz1fKFgmQv0QwW7BHsXaY03fdBIq4Ngy2ZFRu24V//Kl15Qg6a8ja29j8
ASSo1WOa2cx9swanE9ZVb2FSI3ghfOd328+i+G2pNSKWnc324YnQGI/74is9B4m/
0m0CwrXzUxrPNwN/xx54AwDBbWdhT8GzrA60owJ/6oS2tc6YStsx+7iPjB6DB2+g
aGqRE8wrUatFmmXCogxf9nyPlHj9D7Do//VO/4G+l+L2zKcsLEdSDNe90L5e3EiO
8I6Fqo4YddG/fHDnKMcRoXNqVNRWJ6Pf7LO0zdWLfobWCTsRZLX5Wg1FlJxPy2Sd
eBXXhPFRF/3RGENwD6muxFhyxLJy5yb8WQ6n5ClAzNxmpM7MFOJ4rFJ6imqg6Uf7
euUV5S29byj53c8BQ1UTmXMxp7Wr5ACcClD5+PzHq0iXb2SaolDQbULeX2OFKj/Y
sZem794S7P2mPXAqTJB63noKTvGsF8oRDBIkSR36JyPd6jiiaTbeQN2iKBJugKyb
3doR4MI+1klhqoxcKhADIZkTENFG5VSfS/Id4MKMx0Y54T3hKESXDeC1OCAuv3YL
f3/e/PPCgpBBNxbhQhG/oj0QWIdu7eMrez12MWRAaVl4KlyKAg1Ji9mMaV24Qj5a
EjGzkhEHq2i6hr+TT9p3v3gZLsJdHf/ywzHbumWgScz3qOEIDQj/G471RmFX5BfU
3WWilmGKUV21s7TuFeeouE+tjc1erJaFZOLYaMegJT9Ee0lBbmDVKLCikZjiyKi6
x5hYn4F025Y9WAzXNrCvm9TVewWvAsFJQilRqx4VrwAudvNDSr0z6MO3uA+HrhNh
21vs3RkuPnSCvm743x1BNnXvXfRoQn3p1ne83UP0i3yUx0j4qpxQ1XGs4TnEfI9N
aKzaxWHjIy+pPQTLAbDW5GARj7fOUd43sI7v/nZ7pl+GXUp84dYrA75FfnxVEBKH
t2jx1nylvjjMELnZ9D4yL4h1E0sJGGEl7xE29JOa8odzaM2T6oTbcA9r1H4Kg1bQ
dIwFHC8R9gx4InR5eqS+LkhzJ9zMLdIjO3t0VsOqZQvCMQhceMiPthecnzpfDVNG
nea0ddHWJDAE3gY4ycrvQ81eSfdHxU1XMzgcQ0ra+NzYSUof8C3CRGZAw1w0NXQt
HMOHkGgJWMnLZyy4Et4tsw9Mt8az1ruPfUeWqgJRAA4XKHGxfiEXEZEt/N2/2asD
wDQpvlPPeWsTtnajyuMXEcTUx3rBLPc8w/iKOtlqy3FewbiSycdLvthmuXpJY9DN
qSKrqEYajJINzofY1YDHTQBkkjIxxjtSbvbEYUVq9l5YT4fDMSwzcdxJzYdjYym8
NY84Etp5ZrnHEPmHF8iBL8UIahYTy23K5LCOjWYpewWFz9QiJdG24frcZBC/Yvbx
mCRV1uKPYOhX17mIojUuaVy37jtnYwk3Swh9pas71Kmtj1hPoPSyNJNfuC7q39WP
7+sY1ReAqJmlr7AS6eogUDNrWqXK1DJzgEACJgQ7wd3giJAwGWoM+gXfKEpn9wPZ
VwPtibiBgGZENGRrwgx2Q1p/rcjIDygGofZU2CFdZFuXnIZnNweZ1qLl3tLXi8+a
7vg2y9lZcwrVbna4mg8t/PbvGZ+4rj8vLrlflZhc+YDrEqQdI/yi7fnasFLaKeFJ
BqYGft4J4NzTm/iWQ8geEs2g7jVG6v+Wfn/Vg6LmxROm0oGKEfdca332yLXlL17V
Sokt8ARWlerc70VE5U0hA/na0zdxivYDSey45aYT5xXGu3KqusCfoj60L0GurSbx
Wf7Lc9j7A9g/yrV4nYBKlzYRwKs/OMyCSBaBeJtC89K/EmL/DdCuuJFy0EojWXwA
G1rXCJ3hkOCeI2xbpQDP9NcBHIaFpBcH3q8mSiF7nNQoDdBLuf+arMp78jdj9e8D
ZG4biwuikRJsqBRxdvJHsnXxFlXqG4Fg86adfpx5TkMo4hiDQ6oHHdq+fO2llC+T
isoaxRG0JOTUo7psiDB/pcsaW8JklIEiWz75GKfyB/++bKrENNHHm4nHAhMq1cDD
uik56waf+WYRck55YgN445UcHSj4txKtfNfhEOsPMqEFbOLv3yCRrnxn+iR3qj6X
1r8QuGu6t4tvP+XZe/lLHD2LBNJaX+ygPAmMGlnMS6P6UF4JYS46RLgiiOSh2Hfg
mF4uB/orzWyHquxfxLSK42QeR4Y01YquuUFbuJSX1xvkNM47ZTjPPkOLos9H3qRo
sijZcw4tnE1S2JdI+57toeeOPcn9jfMPLMmvOkqFBN5lSV+NiSgEM0mHGQ5kYh37
CAMPQt6DQJ83F+P9cXvOBmJRdqfBc6enMsisBMwrWY2CgWOSIBQvDb/Y6P/QzEQN
xX04yi9MZblDheDsb3fL4Cz8VQjJQibnevYHYESYjr5hDQQYr/1qbf08ncTjBndV
ip/DbVd/rUtc3gZA8oA9Y1ROz3iGeyEDw4Xk/uEXhImusnj4ybcI5YuDj39jMt6L
mGEKvqIX0CA4mvLCRZuuKDODamDOUiEWK1HHty1ptI3IwoS8KhnY0pbvtUd8ab4n
1mkcOi+LeX/g/2SZUPQdUK8e2OCMyL8RDApsssSIl5sQqjkV8nxUQOB/8/tn22iC
WeMHOrKSBzL820uWBMRXgmONuypVwQ0t0wf7zISrPSPkrFTqe8JFAuCh60n2H9W6
gTyTiDUz0dXUABuVdJ85sMfUgBmb9F+j8RKJ25NgGCY0wmo+2oK+nuIo8A+1yFP/
TlKmGtG33bdb9QJAzgbQmd3P5SJX4+56AJgAciMVABNXD7u6p2gRrH+JAMTRCWAJ
uVaJNtvj49e0KFKH+GqkprDmme0THDYv8N/oGw6n+VZ15sSlBxQ6YKWMtLmTV4y5
ELRW/8+ra+qSpBYZOagmMBFPeL/VFG6bhhqI8rn81ap8qO6LRu/zp//yfIPOJ+6j
RH788gAgnAc12s3FhVwBNfmGoNKJ1ejaQ98BsgbGjM93MS09wamq1SAz8G+EnsWn
dBQXsLiHLD6DhSQ9Gpx0CxXE1YiLyDcWslpmJJ55/u0yOlwfPifcsIaQ0OEreW9G
HdNcsigaINV2MU6kQEfdRlyIsh5e04pEwEm6E8Psp/XBgXXDTFedCpVhIWtQZSur
eIgIoW1qHoj0BkgDUAoL70w7Unn575yxGEtYTUz82XWAv0GihQU0tU9kJnjnUE81
jP16y37B2HVUTo4jVwChwQIuGZMk4BVkK78AGPNUopBEWQSaSt5iIqeu8iCDrU8/
Vu1PE2WCxZxXxRDl0uzyQG6g/dpHJl0TknWpXjeS8OrxfDYa4v0GJdQuGT1OClBC
n1SKMA9QiYKW0BDVvKilS5ublDaZnmMaeBDn9LS1zkkpV4gFOAFoDZNtCHXRF1gL
p49KuK2jtg55o+4IhfcsPhKA55UkdXa4XB1inCrzlohRzR5pXCv4g3ZRgUmd8zoh
hyhulh0pWmQKf0L6anT+5MQop/b5XpaK9EN5FZH5/YQajef2WTpX0U4C5QQ9UIv0
ZtyfV7jGsxvwXmARM/3QBo6h+6wuq6cCp/TSaNXYCtKuDaMokvwDjo+7QSVUp0nz
FBQYuFAivquu0e0OgVzNiS6GmHVV1v/lVkdHJo6zY984NPT4ocXF1ozgTLhrkeGm
sqPUBVdF9V1JtE2u2KPXaGmi8Sx4KbJTuvevEMA1MENnQrAl51/fBT8e3uMUvQSe
B70a1G5nE8WuZaz1+lsx/N9goyLTit8PASTgw4680nDPpZ4KtgMc3gar2IshRUBd
hNMhRhA1/CJYgV5D0B+pjW3W9/TKWA1uJwT2KvPUbIxoxOzH3C0TSr5XXxAgTxXT
90QL6xA/eM7o/t6V3bG40DlbpSFYHM5UBp/Z6Di5vKtDA6qwIF61/8ExyA3BTmWG
wW7+3vlC/HeMhSJq3YE/fvUaQH9Gu3y+A0Vyt1/tDynq/bDoPInBsyZy+sD+3d0p
Ci2OdSXu5/cFv+Q5hWey47ssEAJYHlsTpAA2tMm2vYBs8Ks6Nx9duxCw3tVCa3VD
F7ylzZY1gasH7beCWysHePaYK/zTOM8+1gEljsbvtGsaf24N6cltFLDnAWS+QzM7
fMZubwQtve5x1pTvSgkeuAOwKlaaL+wHVTuZ4SnhLePr789PRspN5N4LRjE9UB+i
9A11WGxpR+DRR0kPpQzyezSyIci+Yh4df4DAfb+QggkFk8wPKnPMWUcvjRFcq2Sd
MTyU4dtLngwS4OvqhVqyby1BT/i0EZc9ktXMG8s0Q/bIJV97pjRQq9XW6UMoOI3e
uXmFLTmraGadEEj3pBsqM0cyuZ4ZDMjWU6pBBluGkvIpHuJByRkkN8axbX5NUD8a
kpo/jRYQDpwadeV4rp9C/oBskdVRio165fXyJmrRw/kJxk9EGO1jJ51R2NjAagqx
PlL2zvOzs1F+czRWbQFb+sj25086wYZruSrDHC0t4dmJbsSpsrfq+l6kdL43AlE/
cZIXCyb9kghAOA6TONJmCeEtkbaH50Ts4LBHeoiLDeh2uxZt0atszhSv81Sk/FOG
gG2RFBCINdnlZA802t4FI0dswnzBHpMBOSBQD4hk4RafBhGmNgKbMfKeBBHl0215
uywlPsPtrQSWwROjQwbt1U0TipESxXms+rTz6Ed2HkZUflODOet5SlQ/f9+LmvDZ
09WOGX25tQqweoxdu7Ag5Vy5Hily7fTKHSNtzNNp21XUCj8QVsx2xtxYSYLrce0M
ZOZpl8ZqO9VbYeMaZp3ojsFYKfgK19ikEa40xvbVnVGnwrIPH1NG2Wj7eFipdi7W
rVavV17iTJPKjivNgLRgX+1k3hpfciTrd5xuzTFp2286lqdriLIOZr/4mzJ8gV3i
UoWY6LKcAZ9gfWV5SivhIgdXbGsBDa6MpESuOP4n6NO6eQNKXGXgdih+dYlfpN12
nVNFiF5NrQI1szWNB3rSLicyJ9+P5prGZ1HQ0HWYyNDi0s/HWE3Uq/2AKnI93Vnz
Rsb8HokR/LggVOgTF0Fhnxk4VmW03IoaCVe1V0UW/hamVsFxazt5bmLU49gucnMV
ULrND/02dF1YehmV2jYOFakdImGMFNDrC91AK2lMD/PqClWy3323vsCM81pP5I37
3JmPPgQbXDEM3KWoLuk3C46G73Bo6/bn7YFuJ/eEOd5qPMEroyYIhsR3hIdCA7tK
inlW4Ed0Itu4PaCY0KE6vPZ7yLeWZQqmaBQfleQdFrk4Qh+Em8uNj37Fhfu2Rcil
/ksgG3rNRrVe9m3M08Z6/4q+AKOvf3P8x1EILeLvEJ0sX785Jk5//yXt16W38uo6
MSvoywgs4LFunJo+tWO4y66RXAYOHeOqiAQr5m+LAoS7xoXoCIE2/3xc5LJDttxM
pQQwNrRdIBNMG6954AOuvAUfvSpy4WzDdAG5iSNbjZY6xxMJozvxdh/e4aUurbZd
RfzCnG1kBwcGqaGVJXeESxr0S+KGPizsJ9cXudbZgAKr9Dee6nT2mL6XEyBFSkNz
Nb3tqVfGxrPHrFlHqyc8Zs3McMee9vYLWG9sbZU22/kKrplRF50gvMJLjAgp3U9z
M1FrAa+NswyqV1iihuvV8CgSAni7UHnUaVeXytORNNxsvXvbG5WNpFq9wBx7ro1c
VYUloOLvlK5Qq0GiFsYlk4rrsGJZq7lKDrXuKV9m1K8GkB4Tp9Lf+peXo2BzOhyG
awy/mOvU3WdyYxJwnxIYWkt3cfwKCxXyTdujgivWhP02xRacDvp7FqJeCPhKJSCg
vadkiuk2pvYLhpmz58inO4clLjCqHVwdDOnEdbVfHbMV8v42C0m4m8VKyupZlvso
Vc1Bw6h8iVBYjDP6xqM/8eSdEAPVdkdAwI+yxBsSIRNNfiokj4lFgGVB79qxneAK
O87A5Mcmr7kxnKxqQkIVU3lJYCZPoyHHkTOOGABnwTF+8h9wHsu9mtYAx0Jx4k1r
cK+xEs6bas79NFIvDxQdhxmMUiuKtGuOzuVb90ZBUhjeBlGNOWZ7TsIRYlDq7FCj
Ku0xypvtcubLW9q1bJiu/e1j20tsv68BcMyxXXQzjPIKnSP544A5N4iL52wD1Pgi
wsO9fJVeO6PxmmvVYcmY2iPjLs/ibAmf33JP667tZWxnFGrmNUqLjp1OywvZRL1l
o5ByPjJmSPwahzbYpVd5SxsEZmqfutcy7CRW+qvXomMN4739049rNvFP9lHADCR3
F91q/Ryqhf/LTSOBKqW7SAyIaS0nEp3L829/E5jcXFv3FM1RlOkvzoM84Oa7bln3
26tbgAzuwoCREqY6KSJpL+fNyEPTCAMcMmDMaCeb6g6gtL4rCIPxqZ+gasPR+NxR
hhFhdBKgax/a9crDiRQDGTSZDjlVLztpTKUNKgOsrAX84T0b6ovREk0ODwsa1BdN
pSaPoey0l+pUbfgFOJl5cYO4cHIGq7KDw+HZBGwCeR3ea9frO5AMwuSbdC/OgBUy
2Y9Z7v4UPyz0IpLYHg9KocZDwVyTOrPOlrPDzGmIH2zzEvNjsubnPW0ExXoXqOR3
vn+TAyoLgFpQFrB/XDYRdkje3/t/kFFM40bd8i1XXY2dxE7/NA/emDdXzVSfXtF+
Y+YPav8nwhtIiTcx/dm33qp2r6TcTQVxo00eF9JnTCAZPqywJVo7giCCZqy+Ta4r
MZzdqt1VhoBAfY1GPpwxid2QMtvHwtL++oIV7TZ0M7ExdUUBcYbrDgxYWoePUNI5
VepNtWNvb79TeM+3eQfB3NFVIkGE5TrKCykd1xA0rcZOSqQ6tyxzE17VoUW0QGg6
WqpzHEaJxJov+jKunb96ZbebLhzKnjiGzbADWYj8oXHETxwgCSrWK3evIGYCApP+
L8TPO8SFeY3XGO6k5N/Qrf+l4eABnZABHnhLaanfIVrd1fG4ze+FZdPzwezVugX/
X3mu9mVHBmvflzSoy6gCmuqWuq6uQcrMhFSGU2hyLLD+EN2UqfMgM3i6jhN3dWsN
Ra+uCBX1iFMcISSWT+VhdFMOIUmuNntZFrDj1iAokwMkNVpIBL8EqtSg56ALkNjo
XCrPGQMpwmqZZaoSoEQJI3/Yp/BLGzeV9S1NTPao+hnNMlUo5vZePk7he0iq2CA9
yaY1MKcsrgk2YT/iecKHBtEEYWTItNe93O5p+CWG1FJZHxs5iG9Cq7auYmmyM5Me
7PhWECz51c3TaDEHXBwOU+lNEGx/on/3f9Rh7f91rkrAZh8s+dfUjaL8A4yBAyJl
EbMztHGX8AO60nZYFK2AewsGs6lFiWLnIIbcIfSuKKe8jm1TJLuY5EUd19PQYki1
LbfmdbhfED0Swc6ebUeBZJEmJbrlAJxpUljDO7XVG9MIpGMas9xWswf4i903K1Sr
XDNjjKCLoGyabfxHE5p8yDOqNQaOyPhrZf/fUSQYZufM8NZ/h7acnrin03J5Daqi
ynkHQQduAmPkrZWTdpG8sO3pBKtwQ1VOfvdzvM/fiThZTV2XjTkkBVUxpiWyWzTD
rC+//tWkr/YJeFWztFYUkCHmYlGdidqOhhs095HCQX2wpoZ4EF8nx9O4oCP2Vd6U
5SEFaiuHuyeb55Ca/DpLyZCFlP6kNoDuY1ysi/kXdddtbVBHdKBEDfpJs+F48HnW
WzVk7jT9v0O2a4uwbQPOoirxh7Lj0lMyW5FALrRJWTbo2ur3Hke2616IeqE/uFwU
H5dWfohXltac+mXP0L7612GuWbPg42+lXZaTutB0F/Qn5zxO55cuO6SA9Dh7Cqi2
dZfZCyBPdZXmhPQxcWIrElvDl7Czr238wQNuM+O0Fli3MJOYAzCXjhexq/2QqvOK
+QIJeY91p3SMmciDe/8+eFQvH6ROAE9Dzv07Y+Ed8q+mW8klPTHKU239WGrJyO9p
VyjBXWpjPDkHMBRrofU00BqzOJqEvJmOzsUiF91QGYIgMTQw60DiJ142kuqYhURv
pzBmVWzgkSWMcouw/Zr0TiGbX4Y6XOWUNZkJZdzNBLh8JbDoSDIP/VsRigo5Vhe/
MlpPiMfhpYyKvejsQuBAED0gi3BebiwcnCPoRyinoFs+nRpH2RHaIn2gtb0ALL3y
S3x/XqgAx9YIAztEdSJ/Pk6LImTrRBhk2Ae1/0qzrlwLUWlzorszf5awhF/ey+/G
ORdpFV8i4MLYJCeAZ7KIRMP38FjcWeK46LRK6YplpFxcmYD0pbngnM5aMZ25Zwzk
j4STmRxPW+dN1V9QhPlabdIlVOPdtNF3ShVE4MSbABe5/A8e2k5SQyoBVb1Yokxh
kOz2am64aa6j1rmbXcgdspm4OCKTPrsj6TdU3NaeaOHb4EJblS50edSiDt8hHIuJ
AGpW+6fSJckpFmWPrHJbKotVCr9zgkL5VjVLEEPmHmcTWCa8yCwc0+iRkRRN6wq3
Nm+CkJk+Vd2AUn1CEALP9/nJvCwkRRbFRX63EYwA7TPtHO3chcJgZAlfAmPWL1MG
aIhLJkYdpb7RsfVtplzZmQ6t1NK01tnHeW0FGFcoF4kJVUYiOmMertWF9COdznua
Cll2AC0ZNZQbdAYVF8Ln1tvXHxo7743Z3+FAXb1Em2w/bEgx0e4GYC/LdYzwJ5Up
nwtJCqWCOaCUnL2elzjtmK/yj57R/4dHbcBsk72v2MEiOxPdgubZ1ItLY9g5Hm8T
j07PulAI6muj29CFhuKQ7gFZuDZ7klQcDHs3b5eYkOyxTliy5omlfWrvKrXUldLv
XKISttlq84qwYS6YZW0KuTokcuQSJkuBDKTVGejZIy9hx6HqO+MBOb9ltbD3ah3t
slGZ2VKmY8tT/q6LHC/29P0e7/p32CVvXl0MHEtO4eHJUJ/hC8yJkVq8MJZahDye
K9dJ22NxFQX8gKnAhY5Oku8X0g0ZS7dIufxIAfzDth3eQyzT5QO9ujS4zg6xOIee
OlHup3539YNNod+IsPluMo4USrDrXdb4cud9V2wnFwJb/Do+k39lfWHcRvTHFqpr
093Xrrco8sT9C0tU89GktlR7+KJOK03RFhCXzy4toNR7Cr0KtrpPf1/GHza5njcW
9nSa1SbH+cQredkauKyGPJcFD4fcvdxUJkdISaY1bbCET3Phd3GhADYg7BGLhq2e
kpXJ099O0qBAdT0bF9AJ8jG1SG25RMkrnWPVSogPE/ZWffGdeDTSzajUVhg+yZff
lSv8dcJkWCThrQr8XF16wMhA7gIDtFTLWTvxagH+cjry/f0s+ivm5Xqr1475a2EU
J1UheqVe0x/zAWIMinrb+xCtaBoOR1ljanwdOHjUTWXCkOCcz2U5e715K1XPgT1u
9LASU7PqFnJBWkGTkacRcfUP3cVOW92/zYlpfuH442r4tllBIPy3+QUtpHajnlu2
boE/GnSzSO3bn8Zf0b+XUhmIFrypOQADixfIK8ZRsbIsVl7DeJpG6ZJuKAfOhHeJ
K1x61ewkYa6MwgVaZpzlpPt/8zAOl7sS3Ov3bZ012z/Vh0ETuvo++EbIxI9XA3fN
7AfH9V3oz/WeUDxgfom8DsiqkmmOv1JnVJ+tnFzc5oHWGmld0TuE6aEpZCtZtDem
qjjTnFjwtsPU28/LA3derjMzhFOWscajZg5Obp8Wc9Ux1/HaK04qPGqSKM4bz+fV
oD6bzCcPXvZVBRwx0js3rETvSyhrUJOMptuTVcgtVwUaQPiOkkEfphtdBenUEKlE
fU647NqTDzFXk4S+z67HFxa7+hu4WBgO0PG3/Yef9l5ZjIwY6MiP+aczbcvQNaF4
DMakE4/25d2Cqdzjfeq9cESY9sBclo5ILNNk4ig2QI+qjryklLRYQZsBam5ySqFz
FouJowmH5ZC8fUssQ6BwuoVMOSaR7sgcFIfKet1VmNU9z3d1aC6ZVvDwOuP02pUi
TBg2qNZ8w5IxoLn+srP1kQsBTWggYLOmNiFFUNJfUTm5j3PXVkWzvDpG+QYk8ZE4
WQQHlhH/bYW9f2XjqvzkappwZPjpqW9GQWLT3h2Ar8sVRelAf1ez+6YfZWeLc5+V
iFiL81uMCg+lZqbzIc5+XjvTNDq/XQZ+0z3yt/Si0jZXaj+VfSuMztgX5Qv26sek
BfjTOqSdPyxh9NU5476QXZ1SFuwQz6bs3ZpQh2SYawdBp1mOaa8bhuL/mlNOlwAR
ZOAcgiPilILe3IlzdKN66YL4BETvStnxv5RHZdZF+aRx06O6LlTocfWXCRnMBnbP
0uKJtI5Rm/LA115TsN1QEOoLKyfo98ZrBjKMT6ViRrS3SlhVxFDlyCwvJYVB2vfo
+94fhrJ0U4w+62Xo8F14/xvJbP5i1bFMrw967DYg3/ye1JEcoWoJSyPjAxwvJxhB
zKlQrymEv0qJYcv7lCUh2yYambSyAXsR/Zhuk1TiTDBAKj6X3XO3SLBjBXClJ0Pr
qg8KwlZak3QAiLHIpOQPjCMtIipKMSAuGwZH3G0AwE3wtb8+M6e1XKjHaZyToB/k
AWvmZlnFvqSqQwSb7Y6Aq3hAKAttSfnwe2CS2YRD2UUQxzQPZaXruZqv48SIuFVi
C3rb9GnmeuIZidZs6bTUHOzB3BkMoNOLKyZx95Uh+QnGxYzntG97Cwx+tCy8Wzl/
R4WPEABd4xDKnIG2yNCL2bqZVNlfQac/8+hry+B63PhM9WNKDaT9ELkKgtFqFlLd
+7QUYl2wqKcXiEUp1TDcycPOYyrRs37rjGQg61/QmL/E8EM+uuwQUkkpwzpwwJLE
RWudT1UQY+wy1M3bWOxsHZOqGTTLXDbLVsF0TqL8AY2R1w+1yb/YJJzqFaoX/OA8
VHbR6uJgxt5O+ST3m2bBmChbsX/yNyeQbUJ2XdR1pvSwOlYnWHVW2unJBOOXB2d+
MpubVZLvBN9KJC29uRiDufYmrP6o/sEfDF8zV1nHPj8OjSjtnO0d6VkAuRDhAUed
hrX2KN80nvhCx/hL9V0LggMIHAArhnBGra3vxS/JswG2JN6Pp8BK3/hDIv7DWReq
Afkjf03ybLqn1zUbEqjINDhlQXQ6+t0c0u0Zw4I0WYnB/zkipcUszDGqM8uCe614
AklWTr8tmOhefWJO8lcH+0d3rMbDdt6u+yFe0CfzJkcCjQkCla9KMwSVFmkv5L0b
qgi8IhU6r2B49H6S3zGGWBWdV5O7mlywAInxazcWU87Lvrkw9LSuQxppoTun7x8l
eeGIyBXygCWrrcZYmDF/Y9Dj6U4YYkVGkFYrHiHnJAxP7bmPgWgcOwXMs65r6zsw
NFkjIy75JPLXDWMxpRvpKRre0rQXgErRJZrk2t4RmThrPuUFrTRMyWWXbDkKS+GG
vxxORjjH33Vp6ZOtQeX4xTsD31giFIQfJNuUO1uQ6/f+XCV0/47WaIlhVQF2MiAL
/XXHtASkKWNfZcdRE6z7j04lAg+/4sNTcP0gohRlGVi4eyUnmvDoPDPA+/2Pn3/z
N5smfIWfObCPASqHqPLH1dl6EGqlW7GhN/ux/zpd6hZT0qY+CHvjrDDv3wzqtA7j
gT+qEgKrCsZWgQAHOHxpXk0kF1kLvrxbGmKNuvdSMDLMAMO8XfmRY+VhyzQSm24N
3nKL5/TRzXyah3FPl0IH7vncrCrNvVrqdcal+nG0UW8WrzPCNjBd5jXA2PQk55Hk
pwQoQWGDgVC1D1M3uZ+CMw4EupKhb4gSomSNP6UovYMwnuVACbk8zDqnr6wkcdl7
lY4JbcTkcs4qTrscLfe+ZQY5NvPkJa9y1B7GhFllHHEnwATDbHX2inhVr3SnCz4+
yPpNTW75YAu7Z8fHTmHM7OJhCHpOcA0WN8chLuiDHB7vBVa6DDABiKFM6i960/nn
9z5L11uZAoqJQMQQDpioBRCvGS1Uv02iOlhTpJwu/joWZOU7dGQGRcN01s8A8yZo
L+L0QK3oGEa6EAFompGvTR2QdPH+YakUAdoabBgdVDXXVovQwPmCWOqFDkgj60YB
3/QhELqJ10aYsu7UTB4/RBpKOmMMDqNFeVT3xjduEXlSXozEWMCg2Ggr8uZScuOn
WyqTMRz8dgZKeXTlafQfcTadg1G59zJTLgqets3z/ykXIRWvSyfSWt+ePMr8S/IC
F+FiM0e5oiG4MLAfss9MgrDHivGTUQQF8m0EOu2gSowjtQA+HwiPfeFiJDBX3Pak
Tmqq+yd3+cxJRnKynxdjomhqKkoguh4TSNcBcou2e64K7c8uyogu88EORFWkUFZ2
bWw8z9I80MPHc/tz+cgBPfG7IhVLzUviOKl+IT6TGpzJoLdhZOvFdU6//hqTZJ7I
sMmHi7eh3iHza1gg++Dwx2/5PnG3mX1VGq4yk2DM4t7Ixyfhi/lo0lMSU3qS8mVr
s/duWm+ve1PUVZiO1PZFgIAONEShOjXPYc7wOrVDL/nUcHl/nKwgFBy+f2D+RzTz
ItMzmXw0/ReXRAWMNA6NTtNtvDxuBOpo9xEXcCrs31/f9T6rmbcy/4zCEwmhEpig
40i7JLV6s79/MVxye8y3nEPX9UTtvxRlFP4aOLo+VuHuMOgDfT1pRl89q87pDGfi
njSpH/pDpjgSLtxm8BhtP/y21Y06qOWpz/qdzYfTRtlsTwp2YeNNyOF8NzPqwfrt
TXQZCqbu1+BiASesjgMV0GtsMyQUwql3JYOKLmiU9sIqk/+C8apz0uqaSlGKyFNc
CG9p10wTMpf9nMnxvt2JBmE9XxvpxT8UVyuZYxsxvYijMjfWO0K4LE7s0E8CbAbe
TpTASY81yBhB5fcRSNzIj7a4FzKZIZQGQ+Bces52vH7a6exsDJ5BMyk3v14IvVtI
tedJh4h+kAWKWm9KI+4520PMIL+rnxhobq70tzn65uh7Okrqt80mHT7UuPDbxPO9
nrK/qo5p5TI6bQn6plCrPcKfKQy6REFmpd7k4QVmX0KXUb2HyTBIUvcJbbh1bHx7
/4LngduCY5hVcSIseCDdgK+JulS0PEzesGDpaIn7KuGd+o/PDBMZyBjoB0+cCKxT
pEBcp2nNCXZ6cmi1xaFmA7CtQSIQAmfXMUP5QReGfH2WBXLMp9GIS98hj8351WoW
XUYw+LtwgEBxjBoumZ9qXXO7zx7JjTjst57YIU3vBPa1BlDqdNjaoerhN3c3+JNk
D66ZRa+9WMRGV66wnZoGUiutACGoraD+BRIqVxYBS+r8jsy+VfavQD29yNaTrGkx
w3CjpjXQLKMpuZkqahn78pxGlrnvGzfdSf1mtYDOEJiRGS0VR4MuQV2FlbkCiDCT
znlHzuBWSms9yOZeNaF0dZ/CClXI+AaygVMtmSOIiD/gm+BgCsH20XtEehBM80fQ
RI3ezkJ0lCnwveDQJTGjy+XxjjClTG5avEn30DuCuCY+Dh3jfwnylzLV9vEq/gn9
XPFydVdlvAYEMvXAY5o0FlrSCqZEAit7on+xUsAIYpsqDgGbcV7q3vvuiE9QdGx0
bP3VEZXrVihCoIi5I4EJ8J405lYyU6SYj2WoTnOMeJowZxPx0mE09RARYdzEAWvd
tHprdro0cMBhFOk5SpDhblaCWl48zYeiQMeThJTtBxJx+TEP51grvLjRqHg0qFC8
zPfpwGWM+NHRfN13FI+wLQcbC6/O/4RN974HOJakgB1HDxrezx/dLfbYKjS1yVmI
O+/y6PLuVeq2+OaJQbZ+5XF8gfMU51vjHP/H5FbOA28u2eow90me3QbkT6QZI9oV
eVm2u9x8rKlI3aJ/sNYH+0jiTZ8YoQUWIr+Bj/UO+fn4ENnGUHw9ZLUmHfhSsiRt
P7Tk3ASav02lTX9RH3Y9l59vORtIc5BxLM+lg/3/upN6nJbc8egOXC4a45IiW4tt
Z/c2bla81iJIs65uHlwqI7uNhMYd4Oe5zqZGZA5j40koyj5kXrAUNT8af/vrv8Dg
9PZErzDrLSyWM0lYRZxA2NBuDpocyPKpadhxFjFyZmo19lUO2TQkz06D81pANqQm
Jdu9X6mTBi74OpoVOm18KuqYiiivfdiOGibTkYqphe+qlIuZrffCa/Rgkj9vj5M9
233vAsRkrCqolXyZ/KJGH0/1JR3RcjVE3y0aWpNWYopg7nAGBIVF3a1km3nsZgXr
WoUZXmLdlUqGHGyAWS+N1rMywSUAYkp2dXgyb+xQktEYltswBdlZh23vWJ4m6WmX
QL479wfWKMjK7PLryMnbLIkTnhOJseXJ9OUQCAF8HkGLZW0+ebPsoCXIrU5bfpKW
Fwzr+M+hMCo/cB31zM/0Pqqy2wIZHQ3Qklclr3sJnL1ZedhyhUDHlRJN88lHxNRJ
JmR7QxWgZK2ANw/bK7Kv5mdD5u/7w3GbmT91hbkisTYEceVgMx13267EKqkABd5W
eRRMhjBF8yONMTjWLtc/NAsYnKlLj74HKwFrVXLov1L3OT26OthHajkhdeyPrOOA
Zi5gGwfZ4eDByT3M/DPML+PwfxoNioABSHmcymsud1NsLC9GAkzg3C1AXmyOYX32
G1v0F5DDdGJ5ZIjfZHreGVfv3p9RgBpPCnzm3D2jm/qo0yc7HGnAqfz5qsj9TVkI
oWavzlkWHyPz5GGUlm0Zb85rN8j5FHrmpwGKP8UUowSjETGqo/V/U7TuSeD7LKMH
V06C+6XJZ2PZokvsaiI9BRII2BIK/FiDwynVkYDDGm4DmUdZsiie8IUdLX08/2vp
V1MHWXC1GVofW+/mJpAjM+f1W8/yHyk4MEhEXyEbW3Ug+Ivgn/7+qGQybmYdLAw6
DSFfsW1Dzjltcx+WrLgbKeqWJpU8u+GI/BvM0AlKn/wZTBkEqLjqKbGS5rR15jKX
tJq4Ycyf1ljRCWaAkrdDNJIF3NyQXoI16IVsWMmxLMAa8F58U1Qmek7RbPcNWs5a
+gbj47DsiX7R9gw1JW0s9Gwrgh0iEeG1Hz7AWCHUTjYwgUDaWpGsKaXyLoERh9Pl
86hNySgWQlN5uNmtPHrpSDFMzXZxEgDZquA1+FQnGZoKwT3HtYVLSucsF8T24G42
XdlZbIz20eYMrYCX+vClvtP7V/oF3loh7pZa3b06BdHULO791b9KopuBZad6NccQ
dOm75BNuzApkCgYlyMJMtgsMJixTLtON4DdhsW18CJFC/GhllSaRzKq7HbfCyaos
EktJ5C9KevRArhm90i4EiurhCN1PNC+iYhcF8XcN6Li7GCGnRliezhx1olXG4Fr1
WQe37MgSoKgRagHmDWBXvoS8F6Pxp5JXkyU5ZW0R0h/kSHpd9sh1M4P4UYt0N3LJ
dlYdVkvU6Za2oZoVeHiXUxq9XhaZoCG3BcJZXQWiXjnxdoc1X9nxepyyHwwJRqpa
Z6Y31GNwl6n9WpZekFqJ9qfaRILuNnpzHDYDgXLqoIIHdQFByvEy11P2AcnBijr/
dnlvaj2+nFacI0diU3vU5CanVl9dLF0J7uzFbdgQeLuR3suFkKLIDD/k77+kc4bL
poZfu63JlbLQo6g/lWhO1KtAIAwG1dP1JevZiajWmrsy2XYY7NDkkye0Q2t2Qium
+Q+skmRT5sOLvxQVa54WG6kEWpX5VvWyltJ14QYjxTl4XNka4mSoi+fcaTft8vva
74ADb6FYRGJ7A+EeqEsrzd0bE/I3LVRsxqbarE3M+SWkWcxF0U1CUAwxuxVo1CzM
IFxdA7hdX2+zEFm2yICe2byfx8Mp0TIyqS/YOSkF0tSJz3ppsEszEbAD6XMc/LaU
cboUpBaY0gf3czCTLeJec2SXO+ii7+h5OvuxjtCqeEAW26i+tUYr+3gwFUbfzxrn
tmFOUomqNploxiIJv/HyQqUYy2NzuHPbIi22Yb7x08nyeVbQjS+tnufekpOaL8Sw
BGaBXcyVxNyJvJTT9eD9N1LnONgO6V7IrQnZ/GT/Sollq4Pbnha2B9bC4m0po1Gv
2UdM5HT2IlMbpVJflSXOzkcdrtHPreJotgJ1xhiSquhnAuTMoHhcWfF6MkGTpW6A
29NcnaOcKppjqxXv3ioxY9FukQQOp2Agt89Fz7e72/qYuLmlZWpJUrsfLwt8Mt3a
O7iRlfgRO8fS3OBZUBeRToBHOwcxahDqWTYHRuk1urmwnWb2fbepeOfzMPM5Y3Ur
79cRs/D4oyz5r97rmqbqLRFIAwleCZOTUiF1bydGndbK26kneFrQggy0gUBz36Am
OWFiCGbGQXVi/SaQBdcIi6vaFQrvaozbZ7vPKFmAMBGTanILuV7jn6Nc6A7NrTWS
3+jVrL9yKQR8XRWFZea6Y2aIuA58DobkM38Y10mEHZaryQ7CjWwyYPJcSOycOVGJ
DINf1ZpqEbBUwdvpBA+v7jOZQftEYmICIAq9iH6l0fDp2tc7MPj3O5fGvse/MeLH
SYQQXe8PRMPTLkoU5kBSt0txc9EMeRHUTSsBOBBc32Kr3a3j1k7D7EwRkRSSBuQJ
jbTyZ/diU7wECl+bG9ZodIMpUrHkeanMOodE45krVGvLYA9bH4+xKU68BHVRizDc
AY4Az0CjIM+e6Xo62ALU9QaoGyZvIwx3TkBVTUrSDf/EdTdiLJ9JPVQKFXHTQjxK
yGAW+InEyKWuRiRNXifQ4Ft1g09Q4rmKeEfw0Nv8CFeu+CSDqSY6OgwoF/RkjnPr
hHIcBeO5wA4QJTJzDc/h89I2n0M14H/UJIE+IpkXMsrpQ/UPZuh/WF6gplsA6Bpd
+nITJx2OND8i8nBnMOrzJJNa+WnQ6xTYgK4FBRjgSMQT83YjVAuh1P6HXm4H9IJX
8v0kICLErIATMnodNsbRsLoiAfnmoIGTebXuErQJS6IOC+01mOJo5lStrBEQuYDc
dlhmjSMXhf2uhSKwEPYc23onNPLwrvXIKj+mphef//59xqF4i3UzVFikAiPifLiv
86rIo/EfSTSIExZ58J0vW+vCflzlRlHC/zr0VH2OJa8V0pUusWVbtH1Ju0lV4IXb
tvFPvUw+3pk4htp4wniV8jsQ++JA/trBJloBm/KXrU+7NhgO3pKBFAFdh3WSJply
PJiBmT+D0XR2zozZ4ujiYQCQLZvSr6SQ6I66Z5iuvIId7p5n3ALSFC7DbYHtX81K
CFzRfgFywjzCafQ2PXd1JQBT6rFKfDzmIOVP1Dd5ils9EZPqrihVqweaotZZ1OjM
+8KxMbV5lb8gP0dYQ+7JPeYACdPnGGPqN5j3mlzGedUg6OpLbje662LyJdFNPM6a
9MaxZJHzsec6xKuqYvJl/d0gKfvQa0yzZr6BEkCn8hmXVkKjE+DimlJJfG0KlaPV
ARATIPLmFaHKrWvJj3P3GLVl+EtdtHJhRKczOYumdvuEKH5QRrFv4x7OeaTTKUuU
dTEPvlZ6WWlVZLo81A+1gV24FhJwv5F3Hj3UxCwbjGavh+QA/5ysTP04RQuSGSvX
WAVcoD2izLsXr5kncAJZ0PH8plrG6pZHgyLGq0cyQaXn4t2wTWGPARoW3dUPOzLy
m5D1sjRQFpU6LxSJiVDZFGvAOTnW4EAgZH7w3YBvNGk8oQwdtCr48/opJmXhD9/t
zB6MIAF3B+nHabwX49EuLskBGN7Voi7ZhCZq2T+p5fs99zhK3RAfq1ScxOCeX1hR
PogGH3GMBUYrMT+HNPa4XQAvhsiJcYH15Mvddgdy74akVDeQkJf2NSuXhn0H4lFk
wW24UHRqsyS36hjnAhA1L00A7wCq4BKP2MD7m4oCnA25sgmpv+OHZp6FB11ii8IY
S2AhjqeEwRkn1WIB4z8FFzNaQdIJLtgYFf2UC9Blm3hZiv85XMc9jWala2nbNuq0
UXb1b7zcAkuL2YOnZ6uvGkzVtNcj8eUYfH1lK5EFNiGg9WiU4QJ3SytLfwOSS+LM
j/CJFowp1ltSvpqnUolpEwYnf4UeOav5wIZUZ+/1a0vd4afAeYDloz42QNSQyvj5
f+cQuf9ntVhTpauRrqUSIHX6s18sk7RH5VSQPJcTjPDLmo7xYpvzA48Bic3kGVVo
NUNVJVp1SMWCc8viAUqvDOcWJHy3mhcgbGQ+71X1D0z4OQcwwDx1avUATRf1ZF9A
EZ8EYSi/7yL3iKNm2Q86cpcmc51oKMRKn4Zj7uuI6VuupE/KwlowDcB8f565uKNV
kvElzgUpTTdV7YrzNZ1wmk+JFYpbnfHk9Gs5arCGR9LDhDGZ6BGpHCQXjFfVHGUB
y5iIP1qJLat5PxxqFZkwxfVWKGmhuHvL8wTeCAEv0UC9fQ8DRJaP0X2nLzBEIVkt
37yb/gf0fk6TZadJP9fFlRu2aKgQ3C/z3Ib+LejAPmQuTPEcFubB2putqiYqa7Cz
31f/ToPTKxy/s0E+RP0jFJQAUB7CSnTWbBG7SFjTo2ZLN1vxdo5VY7SWu8F0M+pc
d7JP2SEPdmi73rUmOvDDr4k+TJ/nWt49plasr8z3kWDr6ydnfv+ONUT8+i/DFrMH
MV802x6DYUYXQOmIY5ZBucLIzj7rG3+6YAGYAzrAscKnd1vYxGh3sZijsb3fCr/O
BsQikc5O4xBP+PqE/2IQ/+sbwXMk3lAhgxrvZ7ahGfbTOhrILz+DZvd8vjoHH21H
c3ZzcN3Me2pvAV4MXlN4CbfPFuADmsUoCWbZN696UbTA1J8qbTrJDg8de+no3PiU
bh6tOwmOzes/F1J6BzWtija9z0qa/Xc8f9C2j5AeXQgKXQEco9aoZL29brLm5zLs
QnPSPsWRspNYxI15E1LdBE6G/nFZKyte+TDOTZeGlnKA7pXIY8eQTttjzaR4NeRk
wy+2KiObAEwoixrW4nXgErl0yfyr1fY6g7tZNz1pA2DPxaWdU/7OoOluoqe9cytG
INgYmSOsAjqutHVDzXwQETpkmgMNLt7SYOArYiDAyTy5yXhKQgHO8bwZzTe8rwFS
j7j8uuchvsNUJO32V0ZgfN4QcAR57BeFIAScJ6vIHa8GTSpWcZTIFLqIvP4N2DU9
+KTu94uA9VXCQmp8y0gZg9V5nW8NCJQTygq3+yp1/mhumX0RdBfAI0Pu2k/aWWvs
Q/AFsiDYPlHUlLt8WSdDyEhTPnz04vScY/uh4oh14/J98Ni7+WiSyKVbs9p77pmJ
mWuF9Bc+kGbhwzjiwP2w//ePIFPoalx1G3N/EXDtIEjNjx4vbdIi/3bv3zKRS8aQ
ie/1fUZNc4OJkOfoJrU6wd9nzbNYl2fhe+fV4iw3YEHD/+k389MX1q/3cNeaddn4
/29KNegpTi56r/CX+uhz8BiDuZDfhFTAVVcTEqrKJ2ZXHW7X4AhDEGUxoLE8aEWD
Kbj/OfW7HFX337j5mBWpEXmVqd0I5THOmQNh3Zfqfbu32n8yyZXA49zdCGkTrMQ1
Fbd8ZT/Z8cEMHZjbSYKeAaTllwgOeqQKwIz+lZAhV9/6VJTM8Dvh9gffbAgvtNLK
K7JOuOAeuBfrMQla/LJ2Tymiz/MxE3+wdUfuwlSCtBbhIU1Af46/UhSKogGesGRK
TT79yVj6XnWoCPpajV2MWkgtW5ylGdzP1BycShX02dYtA/AgIyXaV65Dnc2vLeUu
rCq2fvl0faeHyzviRMOYTktkUmk7iLvTg+ZDDm85ENBdICY2txq1vk6yDlW896WS
/RwAURZPFLpP6v0aVySXoy7oq8DNa1WKNi3zN4pqEvO7dOUS0417oCMUnZiTpvDh
XjSI1A/Y7OI7SWcUsWEBqLgflWn057fzA4SzL1doIaWR45q6WmDul0GD1fflSPqa
ykWTKdibwEQk97e4isOTuxvl6sBFP3quiRRYURGFq833e5rrAWl5YZn/GZlt6G7m
iEQe4sFsJrheXcZLuepps5FarWtjIOYoHIerE0FStOzJliWw6VqqaADbT1ho8w1f
M2MeNeokYm475LK5RXIJDeSNC06/psyK4dssY4UHOm//p4ZYCIXMRJG+jle6ULDT
bOqldFL4SE7maML2y6O5rb36JUSnYCkrUWZnRTvdiSv9MuWez6O3BAYBIQ9bjzl9
vLX8nkJ2jGkaIB7L9BiXuUlOT9+KCo6p0YUDpPxkby6HMLqtUTXO9Qs7259cphy8
sLJJzuykEXzWqKTCKvAhcE/cmYJYbGTw61u1fqa3p4s5DerAN3BXbdys266f3a4j
Dux63c0bNK17cKyqpWDcah2xKTs/jzfMjyhh3Yx0fkcPfN+5krfAueyBRGOv9qcF
vAoFMEGrEm6a0z9Gxpw9tUEacXLcgfCdkH5o4sQYYMbQPlq8MSbIhpy1JP+w5l1f
jxd/IN0p6Qzl2okTQ9IqEU9Swy5eItwVEq7HOTLx/PIUh7A2rMKHWHRmrHlzMGW+
lDrguyNnvSX8mXzasP/qNC6dUNPQn9bW52PE6MN2+zf44J13S7SJ2fnP0d3yyPmA
029kzMky297R/qVOeEFRZHuDYW9SQMcx4jZkuB9OLXpzz8QYgRCwuBPSkaQHNlM/
Veb7vBnZ+w6WoV9cMq2r9aI8wrZtqKrI65X4iYZT18kxilKazV9Zn4naCtVT2jLt
QoPMl99k+YmppxfXwtceB0cjsetd+S6NJoiRrfUHA4jewxsn6/b9+mr1GOcTDal4
9GdzBlB2L/7sQEyd6tK+F7OFTFO1WIj7KdehHgrdsFAo25YgAOKDPLu3dnagxULN
PKnq4n0+odOBqKfRH7flgOpOBaSZqwRakwe1BOOmv8z7vMCenuKU5mYtwgLj89Xw
oMtRr6yWLu510mkLG29w+XUlvxK+UAiyp1aw3Iu5EAmZpYyjskQz7SNd23gMinLu
GCdrYWdlC9SLvJHId/NfFCW73PxWPiVBDDoj3/ADfsEZ7tHSy2YNSnC5KLSQlOS4
9I54WH4FYZooud5/fVXdyeOZiJZurek2E2US2xndlv4LdJWgraHnSnVUwU7INzrL
2kcx0lIg/52yQMz4EObdoMbeFk+3Tkg8tDF+tbyo6WBep1cN96lFk0yXK+8tDp8x
rHag5iqOv/p9N5dwPU/dLtt1k5w6S+iZQspeR++4+u3NuR95BRdJ24SS4IiRcw8o
y6V59KEnzgb2uus3xsjTuC7pbxZ7XW0pNAYwqEBwm4O5wkkplxbjzyjmgu3m3MMP
dd7iTjPc7yJaAwIVYi4fhz/YSRYdvbso6u7yDlgDf1alu5strXXq0Wsa1buPu01K
DXAqKQuADbSRQLTBzyUVyuoZuVGbonmQ9mEyRmnfS+3bWX9GuCkLMmYuJl8IYkQ+
kanFKRmGCTmkCR1/fT44f1CtO5tfJ2I+uc3ekwU7oDhvDO6o+hPXtEKGpj6C8CBy
X453KnyoNiqbpHYiScrl0m054pO+cy9YJ5S5cKa9pkwthZuUtn7hJQ9oIGtX7vq8
2fMqSV+Inz0PfpXNoz5bIR4vmyNR5TpPZSVdGdKcWlELZibflzSIOYBRHY+D6CqM
kRXiNSNqqshT0goqU5+j+enPoudjqozf5lyiaVUkziZ6T12o/Z3BOfwWSLc16R9e
Falh1x8TRFWvyb77AYzHuDAzRCkmhjcCuPVAtUzQi3pJYFARNEfBH4A7/2q2YYH+
uFD0VDhUBEm8sPEBDTM/W2wlChU+VG0N/wjNPH03ZqGJaMyKu/5rozMF4PwEDy+b
3/YrEm++RviLNBniY9kv/sq5Sq4BjuX57E7YTgUeddvuzgn5WOdxSHuBn0ebDHZH
WGakLr8wlHYXbw55bHi6kmL32KwWkjfETZOV8QOazPvLcrbM92J1bAI3drP4B9Nw
qrZ6w4WDkvtnIn+8kTmQPk62TvtBL2wOHbQlxecfMtxD9mle4201lgoIc+Pr+naH
RbOl2RWl1AQqLkWW3JG/KcuTncakHwbnoQAcQDt7VEsS5QVZ+wn9/6CChrnUd6UZ
Wu5AMAcKyCZrYo73Ph4olpQXbhvmJIWvq1TS6rg/hNQgQZ1i8Y8FuB6PALtPYW4d
s8sMKYYhrm5xMFau2txCpdn2Wj6IHtrc25zudf5w2OQCx3fX+eewoNCp9BJTDp80
u7mNpTZcoUtlTY/we4n59xN9RKSCbIHqo+df0O9nKxUpqvag0gnZFOcGo9fpIwLn
k7EKBhFk6Rj25hPR7E1/zxczdC60Bv9QM5ffmaY0UOwKk2u7WHWc19azqXgFD3I3
8uuCW+QWYVBgatRPJUJBaxH4j3LGcC2Zw1GBXuQbfqt1b7Pp7ic1bJI+7AIZ9IOq
XQH6UmdtiaIzM8pc5fwx5V7zaLDOUpp8eV/kSnVbrlnpb7rUl+EqZZna2kC7MtO4
EwNMNN4RfQYzRhXQaPM6R4KGnKh6GMztJCyf4vY2ig/X5NC9/Otr7oeZwVLSqJo3
JiVajggDphdhaunxf+RxMegPLUvU2GrXzLFATPkXluf+q9PQeNTr1HJ64ZAGZyQk
AFJSL3M/IeY9sM2FcxKEoQl4T8a5I716JTEp5JF5V5jgbPEp3+1x6z8PHe58dZuR
PTLZ+cZqPrUrGdNZf2WFNN21+lq7igKqRVn7YgRjTL5i9WZsqZMJjnKbGyv+Ec0d
7mvFmKD0m+duCoGltAXau8UFIVWqeKVR9syBCpd0DaJsZSBu7HuihyH2Bx/o07Q7
gv7Z/bIx2PjJkvB1y/YmDeNhy2XlfdlxFxt9qPGCf+dc6IFznVl4Ba4CBCfGs9+5
X12R1B7lpXHJ8GGRrrAIGK6Z6Y96nkQUKwtJqJQwVVweCJkbPM8NmxsW1ef+PKQr
yfviR7NQy7dUgFo9jdXul5mla3ciLR54EX9I0Ja4dX+4PsvsE55i1qb4N9MIoDaD
KW2iQD2dPFW+jsQkHQ5WNwBblBXajRo4SjL+S51unUvESrJVrWQ9VbjYt5AcBHv+
9VNgOdjBZ+YagI+gQbqnKCSSgevMgyo1C+0aPdS1hb86Del+aTQlxrW6XrsgEZ9j
wdKUyp3oXQzk/dSy3AS9WPLGLh6J04i/IYd0NyiLM5JpnDc/CbbBO9ykMuwYj8WA
Yk0UmNQK0czBVLhBhcH/VWiEfUt9jToGb08XH6iqPsIBbvYCbgdAKvaJdYfdBWXO
LQRzR98Vy7tgR5RxoFyLbdYfc4DJx3jWuY+CjFdqVxXSBjgxANbvfAGNQeN8Dfme
1EckjhtIc63wd6pUiXLAKGCSWpMZHCCybP0gZ9RmhToPWe5DBbZn1qKip1EtipLD
8ghMXVRug5buSqVwla6ctqa55Fe2X8AhxqP/Iat7eXhJASRbzn93PH/23TxyVPeO
MpKyr8ZI7mAQsG5m7BJtOZFTlMZSfvSKSOW9lpP22tF85DtH7E04YPkdfJDUMFj8
8h+yz2D18oLZcyzusJmtjICBaLj27VUbHn09bwDm+xlW0y+5jwYiMNU91NxreGEQ
ewsGMtQh6aptYmWAqM3Cr9NXL6fvtbii0YRoMxKRGo5wx78WEOQFo6ZniBKC78Uc
zkYSlflk4on8FUKR0Me3EdJb1V/rCcNysRKlv1TS4YZ4H9SsZ1BipCmuMR9FmKhZ
Hbf/NCRqE5nqLAyZlhf5Zr3bB/YHYLuVIAah3DY4TOOwaVKm1bLi6RVKj2lTVkO0
I3I2dUZ3ICh3NZAjpvcsUqXuIn5Xh+7Mrenbv0qiKnUDNjVJHHZy11n/9M1nW49Y
HO4xgAdWfXH2AyBzg3mauxgJcGKFsRNsSbVCzXdGu4xc4Fi+3wtuAoki2KVUZqGi
/DKtdKKT1ghi63j18GGf3tXA64aHcYUnBgggu4HSK5CTUYBEfOPEcfxJYXz6jNBw
PbXeBltGPNyzy8OUqoVxAsi9rSwXl29lnYPRHxb2pIYcLJ5AQnCJlBeu12WClCgF
dg2DaeSasNjLdMbVwQZRI+j66Nco5DqP19A60PvJ7f9v1t/Ubnuit5J4j9dMAFXO
RR3E3QCHFEUmT4Xkz1WQcIl3vlw9t8uUNAU415LDcoide0P7QoS+9oWHdV0UfNJ7
pJ503aIXK0O15bC7bo/PjYykML39W/N3QMbWUjxTk9t+jhhbdDaQwqX3LHYGxnEg
2KQTJv5dBgcoi2H0feQUO5wvgs9cENiM4dOJ4/uxKyTqwJcxfRtRtziOveG4XEqm
RX1E9+bRMcV4mlrdm8OLkv/qDKF90KCwMtYlbMHU8xmw+cJIDEoBI3aPHg/tp/zt
1SpTYLe1lMuAwrRyEvu1y9mVMD3zMMWv3K43EiaOT6rIO04HLv6KJZ3q0XBGF9uR
REvq62BbKVwGaPyjsYGUVzwUXYuo6kQv2vywPyFtMHjm4RekWGpk9YjxfsToPxsT
9zpFSJXdmQqWVh9C1cun2FJUsjKNBvYy2b+97r+o6Klul63hCXW+EHmB7Sr20kzK
P25k3Z8bzUweb2sA5kE+/BbpQVIGHL67deR6KraBXOL6KN8InNRnmQM6wOikbNWn
7+0TcEJUA49UsVBuiP28O4qkXfZnrcWHz20FZCtTrtjMslUtZF2hqUNIksDfmB2f
7J+5V/LBhkUMn4ANgypdeJOqayzXDVg/woZugNkYuykhLcY772ju4BX29/N34Dwe
nnjXsg2Pg0gMdzo3bG3maOUD6R3+eVntjAxm2K2yFr/RqrHmdSi0rScrFECUGRLm
XaYf/J3xmXOSLsQjBNy6mchpkLTj9xxFmtWbhffrwypKIo7YsrJsg5CTvHZEU+5O
jWLUOFTlbFijqV9gSbwiz1QEokkpUco/9PahwgsJPGnuJ2l3WZHEqusssNomQfyb
1BC52GDlVz+UCwo+ihdfOcRs0r/6cJdwObNZfLyRjR+FjsPgyWsQ1euUrx/lmw2g
taZlY7Zp2AR4af32JUOkRNzzOr/6bKqfpBklvjJPrkz0wCMpsRNHGSczVoklN6Km
epAKoF9CR8tCRqstBG2mvIvvP0Qho+R8dv3YrhN3/iVt5Cgv6F9i2wkbW4tvB+W5
/SmsgV/qpw0AJ1n55i2iEN+lDLLSDYfF1c42Xdh5v/wyUjfsqvLiaeOhYSShhHrk
teokLIgyPCG9WUjl0AS8a1ljs6kXXgTltt9NM/VhEXp5hbJHPRZp3HTxwrZ0GI5l
LAmT85Pdk3XoKE+nLiaThA/f9emKcykCL19u5qUuX3MGApfC/hvYkv+oDKA0bEt8
5tmWyYyT2oIP1olocI7j2zzcMlBeNsEqX4M1I4eqVRPWfjutbFMbp2+AxB4ECXQe
0QpgAEaNvLJcTpzR0HKJOgEtE/qTkzl2wLYHMVvh5v3BhGD9G/pO4Yp+pKlo6xQn
OKdjqhKojtmynj37z2d8s8FFXzgc2TXYacgYTMRbjEYNbmVBbfYPgHcehhn7GZdl
BixTmkht/xPk5MqJYDbk36KA0uqdpLiOXhlfKmBKoAXGKeudUXTbA+JxCKJVr2l1
O1nfOTKy3rrksyo7zasJR9XdfpeIvMv8FfwxKDchKV2faBXBs2cieUoNI8w2h3JA
im3pkhywJI7KF/XjlzGJmwU/EhbJDSDil1+6CiJqIgfguPGxCa1+Y6TxPaFEU7Q6
bMFyn6FHZ7zJQb9+l8Aofh/lauuNXuYiSnNpAOVIXGTzr3XuAtLogzDdwuR/fUXg
qm+IAyGDNQSeRYJUp6+2FB4hmgiGGi7W4rZllqtIbJuO5I6LmGX7QEn0TkXFMq7m
WD80mGc6ya18y4yibgMnuNqI7yK1RpjMo+0O6p9nw40epcUsi+4IeQc2DDPxWtKU
biWxRUGS465mxlCTF+SEWirpJeN0zLO6uTqOguvNC8XOPmSdQoR2wqGRG+ShP8SV
5K6sYkgNoCGFoCDlKYv/uSDwRjJ9hBmLZpYR9fzrRzz+eqvjB5qwO7Rm05DcHayv
+x0ywTiGcLIeSDhIqjrZEn9JE5DtLzv93ayUybSTTsGgaw05SVB7gbbLd8iTStb4
eq6MkMHQN4SHyT1Xix4KgQB792muNM6QNRFHHdNGHyx2rM9g82bT1kFegSyMkrKS
vkfjY/gBKvitYik7LmyWfwZubN4DE00gq5cCHugsegdIcq+Bt6AsVZPOdCjCgiX2
GqGStuUqp0Yp1Q0HxhPcQi5oaP4+ASeh4VpxyXyKW44GQumy5KWOIOn7VoAx3vZG
Ln15WSCKrXYqeo3BJIzAOyTD3kewU4S7E34B0DUC5fQ+zIUM76gJ2AjtAvQbaOyp
NuYleCR1Rv2oV+u3IkFFYZw/MWmwjlDxpm4fv36vW86xavolcdciEsm6QEi0+NWc
DAJEcdZKdoADplpubh/COnE1Y7Lu8B39RLmoyTTmVlJSIBT+Kogta2WKVcV3D8jx
Hjiks4yf54+HVIG3VkTOOHOjDRiNa8m/PEwnerHLuZjpeIP3yOFS4l28GUWTGS0e
yR0fdnPjDes1FHi/3KrW+t7knETU90/sn+MtESMiP1SC2d7lwkwsg+ryz4T4mJU4
dH1zT0o1PJ4+h8NMBYjGfAjP1QUVyuX1n0qYAvUp7KBBLz2Q1EUtME4nWET262pB
uMaBE8miK8PqDP7cVat6fWu2Xkg4g28dHVGLbd+ugin8sX7fSRWMYrsm3IL+5ou9
g8cfa3jsyH61vxMz0SobOfQOtJtvO2FA0rWAk5RI0gobCIxEvojFyp7lPA+ozvqC
di+GN0lxT9g+HAiC/Tgi1ouc1gcudsmBe718/vge2caXNOblln5yIFLUb1xeWHS6
aAisReAhb3x5tCsiQ3sIsTEWeJ2TD9eYTvNqRyxbo5sMTiXCcqKphG/kjUCZI+ZT
ARs302W6h0qjdqWBoEqWhpJn4fuGJ4Mi12p34UNMlsHDrRFBG52GcN2qyocwOuoO
XHdxmcGovlAIjev/cK4rUNL30t2YBc85U3owxxgAPFstX3XB4Lnp6h3C4b5lpNSv
TVeWApix5uezP38PDE+Bxx1sQYgWlmmmXlV790OoEKuvNwLpkOixMTWiCuzWmyeD
bgqwfGbS/0ouxCXN0SCgnSAs89UG9fANTSwNmYrNaVx1o05CbnQkv/1QVbtOSEH6
q1HH64Vai4syDLQqlaBw+GziL/xfSdSu86/dnN+RFHXc76bdDgIVU6ylsIYpRv16
PWxiUTineFjIC41i06vXKaqev6lO2otNsQ2YN/RiLn6Cb4Hj1LTiz0WFGj0nYDuc
UJDhBth1/3mSSmXsCJsR3fMff9C6RaQMtG+NdF8GTRjzOQNtIg8svx+Ubkm7ASvT
UC4U/+I7bSbtoB7IkRzP0oEn55zAvO6cYmVPtFXDVXmzThPaTEDWCxgSJvMQB/Cq
IxCzbX33BH4ksPQcJZP6XEpxiKwcMR59cZCBQcl9nkaMbD/8ldEp2v0luulY3H+8
7+RnTQjR3JaKSlwfTMVAQ79wfIgAzOz20IbtU0f8ZYDRuVPVOKf2kdAdmnh980cU
wSVcyzty9m32QOmhkKPm7uEtei0neGnC6xRIf+iphIXpWl1L83bFgNn6HCIj1+PZ
it97I3HGGd9Q1/XHMi5vVM/+K2XY7YPivHhU/FeqQbVLZi0ZbuVSikLFV0ASxl3R
7wNtpnSUbGoAtVzNSXbID41Im+ad9e09VLq2I/2tHKUnz88sAhdyY5m7nOKr+k5w
3dwDdFmFbTDpvkQxytyH9nIMoQrCQQmTvhFTckerk7KQXpoF3/SjiBcDgX15jZeY
phumMFnaQHAUNxuZBn3eL4m5XNFwHP0u7J9k8rmmc0qnyfq1yVrEt1/WgJrhJbJ5
oD7FrJs4jTIoZpVKdPtd5fsBhffTSg78EjvJI51oUD+8jmYBp+u1xd2ZWxJk9sE/
N2Q/S/dY+O3LdMMMtfB3Tx2o4MTCzvk0klg4dL9Rz4j22ZIFMf3iGj62C5lMFcgp
s15H1AjcLl1YYOadsvrKlfbfbXsevWo48Z5g/awYthENPEcCJl55gkSjeTCoODZj
YJEpGX5MmA0scU2ysgujc0EE31pSgxbGTEhfAOEL8fWgmxfdVBUwr89UYxSsX6t5
ZB0RKPmVG3imwarEydUSdHYxoF9UynXC1Uq+4RbW9saYO0cpsQ+VGwRxdlSYJ299
GIndNOFehXsXIQEBI6K2QOJiLAk4DYimszth/YQfYsRXb9JZ+wshidCbFm/VXQSJ
qm+ghYkQOEInDvfrhdBhAadY+VCwJcBfGH1ibVnUAfwxKBPDD5JrOawa0r/MlIvW
sN2OO/Q5xR8FRqJl5wWqtbBE8IT+mE6vGkjb9uoo1Yj3ekAjKLh42TPRlax4U5VZ
L6vksK8l5+3wHgRr8NWYiE2H0icdNEDrtQbZw9UOcUFbQ+EmHQc+scV3Ljkshw7W
asG4RaP3lBmF8RUUv0XmLadsJ/cEKdkzL38dg8mvNWYeJILGeRbGEx37THwyiJHi
gb3YCu8zI9JgEoXfdB3liL5/5QfIwQEdBzX/2lYl05js4XMcB/HFq0ZDy7dqPXcn
/Q2Boedi47jM7upzCEwgswbxFGr6QBVac4HTisPNFdbcOY1xJCPlAFgRrltOqxtZ
g1oOLncEkUJomcOavlh0SbHLz/DXrBuN0BYlAhF++g6Y5bBbgDu6bJ9/X3UVi7cY
iZYWPo6x0CY1ROXwrFENHjC9RaP1RK7nJ9G3xzWmXfqdc6iKeVelOrxhUIHBT4on
M0nlX2CLvXaSbwOnWrsjTNKtpi9cmniPqLsFA9HqW+/9U7QQyxZhHS6HB6AkVCn0
SM8lIUZQvdBcq4uw4LuNf2daM/jLw4ysuDmxwMKm4URdX3ADFPeXW8oVspr816Uu
xtlJ57BwB+8+newlue3UxGvQSHqYQRLPRsE2T6Sjh/53H2ZxZTWPXxdm1sUrC3cW
alLS8xEDYrDC9ethJVuuRPOROLwKXLiwK8Y8A1yzPmGNTyZH1WXQx5aDUFxJXo9C
pAHHt9pKuv3EpIh+Xurjv0L6RB47dMdqANUhnGdYAlb3gtrLe68w3qkVLIuOsDwV
ok1MUUhWGsklX4z1Et5uP2p3XgJYlPzaptZLxnQa8/yl1NIsrNbsNYaDhOYCAVuv
qC5kjGPdiNV+ADLHp8ohBa6Q39gS22k8ciikbozDIrox/5j8IVmbFUtU9FC7HTD3
iyDqYHLogP5ZrArz4e93C7pZgPz1C7KpUi4rGGbuVqQoOse07I/IbA2ItGVBsz03
rKmEW3IfPEh2egBEJAuICwNDQ5tvAbcMnww5z35pkfwyfVVhh0FbB1wCweTqDPgw
ngnpC1vCmj145geDoSdeI07WXLPnIrkiKKyzpFnzvmmywl/ia2d7Vj7y2EGZjLvW
smWxPGXWOHpX0maMlV6uNxkKmmGKwyWPOm58gVnXkTbnvXe6O94vxmBxiQp70M3h
vOl3e7GRZBTn9DNB/RLhtYqaE/kDgesun1xSgtfiv4UUP4/ednGRhJ89QOacy5bI
rQyFYZWCXkAWDwaxFrtlXelZit5hvnuMCUg+xT0qNuLufL7rlN3CUiDyLk6WBdtv
e+1I4zHII8DFXCxm+3gsLASVQCmHMUNeswiCLPpu01c35+QFlC3I1Z0QXWId0Ozl
Ohv6MhfgDAt2SYJ7IfcKpddy2jUF3ZNBy197JzUkkOMWLZZ+GVB7IV1mfSGCwjbU
q62Ca9+fqTP2G0JvSZXvhkgXGakV0YUdP+0itla5PsXpkejzfNyoJxyAvp5koQwK
vSrzal/WtyQ8ZUgG3nanXp7bCyNzisjbplmAPIHoNAax9SoxFlXVRvgyVH9MrCpM
AJIeOYCvkhisKt+BmeWxIc4oR2QNCRdsg97o9kHdHjVsHuWRtQ6hFfuyPpjBCpmf
oYBvlOm2oR23Uyy50D0hwVcHGPGGM+aztcBUzde4bslKuanE+0hRJ1HH7OhvrJUW
69ibaHGEeOxD+ozQwhKTw49JiIvPwMFvn9Cs13mrfX87wVfjGDxs4Y5VNZtzgq5a
V696FCcagSqCVQYc7aoTBtuAq0RBnvADppozpyTnSa9TQ1MTiXo7VvKfzLq61u9Y
usx+yrBu2vs+CH/rL1aS69XanqMapDN/6h8Cunx8MhoBSSOT6FG2Aje0ndMLpcfN
GAj6z/s5Gvg3EcFJjPjCX4LL9AIpyJO0IVESmOTyETE1jV5kSw1Lf2z6vxRDFYt9
JdyF8LJ6nxyZ53vt7lZoD/UPF9UoiJOi31PJbZ9OJOg4n4xOj9Ke50MLA11hPgMI
jhSK9yYn9pXlqjZ3xbALedmcQshoh+FlC0psI1fzkMKw/q84Zzcql6feKk03oLB9
H57dRoYuKwYXobibxia7FP3kLJgAVZP4uoW+F2XWbdfjgW7MK/SpLi3vLFr36XVw
i2G73FF0qLdIXzsQ4EIgWuE2y4Fr97o9oDBq+9B/FqbGm1TgnQuD05leFX/mE0xS
lFfftb6To00ONMuBqUEX3ZpaNWv+C1+e09t2d8pQIR1K2EZPGe67wNDUAAM+eLsQ
B9IRYvwBbiSW2mm2t50s0LyXO1a/ihh6Qs+T2jteaTOVboI4ldz/H+4corrFz+YX
sQzTKEtCX/NLXrAQZW12eE2bXKT49a9y6VNkcjqMezfnmRyIW8PwiXWSAxkPpYuw
vvIRps1lHk0iBLyZD1n6m20XGGQSjNjr6dhdMxbgT5/8NUw9fe4Mf2F/Of4T8yZo
LDgGXk4D2RzNPh6G/NYL1rbmgUn8ruJ+wZQyvs5uG9O1epTSnm4sqvDNyEYgJwMp
Cjlbw220lgoixVRG+VLBr1pijkWl27Mbiy/zZHR+R8MUk7A8A6Zmv7CiTCulS9Ge
vx93NIZGfj10U7/LYaxHChiVsAYpM2+KOIKC/Mv+BMiPPkv9sHDq3k/nXO84Urju
mEAl1SXeS7n++0DJy1HgWRqtMxMstRNTW/wjszsXTjunRiZ+1MeIivOBj5ClzAmI
SenabGCBAcMj4OBNqncyH2Hoj40ebvSGbG/5HOlgmuNyht2x+fxDy7QXyOo0PgGl
OpTePPOEKTphYh+1NIbvKQr4H/M1O/deRkipiodOXdxkRjn8LFDJ0cUG4QBtYL1k
eNt6r22LVGI52syUh7vUHyAzfCkxbJ45JTKi3Oj4D7ukrvBrbbxgspaNa3MZs12d
B3W23EyQeGwlEBYFyneEjUgONrB3KXyLoLOSWvFDVfFJCL5yhKc+WK+Gg0g0WQ5j
hGF49hKQa7MnJ2SnkysCzl/SRBNoU9g+tQxh4DvwV/vJE2H9YFzCMsSobgRkxBVG
J8zqR5CehZ3U/wM0bZqdyzQkgwH37CWmrwB6c+TzlD6jC713TX4Q3lwRkdHfDj1k
qR0m/eiYK42B4KQk7P6qESkelRa67Xzzzsc//TOAy4NzVWGQ3/f91E48127TIvgp
ryEfl28dc+swyFshrcw1arNCrvfpaqGZSRaatHZ/hUT2wXsUdteS9ktzNCMmWCgA
rP8t3fpDMi0XeTmk7HYSEjakLISdgy7keMit84gTN/c2VAKQSWVier1RKqXI1w16
hGVJ30oQpECZ1vRQYPy+KKCI3LWalYH5pYGvDeR1YnA2yuPHcTl7Nja4YVCIYa11
/6iFQSBrG2iFuznn8SCL5TTPbRrU7+OnBVBheuO7TTeboWgrpse+aBwF63lc+pJb
GMeajKJNLkhW5gQRlfAPclGtqAAO/eOWCIEFlgEx1cCvZp0eHZosXZZgjw+nYS9/
IMKW0zvpSWPzsLprg6duXz5ASblMO0+sn752nzOB137wHyKQrl6KqYfi8A7EFgSz
yn7e9zYyaFwR+nssgmZULdKdi/GvYqzaJC6A9qimAk8HXH93f1HvYHVybfRAZDF6
TebvTAfOQxhiZ6Q7+2WwdazeDbNRwwAc6us/HVT3KtSX8tks7Bd/Vxf+JHt+1R3W
0bvDRBq05yCV2p4tcZq/Z/sil0Nz9ffK19tg5L8u4s7ytyhl1LJ4HfceS0dqSlge
g/iJNA7ecqGZXR+5/1Ighy76/gC6Xb+BzpIw4xdmQcAGIqXqDsyStAF9sue+meIA
5OUEYbqDcA3+ssCKQEBEI8MhkkKhC0eDpqoZtV7ducd1ncDDzJsqKmV+XF4o5/R7
ehAmHQqSZLVP/FWXvKF/DvEjt4tefUDy3S6ULDWeWgV4tLNZJ0Z+F1NijjPKCI+1
Yire6ri0/0k+NAuj1c0dyW8iL3RbVDOBCoSc1jo0EsAfLaJI+6DRXLR1KyH8P1/j
NlK4MGUHjKGK0IufeBzfp/ftlAjWe012mSuTYmo1x4Ei03bXR5PW9PC8d8hLs4kM
Tdpuso0NTwyqbaca/ZLHpDBAY6spEGR9g/Xuf1z5rciuM7o2mQpyeTAP5P/uEyy7
sGl5l/5G6vYYCnC6pY0eDn+j0OdtCfMhyqHllJTDZOyVgNoh9Gbx1cwftH2EQ5O6
RAqa70aUCZM+8oww7pvNc11BCj41NJUvBpkt7j1ndqEwOMMt1OEWVTiOPrCIA8v6
c0AgiQrot44W5khY/j1PPxGoOpEakOqhvrjjtqCl5JsNbAii21Wa7l1axi8q+2vw
CLpHKYKvFv7h0DNRNtoJDrch5JQ15OoEsmSMM4k4GiJmUsgqhMLhJhIzQ6c07V9c
tbO634nnLKoMGSad2J2lH9URgRzPkWP/zJIekqNXhtF6r5Uj1A7AIBH4nLoc7Vcy
+yJUNzecsOO/eZ1jLCOAo/VR7GdInRPAtoVORpt3P9BAY/j1fMGo4iB5kawRuwnn
epitJbUCGpBWgzDQ4ctYqNr+iinJhREq8drxTMEZrqhGKpQ3jcpNIql2dkKNIvTp
9Hlc2tXVpwBJowdFfSpeiHYj7P0AUuVVjrEU4Sz0jIhLfoAjYteJpSL29bEq7Fat
TtPQnAHMb3EdvNXHHgEkTQrFoNMy/3pXv1CWBZhtNogs2mCpn2OY5j9uiJgGMQWf
lTBQXLG9PMoOpG4OOuWet/IwzP1NwZP4xOLmqINYyQBwjwKlpghTuTz3lbn8+ES0
D7Hz6lsbzNxJfxnTXl680ZoxIjz932hP6pyDQHLjg8RHD85JFDOuxKNkp5J0/rZM
/w5jNBDHZBfo20guWSrMJwwJKSgsop2FUbMOxLHigjcvRiRuJrATc/ePkFJXgXxU
KI9KdkPCSr9Kc4r4UoSXboOQ2wAB7A3cABxqSmEWsFIwB8z2t2eiw+NNzlm1kW7Q
aOXvmDzO+ByVsyGJnv5FP5npU3V4MJBU2edHXsTMwrizuNM4ctrHFy2WxGwLq/bu
WOcd72G7HrXk1MlojeLoWzJKPVL5Q8w7DyAS/Rzg98UJVPdc0TuI+sl/HxdbB9BS
qfJtFbtN0S5LOrZBeDgRaQIN8QrhHyzuWTycrhZeIog/8S11We8L7rCudUKTSSwn
ogJdeJtmx8hzCgFpHZjn7Z+bsgQnBcfCBtHqPfc2yZ5AVqhLwYIXExS0o8G73nYQ
33dDeuK0PUvlP0i3DsqWPlRI3kO9nw4tgW/6iaOrtGKTN8yQCgY6UuRf/AjHO3IZ
gsV9aME9v+iqbPCeqKGdFf/n9XWlB1iE2fnyaRmf3gUwGLR2tsHDGf4+qiy4P+M4
eLOrCEJW/vKIAFMAcin/MEbCBQJ7YcXYcMiPIMZKpctX+4jRnZoj24BWALjrN6Uy
ZL8PsoKDmTLNzDSG6vpzlNbKaUfGocyzHS1TIMR+II/WoQ16MgOuyDNI0qE1qqgs
SBljiNXhAuHB9p61vLjrCroTFujVrZKhgnFe7BVszgAK4g4dlcsJBtfB89PZ5vFS
AlwDXj37AwUWSZ5LSby3s0bngIo2u44Q32l/IO3xhSKDOY8+O6+yPMo/s16EFk1r
nE0rJYTUom51gBv2wgjwxV4xzBWzOOhpPoKHY3x0+vt6LVBIzwl6QMSfts3hZ2wQ
mT6sz/qEWwTFR+fyqwx4srC+7lFMGn+XIcFjaUQFlt3A++kci9sJ4kVrvRLpZy3b
YMzW/IJf2pBVld7sNCNdCayxZ6c0CKETtE/Hk8WtRIhlTHTUnru0tObqPixvB301
u/FIXhIBHQxvl0r7RnAwZOq4c9QHKIWKFoiEw3qdvYQFdy9owkKFRYf5DH0TwgBY
LOqZoZ4mBkYzCTC+olsXpA/JdpQoGp2HrDVq09cTM6nFC21U3UQQDKEaXUNNKBOY
pI4Naz8lW4FbuOOMVX5FawM+uZNGqnaU1e64Hd/xx7a7TA2/KsgImhgUz8QeHzYO
eISuysjkYDjN04L7VGRmQBI6ybDwBGEWg95pBionZBRV2SdnKl9zOUAn3vGe0O/Z
y1W0KRCWk+6YuwQbHy8qsQyYgKGGcMKKshrvUgUh1DhqLmpWtnZyLnFMYXZGMqhq
LxbOjyVkXBR5wVCovrYGx+LPHe3e6+Vnnw6Y2E8eAKgQ4FfQv5SyyfdNEhvnmsUn
UE/M5pUB7xN2pz7sVC7XZfS3+ljX9tNtKWKZJDVmL5RtpFv/wlhmO4o2/Kn69EAT
bGiUooshvzEwiHnL/kqY5ivLnW/GwTJYrH6NXTHzwv0IJnD+Urb2rLaPxnbTARzE
iWXhO3PuUwZJnWWWfdfC1CYxTwatT2+LXhfqIhpmtPPTOcNZKA6faKRUIwQGSrNv
+zAc29fB5OY2LS40NhVRrYK1p4OXWEd00URQFjUBufcHjQ63q88LC2k9dopp/Hjy
l2KXQ55fr1BRJulHT1O7E2v9zqdQwOvbq2sKjIJS9s3ToxPJ9BO2oPX9d/pvfsvn
Au9Gy2UmB/BKt4o2/ni942e+5M+T8iqKoKpb9AOq4VUE+YjH5WDseYUHtZv/yf7e
UywUHcCJv9BHhkbCdeSHAf0LJfxjD437FwL/WqS5aMB0eocHllo9h1UmicctcBWN
XU23Lu8aRGlkJZm8pzL4unnvvgo4kgI9j3SsGHJDvXkG4K5v5ol1uY+2M+srLgO2
TjSmrFHLjTQCNvfD+TdGqVRGMLNtYXUfeA88XgBsfEJjSHJrCeDFmt8sZnP3xS7Y
8Y/rI/l5371hRQK9tF7n/qX4ES5Rro9x1jyg/IPLxn8FfOpVpiFRsRgpUjBhGrQZ
6SEvrSVxKtAN150j6ax/1qdD5RBh365GNexepY1dmgwu5XwZb4tH4jxQ6vMu4Nvb
urb9ZqCtsYSFCvdvbBQZKg51Zw6lXz4YbZFHPFrpJ2KAN7hUvg3hPbzcCcY2pFMN
7jSgUIxrACwAThV6eqr/2msBa58THWSgZ7pcaz73LFvKQPIm/XYOlpMWnK3gLOEW
8RlDpP/3voBUWjrHRfDuH7mB77fmHizUIvoc78Nuxobj5Jonbs8JC7HTMhPXBgnq
6Pj6mIbijthb5+zxbByPwVK8AmDlBgS/nf08Jy+TnvzyZJJaGxE8BG1Ette2Glfz
LI1cjR0KvL6PJMGFQrBHGaXLbFWHOwI7j+xEOrjuq3mEtzdK5mVUpJ1s60RwlXX+
B4dmBhaJU5WIdYxzghZm/D6D4JdZcAXWAVOxbLabRMm26oDAj7BIfcMsNq/tDoSv
gUvRAVuMjhBOZtfex/uzDABHwwzt9+vev3YlxV5VGvLMlD3ha2GcERlaLK8ZJ/Q9
0o4JF0QOU6ignOahx9VfJUV+N0nUuOSjM/qOoSfVZ0ZFzpDK+0HAE6oWkuE8Pv53
Ov8hbcrhiw+edGRIL3VPfiH7sab7C93lZ3tSedVMD+QTm4zJD4sS7NHJcnUmrspY
n4adMUWLhphv9etVt3BRPZV5gS3bM10rIOj3vOZZTmqdHfr4wfZNizr/3qrVFRIN
f4IdKKG+KGS42aPrzGwfqngdP2WHlrzxDisJtpIOfZZbBIO7yjSkNl6o0Rcue9in
zORRpqCwfUU3q2XulwG3QvVB8N+4XML7eO82FQSiSZFaZL5YjlcQUoBhM+/obi5y
e6gnwpJR7OjJB4S684VNXiHTowD/ZwnuOlFwCgktMPKAQBLOiePEzbPtl498hLvy
nr+9Ix8Az0f6fmV+IDevFGZaYhCmCyDd1g2Ap7zbAlSIGfy2wLJhUmFVGHvt9WcC
Jv4JITy49Q2u0KYxexVY8CyBBpy1ffq1M3MuQayH5QmZm2UZOEo5atS43ZD9k6cV
u7WYe7CfksC4lX/QfBrsoSLsdLbf/k0a0CREN5stsNJ9jkP6K0QwU+l7wJ94MITj
ClKZFA9+xErMf6G+yxr760FQ9Kg5nMmxB9sd/VQxwgjOZylr/cw/S10qza5r003F
Q3yBGY/wEwFCAmD9rCXFqnVXe7f7yVsuEifqeF/qDfl9HAM95ylYOBscsx09HPDo
w5p+cS5evz7m6WctAVSQ4kCiKnuPlEXqY8ynTRxSzIUedZX7Yihr1Ladfh52DgHm
w/7+A7FVuZt60aEfAyqSfnrWzDanEXlO6vbkbb5g768Qek8E6PbpqpGImZU1WC6S
8VkaKN6ZmAz0P+Vo+CnRAgSAUC8DxyITu7jTTnW3drvr45MJR8rf9ixNl0OCBdxz
0fsngO2l/xEHSzG9J9SsQOTsmPE87F6ScpgwiQYo3y/1EZc76qPn/RyTiadsS3qi
pL+uAAJdKRYLb7HYPiyPUJkk5qaDSNGqCtcJDUFYCT6J5+Erhk9lq4PKOOOgCfPv
3ZzhGpbueZUZlqLP9epalOPkJmy6FsX4w+I3YB8iifXG5OpnXpesI1xCnopFysEo
gX5Tna6dW/i0I0N4jnJNDDeXqyJRW2wzij3uAnAWE9R8cvQukC3L/3SMqekglZLM
E4xlxRMkBqlOCvXXn051olDK/2IveV1KQytTeGV7PSmFjFFVuArKrAo93vPASIz1
vuo490qYC+nRQY4V0bf8zUkLgA8vk4O1PC5Nt88a4KR22UIINSOiS9Cax/leGnub
zNQkYq4PT0H7/QE1XPrVUtZDDwP3H2OGAT140hl8Kw16J3+aN9A+ml9wuy/S/gxw
VJUuWKWXrjY/cqKhi1YCiSoCzVCa9Nf/ADEcAbFbzJcxJ36RHt8LuMOiqHKz2N55
0432pByyQb1xbJqomLsiwV4EGd/CCVg6cqBcJAIni50E1geiwsSQUl3H4qpYWUAW
VSnCJF0zcoJMF/5nerLw+c3Q1r7dYvpth0KVP+mJIAt1fazZKSw02DyGO+NrpOsP
usWcsrSDQr49WZo8XIIeIJk+cM0YwtW+Pf52p2Hrgffy/u1gDOXdZq+RFOlpJ5LQ
HMXO+DqBXkS44a/3Z8ykV+KYwcLO4vZdJ2pyOV6Cwsz2Ve6J/So5Fd+HGGYYeI44
vwmxenEzA+uu66hKKoM1h72E68wZzpxYw1mcL7O7krLg1DfYSc9AqhzEY0RNkb7Y
+61iLdUHLcqg3MKdvb9MqWEiVsLybFJn3AwAckb4FP1WuCj6b1KFUlViDcJKccBS
HOIpb5b7i50thxMzAmYIyJdjft8WL8kkSalYT2k5JqR7VlCs67Ma68xjAz0kElah
pGIq/0MRfIz7FpziJf3P4ORj9p8LAbuO5ObC2f9bC/ovnA3VtnhRXZeZEkbnaIZy
04GGDFjFcP157RgbHaL6ORZoQqn7R88UAh+tzLkCSFWzWkT+K93czZ1mS870Yqac
2jGtXxSaFN63utV8c72VPKM9CBLHm1KWHJcT1RAYlYZGRmrNI8uMVIIMIJG0xKYE
ErK8y6sll/JdVLfvSsrzJ2gS1ayTiV1ylhfS/R3uS5TvzIdLm5C9Y/7mm40xpROz
EJBO+JTi2kOcH40knd1pUbq8nC67bXGfuK4dLjYIG8VJLqt8Acf1bs82Aq3gQVuJ
u3AFQFURFXGWAU/BGlNxNild542mKNLrmEHGY6gdEqIwofxFzGJte4X5IL+pCNjX
RsyB6g9QCEpbhkS9QAM2ktbptbKu8sSw6poUjNTUtQ7THSidjtrUjGIIxXhJxhs9
7cXv7CZ/P1h17wR10sPvWLTPF/rY4UwqGRjW+6PZYlg5gI9Cs2n/Kgys5Kw/MgU7
wGugVtgeTcZAv1uglC/GE2r1+3fimv8OCVWGpHfbCU2/eYQ2TFs36mTebTRmouG3
iRXYTF8tJzQbQYHbvcKR5910Wlr9FujShWDcFDMpKAvLFLsQfzB2T9H+ERisbHB6
HebwwuxTqfPXWOCVBcJKmBvpFj7J6SM9xzPSzt1QU+vQnLEqbdL4ia60bl6LuEcV
eeTa+Sn3srYKCrOP5bKeWXEOqOGOw+vAH80eXxG2SB9aFc7PLoAmgU3c2pB2t9gW
SglKhT5pvA9UEGG2R3o2ddLWSuX3pSmxVzD9t0HzfL/Y4o7cjYGVBLuxhvX6Q+cp
arl1or/huGBdylBzA3PINxJkyHj4A8KgG0heLZPm2qYFppBzLNLptVXUWdT7/IXe
ttAQxDhUlwcx+vXbC4U8Bb7ZDYxbRKHDiy8xA09Tl6l5ISxk5WYCFBjLLQJ+i0SS
nqSLxbfOwJVf5wwTQj57ZIeE/9ywzXjxbLXil0qOTOTN/TWVnjyE5ZPXOBV9s7P9
Vxw8q/dBYCNDKhuurwsoQsUp3ufeCYfUd58Jsa8jvGJ94zbeo+H/fODNcsXv8F/P
OQo09lp7DhABgPghai2UGhIh1d0teHgI4IXbrzBaN+J2unrl+whpAJ19wtlXNquL
SnnuFr3mJPai8DMB7RaZBfUj7OSveHshMnmFK/yZCkQDD0LflEDGZKrYoEO9Wgxx
+PDZvuU7ccgs3/sRMe8YUlzRfN6T7AP+cWFo1TA9Me7Jtnl5gaxdYywSb18acd0r
TSRMfrSTCOePrELxes0XTuVtMEhfDx9/dJiFudPdjSeih7TdU6XNbquy5woTyzfT
cOeCa1tH9brq2OfFUYZgNqSqbdyrqYFEQOQb7I9SnIQYU6pnmWRSiHdXBUE1p6WM
EnAK58oznYJ5cxQck9bRgPmXwjHyeIuDThttSlFY7NmaympjmfRaXU+BvSAG3Ouu
0FU2qxCrPv4ORnTWQQv59yHzZkHIBWsU4nhPQeSnXK4/O4DmqcPAfEwg05S/FUG2
s9Z1iOYv3xTBjF6Bv2s5ej5SlX3ruXr9cWwQGVK2HAQaKE5ukRz05LAwPmdJ2J0I
BSCs7bv9/JI5cp9ejmd5fi2cjNhAUwH7tWebekREAtUV3sW75jwM8V+7uGFjNsst
rlaKu3/LGSmsDGuUaGSc2LO/E8xNbXTG1r8FuMOKzztMutTJcTHcs4VXfdS6FRwF
3DALXun3mzdY13cDcr/xRzOA7B0XtpQBk0A1uEPbAO5iZSGlUvWd3RhgXAUP88n0
Xtfh617kovSpUY5afvMQK0LttS0mK1XffemPLS+AQ2HkWBhNKrPK+bAt9cJCei2U
9ZKyPqISTgCqAdfNxp+qMai19WPc0YJRdtpJEW8MWzC/jZl5pmy6jIgN44yK/yBl
ZDJQ/RPS0Fd+O4/wBQD8iCLtyzQZRBSrP4vxYNf1DV9Mo/r7rkDez3Nn3URIgoBM
If63m5OpjvbEsJgwqGUxinurn2qwud4SNDy45wp4vRnHQCNZ/HWdm0H6IP5ieIVN
OZfZpI0Jy5VKoBUGxaPMoN4AhR4bXXpZxMOuI6toiS03H7BUbVleUHr9gggEhUly
Zo7xRtVxMfmVmGrB8AwtPsFS3HlX1ab3aZaFFXL4nvm97gBooTLQAcy/HltrWk51
IZrYafJEDDj/4Jr+ENlyjW8lLKm/GQfEmQzgjlxCA6cO4/5rDdKts0BBqrdqqKm+
VTR4dv7H7jTHdvhw5TlkDs6bYGy1Fp9cTiaIepwCQDpZBo7vFpn8n1FHS8isMkXI
/WRr1lObhMfeISeMxVfC3tFIkqO5OiRRyF2MG7ihR90JvTdn72y0j8z1Uvm0MBAm
taLdaMgByQ//aoKjE3+FIG+Pf9vnpnzY6ldiWOV6B9wG60ZfFGcsni316dnawTtt
yL9DlvuKnkzBBB30tujv+ds17+lJ9dL2FqgRysqW7gAwYxSi/eTla4AP/+zayAb7
RS8Ct1Tc/mJHXbRQplDNRGJztWg8fm/CCKtWJCHqCPbSu0bpfXG1QTQBKr0adfHY
mrAZUo8eeUNwAhFP7rzBmzLlXkI76p9CfdN3uIGy6O2GRMs9Ko4cgEF2qSytqzBE
o0HvlV437HGzI08wT0KDMoWTTa+UoQ/N3yY3jI5gIaccRp6o6wU/BNT1nHfBug3k
KwcwSi5G6Fr/H9LKbB/8UDUMWnQjRlrggkCkt+rEXm/iqrNFHGtDTI33tCPrQzsN
vYQfL6ksVnePYZEhQO7lr4wuRkQx7bPhTkY6lTyxRu4TkHmxlTSiNTs1Ha+ht5Rj
XLrr/8K0U0UnVNj57QZGHNLdD9Y6FsNYHhV105kZjqreEvoDOj+0EwvONHHeo2CQ
B2DSOyegSbM3WjK1oVkDe0d2d3VbUkYyZz0udeXM7Zes/pzjLvvMosTSYKmJKd/z
h7fkksaAqrckKQIspGXQiUfbx+FPa82OEolxKXQEnfiYic8oX2Tgzj7n3bhyu4/E
tRcqPUcbUfQ05Vq6v7Vv1JU9qFjEbj4LxcgKtN21FrJwUsOTLnSsX2ge1eUnTqDZ
75Sk2XeoJ2WgZmiAxqD0ugBixR7r9WCZOYp0smfdMckVHJ0amhUqSWKd+gUhJtm5
N99f+LSFUJsj/b2HRkoHl+7y1ynvj1b46qRge76WXWm7ZYO8rQhnBACTJbPUadN9
Hpd/dXBOBEf4GgeRp0baIU/fSYY3nwQiSQarRd1fXkHmRvWzL68Ofk5QZLO0NDa/
b1lS0K9zkl+vRqPYrTNlpmC5IUOvFNEAQcnca36XQNLow07G/IahZy6m6FweKhjn
FWmUT50daOsdZ+IRcvLFiFqUenlIlKZdBT2iQhAG0iczHVLe5KfUVCETl6kmjjts
S9fYjrEp3QgOd5OpF08JvaUreTpaNFE7vQ+TFOLHjixK4EdMH0J37GKPkjR/vyTR
ngqmPS/hDT9l2b8S05Tp2roVyKd1axTueZkT45fdxufNPEVzzb7PG8UMBFgVgQ6I
xbo/AqWihEDXAHtVBytWFP3wMG+VTyAEzK4xcDy19NnVLZfU0+Qafnk2DWvo45eD
OYXOIcOh0+WYP/EY2Fv+Gadg5wUAr/npLFnlV9m81+DCfzUmXBelcXqk/0AkcGhf
5EcKtTZwi0jSzJwgkQLbq6vco3GlWmu2GdyprL8Ayi7WkLsbpadgMGiPN9K2Xg6n
6BCWv7xapOojprVuCuEKqDyCeXB4tE2TYr0/3wX82tR9Uw0SI/KN0Usq3BZlO5lx
Zl7nSjYonHSHc1GxqmInyTWrWMrX4+dmqq2w1oC+crQmG9MYM5bBLGNd/Uj+ssPC
yMcwLOKHn91UJYT+pIYcW8r1ji3embqjlnrFhOehDh/SYnbq5hupWCzXZGn7v1O6
h1I+34cgW00QDoMou2rqOzU+76ShV6R9HqWfo25/AWQ37OpTUG5QQHN9KMNhGjtU
Hr80m8L95QRE7Lz7JupAL0Lv559Jd9se5Djyr0yDSNwdmMpRvXkBGA9e9ZPVlmyV
eqQHPZtofjuzguvw+rh+02cLnXOP4ZjclyyNmsp9QVdWTh3+W8SshAHdAto5nBBg
SqaOKLlU8con+M+IJ6hzkrZoPK4GBGtFpHtE4Fdrp6bzAiPa7TLbLDF2/SR7x7tc
TlzZ5fB8G15AbgRAvVITjxLdEy05NKj7EzNhLx8aAonuBZGlVXDAdqsH7WwusI1M
FCdGgva1MHvnxwwQ6Un77+/AKyyCu6s04i8VfqjFjz/QHhz9g3fTN1/ek2zhnQw0
5mEZeO/+SdJ5MO55YRTnhEJO5vF1WNvOZf8NVJaco2DSX1De4ZjL1EN4AXM4BZe9
WC3+47sREOF+7a3x3psJGZmQxXfB8spk4LMg2vMJVg7iCHveK9aszg/fbKe/lBUg
4/s+2EJ3czHMXr3QGYFOfZ3EBbr6qcdmwiwZX2rz6ZNV9uqeGjyIxEgjw3fsbfxr
qzFrjsogbUNHYZfULEYbS3TERCj9KgaIkQ37kVUrCtsspSsFbQAcQQ5i7te0zANN
WxlbVj4hLqQETX80X5gU+y3O9ZTd57Wfej1Kw09Goe2M8FtyOsy/6vKjT/thhYif
JhtZBsXe4mzLyZRH/Dq/1bi+NPpLnHPCe7YIxWEF9R8yGsuhB85BacNmYoRrr7pY
DLujhE4biqvYVtCwzvhf0xo3Xi74BOlXu9cLwNUPE0Urw2qB46pzLh0cPpxg99Ta
PP5/esnXUAcMcg3wah8i7jpQN41FEErm5CwUUi4DXk2QHF41yhKL9AhSGCAQNHQf
lwMf1hZUVXKjzGxAyo6yXkzG1+v4bCrHHcn/nFbJsyxdGIe62FFAs2REoxgj0aMP
hKh+IQqnqsZ1Ojp+Bo3Xw5v183Me1cbMwKJzSwdRIEfBoXLZbzup8jhrvlDbdbr+
D0ZXVsKMCzf1JB1cMq0TaVkSlVdeF2hHqb6Y6JhaFSEV5x6QBYWsNG8Jtg8z1fWz
x2zmN35W7i7I44sbDFgJnwBTXlNjXRRAnQsEjQ2se1fVnNX1xOLvmKrpIum9pyty
fSossa267rpjhSHOQDZIgoTznnxZXZRscHEvrAOqMgv/U5Rk8hJJ6sAVZ5Kjk7DU
ZTf9g5d1xlDDazR3poH9fHfqj+kK6LCJvzziewWxntMKWjd5Q46syWYMd07Vknjt
B4KpNy+Dvr/ZXKQfGwf9DNdz53/4aHs5us/TfY2TVqq2RGhopTmZMr3F6INQVZJg
EKY2/UK2C/Ay1pdaQT1D9oiceTKb2YQmuJUxvEUV1EIQtJgenpura2Cno+a8OqRF
CEfHnE5c8+aOexy82bhMoLU9amCqvU1/qXqY3UyoeWm3oaoVMXbdcc1WCD+A5k2Y
C6tIgAIpGwKuIxDNb/CUnbB+rP6MuAh/ZgsDsedPVxB6RvIaDGt3+FJ/qiVj/hZK
62Q7N+z4PQWc2XgJhFtk6c8WXP1BTTijbUsg1rPB3BttV5wA22yy83CXsE6YLG4D
5U5rD2/41Z2QEst727LEaa/v2prfJXOevQS1YOMUeO0iUK1DHxn/WItT5cCKTrUB
2z1yn7TkymiMFJ5JXwFDg635obDLgwzWhsOOIdk9lb70VdloPflqPYMC9u78R/3m
3xFKYXdPNOC4hrRgE9vPd5h2B65pvO7pQM+AeModWBYtZkiTXW4RBYUscQLg/2S5
LjhNHMY7Ef5wW9DUPxDXnP6z5vMSNVThWVWRbkyPcTKw04rvAB9fv6m3tD1oHC/h
PABf6HXHuDA4kMGyCvg5Ciu45KTnufm4e4F3Yp8QXNvLWLoLJzrEBotPeM4KC38m
CSwXETlGaB6nV8QyL+7CEncpYXAkebYXZYDxhyW+plf8u3GljMsrJa9Z6LLlFE05
3D/JuHvlzriNRtDWsNhxpkLQR/wdBby+5UV8xoFHLcMR/1Er1rqjUxbTlJWGOyn3
84xjWV+UvpzYhvpsQEtPd/V7iTD0Of6sotG/vGZ4Z7j/+1uJRThzcyI01Rg9XRu/
OEdPdKNef/yEbzFepPLvvUuSRxcgYD/kCaBVZnjsDvZtSszJgZBRM+zg69071/75
p6lJaWVUJjS+Xfwyt8nRkN+G3qFI5VBj3X6N3xnPP4GyB2vrtmCMeWa2ohnSpKTB
SJQVMYXQgb6qASnJDb6PLJqBlqwDQ1Rd9qm7TFx+yqaBX+mCVOI9lrm2zmIypNUv
ScQITXU4x5nJgtTW4JIGNZLs2ieOdijHDsILKqZQWjUHZCGtbRj6ZCeKzX4xfUVF
l76uxF89vLDfPI36t5mBB+U18We5oXe9aSoeoW8LQS0HrAI1crAUoE1k3L/dzP6Z
xqQr15ljcznpw9r4+i0YJsNJzcldhB2+CKnHuQTKqRoXfv0iI4vOjYdpEgTipi61
3ALqJT9R0oQgc9Nijck7K7Y3hFS3Kxi2z9iSPuBWDQzFkZoVNMZEsPNKHZCkz3I5
gwvaVfp0ylw+1efL+ylIwFfC3drRvrn+6pSbFjAxFQGKVgZOUnLlwUiv1N6AH7dv
KaXRopNdhmSIBs15f3G1COib2cc3qzHNskA4RHBqgpST9ynVgTRhT+lRjM0lNvvE
Z7qnzKQUZaJN3m/4C5gYD1OY+0151ZkRRivgKfiw5US+Gh/TcVeqfLYjEqAqsZyF
2J/OUnAyL9C3TsJVU9JdSYHfSSvF0GUOjwRYZity6SvDnprvSP85HZFkF9F0fyE0
2smRJ+B0BT5QwQzpTp528Le7hSSu9MWoluYyLVHhYLDEUo+VYCxTWI78TNOLsegg
fneEIIXZi708zc4kSZ4TxRrnnFSS+WtScYv+LPsvuvRkFIgk/LLdtcR6nqJuWd+P
36Kph4KQya0NTY46NSGTWu+i8qm8Nd+wveKCGoEZ/MB4AN8+j+AJ/fTENzOSW4H8
YVSABSW5Ty0+2gV40TZ2VEjivumLQLueRWZN56BaAgbCs+9URtcsF8UiLTrl/Amd
HbmH5nDjyBJqLRcnT5h81FmdoKOtoKAsvJTlUxvAtLGUgyjSJ+bQeKeAJrbN4c7/
2QLS5ufFt6B9m9wGJj3L8wLxrpiRIUiV74sZjL/RlpiMdZTMEOHydf0ybx6tHzx1
/RG+B3aIw1E11BavI5TgMDGaQ7bawlXjco8vxf+v3wjgriSiPZAUcH6NahWtFduu
mIKJ+6jvOWxT66asb3iS1jJca41zsQfL3Rr5DljhZCqUJ8T3Ig3XcKxklblMVLeg
nbWDP8B3FZyip7wiOdhA4h0AWK/DAzjXqKG9HgnxoQMr6oweA+qQ0MfMVSfna1e8
kdhpAF4eROMRovGCb+5FWOlW21kDuGp/pRarFWyZuzMmdU6/SK2EHW2ZW0qDNo8p
YRpnaczvmKVaX3azoh67NCCl5TKOaPCSHwyvCsAX8Cc3181GggyCiyLeoZlw/mz9
1nMY7v1WekGFr5LX6uLFeKwy+B35NWvg8fxmL5D65vW8WNRttn2ZrTFzdi7IayPR
oyJmA2Kipkq8Pe0xt7fSAi9OGcZiWVHzPZinWD7DVF6gVfZaQbRql3Jq3C48oMaq
N0oZs5eMYUvWxaxYgk2VpsCPGPNZM8HVDhaofRrff22b2uCUZxb1wZ8c0FAD/9Qu
0oXw9GDxj8iy5PQ3Sp6yepzUV8e1NhhdaYBTfiH2pMGGoc4lLRnYpoECeS8EYu3G
iVmsGxA+Uj/FVcUrP38VdVG1TUgVb/oFsB0SB7gsNCIk+ci9eTCrQHiKA3W8zyHc
TCd6mn4fnt1M1Ev1xC3tKMHy3ZVOcZk1yi+e1Ro6uOU/qXloBcjjBgFZNsbaA3ad
0L3e6pitAhaDAZRhSLsUCpwo9qHOhrtX6daIQbJx+8PvTNMtfLw7OZCeT17mFSMe
Blrf7O8Pxrcg6GCu3q90upd18HlJtfDPKDfkNnD5ORI00Ewd1yAChDDm9YfGs0M9
LXGNUh1bHdi5SNWhD8XSqaWawcLiT1r5WZaFpkXiWK3puiM/zwUAxmH7j3+seXsW
0MHqqQDzehk0JSkbRzVeX2jAGZbk2daD1CGbfLWFF/Ua3rCgnRowPiLdYjdVEMyD
OS9JdHZB8tKXJQ9sOAafQEreOvRJ48MTwXGq3VsNNZyjZs7t7AGYQcpdhS0swESY
0u7uRvwEfW43YMRSJITiZdjpg64656xZbPQ4CwMpR5zdEDlVb4dkh2pFe0Chftqu
b0kpPj07a+ES2d1LUy5LQWCuI4oeo251AmHhs05A0f91QrKqaAlWx8isRyJykpLH
puKvsJQ1jG52XuBYLpJ/7vXs5ds/EoVOfXGEHDB+rJCbQU4uQdtCtE88F2LqW7kk
5C6InNQCBo1FzpR5MSt+/JExtkuWJTwgrdaykxctkVzEqEz8rdVDFRA68Zy2kZsl
QZuMEiqp2346vESU/FeO9JjGL1AF64StRUCGtwWJ2URKRuzLI+LjR0D1O/GU25ls
C3qJw2FyP2jwAhq6uuw+Zmuu5afdRZvwubQhY8FWHAyr/AfBg93UVIjz1grJEk+t
x0eao29hNP7C3L7l75QzzkorpRVlGgezGaMz4fz7fGtL+RZNc21wokPhTJgNWTE3
LRTrYYLPjs8QK4ZII6HW7HgXF6PCDjWi+akCoO0dQfVRYKFSzqWv+N94VdF9Lv70
cdSrR2reIzrOKBgaa35i3nM3UHtCT4Ht/w3x3tHf2EK+gimsBURdRd3SQBLnogIL
iSoCLUr0dbZANL4VmQBTiPe+JIuoSZ30lTTZFRkb0PkJKTNF+SCLtrLWDXTmjyWH
MvjREPl3Vdfg2G5Ghoz65FmdF3i4D/zgPsTYJLXSGCXiG9WvfarpQ60Fa+Z3C6YF
u66mtQn+mQLar4tAIFlAOWhNYe7nhDx5tVD/rRO6Z4Zj7Y5fYEz4Z96K49K5u6sK
2L39u6rhelmbomH/Jj140wbsRqrSlYpayzbd61/eGFatGZKC9y2tZ1GGibs4UudV
5uiYp+cosHJJnXh9//FRv8YcAQm2WpHU45hEvqAepcgbyxH6uxn3b+H2MGXG9G/1
ujqk/15kGGIAmruxgggn/fNlmHkV0/NLFFclkifUy1lc+aV4B/PrpiORYzd/7Zxm
FJt2YQ78M6i84w2Yr+diaB57L3fjnQFmk4CQEol6Rw1iXEnoKr1ujFRcshU3Di4h
sZnBNJ/kyk5kIb+wRPIcbRYOZkfEwwnHBJ8L/LIQCKiChQ/NNJu6G+PfIQPTXXvB
0yXiYAO6Mw6icgfU4S4o7FA6WEUrWTANkHOX0dy+i0WxDoXu37K2iiMekc57VFAT
AtCXFlK/awYjc+WrKAas7xwaCL725P6Z7xMlSg7hL1AezGvV/lxhgjCgXHa72ROQ
KERFnVYlHJ/Ani06kL6KbXIGd1hTsuzJsgcW1TGGH/WohmggFt4e7hUVWaLQi/G7
o12YszjGrWLaivB3/LYMZPkY29ilISmzZsjI5XzMGKzpPGKkANQ/tCFUjMxWzyn8
ecAxkYMc96+X5szfEbDsUloyE40aygTc1/XTeuOVMFtqS6+WnfeNl/T7t6rKKZVk
kn9IxFLzROlnjHVvosIUxnmKJKwsEqHYZKOfwbjiCguao3DSyI7GFw40HSt72Z/p
4BNeGE8qZHZ3fl8OaFUn2cQtlvYdsDeLP4L7X4zDs6JIR8AXgrIzf2Sd8r1PdjQE
6LAurDzxf/oga3spDphVEq/gXSP/ZLcP2EMfLh3YdiobOuwgnV9wZznmIb0Ycsbu
gI74xkpmvJBCIKs2Y6/Tv/jEuvIXkdeiP4CsONh4BGqtaCVYkmz+QLerp5wjHeSS
rzdvOxbpepFO3EnPh+/nBuRLgWhBaWx4n2zwlkJEboKCz9NUNpmJ6U5wBZA4VdYK
nGtNzNvlHdsdAlgdcEsLl8HXdAOCEqGpreVrDw6luKtrspG4vEHutToV03i7Pd7V
Zi5eJCm00NGUhQP/Q1ybnzM0efQPPuYrymAaqFEmhhcjnhJFVpRlziCwpDI4lK7P
9edC4q5aVAbJR8LhlQQZZJVsLCXUi7zvXbSkgBcik7yrH8F+NsIveAWE3UqCehyj
v46JPsa5Bz7R7xIzoZueynWKcxH2jAwIzFcFymfoYcmOty+YpzL8+MbU5eJ3vK2X
OwBvPSqexxWTyDWGkBhIX1if2coe9uGg+quZyuruviG0tgl7NrX1Rcoob70w1CXW
xffCe6JYYDVFaKPue1Pl+SZchqs56DHzJMdlbcnrdVGtduWltJeyk1VLhKC0Wy8f
2U6+TQoBRzgBN66elYaPX24qIx9ZMAVF96W1pSwRvZXPEv89DUPpt2nKkhI5aM/O
ZHRMWbBfaJlhQuQNFU4vCPSG+acFO8EH5u0Fgwf58UwQaf3BocIzlOvu5WTabN+D
CcQhb77yeKJQR82GCxFoOqf+DZSOeOsghD1fEDVhTDegkrIXcSCJckUZ45ybv55a
khxA9BSZMVC7d8urW0TOyh1J31Ivwtk2nsxrg/bwfpzP9hu4Ayr4G26QP2knxP3i
mSEDXVwIP2LwC8WO7lLdaznfdQA7xfxHD7ZYAGCAhDilr6BZRqLruFEbngJZOZv7
bDt9PvGEOQQ9of7u3dVTnEW2KWqvYCAutdljVnrQLauzZDj0lljmFzfdp60lMpL6
7ZoICk81mMOOD8OrtYexFWBc/RHLhv2Dym5Fo7KtvPBCodQrc+s2yOr8cIUAA9VW
4ciRJkXLdDylrQxB0y/93NW4KqwwzM/sBAt5oSzY3Z9OoX8ffr6fVt7QUjKdgcYO
hMwIwGoNb74VRvqpMJbJLeM/M5PWuGCdlchUbJ6K296aEccQrVPnzAYq/a5eXihu
irnnXIR2NqRDx7M581CQ/BdW6MBruhvJVHJMQSQlSJOq40/JZm7UF/b6Lvd76PcT
pVmmMyCcYqcvOleQVJ51103H3Kr/eOEtb1PPjQ5svQ2cfeqJ86n0re0/UhMNkCha
cZ9CzDy7Ea1jLOPBQguJVGnlmRP9dPMNTrq32HOzO6qW6kEM7eDafmHxPVaqg3O5
Whe0XBqoWPEvpk47t+UjL1MpcV0j07bIqOydIoE19dmObH0uXUx4y3fmL7M4V2Bs
s4C+nYsDFvkVtXeSIHtbTfasHp5m12CNsnCtorBGNDGAEcLC4ejzeKsO0ngsr28W
PYjWs9HtrvgVBUDGox8EgoXAux+c8RoRnd7qBP76wcJgi+TMCZtm8/chD7QLoA3h
UyO7aPf7ksXVvDT8SS5BYxuXDvj2m58XhNsARllj5f3fltgNM4lwBGJZRAoKwFWP
Y2HhD4bDQaXIqPBMe/Yj7D0HZ12H8HaLlvVo73v/owV4SYpxIQvSqVdeEViL1nVV
IZ0Bv9b8IPIj9QZ9dEKxm8ResPEJ1ZW3efjvM3hSQjDKWK34wRuPilKUZM8IEFsY
W1NcrWAZjG6Qg86wWVTl2LIXOgvahOlA7jffMtXuxVrJtpmzLJ/5smSNf9hpfuGD
SGZc3EUza6ac2+8JHRXNe1Zz+dOtVAzqUmtFtsoCCjlzv1DcCUCzAm38EheRWJv4
GijS2J5V6l7MMbLXhHuRZp7bnGYHTGKT9deyE3ckwh/AlLkwBez3c8LYEXrSonJj
AMDXIrzyM5gmiPB8gULBi7QbSuoTffcOFFhIQwZ9L86sK9I/w8/gIQmW5t+3CvgA
IhEQKEzqOqaNwv5NPEuEVEbLSzyEHIGU//0S3BrjtJOrdKrazP60HXgGiQ8XRa5Q
JOmIpfSKQ3r4JUHZegSuVdxUbqP8DRVOYBdz25t4rE2Z5elxaARIXRoLVi4j5lss
GRmm15E+vyJK0AZ8KuqT629sHL1XvzmzKyFhSyi6Y8Msud5BEBl1FSaRdAo6i6Af
GzJpZcFDs5mc8qi7mkeh4KdKI2pq60OQQMhmKzSQbB0aSwBTCCzRD1xy6NlOM6tZ
27NwnpsgJk1f4Ka1GlolgqsRnCdkiFD7GsOfV3J2LcZCEbye3Fgqe3yxJzV6owbv
JioyR2/cLtrZ8o52tltdNQyAD9S4i9xGrdy76lgEYeAdZ2L0kiU569QqzXKu8FtE
rOqZdsjF4N4y7k/xzLqDNRwQPSDHYllFu8t3HRjJCzfZo4jgtmBV+n75jF7sev5p
icTcijJc2BYCC6u/JNGU1Vyv+djWHOR64+a4q2PeMHG/0b8Eu64kwymH4t8uQ5nD
YZfCJgAVXyPrW4UvIgogBmliR9Auqb7ugemZ4VV970ZlAOzBKLJPWOgQMw2ALzIx
hpVPba/mdNTIcvdg9WgxrS1RDpJQtxHslHyGO88XsZ5Al39RUX+RjjM8Eh2epAbK
8ovj38di6HPabST00jn9HKTJkAvSCWBHk99YIW5PhVjtNNuJnDGBt6GC89CtvVYP
FPShatV7Q+86uclZwNC54NJmyGNEtBXW3DM9KUT7MSY+10GcZBP4d6ex8oLRulVD
csufq2lmxX1TAyTZ22YcPQcV1JD7XpXJyrgCqtxc3K6qD7BfeMFWca0NwpT7ysR3
+/QAB6rOvG4ytkyMTGJZWA6Y5TJe1Iyk0EK2AsmK9776VAWRDqvMm3OHzfhEmOcc
UFvT3keIH4HE/GYXHOSuNvNLF9BVGaNAtd6M/IXoMMgM0swKcHlmabreMUUiuhJY
b15piHD5sGI4g649sZ8uyIXSILBF+XC7EcdBBOJH4NlqiOoYRY4olkPUUoClVxTV
vtWCTCop8PGexJdfCZzctkBMsNC+F8AolIMVgHkVS7V7xp12dhUrjTxfwKQy5DDa
MOLBzaqnO+Ajlb91BiWbdLRbzoBHB1nJtsOwrd3XXXINrl48PSGY/QvpiqmX4+b4
DhaXL/LNLEkBT4PUauZCRMgWfte4ip+tk+J5t9aqxrN0Eu2AFBdBlY/gb319ylE/
sU+prrNOfQuTJbWR/q8sx5Gf5bJ6PAPsoFkHzrP1e9MGCxUwADb97xRHZfQG8a3N
jVS0hJKWi++7BhgyNEHX7tdeJna1QqbDtzTUWSo7W5R6XNH/fYy6CReKAJsdUORE
RtmNqdgdc8qJcGsBViDksCigp8PIzJEjyTxuYXYMyLeg/11xRR/7Ob64fB+ezqnG
3KfGw9nkO9hzH9aRoV+VlF/Ka3KJVPmLEekCxrtxWyJVcReezPWYn/A0YIVXPXeL
KDtkUhQi70YyLEh8AUHXLiHfAeVXujE9YaEOBA6Rvg0yfLuEq4rSSO3g9mhiajex
BpKo3RRFgUDA35zlJRubUlBK8WdyWfnGu6ZGpB+GcQEkPSgh6sbfoCwBIJWpv84F
f5qF0QBHy+xZgjgEisxyQ0XEvPOC4Dif2+27pfAJhMcp1s+LIxQhTzBP6RZU+Mm+
p6aEJt8OTOtmgACFMfPWZSofLfOzYS1alD9Jmcwp2y/6M3X4fu/CMS7geiZOy6FW
CmZySges2FfTPBpNFnTQBv+vuuY4j/SoKDt4KvB7dhrrvrQRktx424LWhlXPd3cx
97T4ucY1+PA06w+IBg9y5jWRQ1L+1dt+2dxv0YxB+HySv7N7NQnlQtOmeUs698Za
CAH3qFfEFMEz1CI+iLJz8nRZsuLQqtQluc13bAmQhSNgNXfbCp3ozLAjiY7IP39r
4gU78QW8qp+0ZQfyeU5236Dgbpnfn2U3lkVVPgu3T87n/Mtm0ozV3jm24HdcMqfm
78/IKyCk+hy+IJQCv6QooYhTJ+2Q8bsvwuiw1cJPn5qTdrhDdGslQLHl7uM4+eRJ
mspYw25M6IeD+A1YYk3sf3x/4yvoy7rj1XXbZV2aWWn3UEifWBcNyEtfe23+a7hb
KLvzoWB+20rkT0iBU6jmfPsPqtQnhLFQktC18foYgrUjth6qa7Na1F4iR+lH+4vJ
mdvApzuNIQoDOvAEWD/56ypCdWf4VJtCxBpbZenrRg/Wlr0HJPmbkogm9UlzarXb
4OJ5xW49zRgUvu1c4TX/TWvro/IKNGV+0LYJ4BCxagnJpzYdVhxHgtt0Dhqy9EYl
uJRhnooKbQh90R6/LtHHfHAcxAr/8XSr16sed4wnlK/6s2L7SRrlfKBK3Qc5bdvH
yxSQSsUuJHtqRmHM00KrsWLJabyhMsMrar3W8dPJt+2uisqbOkurrEcLAT6Ujq+Z
2YDUMLBxV+ps7RTgQ3JhPbOIPG2BwMnjcyzN5cbrOmpQrbpdrVQ87ZUCVn2R5SaJ
92TrcWGpzSwk7mTH8Mt5NvxM73qt4O7Jvg/ZJyD7VIYFFH65SDxV8JupXPXKiAyO
ncrOeZRM+WETzsxIK7cZmd21knGdP1DEquMyGJrLbJgGUuTXIpCLudDCrDs4K+xH
hbmsfpkvycWgFwYq54ms7ryVluwSyMlEmjmENoeo8E4cjRkRfvVhotOTgNL+FuyL
A4VDKOxbVtEGNYGTkhK92lb0AiEHqQZJOyukeiP4xoG+wif0uf85OSSvYHiSRwXQ
mPIxmtrr0Qug2Fb9lTN1ROkgnNJ36DNyT6X+9lFcFdQ+RlbCE2fbtCBdWVZipnhy
Ya3eNkIIybvFpc0L5jCCRu6ohM+ZJzRjHjPpJonsIT3jQS0MikkXYZbrJA42LrMl
hTxHpqhhxQZoIac2JoHV+Ks+v1LC3JzgK3Z8plX0h3J9ljwctSDXUhyg2UKie4/C
wCVxKxxvxagYjdD/U3OQQqlok5srbiJCPC/SDc/Kr0heX3KENzb2zrJ0NTOAJJKd
T/9XPWh76CVwzEEWCm4f2cfr3T4xD8LcXdB4+imIRwP3hfL6sBidE+5WLyuZ/sRD
aFRt863Bh7oqUjEIFqdgbSTxziE7nxo2jbt1ihjb+5Qy4qnb17F3ZCvNyZTGHL74
cRA2Nxrr0q8wmPXTxLw3TSyW1+nKKjWGDHq3Ctu+xpMDHR3UOq6rL5MnuMQPRsW7
zkAk1wkRnBauTfc0PNFCucA1LyTPedh7hKsS/NvE23Zot2NCityF4sPNIsQqwCEO
EUZOAncElkfPHmjNnxa0Or4WHIipLpMvcsnaYC1gGPmdvNcMbN9FjMzmGSktT+3/
usv/JzKDw9AcpdD9JX/m9LxahPjLrRKGYRzVNKJVa7elIgSy/4vzQpg2zbypEmmi
4TyjhfItvEVdMCYg4eS5NcfPY24mTGkdnSY+0zU56P4iZwoDKupCflsEaAwCsuOQ
vrsch2YJShBwCtV41OvcdGFMBmTb4zLFgNaJQRGzS+w1l7HobJ8bHANfK05bHL9X
PqaKiuY56Lym1nxf+qJ3iS8JqbGLsQuYUWLqrMueCzZZH61/4695CP+y4hFvszZy
urOjn2BfFvivNHlx/5NvfRdE/z6cIHZNeisoHWc6SVHmARuuupXh5LIPHhFlfNza
r7HRXGHMrjtVqj8oSE15O9QMEZtXvH/stUUJC2AysfMpz8544mIFMti994ICmWJB
NyByYozlLqPhEl+Emuj9Xt47yX9y3LxuM0Xt1hq55UW5jiVsBYtB5w+HFBDDDVE0
ag8Fqh050PbYlq9nRo/34FJitK3wMr7VbwoFRCkUukjmEzC02mF0CkHz4rGwgeSn
agyyXb9SGJ9uJD60ttxk7SYo39KJ+LvrQMTd+LnS26OFDJEW2gj09HyxYRyreHtf
uWi+cPWzqjzjgeh/+/y15jcm6Ig6CwbZwfY4ks+UMcbL/DZTsf/hI8zL+YD/E8wy
9fW4yLnwG8oEK4o0mhxp6iJ1fGV9SGFflkmsAM0EMjdHkVMFaiH15snKdchuM+ZX
DqVX8uiQA81blhShWEXzVtPj92qjYZlPj+ZgEeaQ9Vv+NLZtJg5/vGDalZM/ebah
aWWBIsa7TE87kfbxBzp/cIm4EGyATEVg4AzXaDKP4EKNUOcAiGrOvfW+8rx/4d7T
l9Ou7PFf/Zqz3hWoO4MA9aQRyUFhrYrDYFvptYRqguK2YvPK9pXuCmpy4wfR7UfH
ChPaGVGI1GK8pfpmk3wOi+/fPo2zHqbMxa22w8LXrGx+FBOKZuKWuEDg7RzegLfl
es0STJYBtzi8enHhB3C1zfNUL2fH8GruJPP7QTO9DyneE/5a02YNVHLKSUniLWih
VciW/76ZrJWEQ9EvwVN2QcH2WuzEfZkxEuurYSYPmICfq433PpHD8tOedMfZOiaK
LGmgtyUfF81XXrW5e4xjA4LsRnUOVn/BFOhDW2EvjcEz8yH7xcn+jfRJy6KA6NZP
hT+j55tRDI5AfVg1d4BAr09U1gqArXVHdaJ0fvvEc8aZkAK5I7PwNpplzkrUu5jc
l77m3LbnxC9o7gWuqNHp0HJTcl/NcnljWBJsyoljVr9JqppyBKnrkjBEXKp+cC2/
WgF1p4i8wocHwdYpoLta9/wlMfNE3k23Ct+M3ie20xLUFb748OSg8YEsQWB3Kzuq
IoFvxfPqka2CriyoLbNz6XOIhx2GXPtSQ6BnSY6olFji3GpdSDwdlgKNL2PrQ/IR
oMOQBfQPqWSK/QcTscKBUAJTFh+xglFpnLYm2T/xoaYy/oRaQc0D0AS3MUccmVDo
1du4b4ugUSltPZKds2aUJU/MFxHwzJeb82f6jJzCIbY09Xg/YXHBT27WYShrJMPH
6EktR+bp7yPkBVjRXOW+UqLFNNyWWTpJmntW86TwtonkoXbEYCtPmxM0PrxILLOR
VG+CKcW5QKGvdHMTR2lT+jkqDLBXhyTgK59BdXyx63HcHynCFBN+smOX8Nw8IOf1
SRrSJSqDEoEzpMBTAK6BK5KCNeQW4HiJnemxdQzAv6CtWoPNupKGrPYqLR+XED1f
yrytlt7KYJsduhIlWYCWlWyKFF53CjvjOZ4Q78R6X9xDAPePtnCzQpUph3LIt938
Kxd3ENV4YuqqBxsbomwZ98jZD4QAXqSlUv/n6w7silcfC3BNVIk8CuTSTwo/hwUM
Q7Oj3QqdzNqRfnMMLd6SHrDLHW7/olWj92QUXIvoEaHPQfG+TlXEIpU5DWguwIvh
43TUTncqdOzial+zMO04z/1nnYSQEy4fTFwlU1IyDIou+h7GLrExo60gJ9meJYTg
Tp6jyRuV91qZHLb08RFSWUuXdkgTi9xgXAd6IS8IPOYuoIG6KlKHSAJgpTxldnm1
rcPmYUB7e06Sp+x3Bl8QV7jfxeiWSLLRsOIeCtXzbE0bs5xSPygAURV0m8FjX7+g
9Wluz+nQy0T+ZrIJIJi4OGhNjbFuKpgDlQC1/7atFvbYivcIB0vQoWKmpSKdXQ/X
/ZSDbZiUQn62/uPpJ3tCRqoR+pjhfKssO9C5oZa/YaupLlYsdW7M8Gi4njPlQJpA
1QVwT83JcpXAG6n2USTYADxTe5bhW5HEsaPf8VsbCHWsUPKrNfQvaTySpORcZ4Nu
DBnl4Mu0Oh5qsVMgaewhwllQhdolz+3QnwwCXtJceWCdqUhlnlvgN3OqVp31xKF3
d6WmpEXQFNtTxE4/+tE61aP+W2h0r9+ihtdbqJ6cfVAzUP/ai0ofBxsJ1EzG8/B8
LySlGtOnKorDS7J2uPEdZ6JwXTCLgyyNZoqblfckyaJS3cvE2m/fVyR83aaC9JAM
T+Yl4faLYb1OIynvyxD/nle7YE43yTs/qB0pZBxoNUCaQaxfP5qhcZ2J+QguEjc3
iIPTUts9KUKNxZ/vVhL5Ecs7PlGyU6L8IDKIoSYPws4fGJ8GV7+ZF77EJGckCwEB
USLkxEtmdXR9zjDJX5YA52t3y8SvmyC881y88EqcCRLpLnKis5JYIH8v39fmjQYP
8ZdQ0SUuEUBBaB6UqReqA9LDiZEOOxOj3SLR4pu2OH7fwMkiFzQ6D3VqzqL8kRyn
RgiXj1MfeFqCf0N/5QvRIDtCeUXatdUlCSCQsPxImGgWvauEXxHzTaHZlRa4yrT/
WqUxy7WA9No9hR1ge/d47/V7I4soQxLETK+FRmwiXUkL7vJH91tb6sPvFI6OxDQU
zDu+Sd7DFxxArPD4KrNYDyT3mHWC/9XyL+qLUqglhxgbiqjEQoK5F+JQlMVVYMI3
pLWiOWdyeSzmjxCq1WBCvFuc75thhVpgClDgOeTq6RcWFYlww1pr2drID/OhwN0A
0Ezl3YVjpi7/bJtfzZm8V+d3uXsMBUnZFg2+c8w0Q6jX7cR48v+G0F7u/GlmGLqz
lw3sGls3i9NNxHAreHx50KNIfm/hE0FPAPtiTsRYhgUTbDO/AUHXrqqQCCmNWn0Z
NFX2ililX15NBn2etT2hp0oyLdGRorML1Oa7XxpYfTIdSd8+bU56dhC+9eW9rJ91
zz91TpTD5TmA8keUOvU3AJt1mCUdAv/hYC9HjmaUU4yTJGUFKKX4QBybDZg/F+AR
zfsij8zIilFWKDSS6SIwbpcOI4flPFrwIXO8bg7pRYFi40XBtJ2DKGy6u1/d6Bul
oZ4LO2xa+voq2RbiyBEKKoVkvlSXzAszkZRM2uuCDl1koSzsykTsGCvXmznv6Mx9
8/gRmgKit6wlxUtMJzLz9573KLfg/9SCC3q4AN0A6QTyxnCiign3IJZIaQfR+fP4
Csnw2UB9wW17WwxWyNUmzKZXXvOoDdkk6GpJhIKVKSXSzOoAsY69+TowzaiKrdQ0
zF8K+aVTMAUbFpB7wFt+XNZaslRg6kpllm90Jgu0uVGI84UbIrKadHgdUJbv9BzS
P40QrVs6Ll/bqPm8MOQeFUSHeoi3gFgThIFOstBB4rG0l6CVATwHxj4Coe/OE2O1
Nv9ey4uknSGNplflDNYCUsKl/jIIz+1wyCB9VvglhrzmvqC6blZ0T6IsNrzVqUVQ
o+FrgAcgO9f6NUbGdnol5DvF2i4ZyedJKs4236huCoE5i9JmNowoYGt8HPTfrIsE
uLVhaVw/5XVJsKlKZCcOjQW69S1OXBZVZixmdPrCuA3ar1soOL6bmYkrysQwSn1h
BRwuJ+0kBUHnu6Z2wG+OIdD2fEmFBhj32+sZs9FcD7chnGyDGVyEEZ/r/M4oblVz
X9V1QI2l0nsypYIAFag16u7qkV/UzPYiMp6Ne4GfQMW7xQgomP9zhVoSgWXB1/+n
jxDgUN837gRf+oTKHxi1nbgQG/fEb0GnCJetxDrPjpLsqMQ870gtKk7F7ByGQQSh
R1L3Q9zdlbwAUEJvQc6GQIK+CPap+jTLXd7fb/0Tjga5qA7Q0ahtwgcy+/8nY5L/
0Heq7sLpCDEDlKwazvDpUpBUcM3WOEXnwD04BnAeMweQNat1pOFWf64U6YfaKCWI
DebCIa2V2ceHCal46M2Eo/2DtxTbyu4dZqGGiDNNloIuYlGCmgsK4mSL0vKy+oB2
W/w55dzce+Ia9JrJXQTGCoCg7Qxx80jJkG2gfXqOB+/k7ds9qg1jol7gTjv6jU9o
Bhvx7+5W4V1WHVlXAVRjwrFak4MyS+5DG2y9NEcsh+5ojZnX9dvICAp9d6YLCN/x
Lx0PtlFSJmVZa8JYjl49IrKUFtV5U+VUOwveTC9NYOGQJ2Pz6q2NTxXsD2gM1qsK
fNNo6uJGj5MAlI+fHafn2pqHiKPgtbEH95+60ZvwPTkgqiRatwPObhHuRO05KpnW
pirI7LeK9uUg/P8Fhs/s7bw+lRUUFdQLJjYA1Ty5FtfUae3cTLduVn0DO4y4EX4D
/Mvpq0vwhtPZxnjJGS4tduWDQPsgONmpe/OlhGaksnsOMOYgIHr9/mdTGb8hMHHw
pCVnLf1ICZ5TQNL0dR84v1sqL7r5I+WAcCZMI59zL+iEsjnhdpGLuOX1tOWkX+mc
2f+DD4q9ohjQbPhcUU/xWKcx4Z/S/5YlIEe7bYfcVD3rgHJCZfmU9nopQ7pmUQif
if/nAimxeFvj1aTDg3OINowleV7sqmg4rCFzqM1W2AnGEUejk35EJR962FU2Jbkf
DY/yBcTp7hzxnz1WA73CRsYOsdfPygiIGJp710QBDTT/AQVdfy3gmc/PzunVYW7W
rTtMEM1uKnfmVQs/UoapOisYzeru8KDORJ0rk4DiYw0FnmR0EHAJXNwlpQ4QIp6g
i8G5/HRe7yAOTSmQvRW+pgaKmqZkarXPIk9yq0uhYESy06PQX5d4QVLNT0/FLDha
WfaRWk2d6vlndfPgguYKSZCNeXvh0uWoLEYO6jUsDA+XoUJ55yAE8z5mqmkJzoNF
JljFWsujS/SPTKoLTNhNM9J7v+MkvNhVGC+tnwjyzXmMRazGVaQ9NMhHSdGMsgyA
bLTcEMaGYiHTCcYxyDX5T4WrTfhEFeF+FyOZB/Fwrm1+bIn1pvzDSo6R+0aV+hX+
QpUXZ6KNkgwrmg5CjwBIXH4RzRODpH2u/Y8AI7Dt5Sl7/1uZyzcu0kEuEBgazYOE
ylFeHQxgl9LPI39+2c2v55AUwj0kPuUP6kpHQFCsHQefvBCu1AgEWZpRBu7TJxVn
ZYDGRBXi5Ex0vE2vLueHGIVLL0lhWe1GYRrckB1mSX3MpzxhUmVGT4vkQ0VTROh6
78KuBdfc93tfIv74/gdopGAWWgPuFwGeS1WfjvFf9f6550wWLfjemx9m6s3McuwG
ov5Gvy4Of/vfPNl3X+zTxyd/QKI7XON+Wnz8aUXdCOKlrge2b11qRnw3YEEBKtGa
OlHhn2jYOs+ZEvvKr9r4f7WefrHOhpHM/H/gkA4Njf1woKnZJvJJ1SzcAq+X0FcN
er6dN/vARu+ITsCHIj07zaOoILrbJgkWSYQXaWFg8HXUCdUF5Nw7cKVoTEx7cKZM
vCpdVpsL6Ubcz/J+L1vo5CWWsD+KDI0RK9vjj++T4DqerRszwwf6ySmx4iEqjspY
FUHpIG2ciR9WCro10v9eHZxjkle925UquuELM79Sx6qm3rCXd2xEM9dXj9HF6NWc
OHXpsAUTwElz0d3dUsXKGCUMFiinTCK+OJrJq7jc+T6MJWYrdooGnQU91TiW0mVw
hLRWHTMl7zaNcP3A82XYVzlhgh42vegwPNkT+D8b5AKGQvsUOKjhwr2OBe2Q3GM/
DumX3j7bxsi2zdKEhLTnPZsu03yDfJu3FluogatFW2RNqtMiL/EguaIuVZR7kgn8
VaxI1lI0zwvwDEfFs1ZPA9yjblig837HBuPuGvrXnQZ9Wj9J8JABowQ3KLcccPa5
aUtae5I14OuDmnCX+zC3ZzBio520GMj6hnDgcirhAxa4BRx5wWSPRGuTYKlVPZ5m
dGlQRr/FfLRu0MP4kuwUKSswLKhP2tBcCicIOn+jYSv79UMnzpQNnrVo0NNZjGX5
72Fy9NwWTjb4yI7WXkI895BkP/IYfhrKhygZ1SEaWl+kOm3Zh9npoH09kMpKZ64z
EXoMAklFmogRa5tHTGHd946mWvqq2auMA/olkp5scz+81p93/kO2i4R7/mYxPGi9
XQF1MwoCqZcVJCh014pawhTOfchMV13xaNEvLW5yPIMjzvwnorMjEqzO4dUwzUt4
CCj/f25U+OOsLhooxGrjZ3+LpNQhYCvbSaB9DCSVwexUJPF/lwJlZsSCif5ZzZrr
D5jRdSOSsMj7sgNagafHNViTSbGpbHLt3fONHKyPAxMIeb5BD2dbbZLvXi6vS1ye
b9ZlL2/MStysIaHXmeqIhu9M/pTgcu7gHRMylUn8DIOe3gjlhDfdFMrSrbCUBp1m
NRJD92zdHtRud3IkzMDkBERGdRITCgfWWID8wr10JDx4F0fX5Xek4kSg6l13yIme
f2urOIl2gIyyVkX3X4pVUbWvXN8RMXfR4Vpph6WnFItBW41IQFtF3LpINm1e77tu
6nMusqSI6BY805OLAioxMtO5hYdKUj3H9gY6vUxl0fN+wLzDXSSl4GFEgk4RfGQH
pefoEUXYl3DNnljYuK4VtlHwh/WVuBuluFMhDLb+LO/uHTCgMv5xdJFDpmdbP+93
+i+lxRxbKQahFNa1J8B5sT0Rw7N62eRolanDTPChhmGw6O7kr2UIGgOaveNcqszI
NGWJbZODwWGqSh1yH8ulzY5DWX/YU5pPyq+AjlpdKpo9+q215YEzPW3pYL8MX1hB
VqVWOC3TUjlRtNtSxIKPnDvO3sHx+ZZkzqZqsf/AnaGlx3gGBIqIUMKCZOsEP1wH
h7576la9uzK/rG0iNA15rgIdIbacUPZd/WhmrFSpSdA+SrVPTOYnEL1V4zIqugVR
ZcXPVeNghGWC4tEG8JRziPdAqYT3HeC9IcLnaXb2Al6sAPoL+PCrBEBqM63iCxX/
KClf/xzOCvTpU35N/z5cN9zkNuKqYLx4jYHjOfyL79solqDxUgVkAMhegIc3srqK
iO+MyhBA5dtXmAJ16BsABwplHA/HCbL1eiYHRff6y9nGNtYijPLWbdHO0B/NYfAF
YDCpFVTUU33ZDAmHrMjGEU7PStAr7isywE8fNXftg6q3IFrdK7sfJ7C/aPNDvgL9
PZvYx/muF9gzdCsijB8i2yZSmAfVUhR3HlP3kMbt55KPXthquezAbJo9FmnmPsrq
5LB2GNqIoolWr/NHP5WEY8qQ5WW6Qtb9wVKy5miEsYDm2Y5JjtTivK8gM9YGxcf4
ha46xCs5Gv2Imh02Yg7Yj2QDKor4YlQ+mpE2UmvhGq+ZUgOdYKr20soHH8otuQ1Z
f8kIwb4W7RzAyyHSciyBXq6X1nhWRsChri/81LDmeoX1E39lz7O27qTJuuRLzKwv
F05jC0VM4C2UPXBt3yyA0cizLEeAYKkOnyaEx1LtSvA7TF/D9LWTH73IbVA0+UL9
2yH4sVunq2lBBKKfx/0W2pAi4DK06g2Gtt+2xdYmsFBALmy+Rv5OA/RMEndG+Mr/
mAFadSaVkEHFqmY55MAaosdEjAbOgi24/DocfOhKRzSMkP98CE5Z032WzZPcz0x+
qHiNMOhKJ266I98zdejIBO+Roj2iD6xHashIe7jYEiaXAn21mZ9hZM5E1hj9Ne81
gcsDqdfVsvcAv48c2oDBbKSsUxUM/NdVpKjqKCVolWp4TiBjqIow077jXM2xjZR6
X68tRpiEmZlgA/b5QrCE64hnzGaLBxQSFWLEdf4UckOoqTo+IX+zXctV1R2kSZcU
WBaSDc9ZOBNscvGwFI77eVw8sTVenilHOheyUu+ErXlV8TwdlSgyi9ERLxQelLXl
4nwC5IElmdFikb+61goaU1J/Kbm6wnmse/Fb+A4guk/jkfqOf/iDvFH9R8uersh0
uzBksW3W242Z2YnNmdrmKNuCsYiytVaKl0bEi2OXQ70Z+Q3KhTCHx3N/o2up0OEh
ehpf+1gI0gvt6+7FfsGsYpUtRpmsCxu1V/0ZKMXxJfrrpPT5XIZLx/FkoXakN8+z
AewDhnhjysJvQzo2VXsSv2at+bJLQMhw3PuaBRNH7X34H0FT0heNxVAdot6+gnTS
ZqX9LmakuiGgghFvR45YIJmZMdcDgUBnrIT+Isyc4nEAVIaOFVUgIId+F4EdLFlQ
PNpJD3l2mZvv4AFT2ipvinwCYBXgJUTtSlOVvtjaeZgbyWx+irFju8CCXPvY+gfp
EhQwwSWMatd8JdcdHGb7AmP5RQjh7BmZPsRiER3wPxesfdTkycEFpW+nHKfVtSAL
j3HjNPZNBLeKwHn6cNLXDbuztRP636tQdzWVoL//S1ZU7bCKR6o88Scg6kgP6L5X
AuGAxqq9gs0aKGU4ah7TQd82ZmC3K2HGeLTgWWn56OTUyQnyw6gC4BN+ocobJW6M
D6m7Ck16AFvnnY4pUE086MFWLKszhiUpDC0bEqjy+Dcy59YwjwvX6B7oyajREo3D
xPlNTWMfMzsvsmiVkwxqWDcTudzDxe4NKeWOgSVGS1k2VS6NfYAwFIugPjOlB3qA
7o2fUiDBTP69/OD05UM+P9f7zipbiolPyfpjonhNSptvCZ74C5PXvtivwYA5WW6C
YpURD7s/WfE+qWnOdJbFyHjjS0pQxCO5d+0znHHbXkc3IRO5PgBxwbqX7yp4EYyh
E+yWM53ZTkBZrxlPbKRiIjRvVNUDRAOhZ9uM1zN/Ax5E5p2G4ExuC170dh2KWQUn
MwCYA6Dw0oDXBh6gxmEv8B7xx6o3By/4GKMISTNtYByroDllmbWT6/Lm4T0rbdzO
e3CUGquTmaKHXSi+RebO3gNlc4AI9bwYbw/IQgJ8bhX+bT338yCMvBcNRVqAscTK
PqBf39HbsVsHd+tEWbQ5dikEZd7SX2v/oKCgprcCRK2d4jfW3dDydEMgyEMb5sfx
jbajTbr34C1daMUTRFUbiwWPIpi7MMzKGGULG86roQtdok7I0XyCRZ5FLVxfPsR6
w+H1Tb21gAADcOdPqdYWM8nITtCyREXLYv56TkubxfET3dSPdjH746P/gXsc8jVE
OLBVsNtiJC1G7vtngQSsQixUjPjte606DeT0+DmkDy2ZbTFnjVXc/XzpKOSRUgDj
hGnGPRrJj94WsqBQB0diLlfO3XiBclCLQwIJGAew5VsWYqDOc+XtY+lXIsYSJ68w
cFmsN2k9XxHvMYbXTBoHCz2vx1Y3PnWj9fS4nQJtzvGC6Xz/o/CjRcxDoKd/0uNk
KQs0W98TTX3FgID6TjTGB1e2ormT06MoAP92xbCHalwXaLG4DiNq7RSZ2WYzxEHj
uREq50Mpzy6OJZmo2T0vY2fL/7iYScTpiOotAH+GkfjGQChgNNr1NscjeT5KEr9T
+42kSVC7BxBOrpiNHLD+AW4kjZuKf6noWws2tEFR2FFbmPqtv2wyHqwgB7KGWfnc
RYMAdBt/348wi3BnxlrwflEgOngiMQkXmsFbA+Kz+yVKxZMg6aNJrqNFkTETEQ1I
waPZcAh2Qz86NftcEGB0R+b9DG/W4MuzuFnehLFcEqFzv8VJiizc4N0/FXoiO1V6
IHf9qBgUGekA7VcvuRyjN6UMXdv6VQgGFxPdqyaxmD6rDt1sg0Bh4X35UD2mEfUO
Gom12LqB+uqKfPQ5NUXdlLrPGs0Oa2icU65dCWIB6fzM1vkgHZZxV8FWFUGSBjkH
3JWYraol3voIdbI7sBzxubk1w+qzYnXGvIPX2xnq6ty/MWAqPPrbBq0/hFaSkcej
gSnZ0s0O/suFUITg2ByVpCTSEHsEBqJF6mPsL7IqBSDYRFSYvH5p3PoJxk05ZWXr
CAn8yXXtC5K08HWc3GpccJTny9kS/JEcyUEbJkxjM9My8OKQ0r5ZJkcSIlN/+N81
FNmn70sGZFcMPVyku4Nb11sARkvSlXIfn8dGVzEclgcuxiFZ6QkiEbw+QBxIHepI
oIHkNJlIQYKIDIZYGPJxOSef0X+qkMzHyQu/pa9phz12rXI5LPBwGNFmYHkarl3H
cBFW3H00bxW9XTiKikAFnYc+5/j8cz5XluuodMjQVokbq3heTlOis+IYZ6t6XOM+
9HZhA0Ai6rcITKpL5oZmIKuJKuvDVePx0c1mKbtpsGtKq5WAI5kKUCx93I15HaHV
nxuWTAWDXAChVruACk8dZDBtcjMNdNu7oHb+W6S1EB82o/vD4o9yNPRMyO6XFNHT
JN//XGbCd+tCp/BHDEmE2sL3P1Zg1+cMNwwhRTR+8byDLFYrodJ6UMw8B5ej+tM4
b2Caj4i0Q0sAkt2U8wD4yw3QnLJCkoOw+rwW0Sf4KZNkrCXkFX9MPCGhyL1z2ZBg
LH1QMY8PJo90uNVIfFaWpXqPzCDdYLTo0Xno0qVtTQ78bVnJx0DKmT0fJtOfM5IQ
AcbDALi2q9vviOoqgv0gf/OCPiBQUWDILLCttE/xQx9MkjURuNMDEEk8rPRX1blY
Zvraxryu/AXH2XZrn23AbWUIP3WFfdcRV+tAYquRLzqVm+cMKP+Nq18OVPTMeKlN
OtcmX+vjmaudJ4ZV4hkURf+qChhHYJU1A+qMw9+pGRwqxrGqhLmUcpBCNqDN1RRO
K2xj8bhRHnRxdFm6TOHJrW2EPhOrqEnOabOJM3ui8zDFuPri04Fs0BUxCSnmOfr6
8gKtiEw2wBqWpfIi5K7WTfknScCYBdFHXeyTGjJUMK6zj7ret35nXCiJxHYo3bmC
EuCvsjKcSye5weZ/yAf1CQ0vO2emjOElwbDuOsr5TIYxVu0esNRlzkGwMPP0XqRu
kVKvK45Z1p7H7t51C1n8RTKPUsI9YAv8LQfsQFLY/3R6ggwtxH7sehJya7one1Qt
mxfT2qnr4alxw9ztTqbNfn0VVEgvl5S907sPad12g0C4btohZGBF9iY3yuTbhlVO
sRQUfhMEnNv/ir+J7x1oFTqaBgG3SScp46c3Ul14EUWd6evpxMODbMZFojQS6B4s
QSePPX6+lVQ7TC/dkDWrYimHRqfNGu2BnsKMVWCuZrI7FoiAFJpcb2wtxk98Xolv
RGxetDHgY3nz2SAUt/1WHcO3DLnaVpS1N+2GmOZwtwfxx2iZ/2Mrtd7pgBqsjecA
FvOtfwVn8G2PrXJ05ympGQWQCDP/9PoZK4brp1Ty9L9cf8YnmMcxzHg8n3mm7ElL
ApKGdM0jj6zXf6MeGMPj5b+gXr1/npPqJOkWlJlo3ffW3bylB5nsVm5eC7vSW1E9
f9qfoLjrVkzwQGrd4MFkbm0A36akW6ysYl/0iUngCbZwWsdRF0bMDcU6Ur4E4cmp
K+iIj1Cl38NHumYtQKVwcU9u8qZBq97RTlupXxWxI7/Ol98ga3JweX9HKx+7EG/p
HNxACndAc4znXnTD1ajkuWu87Slv+fzY1+Z1WDw9OwBX+mxVr7wqOHrTP5aSgTOv
IJxmYbOlKyYTBbDXIp0MnqnK1C0dzIYN9HYRbdmjg0k53i7RNmrsY0JlDe7gMTyF
+kaz8WNTUO6iGqCedyBmsFeYq+wZpDj4/JMLo5pL6FpUNIp6mNl79apoUhG/kXn9
rKTljMHG3E2unRTktzh80kGnOmBSQwSCku2mruUuY2DUq/nAfOiIPdUQuuDMpU5y
cYYOMgKQB5QxjJpo3T4cDtUBb9nGZn6ZXXSjrcKsrfSR1MbrX40kxgYW48T191/W
w6GWVGLhAw3ZJN5/FgVbulkZyftpUcGz6xj0u2eyvrYtXBZAE2jKtRGjvboCsaFg
riwqAhHom8TCW/RuDWL5rwXmoes5m9PZ8+tPwsuQf1UFMfnBAcyUPegEkd2KCuwQ
LYngpPHvE2sXXp56k2Q/VBUpeSAMkfbabyoCGKxn/gvSP8MUOFwCp8yqjZ6BpK4w
Q3mea5VTdH+HkEt6acVKdjU0u4IzATOL1SgdP0QBOSqnW5L61iRTFK1Zc/EojfCc
Vkovqmce0xO8aFN526mdBUhLZN8hwY/vSMdTpiyj03ff/ajZw85QMW4ZlWMQyHQg
ZEfkduHcJ6GUz673mGWAywJje+6h+EewA5M5a6bZ0fOxpsx/FtnR8soSDHi/3Lxf
XSJIELcLwxfyedqu+PSJE+TsbxVJVB8yD0apbYzS2hlnv0HFEdb/RTyVcxqCV3Ox
QqX9/0s77XCgiFSdRLtFXxib1+73Rlwfh21aY/XdtCguMeoQzlmn9jec+2abNTie
HpkLyYgfqh7PLBGCDVQ2F1N9wTUEtbKqRX92IgH1GIrM5nBfRmvctQMCmISVHxMB
WdqL/piMveh1sOMX3cE649a1n+CD7iJjx9D79Pt+3biDWRNKU5UgxDgAPUUROiVN
c0wFGm0IzcVu6dbkdwwnQYXViZr5z5BqUMvOfPFftD3FbUhBhwogdntqhRifA3aJ
fbt+ulCZMbDocBk/T88a1vgBx6fDZvycYDHAZwYARbLJ/mRBoHyLBbT1f75y3ZfF
R5IAZbyB4lgS+GzFO/EGnZaPowA3eAdWnsFRUqMqKiL8eF3IRbePoRgXz45QmluV
a7I7ipkZFKpuVP7KG6yGWO8zLmJ8zNcglZMTr+frB7O9Jvw/tn4//HH0B3mtYe/g
0DscZKVgNob3McnJbGpA41yDP72zjpORUPhv46V0sbLxyMmbbu1TaN2fn7DzIJky
RunX72NMPCKFmrtJGzlnFKSXZ0E/MQFcykBspGGVq8Go8QOTmmB9WLS14uUfxIdQ
Usoapi+ujdAYZ3NFUrr8t1cNJtQAm9bLWzKUnJD9jFgKtFCqD219Ky7XjPwN11uZ
aAiXLNX+wU5+dv2C+e4WzSX0jztdNlVmuuXBa7SWibirvX1EoFHH80DWoovdAUJ2
Bne6IXEYOXimspUnaSYvRQsXQO9iCKtnd9ZCT2kCDHlm8tiLBLX02bhdWGfwtUUm
JhY7/EgTQBxlU4EkDpzDiVhynaUzqJIGPTy56wyj9fYGcbzuWUybB03CWFtDppjK
ygq+al4cEG2USMwNcs2zWpEA72mULv9a1x6xDUHo3L+NQlKSr/EzClisr+d0b990
71V6HnDNhhq4nAD4bXinwskiBSW8d9PucchrT4U72Nc3asI8P7heQFJsfOOqSr99
NFu0bCciLtL0biIi3uhVnPRdmXVYPu4GACHsILZEdsVkcl7JnsxwXGBDZU0gGHk3
4k0n/Rce859cl8w4FVz5UTvRlbNvIla+KQz2+DVQUF4vfTn5wLMRh3OAyMr1HRPv
eXZEYDiABA6ZJnuyxbratTMek/N3Ac3EUxErdgaHaftbLCrk3TePbe7Cu++EYUIo
Qjw2B1FtT37wIO5t7MghuFpx4iblnycCfz2iqwCf4BeCTGnSvgg0HNABoubQ+ZAF
4vqyDYMW2s9o1F94wlIbo9gv/9RT2W6ifxD30/bFr9EDRlRzNl5/UsQYZSkzQi6J
R7oHUFAIeKdvpiEkUhy1BMNpUBT79FGmMTGZTg3Na3F7rBS0kQLoru5Q22d8m500
vx4LalaOXd58irKqTFUzuJihTZwRX3lLvwESDmhPcBzr7Hgzay92fS82jdwF30iD
6B/CIMYC652C+gX+oDiXiCABvSP+hcJ3N+6Jv3HVEwRz7WHYbRccQRG0OEgmPGM9
2tHfN1JBng9gtUt2nmoDfiLszj4oljDXsCIL9j9hHdz9ORyQ/X65fzUtcR0LZNtv
seX/m9MfHHwiE2mNwflSxxrUGhiIfLlBq0/TH7y70SCq0NnNgo68mVfyH8qr369T
W/3vsAJSP8u3Y24lOpfUQszpLFHPSePaNFKfeS2uQDJBWjJrEtEcRm5q1O4IVwot
tcNNzedVywyRjE7wA4YBDlSL+b5H+JjJZRritg8pEn12WuKMANELR8tgVdNRJw3A
9PVtkC8Ryfet2r5VbODSL7dq/RJmA3XW6HuudFp0DWsdvLKicU6GJxB+I23HJdRK
BUAqNcsAbwPq77P0VEt5UOa9XF+yL/xJT9leWo6mkOzyj3D3Spmf2SOgV9MoWsn+
0VEugMHLcxGcYCPxYW1ShB06Zu8Lj7upxQnrUeb6lrTB/bNbpnRmqKmC8DkSHxA+
zpw5KRRCmYwCQUtLMSBydJZUF6uQ9K2YaQFnxzEPALOJAb+W8oltTLVAmcC3YdG7
9kUDx8bCGFqT2qS/h0TghFiNM1IRChHbnnh+xDEMNSlBhge+fO7/aX3LyrSIwwiC
Q8WhyzeXtLqtyaBKO/6pDQKve5IU1Wwg9ieNZrmkWHroILv/Vm35nYDdlhF4ZTPq
WctXVg0Cd2UD3aVoOUTtS+0NvKCMKJllp/4udN4PyEWQYkIjWnadirYxs4hR45e6
3Xv2q3TNVg4HsobH0/ljGJrwmZBuY/XYD2ZUj1AkWYZfIvS92HpB6MjfoxpoOfDX
+4DP9nZmgpvXn6iW+9KYASmmxHzpd8EO8F0a/fJX6wH3yTiHKltLln3SuzbVuYOu
qCkgGrIwM8DfI/JbB9cLuB+hKyTR5gyxDfETXKSxZTAB7SjQPvzwGkgC8/589ebw
lxIF/Eftxz8LCy/2zG2P0jXroQmYBvTjPI56rGi4C1xxuTOGyqMn0mLR9CNXmqdd
+sBtPmIKutgLLFn+7REMDTu4a//QhQThPPiPWH+68BgYJEAxwbT3uXHNn7TOaDxz
q0/VQK/3UBW5eC1JHekkONfrVrmU3zwyTKMYJipcLvdP7KESC3UCu+r1ogETCg4C
ayWfCiiUGZQGR9Whn69vuzu2xVrEmdce7PLSDifeG4a6jk2bog+YN1fktrRXNvco
gcWSATeMZTGycxolx1Hhpr9gdR1OEg3djA2HTMLh4YwdImdSMIuyxQrVKA6MNs2+
Tx5jhmzA0LsN8Uf+BUBJ/+8w+afXQ5d7wIsCC3znH+6rFav+yzwzIEWphi4xiEUc
LUZBlbd/eXM/gRXkfYVw00EFODz71PIQIw4AyfoJZjzh5kdMlS1wkx8b6cv2uJL5
fcB1psSWnlxFyQK2N/P9VboR8bigtFb80VWPg+glw+TZWREOEeGoAs322U+U469p
SSL46yy9a/M7JHEsBIEKrNItcQQGCtcXIy68eGGbuhAEdimSn32g3mBCLywNWqPA
KMIlEKOzABXZBvw76i5MU/ksyr54NDVuBHtU9BnKabZ7xXTHHF52xR8ymwC+BHvT
q66Kbq8vjG9eTZsYSAVdBEywGpY2aBwzldtS9Mi8FoZAwTqcH2ZkIXqHuNKpC4qD
K7h/GBaR5nethG7y3136DZkF/ZiQ+ECStOHgB11LHduY7oukpnvsXQTzr3TVPbmZ
YrQr4oQ8pbd2rdW4B2/psGftJAEmSjXjeVV39WO6VcSpcLfHBGVHUColYOJC+GXQ
WThZi03LkXDL+wOD4SP7aTtMgClVScJslYx7J394l65RwRjWpD+X9JD48ycUmW2o
IGEvsTShTCg5WOzj9j2kVzqphxWNLIAIqzMeG+R+/A3RHJgeg5inK7YibXU21UBL
pT7t0Xc2rfJsT3gRiMfBisi4xlsmjjDgTiqJEKbkch+FOfIojMARUznVWKV1Aux+
YO3yUgYXdjr4sYwhWnKAYOwr+LKr6E1aXYlivmMRKKrw7aCOT0Ykc+hOhJfvOu13
AqX6XXmiTiNuOp8K9Ct3YArCWkBYGOh8FMfWCJM9O60mm1BYxUfPJ66jqvFA0k07
gOH8B6+oOTJOvp3vRjbfZ2ilb6tNL1gAoZF00iY19ZtGEI5m0rlSU9tM3y3YwUds
TLcbJyJC1kthOAePiTq2mZM83XjwFjqL5WkumliKBgGIZ6SAf60htmyspbFlSwUs
a1m/IclZjngZtany695X4rECrEDMqBlbxSBBTwUiNUBE9FOLNivOukGoNkLJFS71
DA1FSIIu+8S7RHix2N+3g2mwh7JBVy1D0s7qJowEvO9pZ8SZJmKXkkp5fKLR3ycj
/lFYGp++hogMjNH2KoyfOd9Doc9TuqrXMVzJEBP+uCt7OlVY/msHU9Eca7IMgPJD
OKAX64lXoVxXWhlltG9/cmD08jOeyI8EseuO+jSCkgyOO/ycjK6rK4LhpcDGsK9m
Vt9Sa8eflEoGd/ZWT4WcVxL5m9/g4SYv2xbG5uFx4KygjY0GgRHpXLtrQmq59YLL
rkshkcAIAIYq/vJCq6cSpYzvqBoNKTK+30yd9bgOjJRpRFqOvQFjrlxl1cRJztxd
QKt0J3LVme7rDThcqvU8nH15z+6Xg6PD7B1tZJ9+qC4xsC6S5yMgkUeUDvkGHnzL
ZcQ3IeFEc/EPzQT+r49sliwmZXk16CAUDXKQY9o1KP/y/Af/RkrgxIUKCDMOUmew
d/hqMldEp/iSG1b2ODVfCRFipOkSwNtJVpopX7fzDfQFsUC4qfGINSyERxWBsX8D
KikfQDzFjCXj78qOXeZcZrNt9FVZ9L5yMLqrvCvB/s5AUAEPtd4OOp2kBnixCrfR
m9LElXN3dvAbpfY9/I81//ERzj0QCB7hbfMswpQU+OxkV3a9O6x6lKMRBHLiGBfv
g5ayumytzQrgxftAQdkhU53DI8W3ib3Wbd+J4zf1UbEt1zo60Z18s3qSUHMLhyNp
nidtn2Pneszf6ngCT54XNbQwe5zFl6cHw4wkNrdQWg8Xl1M0FfkyMFpFlSXXaODE
58dKeA71ZvSAXyyMWzbmeeSGAoiw/+a4fTS9KqJEWYQAFd6G5iMEsn5FdLgIbXYw
O3xsFKqjoUl7TMDwZmWCLHbdp8UVICk59Od4bLJB2sUe3vX0kQMsVXyZHGRMgw5s
D+HFJsOJLBR2dL9Z0V4SPcEqI5M4bpBFqPnwli2pX5RnNJw9NxtuBiCYhTP8pWE8
FCatjSo2ijyDQ4AVghQtlmbUMqyKs849Vx+dcOxApAV1fdwQpSlPSA1rqOz0P3t1
M3HJdBZWiGegKywv52SzrBEkcJ1UXgPeRqI4E4+qzWJWjDJEZuz94rUJwYXXcqXM
nWjN8jUiWBxECk8ijo89hha+jO2LMMPTGwff/YXvQ6kD1ZSiAFAZ+flFLwwUitHJ
Ur4SFBrTKsIwWBdljawI6prGhoooRU42y8z6IcKIXyaJMdStefL3hzSyQ5B55a58
2+ZatJz/8WhfyDmIAw34gZeiA+mfjBrO8ef56L3l4xOLghh+Hf413fXE3IzC/S7Q
vhYy7m8W4KK4+mtqGR/eUFFLrvuZcPNCWuwJNW0ctSMWFq6g9RITATh5CydgACbT
f0wxyYxBGnUGdAhiwvTVuM5kbAO2mYSjKOb3C9k+F7kgvb3qxF07+1GzeePc9LYn
oxtfCzLpFrVawLt7o2RVhicAzYkEgAKM5dYNacTylUOsXtGMNuRl3XeJqLLwkQkz
eYtcgPjuxrSqU+kPVME0znVIJbGPB7Vj3an2JVheen3bBOtheliX1/hAtdRiFYKd
s8BBsmdfUm8quFWEZ/gHT8T0vTvFYkRkjAuvXvW5H8QM+uzW/CtfXLyOcMyD3vpO
gtX3ouNHIDLkRufKRo0Sf8REWKuphJ50VlRS/WkYQP07FzMOk3/C53VpfbdiAIkQ
9Hl63q4xlrk+DLci3n3u3YtSXubICgQNFvgpLd5/dVt/ewObiXdbxOQX+LtaNdZy
TXSD8UaQxurBp6LIag9Rk5/fB0+n72ol6TJs/kCT7Yhk+JQjGkP7BdwA3bwkosfU
l3THoBTOhK3f2WT8iTzAcJZG4rnWXVV1WTq0t4uM84/mhnBOqq8DkKrrkGUdh2sV
TpL/9gPaiuc02COxPFR98K7ka1LydOtQZPzOVVkB3ktnMoWNSXRJMqS77vbVK4BA
8iPRf4mgpVgNeMVA5CN8OElmhBLExtwhOCvPaH3deoriwBh7Y6gjt28gFdlr4hkW
poZBwhXipoJ0YtcMGWAoN46rOoBQ4M/IrhTRI9T1Ps30HYngq1/p9EVR5Y3z2W/l
8IglkOePB9lrdQoghIHHF1QjoSg8L803LeXIOUsvRO5mNRuvd0yiAFbI1kAAQh8y
IHqmetrzxIMrmt3vW3thNSWd52WLw0RYC04arOMeC7aBQvT7px1JT3qUeaP0L+dB
v8ACG73lN8Tr1c6WSgkosdI4dLktB1L2XKPkM/clhk9JUeP87olIyw26Wrj1/5BX
ESmclwkcgpgB/VpssBWNRQUs8UboO2Wb3WYoEC8fEsT7NNBofNX0/Jax8p/+YMpJ
z/1f4dpsOh+PTuRJB06e1gGk4BWA8stzaoAcg2Dj17e8L3Xc+Y4cO7hYMo7aCAsp
BvGmb98Gb3lLF8sumnw0CikVf8LEXwfcKA1gj6p7Cf9w9WBxsVXi/vqkn/Qs3PW/
RdpmjqaK3C1ALF138PGfKGsySlucGFfTd2yjAe1s9DEg0j+YEP5E0pINHUiG4ADn
+nCxuAd2GHj4QOOSExpgujT45LMJy8+1UpYV3GtmFmfOpF4Fl72CSqBGeWDUbr0x
ekzdYU6w8Tbr0vwk4a9fif9VSRdrUgNetUIjdtZKnxKiZGQK+pFOI03vf4s2oHVY
TZJTyinzCz+v2fkDJtfwxi4Unc707QGTihN0SalOONl6EZ5+ptUETDSg2DJOmzO1
sqEOaph9tAMsRpnk8BJk8uRwM3lm0mXZH4tuIh0fC/HHlVofyDRlb1irrP8S7rhV
a0yO/BHRlSWyj9A+UTGHCSNrZFfSHym5o3/WdmMWmrSjTRMyfYmWXtFZar/I8PVo
fEpq3KdpLVXZjC5HfMssSI2d4ezuGCpDB8TXwnF5SG8wWmpjNlu85XXFrMwi/nut
vugyxLDKSZNrpffWkQNahGWcSGec9wrTVi4viPEBWSn2R9Fug7sQ1T9pikh80dKw
CAbDmexPe/w56YiyOmwBjfV1p3W5iB4H3d1nm89u2HIXqpda2fMRGkckTjkWcu+j
QjO4cqCaTMYt8i3ZnnXWKMOfp2H+/HQ2tXIMuc2XATx0JocNwCKtHebi+6HixuqM
AyBd0YOZch7av+iONv+BA5WN7bRcGHWFGldC+J6pvBkMTYGCnaEfdHCSEbwwTbX5
mennP4u2Ewjx7Y2og0q1ngogYZa57n1D2DixTHDEVx2tASS9+IH1YaeQxUFJmx+/
sft+Ya4vjjAHEcq/sLuKOrpOtnUKYA5S7LS59aNhVIssBJ9x4IAGrnxKYJoJoYE4
IgeNBbOQ6gMboK3scoOG8xpPhbhGLnGf2Wa8yI4snXQ/N7Y468TLb2rbZujx2ZQ9
1L2teAICg5jpfaXtkPtN4eN2qIIBDv6qrJ77nDmopJXS7QKInqUU9PbgOAH8re0y
dzjC8INFWRQerVNK24nGkbCmPkFqkxf/2OnEperrN4vMDDy/4KWl3XVJRjNTHUcr
RpJEVP8WcLDKpa0z73U8MtqUSj4qo8lofub2PRmjm+I+OUccsAu3S8Oj/eCHad/T
ZUfF1ToTzlkNIzU2nUuq+eyoQwYUS9jAFaWpJKbHLFRoPxzz93GF2mcy4zGxjJom
F6pAbu7SN+k78Am4eTTHkSOr30IsGCdYG/UKsjYQMACWxKVDsq00tRobLjsCD5QY
bSd0rtAYZoORqEI2jJoKrFI0hK53hvxK0roYrkV9Nx97qUykEEFtuEdIOGKamP3A
sfl73rOZL0lq3ms3lbuKHjIkPrs9GbUBvv/thRIhem/WZQDCO2kOypRr8s/cJXxO
1SMLbFon+mKH5RcQjxe3kGVpzO0xEpR5NLHhlbd1t49FUYOJkC/0RdbkdozE3HgG
l1H572jkc4NyhC53pHn3txJiaKDWZvqZqPYSey25iJHjRfpobok+2+/8dXa7hKLC
t6jqbyCOjwrZl2Y+y+gUzWv+9JPpUuo4aE3UO6Tw8/7ZDP43If5jEPNgEd4GYdsU
NL2GbLrcKv60BNS8k9wrN6wAMXTxsX6k0XKsaBPXK/z/DsJRrO7oEyYejcSBQdws
B4ONsggaqhqrO8huvcfpzRjkXh/3fQIflEin0sASrIbbN86O8lT9WsGZjcUwL5Zy
UrxU7ivL936hPCiOhQcyfdZhxo+/hF17XIZ8jslNeMPmmUzn9s32V2U/JB60cWJY
JWSVeb0iSbgI0QwVwML/k+OeTj7M6BggwmIxO6c2JkuqnUG5MVB+z2jYC8vgt9Ik
y6G0lc6goakHiXfOj9GDlr42SJ6MeQSSZmXJP1KWEROSp9vSNkfq+3bsAfCG6UhM
deHIiK1cM9m0+cDUHq1c6hIm79sFYJtKs2qqEEEVHDYbjhBxDAO4kKDgKHUM2vIB
VFmSMCs7Kw6ahUxskPtHRWiZB5P6z8D5bijZFZ8zUCajPt3TY3xuoX/6osZVAPtd
YAmgVFefQjT4iOTh+orKklhJkOi5CBni0l7ZZWvYEvMHmyfVKN8IglobAINSKkeR
tzopoMTIkAzaInusnisG/4XtUDUVvpn87jkaGHF1Fo7NwmNKc+nooS8iCkHE8CDI
C1K9qrS7yUAP8ArNJk00duoiOd5baO/JWCLwlJUDDAK/TK7wqpxTqDGATxM6SvVm
9glCsCXYEPtzV/LTJCLKqVcViSwG0+vqBvUG1tvkWAdPgzc/9wo7/Bcmy8V/6ge0
HBHSPl1kvCLvKaQyE3fBCadvKuEtzs7Uq4Y435VIDG1Yamh7sJiGPgumQQOmWO2J
VLKVSiDo+qybmOHggpnuuloNXr5khBq7FcrMa/yQULX78e9Nn+cT4MXpYajKELay
vlo6IcxQml5q5RlH5r9yK3OsV3c8iE4GWBBpmhSwJdwoGgc/3lT9l1zuq9qwdRfJ
KULW8T7S1mPVtT7UnHraYQNmw0yGL9F4g9N08GDsm8bezaDwyURIczlu9Ricj6HC
G8H4CKq45rz2DuprTiTLohaKoQbNn0m1dT0ByhJuNqFEnW9Jn0LzIg/+Iee3vZFO
4nr0ArVQlZKT/WY8RBsNUFFYvrb2QWfut0x9+Np+vX7g85XoSAZ8Vy9vRtZTK3YN
8msiilV4M0QvTYpYdhsDYu0+tARKw3K1CRXtAQTvd9yphNN9KlQ3gz4EPCwteUzW
DugCtcT6pHREkpGwZSW6k4qsoATSISiXrWxPIkkDO3jf0PmfzhcLiEV/laKlQuL/
deY9p2X2aF8aNraIcpNNl6IbrqYhp1ROgkR0LJSetBRsc1gEUMMnUhTqb60UxvQI
Yow+XbjqsiD0p2Nd5RLBCZj17oHthvnbFO9T2/CISVzTQcnDkIMo78aCRygfsN7Y
Hv9SKdoCJMwYAIbz2PUHU04LpiPPwJUgghktIoCHiSxhyO9huqPLVuTuXjFJZQY+
+6flFyasEkC3YBfz7FvDUL35Cdq3BfgImlf5uI2zCojhUtkw2QYbfMMKmyxl7/Qu
wH2I9BCZ7Ux2C6V5qaE6CwYT9enU0gBTWqvmnlJbB52pHpelGfn+vRijuE9mNuRW
4zXh5ujuSgrO4EekybcyKdGl0tOHGAtbbjBU5M12Fs77HWUK91RfDmUuwvgkOFC3
5+JEBKHb/nCe+ytm96HlYPvEwyvCRtH9eDquIPl0dIQEggd6sdAiqoWJqQGVgsS3
uGwNdelX/qv4bbmAlSfvruN61u+9ZKl5WmnYZwYwrcWpw9LlJwQEnCpWgkaxveOz
DMkYt2XTYmr4bcTCxcQiQ3Bwp6d2iescwoimTfWzS8kpOkIkMzN7pDrQ25/oxij4
/F7czlXAZ+wj5mLW0IxNMmpPRDbEpmWAVDWQrpk17cuM/RKjbA3y78/wWTf20L6s
z6Az4z7wa3/Sp/3ygX39cHKji3KYD6Q0nScwkPL9/YrGjTT3IFhuSVILaWFsY6Ay
NbPcWrD1+8jD3ZCsI4SUPf/mrcS58Ek+rmwh0o1UMQEOscli/1CxSTyqYUCpsC9u
yLS5ZXaVrsrEDXwrkDsVTCdtFFrGj6AuXLq5ZubvjPpbHOBaA8AQORaZfXafnf4R
89QhP3T3iHZm51DLtyvkzvE2nAszrdt7ws0La3rhISYXaqf6Tdh1XykJnqEZE4JL
E4ZaWw/jFvGzOVIdRUWr9b5/QpjiyRfl41kHgt3We4jWMMmi+X3DoNB3fqQqtLM2
jy8DBV9IUVmt0xfn2BmTsYU1Gtcj2iDq9FyyuhP+zFr4pqO/6FBsTzGRbp3ab5I3
EovPvjNOJeGq4qPc+MjGb2JxBSg3u0NLtpg8JXuMfvopSa23OyqJX1dHYc4A6syl
15O7zRKwxA1rt4dZrL0gm5ttph8C4rXRtdet1kFir2SQJp087145YkpG6nrBaWxG
c7nEvAN663Qob4XR4A2MEtmwin9kOjZ541oRh3L2e9Dt+4ryitOsp5e150MYFEMB
0SlQQLs8PteXpWSi151ZCSWxW9uF5wZU4eYCcFfzNbGZExfr/IcVFwCxMqxagrre
RNo4f68iyU3j0QN1mKm2kQwasyub+MysR5vTg0yNEZAn7aMHVNCP9tSbZj1AUODs
P9iCpSzlTDMLdg7Mvngqq4G1iB9pMAwEBYmvUPdphXF7POiQyzdc6rQ7rxjiMAVe
xx5NBaaGTm0aVsm+4Jk5E5XoeVYrliszs+2yf9jlNRWfIQvw9jZVSyz7J5rGCsMG
Fn6GsNR+2db5kyrw68KhXrGybJIV3/nbynAm9D8SCt9fJ5irN1sL2ThWbRpEIwBc
GLPrbmsNzgtJY0H/siVjZuq4itSYJli2mg9IloOt9e8AkNkDbZgsU79kYb1BL4aP
lYRO6njS6x41L/OnWEYTAFe0x9p21NJrku3It57L5CCWXW1tw6xdzDaJquBTPiFK
aLi7OrvyEXLIBF4oyMQ0F8vqfDpXCzqFgu4LkNmW+9Y5KOF0Eb2e9iPRWl1bM8ZJ
HUejFMnNrzpFdyzUXX7hIIclXB7JTFo/zzrYU1x7pMJbnZqdwIQ9hbiLi8Mt/Upw
qePIO1I4f9ZPLoy32hVcp8azTempjvTmq7+82GzXtI6Ajmgq97Xfw9ublYNRhVep
39RtrJrb2wM43ZqINQ5Z++YGugI2mr4wcnQh4HT7AQzRQI9ONAiKp+BlnNAhYgix
gl+3SFGY0qxXVGNiDqNiQdpv87I5nhK+NtSa1qIf5QbRyWaz5L+jXaYg9zK4FNxf
z/LxP5nFtcymisQfb0R38Otz6Yu3lSksIaByeZt4iNYLwm7WOZVjdDwRFBIQp8Oz
PTgMlMouuicS7nRbiSS0fFTsG+7JWFAJBxo7BkkDwotLQq2pfIwok/90OSW9d6De
gdCfqo8iupNywndAhmyU5KLsdOQ6gdojsnQqZfz3fJkN4CKzs3Ed4pD62BpTTDtm
TvNvpORWGN2IMCgbvajJzRT1Fm66b18hGp64aB8o17e0qUE+04mns4We9w3rOwaj
YyH5bSy3ujZLwxcIrC0kEuvF6EV8FtS4DRooPb1ajvuzpLmtfFhLJP3EBME3RkLA
rQsjrTJshnZGbvCjUo4fj4jLf3OxRjBcAjAaGkDFX55w4kvEsk+UQ5hBPaodnXs0
GkHU6h6vxgIm17L2huKvFZ1vNFUf4tg8ZOABLcPmBR6d4Y5rrUos/gsqteVnMS1K
lJPLDX4FuvcqWkGLij8diUdIq53mQRPBGkEg11HAx+R6WE3SiC4Jm0N+bten/1zO
ninRQSoTzMudh24n68/1x8frLeNDQjCCCtczfNPuf7mkye8OpuECxkWqgqKCnzwk
K8u3JDn6T5eReu4p5zviMNohb02wlVSlSA1uTaKDbcwI8kZHCCgUe3q62ta8v0sa
UomyNAE9uDy1D5t0B2pM8FYe1lpFTq9vpdzt2xeH8X8q92G6Cz85EyDjO91DkAcZ
CNzBIOssO2UsNtGHR9xEBltF3BJdQKJTrgvcFurpx79FKDVz7h9oWqWCYC2JlCHg
NEMq4TFKKjfQ+s7aQIvPKUMukt0LgxjNno5sQVlnxgXJHBgwv+6EcZtMeLAGB7kj
898ZE88jYiUuC+fBnu+LmY6NOQBN2+F9SzlVNOIWxGqG4VnAmZAt5mibT0451446
0f0n2qv9YRTOM/TLMvlkgbzVzjC/59tMY0j6lS5n4kjpRNVnJDPtr/eDoKkICBg7
D1wzqM0T1KbitLU2hTNc9Jg/90tW4YFviOvTnJH1H2vO8NYcD8JlGHOEzIkwkp3z
rBWblsEKZfrTQCiZf7RzEN5c0fW26lPceAkcba7w4tGjW0DwetZfW6zFHFWaSVJ8
JbUjCPHopCqO2TKgJHztmGfPXUgE/i+9BBW3SDH4r738D5L0YdJ2+g3zt9P9MSd/
o7pFSUs5S/XghLnt5hI/ipLJIUXFskBJgBrziRYiFsVDClKh5EEYCznjK946JtWL
qbsVgjkN2ipkRqfnEUfS5TORGu5a7YY19v1HoLAxWXhc9XJXXWsjDiI/VEfHUP3c
gMKxStKEcv0DC0Bm6ezCJ1a0CUIRJ2sYv7uW+/yx18bPBuLKOIe0bN5CYD74l3kQ
J6Hatk/bfQhIHCCfV7i7nTE34QSeqZ0N2/ddi64R8h40LYx6wfvhUBVq2QaPn2hM
lbLcPnaDTbhKxJcM9gx7fjNhHRRwfBHtFj0kze5N4VuCMi2+yi77J7OHomXJ+hCD
LP6wWRFrYwSrgEHWW7SklX1+RZgCCElstY0msIMcp33e3nVCrFOpekEb1iSEO2n2
Pd77gRAQt6LbHyTot4FogzD+V/FUBF67DIGT353L2aKtDbQf9evu+Gwx7adcPFK+
BE0JhB3j6aJgVqe+eDf6+qCOZbAy38FW0eYo6sg6/hbcIo4ddcBVrnFpSP76x35R
kddjvW2aVRyKNTL2lq7W4d2fkBVdMfOKwhIr1F5EDjoYQvO6bxZUUp3ys+KdcibI
nOOrSS59JxWrNtEj7Icw8jZdxOl1pzREm6ThvCp9Jq50nUqmnPtVKmPpixzKyVwq
w8LZzbt530kuxQWdebZXtjSZVKJi6sGFUoRQIfAOo8YSo2PIHbs0LeiyqJ9S16md
t+/pPRb9EDK9k/O+tTx/ih5McIg15sHHsEtdfB/DVHgxpmkodDHlleH+yaOA4shr
NLypYDeDDKwp+wkl0AVTSI1KpVwynPsUVtIZ2H6+qlqKpkM6ydGOcwKj2MtbQstD
tAkXcnnsVBlhZdDwqKuKjovrHGVQl704jWExfF7pg60CJZdp0WMkvo3qJUxnaKw9
2mQApwg0OtMhomFEj+e2EjRgV7yH6CV/YpuCGVhduwbviWyShfSgxRiH1MjQ3Jw0
uYgGBTGIqcvKqNHcqhOB3QfoV69AluDp/A7BrP866Ju1Rv2SjShwIFc2X+NevjWe
8cghwddoqj5llnkAaaTBPzSNKE7xKBu/i/lCgAQncdNVv8yftV/35InTmkpGFN1r
mWx1zrG7+utP+RwnVC5IoXpT2nfyUcTbOjH7hg2H4HC3XqEGMuvwkWM2QFOAN0uk
h0RM+a7UkpalcLBrsSdkRt7uFXJ4L8YSZtNf+XGRFsBI4egxyCDticaS5rfcRitn
oB1EXnDuv/8uDEWofGyR7HkzfTaIODaIEtvbIy9UMLI450vdoF1rgq1YMnR22KSL
1YnYMtT7YC7G6IgD4S83X+QMkJAIs8KSatomIQxM8GI+nY4GZ5oH2Efwr7LDRqaI
XmoN+5bKimUjMLfagBVkKkpwynyEa0O9BVZxVK7WpctCBMI/+ZT80U8q7Ydhxt/N
wxGnVYxOeIb6dk9qupotFk4ON+Z3PeaOfBiY/cgpv0tvCGRzJGlLOeYGWkNqFhfC
W0fwgOkmTV85uXiGOWwKmRV9Mr7sR9OqqTphByG/xS770OCWMtSbOxmh50W03mqo
XxAO1y34qDk3A68A4WoEXhKy34dEZkXZmtMmeVoyUhysjl2iWTEXcsuXLrwb9Pxu
hmXrgnzTCdAQMWE0JvgxCtFFMz0tAmwXz5G95aaG/3Rf7B343rqSXeLyAj88YSTh
9Bv4sGgOVLgdqJCPDwJF85Jj3gnLE513JyF8jlXC22UZoT0ppv867v74oxQcZvIn
Yqt16HHq3LJrfcqKTYM2Lln4tS3cUHylVOWt1+6ODyQ+WH/sZVuID/bs8ypzSF7v
avV1N47sk8EQ9EZsv2Px3S6qOpgR1jWqrw7lG+KMDYGUd8AEKBVFxBHkIpRcTJ5Y
Zw3kvKevAzrx/W8EgC5tXIIz6bbd88ckc7SNJxdasL0SMdmZELZrp1ZfyLk9BlXQ
Cpf09HRZSc1Dpe9zrE1zd72u5y3RTk0Tjv0GcT5aIk3MH/+x7CPSdzwNNNHL/cIG
BXUGLskkVEOY5UykV9lF0y6ziE7wn934cHmel2Ww3LG5xzx5plb955iNLhBqCucg
hFLHJ6RrHslscrIFpiHD61nE6JeoZCKk3lB5sHUGHw9FLUvyCJ7SqI6r865saUls
Xae22dyOLrstItDoGm3nOEu1paJC1p6QOd1F6Kl1Spyyx9TfaPcgJJgptDMmsj+O
WetfBF+NMZzRg3hA5VIwzayj+qFy8mHxvSsR1oLDIKJff21xzsulTvlEyKbNNwdV
u9O5GncJeC0t+MMwJPCSt8ZIH4zzL8CAgtO6A0wbsAgYIXScUvgVnoJScHtTp08q
feae7XrLAb7nCEbUglw/MgS2m7A/Hlrj7PTuM9RwksqHU1e58kF3WCY2S8Lczpdz
H1tyyLNH7+W9I1ssqDTz3l5P6kH5MywfrdFxSlB38NdV7aulLq5qk1AY0kKFSL08
tHKWKUT9sDnA2TeRPL2e7aR++dkzziHD2WLcQMfUwqG3PnfcCwDBUmhHJRcB6WDz
Ff32Jj7XZDqGTLFBCBMBzFGawJiKsVr+7UI+vU2Ep5mL2Pn/oDanYtC1lk9Ioh74
tP+9bsr10azuXFGOHe4e44668aHT8B1hZ7+mqwPkVqX7+q0619X05A7KOsgubTJs
xxpZJcHQab0+lzO48/SSULQXXgGcw5/0kDo+9q4HSj0GL5FL7sqsri293OlOtbR0
biz663YqWKCJsdn792ueRFbSkKqqqvT/9NbfnGsJWnnoZgoPr8AZP4wTXwUTggmI
Rf7nslidA62U5B7qI0/IfU7om2jLirB91Rvvwo1VMegdx0l/+rEqk1pAxp37jGPa
/dupxGawQLYp1FB5doTePB9p3spS8FfCO+tgXS4grsNg/W2s+Ai/iywKlryB8JKX
z7u3djCG3JtB93C1+Mr8lTdykdhZFAbWrcHGsPyGgCPzQwL4AJovJyrwBknYZjkh
dG3f5Mjc0hp9OUqnkS39oI58E9rhmMSTZwPotLi6riGk4AHzsxWN98ghrgvd6m6Q
i/WAopkwjoe/jXhgMznVwjqARSBLf+Fc2NUoHARFHsp5znezd/7ywhZ9iTO+wDV0
sEn+7j7Y3MpsgN0s5092VLcbmVyOI/r/dwQhELP6o+44E+8DDdDEKPhBnbB5C4MW
pz45CEsLnAFtV0sfzQzRkTMJpVkfCGyNlIDSa5532dgF8X9NX3ya+2aQof+jJ26L
+HNuuodhNcsQK/fqZ7Wn4e8F3zR2uWxjdLpX+vrI0d4pL+vpV4OUv/JBC44DEYuY
iCHew/m6GIFt99D1fkUOcbfLDELXHQ/fV79bp3Q1Mgy8pU1frfloQcDq4sYVdwda
lYJUOpvZijEKB5ZMnprizQKxEGnahW5I6hkZHB+cLK6YCBvvjRLoB8w+vWLHErxl
42GtEEZcWEzENoN4GTe2ugo38bIxXXZki5LrJvvyyAUv3p/WZqdDPxeblXJvJOqY
l9+ZmTpPqcg5spE2W8lGgFC7/Sx4bbYjIoFSrBHVAEmZBEx9j3jguf4PM17zkAyb
orrHoeIK7bnYG9RlXHgC8X5iQZm8AAOoDSpuJ34e3SoNKo2gx4bwZ8Kg79fVCZLR
QfJ9qQrONri4ZRfv6vlc/Vg6+q/KQyJZYXxz2LSMnbyZLuDgNQ0I8cwdHNKTvEVj
yboplkUVb7othFnsjAaeLQ1YjKX/1SvT3fRtOeOqbABmCL50jUeclGJzlM3sxrj1
K49uRzSQn3K7ju9c2oB2dGv5WcyBjtyQdgGqa5HABTWdbZY8tHMHuTQF/gJeCUUZ
Agu/JNnszUM2IplW6Udr+2lkHmRrHia8JZIt3j7pjFNc4l8fLGN+AtB8o0by0e/7
qMPO3p19xLcr21J8W/W5bhI8+cmmEycXPKmo/Wg9lZB8rfgML0UG+hcv0+E50eYQ
w/iT9JNJa/IJfEKQ++IypJ9nzjrDlI7YjjJK+uGnQv+726DUxv5dEpz5ERfUStwS
G5LqcUJNoYWOl50UndeC3ONcG9wiYNxQCF8HCAMumH1McRQTjycyvZanMcJn0LCa
dy4jX7OKEBtg/pM17+ldhA1q4lLkQRnMoLFoWgI5rhjrEH0QiIGePvJA0AsBdBSv
5REQqYIRtRW7sICO5UGPZUXXu7A4YvWIUr2b9wplsXbHonOwToXvyT3Yzs9W8/D0
uVQ6MxiEhbCwpxzeswPsr8aTUw8bo2KMIqaDAUDE5m0wF2hWBTVb9NuOyDRnuGz2
95WEclCKrxxyDK2wzjmP+GQkqY4gbRMI3lC0wKrWQd3axjClU9ddKu8DzSUGJ06L
TmuFpbFOIDEB5gF9alG9vn/57Elk4gXew0QWisdcZyxKT1JsXPHVeTxyjjNUhKho
pAPYN2P/kfReuPnLsro+O12yXZIAlOT0WBwgT4Xy7JT0yg6XOZbZaLP7np5Y4jKr
s0zRiW2vYyAkXVHUuXcw7Gcdjm8X3rOKaX9CR43be9oWVsRCzw5/P++z/GKKsS2/
giTeNdVYIOH+33vrsjb8sXKkLyPPezYAcoOvS0z3yv2Rtpar/bbzJFacctYq2Tea
e80L4LZsfr7/PzHQxlgp93tK7JmIYj+2kyHvK9mgiOiVgZHmPaZcjl7kaxwWbNOm
/pAAb157MvQyXAZCSdcTDEuPOFdUM0+9V1X6KxOzxCzaOLGb6986yLRFvy63G8lu
C1o96VHsWlrS1QCloEuX5iKYQKq8sDOIk/0ZavcO5YE1+VmU7MD1RyOjSE/HTZh3
2WTyGmdplAOziZRAGdIykdb0a2egCNPTK73o4jmWDnd4bc3yl1pa09f6g6p3U52r
Ar0dkfdQvl/N9O7wdx6WKnODlJcrAm+e4rOYmlVB/t7550Eh/ylAfP6StGYh9cEs
Q5M5CCmRGI00dQDtkBIFc5leBySomZsiaVjUkj39JKY1ATtB80kqRdTrs2SF/Srj
cVFIGwxq/NmAxtg+n4sonJszfEJvfcFWXvnnJB0WtCTbUSVxMN9wz53oXpcoLJaZ
8oCdyj68ipqi4iBvQ/xQyZIiBi27Yn/Y1rdHzT+l118xrD94xZuhqs9ZGykoGdLr
apcLKotL9ppXRDvVXKV68raDQTDDut0xOWAaC0FeOMLltPe/n2LnaS7wGtY9aMDs
pjYyMrVQPQwfiy+mbVzaP9VGVXJYamQmhxiknZ3XI18mJG1U8derqxA4WeRXOPLn
YlheMqKA3otd3wvw0EkfavWhbzsm/Rs7UiLqb2zPJ0IxGVpxuRvyqbEFYBR5cUeL
piWAfTA6SD7sg87SSZ766l2VtOdJVKUcagTehD68Y6TUjM2Lka8lDnWx7VId+e5A
JcDQEupdsQzLKYyyZ2aPmJ3UsTdULXmb75U9L0q1RQ9YLllpJJAasMR4DIfdSa7/
l/4AG4upMNBM1zevP41g4UoZ6dKZJ6K3vP7vjN54mRE8pW0xQWgnpQ1UJIi/FGrQ
MqTBPxZx6SKFU7TenGlWppsFU1b9qzRt1AVadZE5Pi4pLNkHJRE7O+NpAIq8xq+x
VN0uuByopC+Er/hYl5lI28iHkYunb0NBPLzo9Q9vyUigtYsVba/fkEgptWi3D6z6
iyS6cRSZo5do81MQ6YUplDTvaB6h5+2dV66WHagOfi7zmHTAmK/F48Dm4NxzM3nx
WEAYguWPY6WOiR3pMN+NtKnwLnP6jGcDWSPWBuccatN1rpG66pfhYYyaQr7jaSTm
Fg6g4gjVpnGJwSwdPkl+Ui7HSyRs5fZwUUXrnA5zhtIYoPd39Rb9ozAPMQGblxhP
eTJoLMykCbxNpdxQ7GQbzl1qUms/RhAHhPoYLhrE6EwysIjauxINmbk7JSkPt81n
1tQ3r7i9qAL1bZXHtnqq+JWjjFvevNjCyyNra14s3yLfItTI1iC252OBCGggSHkl
SNfRWBfexQEpKgcYTA62P//V5joqDDG3SqYnqQgPDlF7gUY+2P69Q1vNjP84hNdt
oHpJlF0TPS40Q5wRTsuqROY98S7IkXYPU6PVkSgLq5gGQJ0KHi3MIEO/oqd9pnRJ
ePSOzI3EJTrT/83cvHjLsmWIME+cX2na+2hQle6KPY+Dv3JlORoe2hpVwCB3hSXj
lJEtPyMWzbHibXLXbtWuLaWWCcmwXrZXyNWFxw1mnHG1gtVo1xS+FCBfcVEuSZx8
G+fVZ81qfmRuPnkHIsFCkZ8AH9bJtq9Mc7ZBr5f6ZgpcySI65wL4bh01apOegrqT
U6Y8C3Z/eo7pAfOVSI7A/DyABH6h4tha6GWEPGbD7dS4A6v/fs4xV7F2KIugP+Hb
zxNW+YEhhNLlGy0sp4UpWGDTV0fnH5O5AWYcw+vw4NBDR9Vfcu+Uvk5t3w++y6Sm
5gCe17WbGCfKplWbe9EgrK3AWT8VAVoQ1aw/t+N1M+UTVM3EW2WFOVK/wMTdNnUg
eQocTkqVoSw7r/eFsspgRnol1vxcOOsT6/RFV/bmPfoqW27t+R1zsQdwo+0RgJVo
379O57AOHuEXN0Iz5F1E1/EBQImzEHvtO+eK8qCmQeTOx24x39LiWeAekcU+pRQd
vZKVssxnhcTbTeG1mHp4ugAhK3nKTw4ID9yexebIu0TwCGwZJ67UARac0QWzRRE4
h8i0f0L3Guj6nkw2+4B/Eze8VSail/4td2g+O5qcIGPuXndNHqllqArBXMW75z91
wvvroFQ56lblQC/oeMYDnBuMOcU/PX1dp/1lebbexwr/9l1S4a0dYHHAms/K3/M5
KnR/XDH6p5WhEVT+vmu/fXJGMb11B72P+C69nlW+O2wFMaWn4c0ESOwMP15qyvXZ
jo6fF/SIiwBOkJ1RmHHNIpmGnxCxtf2QTPiWKxW9z2rFjclpuXDKMGzBe+LTYPOh
QnlxvUpOYyWaYKRp9fD5BC0mZ8ot3TTDntAnU4frI+QHvrReQwZPNESUs0TXBsCi
f/1w9ezNJLZXcyhz0l47Y86mvQybZHzroGpgPynGTOsl3evXY1iFLrhHjLALvaVP
0cgOp+GjibTqZrIIfnowmaZvweNwDUwizZo6dRMdjBujSbqW7v4islI6wM3Ap66g
EJC/Kj4l3fbRXfxLI5b4gjNPvTBEZsIofND681d8Kjf1kQXc2lPiAwF8N9Wzb2J2
Dv/8UAcHXSpOJjEuonQR7TLwMEFd0Wiegrzw8Nw44S4r2pQGNnI/7jnjY2qQ4F8f
5McIjZQ3I9xMZOTsd+JasLkIzU6GDo0e9Ub6pREg5aNzx8gRBqngp+yK+7XoV0Wt
DUN/pUEaP4fvrKe4BmEIEL71DY6hjYDVTqRfyDZvbG1KRkTJbhzbF2uj/mcGAkjJ
bsaEyG03hS1NbHQ545tc8964SwCS1FYCeE+I3dleIsHP7VzIxfjhnaIN95gcRjdR
GAErKTsjbrZxKPz1+ZZ1vXMnk34yTl277MbDQ3Y448gnMAJeMLXs7e1jgZMqXnVC
bqPs9eh2miFObrL1BGDrp68uJCkafzyNfMVDC+tMNQp0LRjOpajOEn4NQlKknFNZ
dEPMxfsp58EePCWZy3EYr0Gey0QUIKIuT4cozB21bsauje2E3mwfAuNXdA5ETZHT
kE2wXQz3c7tpkROwX2b6uOYtBAECk4vidIE5aFv2S9Asx6dOYmLus7H4t42PXHzl
EE2JqT/5Di33bgd8oAzeXL+bM6bL3R63gqH9EvYYWofJzw8pEQaXKvxy89JAshbA
MH049kirHy45KQhvTeL7lQLXZvwCae2Ve/VYf1L85cEKEqfloHCpSZovZeBfI1Q9
Cv9fRetW8M7XXMp5L5R08pXCjiohlv1BbKH+rjTiNlJG9lPHhCXWb8+9xum1OBaP
q8LeIJR4pJCvSvGfaz5rzbglqaP8oIUjnP/Pn9AVUXodm2Tg6Aw+POwlIoDzBd2x
BHEwW4Ivx3dGRNHVv4tZMdAf6xnaRvWGpmj+wRNNEikiL1Sy/L8YRZXo2eKxb5GC
ALvVFxAOkQ8HV28zqCCNA82WgdS4bjOTn312T8/0qYJ3FJeGb0CJT04ciQzA3CMf
pZBdCsC73D5ybiCuZQsv/GbfXVtYNuNJDJWeuqUslHhf5mGlqKHM2h8rz5Bvz8IM
Oqi/QiHBOHFK/snngZgVkNzMddYlHlZA4f1n7uPlbDyd1b+bxvnLEwsUkl6M/ZAf
OVcl3LgZznVtb9nxXgu2An4USrrshigsFp0/z5OuCXnTx+XOO8loHqqAtve95rSO
lwOb8Ht+7m/upuCcoZM7EHMOYZrg0Opje/yM+O8cio+Z2cd+RB5L+CBvcZAjvxgr
+OKT2hVp9IUyBAc2eX/6cap20cjzVzk7t2ciKYPy8L5z3s8IpCM9bZE390ebLlGq
9Zk0lE0LdzwaoUQ59J88ZGeYuBLkjHXQLQpzng/VITnERujk916bfX3FxbBAgu0r
F8pHgTCIwUMXdyCCUJtnzA1I3TXCPNprnFckU4irgWz38XQfW64dtMzIvL1Pa6LP
rmUiC9JvBU0WTZ96+UFa8Dz8KjYg9UAAtQG4ANbWZ74BjEGvLM9Pwa04MkKQGKG1
DdA7iygfIlOzyf/36bDjvXxYYIHnLMJIHnyyMjt4vhcbPOL1U1Ir7m7rBTL/cWQQ
j9X9nLu/Hu2lqmyF7S3vMg0903rMT9Uu45bDfQpH7XhnB1oxG2tjhBxpBfPHC/VP
evMLVTgugffgsvkZuXhsyIxVy7/IEbiYOaqaDz4p9/4zmrDWaF6C2TA3C/JwxkqE
TCqeDoutptphIu7c9J3ZcBB1ekP8eo2I6tEWCdZpbk3gnLfEB598g5fb9TKzRYhK
ev7MMZ1SuN1bwHWOPGEjHqvLQTfJM6Udaq4GZ+pskQWuX9K/tmk/TwPk9aOZWtND
tTEt0oOoHKqm/jWG18Gn8//jgoYsawSnc4G/O259sH/Zoz2Zaqa7QpMypyB9hhvv
nZFTZ2tCAJcx8xogFJPTmH1dXU2nEjwg3y8ISFbV3SukRZuJn1t9hdlo5seOn+85
k0KRBIWaH7T5PES5m1a3EsDZmgP0o04kuwl6muLNsfYERNITUTB8J8Bq6FF/p2P8
fIA2Q/Mq+xFr+pC1dtFyrNyY/cZ9kc6eRAmHlEc1drDqtCoVjroxM6P9YL8BPgXc
PE80YSklbD65nJwB9AKy/pUoLUxVz31uF74CH0EmBc6pHdHs3whHD2OLe4Dtg4xV
8xIPvdWHCKSddV5G+e57K2w8uEjPmE0dzv8mZ/VSZgrp/7sV+xIjxpSpZMXpShzd
y0IMTmmiVa04j83bln6FusciphjmYw32lGTN6/3rd0FTL4lBxhvVlQeRZI5KP1PX
XOZoMkAEfBpH0NWQh7iGawUYYpuNasG5MOo5q0zzWq4FWr5LxMN8apLgGiCWJip2
djGcGcOhFYWGTh9o5FgGDoRT/G2TNndnxCGh8c4TAnVhdcpZdvAmKWmKv9a+49Xk
4IxNdzuQgpee4txqjfl3bVQ9Eukz5Oa2pv6IrDpLdbWWfU90JTnT0m2BuYqk43Ng
9jtAemMc8002+s6R+iZmrt0YVwchu8PvtuQJdMQSmdp7qI7jWWtzyKA0xr52Xqzh
N27JEAd32OyauluSjwI4s965JIrJCeJDRMifj/d8YSlKN095S5pGya6gUwxzaJSB
8d0533tNXQ/eNqkh4f4oBN2GYqF2LnWuQLpsK8ek48jSwJUTH65jLjDC5LBW9Ay8
6xPMB8MA0FRsG0VEL/1fTnfSFOVBFc9i0Iqnc7L7IAAsPiHToFVdHnj8AfcJ2V6u
dYWTHTyZO0jvF1Fp5kjSbhAJwk+RFSpUE07Fcpx+PyAeA32iF7uNSOhK8gOHbUzO
1xDrhMgts2+gGNKCeV1qhpKHc8uu/amUVfE0r7QFXtE1w3z257U7nOj54gr3nvaj
hzEBEham5bCtjTHzy+nEaOqrwtjRbpZjnXfAMBBRhx5IZBYbP5k2ruA0b8lICxXB
ra0lqHaVAdcqwms6BvU3iWCV1EZNao6plsesIWxhb2ZoR1oIYSxqSmAz9JbtqqaJ
AKTJjMViQePcYX4XhXk+qYW4d0DNnkW7VnuDXIyLX4RTxIyY92fN3yq/Iz/GAr7v
mQqcHGKRnAhRF0bMk4ozOpTvTDmMs5BqGO3ARuQmA9kY+1oyRd9D1TH4BzTogr7A
gi5qeMJQEcy0bTuG95D7tfDC2rCPqKwhjKZFC6GAE8c3j/tbHIdByNWD9Pf3oHKC
OETDUfnpMdP0kVXJBYCu3I004dETBXhCtgBc7Riwceh2aL2bq473lYxOKMAA0OCE
VtCNoHCpNvWLfwWSg8BEs6cMmV5Bf1E28TIkaW54hO6XBfpb/kj1BcoeFqiVFJ/C
WL7MFB7Q3sdFwB7go+v+Mt88ypUK83yCfzcGf8e3uSiRBfsC1Rzih1INp7culdwV
gGbfZjQzvPqzWVIwcOoA64OeHii2gfWJ8ak8ggWINdo19V1g9jA6TpNia0faEJyz
mz+JCWcI1l7HWLYXvnXv7Z7qPsZ2lF6qrTvaqZhXnMSVnv91JK3eXb19yWjqC2Xh
uvXOsj4em/so1qg5eqrOol2wYhcM2GagRh/H6OAI3qxV/zQ4wEkjpov5SPJN5m8i
hs5SLld2IvQY9EeNjtziix7TRobZW68rUP85Rl2yGetcLZ7DKan7u9TpRcumlj3m
OjCiy16VxlvwRyrsStqcmf60A+Ei4wbSq8qxY5f6XA2qFLcMBBJIDu1M97pgufBh
MNT6g1cNsHXvh3OxI0EtYXxisxkQAVmBhsne6yMWCRcYLciO8Zi3df4QavIVN0Fc
wj4os4ryShQk+15TpLKHDqod1n556dHq769l39Uv5cX3jCHNbfUI3S1qQXjaXzyE
ZkskBrDef0l0XSKHMJI+zzF+Hr5BEysYMJUJge0Yh1Yjti88YsjkC12XrgEO0HmU
q7kUoV1QYyEmNftVgOzz91OknDlKfljSLAVqNqyN7LO5BadDDsLeYsFEZVC77vl+
CdJEDhWl3EAxKATIRZ803NSOzcVVKoPpq9+FpWpj8irfQwGrbJFGLj2lSOKz7LVk
PGEA4C8xMkm0ouawUDUEuJndoTjVfTlzPE58Iv8lRiQzLIoX0clg2jlz1G1i28bl
05iFsczXWjGGTwstOr29QThjGT0sRNQFfHlO2puCvfM42nAU7s/1tzXdpXtv1nTt
c6VkE4X5QWMD1Z5qZxkXpMhzEV+oYmiLB4kxAFaEsCLhNaKj9fo8Dh5+9FC8y73D
cQyzJHmaGuG8/LPAAUQA/l2ehcrfsHAfPRkkkP6MPvG/DhbGyQTaiie4amo78NqQ
eOb8SDY6ZRk3PMvtXyRYvWkR4+A54RxYYBZ6Lkn6wtfxjgXYZ4SFNBWdbgKfaSk1
AujXTWYy/QuRqfJFtV/fPxOcay54aAHM45xovp4+GC4GesoKNS1zDjPOck9l4H5f
DPiVIP/Q0AumhUOoGltERLc5FryiwwnCsv0TS8/ISOcdxhcNV3vmF8D4JoLyVDfS
X8jEFNRicX/9mgka+SfrFs0qqJXQ+Ff8IO56tmpqI02uc6l7x6JpwHHTDDWvafc7
t2DCNCmNjK6NayVWD3aV8QxKwvrapWHZ2r4XNwPD3tWjfjK+4ejadzPXFQu8aOvl
6vXkiTW0eB0gx6/uXck2+40hoC0kYK/mB/md9z57rA7dehadg7bc0ow9LrSs7U0g
mvcWZB5Rcr2S+iJNMjOD8lKfXqV8cyOcFXvKwYssggFbpK737/nOm2jb1SSSRbeD
VmF30WVfUz3QZEH53MRivby/fL4U0rQd9aidfaWn/6chUqn1AycxzozremS0ti39
GLi6O6s8s8OgVAKgPq6u1CahL4ten7V2MaxtJNLR+vLdzLAfOUrVKtX2Ihs3YLX+
VVhF6pBSEm8GuSGyutdAaiF3/Md7Qt8nltGtPa7+PpMkgZ/xe/l8/neV8y27BcJy
RBs4qST5p7xBjCIbv4XMLShMXWP2a4oZcegNk++eOPRJPMsSFWviDctSMlBun50G
sOjp1Z9lQ4TInki1Ee8PGeFwu6dp//s09NjIuZ1mrfjKSJQ72NvrLZjZ5Uq8Z2x9
jm/0cGY7/KSLQ2Cu3qHC1MEw355pu8V3FgEBS4bDeqEkeO1KhOis/GEq+HzAUC1E
Pa91+IqVG2ozYr9pqpuwlNgcG7Mc8Di7jybuchX+SiXUBnoxhAGP+xv2dfzxCRi6
tPcSZYZdtWv3Q1BAMSPjvRH71iRdrjVbvKaou5Akqc4hrGi3WwxZtlmfosR3LsKi
8izwOmyPCSbvSxLqlGlQrY1pBMMLq9f2OhvhiIHDNP0+RSpVJY7AtDCzwP3huvXX
6xlQU/+TkReOiF37oPBSn10aNiTEvu+8nrP9Q9zq841UjBBsMdhWQtYhQBNh5KUp
kaGWBiCz7LZI9oTQGuLUd1qXZI3bMrCQ69mA+tDtO0v6ttv484xjfS1vY7RcbNZe
1OKQjdEW3slXVEWtjmbllAvQXfcN+80Ef/BPwAd8JKd4YRad6zxpPmUgcmhkfyN2
1lS5BbBYCd8GFcsrkZKqorIEkTQzf0lEULzH8lqn/yc86V1aGG6mgy8fMZsPIQAi
IY7hwHWKms7t39Xf0YMj/jHszcw4dJ9cyGIKjNF79xfyTGzUQOWH/iv5DnDz/CbW
I9JtrXmJJAwTP5fNXg8/agqxLDHuRzsaOOyYhVrvAlMl08vt/sAa/d9y0Lalys4M
kSCodiM/ckZ8PUTivUXddnnURX0jHPvbkh8Eqx8d8TRBbQvif8uESvPF+clfYQLx
Z1+veTJNz6JpMAd/9sUljpDepkgACew+E0u8577FVPk/+JkzhlLG8BFRftlvofQ2
SRzx1Vc6qQPmnFMEI33Vq/S3NFsjhi6R1Lmk3HyRNSs6tlC/SH0pBDky9mmdgatq
g5Dg+OGZ457u3lOMWWBeu9kYFGOxJfL/wHc8C34cw4bkx1uGoYyKYsVeXL7Uic6I
jSx9p2y/D74vpYHmPwE+liWKX5MQN6v/8ViPejpIF3I+3ig0OpQBedYhIMKX9o/R
cxm3PMUEhnlE520/3y72CKjKi0GKky/HXJPgy8WVLX+xhW6rQKPH38uD6veWCTeh
TYbUFuXiJCtiAiN2lRbQPgmH+52zB7x7VDAjEEMxZP3fFIHS9tiZ9mwDRejEA75N
jvoP5eP5jE0AXOIMTOEM3JU8oRYSR6RlA2fl0tN5X7FDwYdipyYDudKC6iq2SzMa
AodBfpaLzOVrd2jlWN6y9ke/+wsWipFEn+TffVsrplStI4FJUMJeh74u8Rq5UVju
PoNi1L19ydQd130ROhmT6SQPmaqTCHPIH7FN5cTVHf+h+M3mJ3Vmtep0d0+ma0QB
w/Qd0u4h+cru+3uPmJrlbq3f+aWCzoE87pMMpu/MO4qkexsOrOb5PkhGM16AB6QH
TMBOBAQbt61hlws7DaghQ57H1AE4EAjrjKO6vpnFvuamSkdQY7Bckj2YVElkO4ZP
+M08JweBHJGMWPgWvR3WwEdtgPlnFnVUY4oFVFC5xGf9AkecmpC8IWN/RfN13p8q
F9M4AyZMccJIIl0EEnfmeVQjl8nt+6l8Oh/hpYV0Jeum8Gqegscy0F+5AJ9ntuqd
EJPy+OOZ/bc8LRA3o7rmBIOBqOsodncnYgJi5M5va9DwZSZoXSulN0UhYcEbkJOa
H/9p3A0xRAp6dn6o5gPNXGpwObgJNBGQRy3RYfertACtgFcYZ1BV15zfdF1Bt7nA
eBRMIvisj7gcdfe1QNlLMwGO6EckJ5ncTFSUBFa4qbktZzLVyxnAg+SItmXQ89pw
n5S15TSEWJOnrIuk3iUymJx3o+yQXuau42YlrHgs5GJHXM7V7YzrFuGtbRwszSHs
VUK8YG05O+3oj+tLULaF0ebV4Tf3HNZBPPWVIX4LF+KDE4hjJzninb+w6FZo5VZ1
1s6NfNwuksMvnHP0dXQTQd0Mp3s97TzqcxOAR2FnPm0uA2Y03NVUFHDc287Hb9Ei
J5kpachlNz43Pl2CMDglGfJypOIzL+Rv0ZSQcS7YH0yBRw4c8hFTSvMdUKafaB0l
jdUYU5/t8P1tTVy/eZJJ8B2IAG2V9d2VLWLibBnoIK/osXv8CLaPFvTt9RKfV5u7
OXaa65tvvz/cUWop4Ylt2WgPXkoMhYgDkEv+f2yEPSBFiDbCC9yXQAw2rkCpzE2f
26gcmiH9rUxn9KkBsCYyE9dqXAC+4a4YZP/g+qjm9W9VUvBVF8xF2g2hI7SMV2Pm
uYQFhshElgsJoVOcPe2wFNt3wM2ZFqnML07JQ9o4KqJPZE68W1/mO7VixNygBXHr
5y3YTsAf2f6tjp4l1OVOT6rYYVliYuq+ieXMgOYdr+eDfxFSJWpck2W0yO9HUloI
QAC3LS9Pkyb4p1WXRyFcqySdBvcbijgNtofwan+8AlGN4zq+vA4xUZo/Bc8vHJTO
hGJcC6on0VXUZYzHM0qzemQ5QK4IMPKGomZKbD0356T4Ge/Nkwle0/eTCTcpKF8K
tlLz1yrnqS/QTe17V/MYkAROoYEK55shjQbC0p6tN8cz3oUnSpxGxc3F9IfM/ILM
YOb+ZmsO4wNgxOE0EABgO5z0zhZ2c0D9/sxqBw5Bh5yAU3Crd536z8JtdbOWsL8Q
WNubQtd6zPCOcNNrJnvlGON6Ls9u+PZ/E7GkGBycEoZ1ohjI0EmkelidtImwZpxt
CwlrJfj2WH1Gay4yA5Ik4pLZBlhVRry6aE1j9UjFbBr205BUa6x8CMNYW1QWd96t
VsuJ/CYXfWX/1t/+sd8efl+266rrl+xhYes7vGPhl3rfwpdCtnO8Ux8mubWDfqe8
g8xXbuiAlZG7htixpl4pVQmKmZwhpijvbhcIxA76ztGf37O8uL48YeF77DxZM9zZ
vG9Ybq2y8FYlY3ThIo/ju2AgchS0xDThWQQ7DwobVuLzS1RljxEJUcGBHNjvXg7j
WEexweMvZP1z81Syip5kZukQAMi9glbbOHtEMq9l7dIfIJ4+kUptJ6HUHutkqh9s
dg0wdAajPGF+5B3wpq/r/37kacw83DQSQxOcLAzXdSqfXXxS1NYouWe6Uxcsebu3
vbzDfmb2A9qf8m3EH2nkzC4/zNntpeX3Tf/gVDdrhzWClcD6JNO6lQjYrcUsHzGt
rD+dgWGxzCvbq+qf1k124skTPG28C1SnTiWMKrD8D8JUsRcDjc1YFSaC/hV8fs9x
3ufpXUr13u5QCPQm8v4pq+fUVj2l0OjUDKFY9LBy3jAOAmKK7yl2oO4jvzlURBSU
ckWMnU6PiDWTlQbeirnPRtPVZs1n0B6Yay3kXQTjAsNbdxFjJshccBymUN/YG8s2
wZH9LSC6v9OFghvBmRNA1lUGy2ucugulD0X+/03XkXcUws2ZghuRf3hBAmYiPrBS
Rh+6H9bcsvM59FezMw7rZ15VGXL2c7bF6JsMiBb3JY54oD3/OZL7hmpYZxAzOOAx
cCQuRpB8hy/z1jB8d/sNCPuaKscxuUDKSXjiLHXyJgo6Vdw6klWmA8FLn20P1ick
+YoASur2S5hBtr4vsoXKZXJeeDhMUbV8JZIjEtd6LiotPAzQHhaHV6LQyyBAag4w
AoDYiuO6NQ3VNrFkCHAxp5LZWh945GFkE8Ac5eO+n9xqe27wveDt7VaLgJLcf/NL
1ACJi+SbqG2nXCDFsuWcEg282KGfEVgwxInZeqBPuIV7o+MBktL70XjdPjURdd61
SmMXp3D5w3bOB+Fa4bFqMUsoNUsglVKmr8bKCyb+OcAvUlS7XfbLeFdn/JwqpPe3
44eUNCeKnDsyr4pqaloBdk/xkx8VIcBZ9kHrEvEu+mU4cu8upoXV0qRom8cG4JYK
1EGAH5TQeLalQpVohFsxhzorvMBg/KoWCVsAgcoY3vMgQD4om3F+HHs5+DTsFSt1
Z0fVNhBHQaodeMDsVInnCtyyPavHbPvq7zM06Fs43wtK3hCPOwnClZjq+qsljbYy
tr0RyAi3MacJd+BU1rRY6C0uHq7ZmowT2MdaqbG8ij/Fzv0Bc/+Nj42RR0yfad0n
JrcQEPpFq35zEvFhKtA+YnoFS0I16AWuc/AlvU4quR5EeAQSe++lehpNK5PrUOwz
OtJdVLXVUbLwVpDcpFeaM+pB7fZn13/vzQZcoQbufP+rGDQqoHxrtbHXzEasPxZH
McfvJRG1RwiEhgafMIH7o2Foc/xtl9vYG14P/lUh+6P2D4gBvfDRqzkn1Ww+9gM4
su13EK3w5NOveKXoHkAV8szEwwhU9EGHq/LWx1ICLDWCTnylBiQu+qcFdVNPc2/W
+1I62pOABjZ+aTwHlWYUlOdFNo/+27aFbxU+pttZ29cMUyn4Pmj54CXxWRmsIdEm
oPw8c/qhYrC7mjwhztQqdahPJw4azc7oDDltTk/X6titpeUzrGmT/s2aUnSRzyrb
7zm7xhY9yWlWt/kWfr/Gwflz/Q0vHnS+6UIIhV8MFYilRM3T9zdExbwPZMFhRJY3
0GiE+LFoCHXZ8Ed2i3Oar6lg3YQYuBMmScG5oGrzvW7Py0Wuf11g9OJrhjgL+2fM
PSbgAqxLfOBp+kS01lGgjc1MjSxT9049hDjkUSFUMsIICalNBBlyHulRKtHMQ7yv
EcOtEReDqtggrxOzbwJZhFaFDBOK7MOWmAXqaSOmBO2ClndcXmvvfO+JXwBwi+XO
bnYZWf3Wjtw0NVf1m55IzCJEICVHXJi16hFSXPY+dys5wGXF7KO556hI3596CANJ
iU3Y1zlQGmVpg4pn+7cuU9EIuMAdQlQf+eLWswpWX62LZ9MjSMbUpcklKQgmHdZI
AWsBLBSozTDjuEsba7jvFLZbfh11uZck1s4VFyFKUyIoIsIMBi8wZjyhn6Y7NfR7
PGhWR5iNJ81BvICD/a1a1ozNRfKzDHCNl3DMQLc5mpJzXwFhtqjOo+mNTuBGLbqW
fts6uX30aBKuC8vUDh67LdafTBoUCGm3y0LBu2n0KBAZqJR5xZshGfwE7elWAYdL
mYxvv/FWr2i/oIBOFoMpLp6LSYkk55ZcWGXVIcp4yS7tWiXRPoIIqpB1cD2x0xwu
EiSrxIXTtFbteLWWoY53QteL2pescpLw2QDj/vj/m0e2dXT+koBqwZoytjELAgqC
IFA7tmzbM6Cl8hPCWlyLF6EQb1ptb2zcK6rzVlMR+qYRPGvcwBMY4Z7KqJAtKq1K
hmIIzv1ES0PFKcza3kyZ2mmMw7V3rmeFqZaUmWsP9oMpourBaNbFi/0J8ZiwAEg/
ChL2xG/sN+in1UfL/SbJX3vgVXQK8rRXXYluNgkRTVkTkUl0Jqzhft0QJWf029Ve
ingSzR0JBzcfagGLTMxaHIgTEF+Gkfx80kJ6pYdQY3tJ3Y+JpdrMbPnbazK8PAVI
agYF01X0BdtIQ+GzM4IzEZtmvATQG2me9fpAwl3vbME1SdOGkXdsu/qwenkNLPWe
+0CCSQqNgggNi9nzh+pA6Q/zdMUmf5ZF5h3vgAtdvjPnTnIgPrzCm3hEbH5pX7Xh
QAWJS3GGBBK1NqA6Nbwkx7+5+bXHLgG9hYCzVnNtm8AL+seb1tJAV21wLAq8df7h
4irHI7d62iMstW9lgffWFwsHZhwv512EGnK0MOsSQxmLf/Rmx4XLKTuTUlRPUVnj
dlufsnMdPOzMzneN/5AG/2eSioQm97TTM3gxIAzm6O23F2kFKm44UgXDTzSvin8A
xc6cqCfEAnSKBNvrasHcEHZ5jLxGEHXLEV7IY391A9AUecIyi8qqYl6mS43mBlPk
HaXCzJvorB8/VtjAL0WyGBsBpbVW4jaXJ7sBL7SA4WK9xDUd1FbkjSk+vsq+RTcL
xpJYD0B/GGelfHwdRPDsSFUJOFgvQuG9N1mJ8McB1Otsk1p0hqH3RwDOEgmI0FyV
jTviI0O9Hm8f6Fw9AQj2e1aq8s5xuY/ZLCFmOHwJnfbefjuvGsB0ct2ZjPuofFyX
2QsNxqqEUX7fOTeJD/j4DNiORAKefus9RVt077HNdLCuvr18i8sphYA+ke6v56z2
yIRXxyodAoqiQQ+hoWOj285spg7rLAaspq/pePukbcIURAeimX0eRiIVFQEU5D5B
Ukcz3qEypZxlxMdk/XH+R6/aCuSUNHUZDl9wJ83ljPazulH+3FhyCpzAtCsLQ9OV
il9IgM2wpkaA9xZ57hu7R7WDiMD8ZuCHhne5M4yqxM6sVOsv2A9EC5vhZbUVSE7s
2swVnIvV4pWmySlNsk0b4N/ag4l3j5OWMKTLnnIsTBjlQmTw+QDtX+ktFFJspams
MZkA/TEFicXlkV3FllN5l1FgK7JM2kgg+sKPEbti8+urDzzYSK3lWCucwg3F4S3x
GTcYODX7ZlURIqL41umEg7JSDo+ZZAJqQ3qe0Qe66A7vOOaQb0GhlkcLLz3o17kZ
slir/2vzp2iji55YpRZd0GUXZryqFXSrd0Lms/fEC3zBOFq4onit28RzK4O5OvQg
zrjYqFMwN7hku+BA9MKz+rwckyf50TIY+QB62mr6EkAMKQxRN/t1Ro1EAijmunIG
+X7ptNb75EcTIz6gceyTbWdloVyuln8wdnTKypyAX2hsE8bV5Gnv1ZNxhACG1+lB
pROgPWbsF80Ym61SqyxPKqJPPoxhX0OvcvvCtAVHt2RyTjb5Iqn6CvmDnBuTLeKC
aK70f9HlOuZ8iop5q22VeT5IW8+UMKRb2lF/Tgvp+cs4EzpgT5Ub2whzPrUJMbB9
AwQIr2Z5me69Sfo511h4gbAX49WzMF+QED4kWyadbJELdf6FmY7z0DfcVCgHGJHr
4LowVXR+3V+Nr3Y9PUN3hZgJfZ+kFx9bKln3W1sxFSdW2wtWm8optMdWxoZwgkCK
P/aRzRUv2G0eedQTMgsMDTHs7LswIEd3RDLbiyBIFD/2FJXvbVMA2F0H/dFe0drv
TY8fpqLSY1xVIUEnPwAxHfcvhoysf5m3laiwlgHai0RRztLIrmPn3XxnsFFojs/S
hu7b9nP1sSt0i9y3y3OzZj54r9wC5HNw7yDSFBxAj5ExVGvZzzMkfKECbMyxHzPs
8CI42czsKKq+3siW6JKgsFHZJPla719pbHaLtnRkUMrp9QxZ7iC5pp8nLLS34J6W
QHUwYnuQ7ITDWUrS0L8jeD0dur0HRvsu1RWIPUzmhQ18+oibBXH9s2eD9Ri48086
/450U2DJpCJj0ZHKlNl5xeyhzS8P9+L0IWhdRkrlDJCzYFEXsJ2DeqP7xiKO3qx2
pgl3Wdkf5OE/aYmBgFtj2brDzSC/VGJHyf/phXvxPqmToDrG++dVeOAMvLlImNmw
Msz+9LsVNgQSk2wa8gjn2cBRaf4bg/Ckl5KlMPwNz8P5cN8Q47fNBhMHk+fEzDe8
9GAZKa0+4bGDgl8ji7Wm+NBmKBsmVuSRrrSujkC/3D/wrZ/xROszragaRceh0g4l
XfTzY/wfwIPuPrEFxh9J1IX7m/GjJICrXLOLNeF2phdjGM4XgNZe72fNmgcrsw7S
P+LhckzovqMpmGhTPhQddekOuPbOCHpRxTy066Yrl0wRl+Pl6ZKvV9kwheq9morP
d3XJF5dFXFi7jnoyCk/ju27HKcIkGBJiHDcjznDgxtrO053kGlEwlndRih74rz2C
Qs82g/4ACvq4PX9Bz3TkDL84+0CgRkAHSNRgsoV7oR4ryj+0Au/ytTprvOrJ1SWK
fT8gOr4n1Kl6YZMZWoX/6iH3ry/O6NgnbzPdlDIIE2Q8t0f9EQJH1RZc2nkyHheU
QAN3+kdQ06iFIUnWeJwjIunwtm+6cIFhXYe6A+pkNQ1lbGeu/GcLDFXGw0XjbsJw
0DJbfqmxzqY/COk+0Tg9kdeyk6OGU9/ZoOVC+Z8ZQJsG6eORj7YQzwiGXeyHgVPk
1VCb/7zT1MdfFgy1s82O2wbXAcxYdpfqXUfE3T7IFQ7kgTQLpSYGesbdS7sz1Yws
NP7hTjeiCR7ysT0+NxrhPuXnWnFWx0yRuk6kLi7WVD1nVdS9lulmSs3Vq86N3SOz
rhs0hVcCJz7x2liuLdD/TkCzEXGEAqM3sW05PqplBrPNBCKA6jM67K3/h462F22z
VgDq7ISwKDgkNgjEi215M4NDO5DZFT15d/OQVR4ITnlmEqtFZy9eW8CXWWvfB2pw
/FAXaV/9DKS50NLuelvGyaPQ0w+EZ/Q+CMBtbINLvdMnvS+T3VqZWN71fD9yCk7t
D1LlJG+vwAhWjBE0QFqZe8n6zNpNQgw7FqJjdBej+Lzrma4ggd5BqJp6tdUESHUl
98F9jeC99RZUvmd4nxrjH9Tx1X/zMI7CovcLU6K64g2P6Go57nFjrHsxe2ZPoJCc
6Vo0Tyt7tSAr9kaiXnT2iYP3WDTszwKp3P2kF/O6NhvoBaqx8noi5h3j8foO+HOU
dZVCRg3Knsog3b3hiJlHEacWiHUV0F3KQJK1/tRIQ7v6VlYKcrRvmalAW6y2jveK
v8fXo95GKT3tgQbjeRbql3uOEvRxHoaVWc0URa3mEvyzhivx5OzzF8amNNSqpNHG
9BhuS+c2QpBlRd6qUP22iMtgdFChL6tvWIRvAl4Ryo5AHtt3MwTut49ufeMn5j0b
HRRk6oNSNyVbczCZEfaZtORVXcQXeXgOACALsjgDgOkOP0/ooBl/HR8Xd9bUYN6j
IDfrtwofgVYoh5Dnlh+dGvWq3pxXvdZEjLfFbVrzXKxqGfTtUuASkKnnIewYDISk
AW5DrLmq+6rVnuS0sOU5pcFwbblC9AVH1W5ih8M5p2DDsm2xTqR+jc9N4KAjfe8H
evpJ85yZwE9PFDzIeXzLseT2svBMrAfDm5Dm0l10huRxW47Z/rRpQJ5qEVMunTme
cFBXi2L63IAA8nFByMXbYIUkplilth/JVQhVd2BeVQ+e3jUXeRs9hOXsO7QDjHbh
7Lf8twn/jV4p5LnlKlDqwRiNCFRvFJUdMpMvnjX5dKJYvK0EO/SNcRhNah12FFZE
5b8bHZxuSKB9TJ6wfPp8x6rFTy+wEOEb79JZPGnQNMsMXOftmynETvt4/aYdipTD
6cC8vUsdhhXgiJxMsERoI2n3qRMZsxEkTdxdZWP3qkOhnMtWgJc29HH6tTZB9dnY
5JDbtl8syqrP/1W7jeW7T+NbC5sPjPic6bHAzlgxBJR9liiqzND5ksQnHWBwlf3Q
2k2akp58XXgIWJBq3UH7yrUttRvjZ05VKF7nrIxjlJn+gVhgddFusT40AR3t8reZ
ZNxBH70NhfF2fQdkPfcj4+19xSKWZiEaeTtB7hBUSBp5bDJ11f3JWXmADEqBVChO
omuTzW2iQLP0fnWRy61JZg/C7HaRZpgl9C9FmtY2yRuTZarsVUQfO/1kJD8RAF0B
gOJ/D0OLoczomRbdMxaKcwdiyXy/to3gCqzrPrSZN7zeU6Vr0klNBoZcgYYu1Uq0
nE60NM3cNiLAJFdg6dXVdJQdxJtiWoKYXU5Wx/t96TB1fZ2ChWo4TmSld2EiMEZu
6IJYX7oD465ZQXLUMpRNzh/Qab75HUouqLLRv8Sk0cM31XJH1AE654FWIqvo6s67
wYFc27t0cNV6quIQAXT+zpkcukCmZYqrKV4ofUZnLlqQF2UiJ+VuaDnTP5mAVBnD
jofcUnvzJsKO4O8Mh4jwSvVC4tIlnJd+33uJQjc4RoIFgWHGdS9UEd0oL51oli1+
U/zAFah5MR/Nc3QIEE+GIT/gi13LQJ6qLxsaahPyZy4z6Bglkv4++T4G3aJJajQT
xsKGXjCL35KJ2d7VxOzSUi5WodFxQbr4yzRgGcLS3Wshlee6zgtC3Qo/tBA+SjC3
39jkW/8lY3M+MbvA7yKYerfyqNBC0WSJnlk+NhLdyW2vsru5Cf1QYPX9xHbyoPH/
Lsi5z5Ugpoz2idgOr68F3nqaAhcN9I4G7Us50jZDGlVQcFrgvvpN4nORgJU1VISO
vG0VZJLstMWkeVCVAmWpE5dEJ0o95W3oErGuihga6DthsztLxaTWauwBX+HEEznU
kFrmtykXjqoXR3hfAMHSDKyXO0JN+KtrTv4AnNKSBmUetcWh48bkxWkh6GI6DC8z
5No5HtNWK4W87qVmTP4RiFztOlXsS694khael+ik7JJ4z1GNlKn5CpYxR457JWWp
9YCViF4YcWfZIlypo8v3m6x7sje/Kq4DV++KBUnLppCnO0UC2FwCu+6500bfwKws
e507t4Vuv1E0C85WcofCsdR1InOJAhSyGMzmhK4e2uvtngrpkDLOLV19i7+V3U8R
bRAPEpJGHsn+0C9MnXzlnT+ss7fkzTWmS6dZjGKX4WOnpToCHL83xeYreuJh8T5X
mdWNYKW7aXnxgUWk/MWzHPdEqaKVB4Crf2g9YCQgAK2lwyXShIdFZN/+bZkAamTb
6TwfMR9IzgG43B0+C7KeSGeG4Bc2MwWSTTTc1RrE+jeYRQp1kG9dJhGla5XK3XIy
bQiCuBfil+COCXdPpSkF5aL9//mHGN5skCK8huyqBAmqTLPaTdBoq6jOaQgOC5ta
7GI/ThJel5t9J3UB1LAEZEKdp05eqWkS6GetkuOZj74PmRD5OiVkjGsQ9m3qsjY3
/pknHJ4y1emPkJP57DswdsNy9QZWdu2FSG1JboaFT0QZE6axNd9q0wY1R3phWJWY
lvF9gujwd419qUGgypdIcxaWdQyo4nuVHx1I+eV5aSM7WtU4ybrwKBrFKrJ4YdKK
fOtxqTgXUySmEJ9dkTVDxFg1J2wYWul/M54MjvbgWpHo4d7E7SYnYcB3nuXpfk7B
mbOYiYJo5xhRNXm782ETWSwOqUmfJoIT83saZwC1dz46PcZR4vACFTK64iezxFIk
iY09YAVrUOgwtlfAJb71Fe2hSRA6BS0PrIxo4txQrJ7i6vgui+LmMuh5fLxRsTcT
A4ZX6Fb+n1+C/2y5AqM0p6CAa6yYLCO/mgzNhCp79KdrAe47pqHez5EEu2ZVrrjr
gA+T3ikvQPzJ42d0iZPCQWJeX71yc1NNp2FbA9x0/Ewen44jdUMubcioORd5/hod
GsiAYOPrh0TmgGKENoKE6VqKjiaLiI9DcZRW+x1vw/s44d/IIAFa5w7yIZjgv5Jw
vyWbhTYlwFpaqt6ej3TvNfg5TtsLzRSBU8GuT7KkDuwaY14k0JJrt8ij00ldfZyD
JddSDkAPx6WJbaE3mLyIpZA12bzMM4of1nDoeENlxNnYqrE8DXZqBk7ExutUjvjv
ozFsN0yAnYTv/TZ0wEFyF6t3J9jTvPES6UM/jgMAUHRJKd6UFT/2t6FSy4kp9ZJs
HL1BSDZJ6CnIbHOXHttq/ICEszNjR7dkjW5z30tKSyZTN9ihxIXBE6YoTuvW9GyA
vZ2OKwTf2HSFMOhJc9JXJORur9pvxA6Sj6ZSeYJMQlr/FphDInGvt2clijXgZHaH
Auq4ScVw3Q0Cvq/2chvmuX7G/UIQ6Q9YoiDek+s/OP99iaFYfbuekt0Q6CoLy82a
4jOzpm8SUW4toiiJVUEG9dBeEgWy2Rrghrp4DnvRvCicbEhk18HAAjqJbJPSDNOW
2sapl8iwl5HLG1Ee/yOTcZ/ULGDALwT8BS6wMbjkWh63DoNH52ZkLt2FQSzC5PH4
hHJmML5fAhMUvTFcUMd6EOEgFOMpPdHBYUM1tyeU5f98A9vTP7YRQmNmza9oEhC1
ukZ/mci+HFfaj/hu2rPE6mjhFA1LyMKtWR/KHCWihFGoEO7uN+DB3SxEcQpA9yCu
nc7D5DMx1adg19pm8ZlgxXztDHW6nomHxAMmPYWrl6aqGLqaEZFjsQDuhis/nBCo
AkDFI4kEdS2iC+fqxUFyPFmE1efyuMXMFeKkFeUhQRwgsLGEuF/8iUQo0KLoGk5X
Y6zCaHacywRzkMK+LRxSyWqPdBHItay0tNxuooWEaxWt6mVD9bLQuBzz54/w21Ho
cvMAing8gjeEBIxXNaDwGDOE9HcgEV4x1ub4dKOgmwgAxeIVakYMycGD82hgvqEA
oT4U8CZTMJY1xMOprrn7IYTUefIBvDn+uLKLK1qkXvx5fpkHgwEyq8qWgY+VQSIX
IYu0fdBaR7vfLWxhK9Y6giRNPsXQsXZM4cshEANJS0GMt1/josrxa/foiXrGblJt
+CEd072VJJiyvNQojEBwvikrNZH2+pNIVHvLhKnin0dLI0DDt037m9SHKpzjPeru
ZF7SmKN9sENIPDHDNP+xEot7HV+h0SWrMeDetjryEQesrh3Rz1ZkEVzQy/IO5aPc
eAy6MzfG9PggIbIe1GiuHd/R+wZ14r1HBJUZ7Hc0q1rOwdw/RkyzABl9Ma/V3+Rz
8vYLDhzAkzQGfAxHm1DT33S3+q6wwmk9S0RjX9kt5cJQmG6htf5adaV5FNFo53vj
Jt4avSC6Df+1YLEREqqqTuOPCP9y4XjRFYd+F3hCNxTRjnqC9QHY1JFf90Ous0gv
B8SRUNOhMtcBSAqS/a6S7+R+DpfvAeRLKfXUa1oReevYpcn3gxj/MUWmBe4iJOna
sorgTeHyMoNIvHXE/gLEgG7V3HnXsjMlMkqNVDYXeLXyH3CSnxiVTVcjA3yUlW2J
J1+9IZHWrrm55B/IBH2s7ZrJ7ndfUWFk5Vf+Ng9jIHNnoezTGCpLGUiDQizMpRjk
3OnKybNEVbssAqzG8DDE+F4xpD4FVYB4zSso886f1R9+NNdAIMXwVdM6AZXeWH5P
4iGKMrzBu5tJwqO42OgA+vUYubOl7NvL6GYrWvGN1K+IWfPccv7Kn+b0REELKEoL
b4Ruh1KGJeHTuhbve4srGgQko2Xux7zIzsBzBJRmx9NiB1IQaBToTZv4j12Bv6ly
7wasohFFclZAotF3+5bXoF2jG+KYa4enS/sBnXV7Q2G6CcZ+6epqjMO+O3zRzqSu
9COzhwC3JbcJ22gEm/gn+M6pn4enlGhkBTD626/eNXjHldLiuDojPu7dYjG7mgs/
sFOkV5UQmSCHPiFnR+fUMIUEndJuMceEhv6yCTO4L5W5Lre1wAWvPzHmW+mGCDCb
vnRwfqfn++cnt5FTQV7soYwQltO5I0g2cEfQI9bcd2Pko7lkFP1o4lzA57Mb0yBF
buwcvdaSimZnQ8ZGghaQSeM3V7Kmpnt7YpmjAavY3SdwH3k87s644OAD6dYaQBj/
7AVs5C1ES0pUGKdyH4seQMnXbu4fhooT3lSyh3+NQq5/WjEo8+IBU0GkfZJulsju
nQ2xpuUb0dAZ5aPFt4p8o08HgDhtTYRXtrddDokBrIU2XQ+iTGwQUOfRWVpYM5Bu
UcONluv6FMB6t32f2S7usTItVkC2vKdg7EgltySYYBB2SzRvMC2s5clZ4wmOLaft
y7/G7iYujhLlZYY9p+ja5eWiGcmdMB3sauCFxRoapU7EI3ehifRJQIlWDYM8aNFu
lHd4kqQQW34ue7Afg2Nc2P7UDuGnyDxM5knE/r/5IjCZRT/O0iVYY7/Y+70b5ZUn
o8q6HDgskXWukEX/Q2uj9v5Tja1S2tHhGBYEJJlf9+6dgQYDaKZStULAjqL+w8Xx
Fu/c+mMondceLTRjWkv6VZN4Zntqr8pneKCI8WydKGTUjnfClZUpacteQE86eeeE
I32ENLBDY4P5v9KrcB0h/sT/rryoigUWcaYYubLFBI0CIgzuxN+qXzK2lq9Io3ts
v7e62tpVQRkvYSFBv/CACIVcnaDOp0II/Px9XghM3zQya+YVYllQ9KjMRqniR2SP
1k9AQl8y5x31x1GGb5ywlHwvqC/ZNTU6HYJms5Yp5+59oGUjEnkhy4xHi4a7dGE5
7yg4bWR/25WGsD+hbTnq5A/RD/NSzLZ93+/5RjUpgNkoEnhZ2mgXKHXn/js5TSGc
DckOyrzs4u9xMlQ7bFx8DnHq1xW5KYLvNgEhR2lnSb/Pelm5bQIKOD6cZg6HBXLT
s92Sb1pdOrfwFSsanoKE4L29sH0JcRiUVeoHdBwraL25tuAdneOiTM13Lho3Ede+
v0QGtX75eBcudIKU8xfLfqrZonDO+i6qic1yZEeL1v1pdFW5K4DXswtksPOoC72p
uqDYlUzkYwn5e+cNzfz7vrBjvTq231Y7o3PJQldBwOZwKksrOfMcKRmIX8tB2xIW
YccKQq2AOD3/uQac2Z6d2Y2r25ZSUl7fltSiOF3FkEKnAyNaefxLUk3/HDzvLJg9
i12mEsd2xRaz5Dekjt6D05en5w0HvtT88ZA9644KQ7ERcTz9cour3iUmkSZvHH+i
Rzul6KcNVgnw+Xdz+zqviumFtHsSfRAbV/wAVSIVjmLurWhkvgDHk4emq1/Gbl7n
wvP1QkRo+x9hEi1Qf0HHPE49+w9cLD6JtxDgWaRn0yVU3BskMvKPQMZMAihRn7Wg
7+AS9DH74/qPD4t1HAI3W6HOV20ovLVNun7cbaZqd7WWQwCamRD9EizETLXDckXe
Sb1XMMWXUjDDSD2Uft86UIwL+JtE4ql+EuDytP23+aQX+o4YVKWKyenujhMrbeGg
WI3Azr8ZkpM19Fzh3DNPUfePktHcyGjhPU1RRUcVWvm0uJTnGMTYsEYsTFt53oWR
6fT/8DyVBerDg9yZbMZrxovZzgEf9hj84yvywI60vYtwDKX8+SBWfi+RnOLLFblb
xjsNA3xWfnYRgOJWzYyXp7JC3IBEKRilZQLJTDFvlouWaN3eXtHxqKYpYCz+Djr8
iDnhUfmA64x2kt/0xzrezbpyTY9VamLveRLZS4k2mM3RNG+YyQ/7VbTc3QAS6M8S
S9AQpsMV9eiXw1Tf+LU9OAav+mgxkuqR8KwpxuhoEIGjr6daoocUCaqvr0WgMiXk
ic6d/9qE+jhz1oTEUvicOZro6PCXG+ghkRhb166HxW/tlbcgsqmU6UbepPRVQ56u
BQcq7YSNCHaVnWyQcHzynL/4yXoYpDtoXQKQ0OSovmSPtkBGRBXePymZqfswG6Kl
W5wGwllsDuZ/c1OlhX2KGrGAmZePqfXw+rusfwWMyIhRbHxSkb7u0NwABuMQrQZ1
Vd567kiE6P0GWD5Xve574Ld7uXZ0yQZWvHLwsZJvJcKaQ1C6o8pPYn0VK/nkmdzb
aDBBqJIvakHKbYOGI+zMzAY2/DX5GgRge9rO1//VTh7fDmbCH/FNfxK4VZT9c/rN
HK3RQxXAV1tHBaw8gNLSfr7GDRnbGz4KO7uzovNYT2CnD/YWyMceIW9/yQy5Qaau
BFXlQeagmloSkUfMJVrMNeG51m+Z1lm0lO8kdFycAH3l+nOKxYvlB/ixOccnt/NA
j+08OvKcSWsHScQxmofBkz94nyx8+p+/L85ZSObF/XmCEmKMrs+bqWDwPw3dSDHJ
wKHQcgnYNo+5PMcmNHtu+EAc7UIU8va1xMCOCNfv2TSgg9lWrV0b7NlocZvmT87x
uhoOsgg6tvy6QmzyNutgrK0etreQH8nSPIYqGLIULLxtiC/ZfIfawjU+ayQlOQcI
9WRdyNf4KcOokwI3E3Yt368ZVlQN6iuYOtbHymsPvlqJAz+mGnlB0U5prb1LTxEQ
zebNnT+K7xtEybBnmprfh8z/8XLX9UcM1KTpkbr3gbGYbqc3oQSHdEcUQ4oW98KO
SHARoU0BxVzrG7iz8JVrk7N99fRZkirCAk0yBAVv9EcVPjdAo0EZHp5N2MWBaZh5
bDNycvg6fXdY9WBGqalHFLRHr4uiHJfQx4k6ok8UiXQnjYFLmVEJZlj5fqlv42q/
rqzzUHePOctltENmmWAYZx+7qtbPAK+6aI7ZT+iGOe8E4iM+L489dr5uY032WgiU
1NG/TPMkh8f2hql0PpJRiCmqI5mkMnaBspDaePxa1adYIAZkknRAdDq/Y3AJggFy
rt9PBWrUaGj9ldaGWLuYH4EiGFSgesZJ5gQpFpynhssDIigYuRFQ8GpFPl97+ZUt
TxQZwF6naHMnxXx3mh49dZkpyupxmuFuJwtfcDilz0HowzwmVrEMbfJm1FiCXqJt
Dsau+BSjcRyEghKsQFc9CKNogGiTjk+mzJ5xd2G4ZuHybQ+r3i0+Rl4wX7w48Q/H
eJSOBo3adnBoe3vU49+uPxUx1VHXlBl36v4Mo5LxziCCY3h6N0R3KdzVBS4pkJUS
Mh/hZzxPntqbEb85RvmMayv+m3uOIGhEutwpNplRuxTDbm3EkeAJIT32/KFbmpMy
RN80M80Uv/k8Yd/SGMSq+TKPt59raLV1tSWvoSbpGlMd4zcKTbPBzr7DnQh7qbhA
wef+RWyfvbR/EvRBG0UnS9+kwGUsFL1mpT+5k+OAxR8wVP3EiVcE5a1aomFUq3YV
Q8bzKysII1VDwydZgJ8sKMVZRnixQWEAW107KcTv3T/NxjVZ+Bxheg1f9JLAtQaz
J3Ri/wfPGxiyfIbEdhqUkB+ujwEbaPMQCQRiQzUPpE2vIMOzTElZdtvSVpymamyk
+t+jMrWnWrbyAyQAjXq0vXtCJWRC9TtpPN1qkyZgqzZ1gFFBR+dQzYKVOeb3lLio
LBTXQq+GMy49XX/bDHN0ogsX5qwX3MNK52fKf4eyz16RVM4k95dEUuno+SVOHmQa
lbz7WvUee/SNALdko1raYG6ItSJbEJNrTjkvJlb2tmwVBgxlch6no6+zQN3c195u
9VmrvoZAVkkdqTATtxoOBaN3ymtNABsyxgc8VaJduAfCwwQ2vZFM8vzgt/L/Bc0G
YjGMJ/gDDVHedy6jli3reYE3S3eCnyaSQ8iFYCkyR1/KvVGXtM3UEB+l9WMIxikC
NsLwEj58HJXeNt8zFF/wsew3K/eJXltGZ4fWtF7uN20lfWqsJedi/UXcydfyYPSz
BIrFPVI/zHCJ28nez40Fh7/SX03KSnfctMSmrrnI7evohlcJEGB1mzPZkGSRxFuy
JIxrYOYuZHiQ8fZTKeYMPKPVUjtzpxt5Ad3x4CQpi+JZfxgur6WPmkAUHJfWVqdr
0UJZ4od9Mj7BS3b7pfbXedbiwZVLKcKq79BAQjTbswBzy9NTqaz9ycxdt1evA14C
yTfyIq9oUAnGP4XdmpQzH5y2nNXnFvnFRH3P08wPCBVmjBSQ/hi8a1ERhUopi444
9U0sMWcl1ISBg5OJMOkB/g7Q2TLp0TjI3sThGDCmcXcMm8cmMiUFDf32xfOxJa8+
7Z7tB/npVqzdtV93EItkD5lxrQTCJCBwbq+Ivw/Xne6v6VOwalm96wPxq8vwnbFn
ddOUVAjUVJL1YkMOzAEqI/YVA12yHoLcRumtaIAe9UXy3d+Xbg6I3dc3MYBZE2RR
WVReKlxxvbFe7hNVEKBTooR1lPhu332mHBRtXub0I7LwxcTln8/ONpoEt1ycP/3F
VsypayM+LKrIc2l5IlRnDbAVPPHHTY6S/R+ro+/KrncM8P3Q9QquvMWONw4jQSZU
ToM++I2X46rZUzAyf38uMcI/qAzPvJGqZJZIOXQXNKVAneVGCFwqF8PI2VueYyoV
QqK+BaoWdZTur17NF+JXk1g2U4236SEBq9zs3SzFdRihtH1FiYgpkZQvhAkLbbX2
IPbBxjFFIbnfghXPy5Tb7uZEgoz24lJ9vRtlgOUMlPnnzebnx2ccY9l1stkC5Hph
CloJkXfHojVTxSavzNTkkb1oyoH0QqYrmC6IisG34xQRdjk5Y40nQGhunM9k6EGo
HIuQoyAVK4mhi/u0UFRN+z0WbWousG3vn4RSfOde8ZTY39oFrzAtr1BUHJQiTqqq
fe7uwoo0d7naElAmMShi+ViIQAFqSTbuV2uDKQqtdUwHScQ3V3EOloZapUxLfLIZ
rUPzX05HZMbL5udIZs9v9iEy80vFWUirGZJeEhtAeBMkFuPr852+2hcBeDZyI42h
9NsEf4K+IZIAVADWpmgmlH/vli9ebVeIDx4UhxFQdKWU+WUlppi0qPRD3m1TgM1A
5C3ggqtHlRSxaeg9meHxoWvr9ajTpIgxek4QwdF2LZfrhCuGCAE4OtTPxr4vtnc2
z7j1ClciCsgIDkWkk2DyqtAQZVqQHXi4gmDL+wTQN6Rx4C3aDWgAj5tN1G96nh1c
4FPBQFvyviZasrvu+sVjHyh9e2ID2+mHQvOVyzNh9EvG3PX4asu7vFbsDzfW95Wx
4Qs0PCs6zEy3Y+qIw7O4wU+bVG5XBnlEnplN5OY+WUrWJ1cu0nVmdXofiGLU8ipd
X211pQpbo+DDdZCt8kDQGwFCoNqpbojIh01Wm6x+hxkwYOugLmQrcP5PB6t8cCF8
NkLCvlC8RYKH0vmxVBsWkVYssFk9aOlEL9ew2HBHYMIRT+sK97nXQSxEAPUT3FQf
90Jj7/kJM7UfDAAgw+Brquc3LPmCD5ojsx/cFiHN6QEos6Z17U/7Kyl42kBYizfy
9ggraWumoah4x6sH08hFd22C6OQHC3yLc5m9PbA6YoQVkdqVsIuU7K9Il992hlh5
2kSOeq0TzYgsYohlskKRqVv02wOl11QeKfNPr4DkiR1Asbsr+BbsmjiNW/eddmTM
1mwhIt7BzWAD1aI6Lr9I6rV/pajSDTixkMPCsSdHu6McoyAUsjRAQNkP17y468/f
CQk40RMHG35BTlfxoiYcZRxdHYplrbQgoUcEOAJdUjEquv049B8d5p88Tw568fFn
jRNcgMvdVM3oMnaGkn/GDnRIKy/dsNsg+v+rrWDVW9Eda4FkGl3j6zrxUNvlSMqw
N4xWQYmV9tMQOmDpq7CAAoG9VDM54KdA03giUwVRCYuizaLij/+V5kUE+l9LYSym
JOLy8alJlLTM22gm12TImtY29WNdh6YD7vBpEX6bsniLAjFP+EGab1v34yQ2l5cq
YErD1RD6az3CvWt79K3vD29HTAC2qBcCGhJPGd+PTb+n/g8WKM1IZTZNhgJAO0BY
ApGutZqnyRTH8WqortG7nUo4U+cG6hbLzN1D4vkqBsXWSfmPTIWLs+cwdluhWlGk
fQ8cHewlQApoMLr5dN4gEf47RLUo/L+2tIBoNf5WQq5vNzM3/lnIp06NKEEX34KR
Z6+OkhzENSfwy/tTmxiQbQ7MzxjeV+nkYdZQrGx9oL5NHU9vvo+BvsKIqRQDtUS8
mL3TOvwaCL5ypRVC4QVw0SioCaXePftnz+aTcZKwWjvutp3Q/4xrT8r3ozbHjsDV
xyJeuR3CshpqGe5jCjPgbFUfhKbYv6Fq0sUbEPCTpP22sqzVlOwQ+Wt4bs67G41U
3cRDiiSU51OJ+2WEAn6PHU5jGHGX9B4+d3fIBD1tZ92ArSWkBvTMTpuKLZdZ/fU/
2FNhqi8k18rWRtRCQD4S+Hh9tqTOHqzZuj22A+8xjLpvQzTzKD/2WxAyehp/5S7Z
yuHrnMcRP1LaN3hvtvgX4NCD0zvttRuvOuCeeAI0uMIAjPJ4DmT5MfZGeSIfmi/3
NBVdYc9XuanatQ8BmYsLMVzyJ0TyMjACSw9RsT6iPEp3ul4WUbY0nsrwlnDNunH2
Mz5zHgeViZl7i45lWq5XSceo14iIJciTiPpgMlyFBswocARKSvJGd/ETrWUpkKdY
4Wf6LSyxPR5FdsPkMnthmPTlIBYjO6jDkJPtgG/FpTsRrh12zkhjZM1vo+LfO63N
rZF2+cAyiysMXqNaGHwaZz6Whmsx0276zdaOva3KRNyNvoJeEg2rtoLTsuSHcTH7
6RDZQsJ9KmfX9tZpnmTYI3nUL6+c3Huh6KrJ20gBsq6SgdGzJLq6ctuUITjdY68H
KZ8yf2+yQVAJQnOGYca7ZbQ4kLoDczr0K1kZmfcLXjv8+6s9wH0+SctUBfx8k6RI
2qbD/m8Iojuof/NjpSEPgQeTUHG3kL+Ty/1eR29r6GwlEqW1bm58o6KRWi/D+JZ6
xCUtQeR5CbUF8p+lkVjXU3aUa0CEe4krsYx8UsxZ4XGplWBKWJxEsY7ZCNIyLMjY
25KaFklTShS/p3ei4AHdgmAScESoyp20//EgQEkLNQHGEmlv5jd1r8NQZ76xOF8p
XfkOdARcXP4BdMADmyT1AJa1MGmcIxAiZSb6b/pxowJ/GTU4Zwj0xuN2qATG7JWW
xel97T+cJ1TChbOAVztXyc/TRVuxEWG3+S/iXGo0ADK5QsBTG1yCnqcgCA0hqLIn
uYPOYjJHDYWImHSDjZcWPDEH2UG6kLGAozxBQtxG+k6ZaAKeqEJnoRXhPyO/J/G4
r3Tz53DJedYPu+Pu05SzjW48RQJqxb0CzpQMSEOpwhDz+3F5S5WQxo7iBCIpt69y
CETJVoRrkT+l05S+8SzFYolpu9pQTsr81PnPxcHXhTl3z4crfoC3rF++a3YHh5TZ
EIq5DooevYobKNo+hzJqj0ynjGol2Jbr1TPPIBZ4DgusYCEVOijNtMTTjAIBv19b
2imL7UVIWbkqCnBMIgxW953diDnOcx1FMqWHLm9jyICHR+s5GtNX99OEZrPyltWr
BKl/Lu6yo+llF4Jf76b8a/XUIDKq77IdhxJMk7uQw/yl7QJRywlJoFwV7K4zSBXG
dq8Y0tYxib9Vq3Xdg/YNNLuqT5UI34caSxlLf2w3t0DaxgvoHTnDSeVMO00wb3HX
ybU7SOGdszlH8Tr5BDhr+84cBCXW+yYQeHxNWQwvr+Unj1a8GFz8jda54YHC40QA
NtRavwlNzEgKFl5judP6J8cECGHaVA5LS2VDja4b8BIbY7BCdIkVS28O2/fGu/Zg
ntmME6UhhqW5UPULJAjoIXUz9RnQ2T8J8NMDPlBeOOyiG//v6hEg9WNR7hpnb/XA
D8C5hRlmmXhaooh3c9LP7cQJnKC23rYGgkBpsTwEemBMoz+XhSeMXTkWjmby8T4t
i3c5HBhWMeAE1ITemgpTNRuyM4m15nxKdq+UG8fI62JzoV6As44d6H4L/0K1+8tR
QualDqVLGsVmnK3Yl9NbKYLql1dL6AUvC62jh23OKZgsCOOqPBvr80ZUkQ7vpVwx
F2/Ms1rxzOSiLskvM4blzdfD9X/3lL94Ppt5SZxh2CFlmt12kha6JfvAVKf+kHWf
FHhhjJhHHLzY84iUGaWhuhYJ3g7YIOcmJAsHtHY9hZ0FM1hkNmt+7oNppnZDVMVL
Hcq2et9JkxH1NxmFgcE3LF/2RhKmzWu0CtfQh/I4Xt07YU6f9poLYwxMBnK/4/dp
Av0qY6Wu3FSGKQo3YnpoyKXK3TE1HIcCJygfKWfjGu5kFhSb45XvAdUMKYWW2JLW
69z3y5bpzuMOU8gsp0sjgX5IH4C+aVio2E/7SKE0+ZI+eyUJx8ksC9PW+7RPz9ZN
C7Uo3DXSNqAZSX1ULzpoL0WuobeCFCMrPJqW1+wGPtLrkSWqRJLJHSpabaFEJ2vN
2sFmDwYgOy1DYuda39Kb0nYF0nJn5wePrfagEcxJ1VahAiJRoQRyV0b0jsqDQQBr
0uehhd1xrRrAlyWeNUAtQm+kD2nKvYVIyDdAAOyEZEzFevvcCF3pcopSHj8frEga
UKBHKeHDMqDih7jIVjtdSE3QRjgpByN7QrjmsPb6e8doO/QqK2EJiqhY9kYf5BwJ
DaJqUj1e9Dn0COGmj28bsvv471mq2erXUw786w0QCF5lFxRvkzGymf4Rhnr0GaGV
Uz89VCSZeHG5u95u8bMjXTpA4KoB9sMMsOALRNP5hNanikhw40X1HLm+jzHGpQzh
+7SIoNNpqbh8qShy6w60dC6UCWjNRzHnICFKvgg2wR2GlT6PNysuzvYEegnX9cEi
k58uAKitBNieF10lx0p/RUU/RwZDSnhd+LsdryTXFeRuZaTm+d4xO5Nd7S2rQl/N
1EbLhs7f1l+p7ws8SJGg7PBg6qQAbtEW/09mSC/tS9zxs3ehg5mmkbKR6gNakPcs
ihMcHQCEu71Q4Eb7Keiob+ZSg5tv64iB6leO4zIs4lZsQxasggDuu47gP3S4xMa+
7Trpa3ECYymggeRDUhM1fnEuX7smFdpVON9hXgKdukHeI/9uOrZ84HCatH+1gc4W
1VuCICjBsqmBuTDkJW/cHkJpd4V8Y1x6EsiIXcNfcgqcY5kp2wKlVfvYjCE1yDhp
yjfkmNIFbYYlN2wurvGb/oDFJcXN5nQie7F7fglJggltW6kni9n1a52Utsl1z+vM
cSY47P7koBPsdB9uFHTGwhB4Fg1msGGHWnG24539G3kf+UgeYBHUXubXs4DHtqzR
yjUEh0EXRcfCJYWzvy34FKpOS2jHj4ooagcuIOAd5pp5rijjwhASn/+mvM4Gd+k1
t7pT2ueWZ01rNndUO0ZRgqnEhAlPGpWSp+aon7VivThRQisIxnLUfGgFO35OFvml
5gzae4zq8WnAoL7EkVzmw6iMxLAu9nenEi9dzR1Mrky9TshuIeQJA1/Lgb4rywLI
MwBVWFmMfd18K3pDPOUeV2HmvD/fxblwoE5Wt901BumGz2oLvXGk04wwnfsU5P8O
0gm9H8p6ng0CFWaIUQbNxyPsZCO+SzbWl9uC2zrotSe4KgSE0mUfrNAQZo5BLfKF
Q2jYdhZDlIX1FEyNVOhb08YIlsGiJK2VO2dMg5n6uM1MVV6pZpcNoD7IEn3vh2wn
8+WJexeHmVtBF559kg6T26blLh+qPnsckzF+E6ejxCXxjf++Q/i9k2YGlWM+Gl6h
ShlqzXqURh9sb00Y2eOwMjz1psvwlz7jpCWJ3UhAI5tyRYy0jvQd16fzFjhWFRqu
tKcPOHdgxyGEbAYnXyfbb8Nwck8YZp/knH/RD82AmKXCmLgyqJfmlAQ4ggHlqUao
IRRN2qZpOy2/CPWIgvu1F/favBuYdUau+YX4wBBJnaXegcOw9Dec1TrJb9oGzun5
MKXExRj3UhY9wi5IqIS8emav2mzhikD47X8hpSkpLUQSntZ6aq8llS5olnIyK94v
6H+BYF7YHbTPOzm7dRrnUqpUfOBUQ2rdJ9HmO3r3yfJwtemBBepcPbVroyj6lqob
us/FPvrE/V7WZDNY4Lif37ZW4pPp0n6NUbPv/n7my1rpPiaoQDCYLQFgzCGhkSIf
MKzbLzcjTUJ30f/UoU859KPADa9pR23CGBW9YEK0XgV2EXye3Ro+gFh+ITg7yYta
n+dg1of5FJhiQLXaT2q5PUSszTK0hYrflOTIteLSDgpEFWnkRTqVNkLMvH6VS8qB
vD2xqNosZg4vK30COkwoIdw1chcpkStnj18+wEmGI8cm9c61iJdkqT5xqWoTurm5
5IIhogyQmP0YIX/OtLWY6EpCBUgqVLGY5lZMMf7lOTm+rtiikfhk1A/61VhUbmAq
80o32Lf3u1ifGjLwgLuS1dwdD9aon+Dbe3ve8MF7Wl0o6p4s0gsynUwm51CegU7e
36R4aPfNVDGyfWu2qmJw78jY8t9DcoMeMpr8NEW4aNAvIIK6s75oAv8MHWEggLFW
ud3khh8TlVe0SQT6zG0KjnNfxo45zgOULCfo3eVHO0yYESwn5X6ADtfYODz39hKQ
pv3fGr6D4SPv2EFyCOH9YqtCJG/VkNYxu7+0fj83eJ1AIDJgIod4SfYTZLXyLTT8
25fPhue1yAaDFWsEAYjRo78PD3fgSbp/0EBmdRNiztPcSiczsR89nlXoOkCGSWqY
dlz4/xxwUm+drXEceooQTAISPSQ9zpF9CTibhYFyOwZC6Esr67IsojReiZJ7YwqT
pGzHwPggKPm5bUO+Umi3owZ7VpmF44KoF0j2J+8kQZX1Ld5RLDpdGtl8X7FWdJjT
apIUgTumKkJfoA2VB2Z42udO37E//0ddoFeVelTNQGm+1iI2iamGCK9lWOIvOTA2
uYynnoiCuiUpApHWs53ctJoeqYfBG7NLTCp/1LooXr7IKlTx7OzzuCIMB/DqvFyI
Kg4tJYxgwTBxIlaA/SH3kTrsk5yymvkNJdgsNq7zw5I/yw64HW0cyY/XpxzbYsir
rz0Y6qB7or8mH/Wcc7271XsGUrpeNhjHWo4CB61ai3SYi22RMnQWYUvtMVVxCUZz
Pbme+2lNOkXeFF34P4lA7joJxf9MNAzxPcJ4TpMbZRnh0R6KOceRimM/FBFbTrUW
Ogqd3tiq8yMUwzHBPyRPhkS5bAtX2Rrr3EEoX3H3EkFrkFqckLgUFFcFVBfcFRvA
5aFRJ3jUlK2QTDz8Yn50jz2QDB6Dxm9WtPYWeXgHf0wx8SayJKSFjev6Dcogid16
L98VQesa2WQN/xpabHm/naE/WkQx6yn577pSESvFy31Fl5Z66C17bKRRPAh/niD1
7egDQSuikDwnvtmJi6hitcCEuSN8ll05jAoBzdngbHuRykF9halFCUlj07F7sHIk
4lDdCYAsCH/A8uS1qVrR/epqKOQTbkk5ez63wpWXgTzMZ0qLbG7sXkrrB6mBh0Qv
xuaDPt4KntwgOEjB+vBSVNrGwU+PulqwXDj3d3yPOGCceDVy/2GWHSE6OJCTURTt
197s4Amg4yyi2d+tV/9ZYzrm9FmXNgARPkvATgPT1b2JIdDP1JU5PoiENwZPA1rE
m80kTmzc/pOAHM3tdqJAGxYwaggCTtnpKBB8QFhBWMcuUKn2ZJKY2JGIY0qqAWpJ
dTC1exzJLBFxl0VckVIWhStOkrVQGrXA4fpBZL1DbGkiqnS3YaNpQuIJ5ov65gti
eafLEr2vbsCKmfaSQWB3qNNiDLon6r3ce/gxvt4e1JSanmqu0wntd7DRlYU+cqYy
5Eye1ee3BiN+UIj6xsTKDqPkQ3FusLQfLnZb3G9L8tHTc5eGk0mnaWvz5RcXXDEO
67sF8u7CAvJ5kERbfpUsKzb4ek9juggk0LrkkuvfFEDXU3rcye5PfVozUUBCuStm
DXxrSXwcRW066kfwn5HZCRcgXGHF6JjINRAkxnAk8fOGGua2q04m4v6YvZVucYhk
vuA0qRjo0VMP/K7VmlRCoS3E7EwPK2nFZwULdWsWb5XxkXUUkaKlX8ymQk6pY/D9
6PGjaEQ7R5mhF+k1mAvFAbDwk5Qt88nTXNiXUOVlmNTCAxC38VpArgJtP2Xlpxbx
sf4Dd1iLyGkh8qSkByBB32HnIw2Mc4lUM3+ZHjNoBLwQA+8H059Bp+BaeS1BX6V1
lwGKsERCYOswN2BCusI1OEK6necDfeQmKQGUqRqut8kXoOwkd9xEGc3qt+9FweMD
+TOjTOCgTjyJyaiIT3tL33TprDRvEacCdDVy/0gadhyb/xgn2jpo7ENEurju9Gds
wKoa2jWq0iw6Yej1S7ygoy1GwBNpieTUctfs/N8+7LoAqa8T6mf6WC4EdzvVXKOR
PNESqHRQDjn8TWcIGNj6/BsS6CG5dv17ey/aQi2dco2xdw28zdx8KLvkWCkfpZc5
ZMXtjOH5KQwbIzxYzlT1Ev+iYIRZ6x016daFz5PdjFjyTZASDbYGcdFdzHqBNpH4
RWfsg/HLDAYaVWvW8iNIKVP9gNz5B0VkuBp8XfFNRjYYhfp4sZ2MNoBZOia59U70
nxIiHp/8MrMInnAckIKaK8KVNCmCI6PrwB0RItedVaq7m9dq9rABA7FdtSFFPAxQ
3suENkZ79jFzBZBHYa3H1V5MHDaxlAR7w16jzRQeRJrsVcgSF+EWV96s/GBTjq7I
6kEjaAZjle+LlR8smbRuaoTSf6d4q5UKEvnKScLtLBP8lQ08meE3OcQ3OnxpiW9V
X0M92GCpAoM2jM/KNeyzzUH1p9q1N4+iIuM4DkbTUalF+gPLkS9l0P5+OTAOUyl1
MTIEULIl08VZsocNwdhOhHkZ857Dci6Gj0/SwNAOEOsOXyNSOMufEZgSQbiSYcOm
J6YQI8ex9lVlZtnW+seyk1HhwKoCHszdyOu01l7rGo2X5LIcYvJ9kOU6ADGXkCtO
WxV2P2cb/EOXa4u+Z9HuVffXI0vYWWG3vc/D4QvRNhN1KLAvjHz+WxKsa3ENrME0
9ygVScQK32wEnLx7OUI7W+qpFpo+13Ibudn5mkrvpTfzaFz7xS2g2b/EiArQ1cgj
+F4CfuSW/miFpkv8tl3+B6OrYsdPzmrFVwvw7uRvRr1yF61uwmu59xtjhmDfuEyE
wbM37kFuHvzawl4lNU0kKuZCZnqKp8aANBUwcrKrzH1rzMMXyARa0OZjLeuocFiI
th6Ptp9VGfoD5KUJ9U8nJiSj7DH5AR6Qxi/0cxqU7T8uo0Y1AmFMlp4wKaJVuw2M
o4WK3UGdC7qC2EcnSMx/ck5agu45vBcnp1PXzhbP8hQH86CmfZkFD6t6edSPDh3O
1vGExhkz7XTP+OB07KwLZcU3AQxIw6PiHb9rFaODfHahrPA5cmx5QiVVnmf2q7tN
JUNUCCqD/fCVLbIcwnPNx/qHgIVZaEaDfSy8eMmbnOYl6hAzfOFK/OY/NU6RPiAv
F3oMimj2ihbgMJWQRuFx+MQojp6ZLxGPlvfCxm27R++eRJaINL9z4/VIKwuD+Lw4
SWa6k9oUL2AOPgLTFOvNzZtOF+89WcbmlcE1YJ71h1dj6lESPqz/VoDUgIlut9wT
JJb7cK6T1lFP7XwPtVLCtHCi5C5TFVJgvby7w5MyJb54r/q9bkq5vwP5acU6FDhb
DJqesJGSb2ufWc96PuStuzET4l5JWcppdwyACaYrU/2M3gH7EF4Ze2VkIbjFhc94
IwI3pkxkoeXp1cZLsnyLoTgQyVHNj9NYJLd1Yd3IABOecLcxyzvPfneednaF4xMg
Su6FXAts+C026Icq+XnHqObIwvvOcpmg+B7zhl92rqC/CqZ9+tW6EUieIv1KBon9
37Pqh4/WjvCZv8qGULlKpGP3H286pdpqKV+6GywlLn8ir7PN6KEoL32dG7T7Jk7V
ahg6TNo9xsv68RyZIqDMA1fQV3Sb+9WnLsGhNzv7TfQW5Vsu5/dXmM67IzXJ39q7
zoMKEO5lpBSCuRBViq/pGYZ2usywI8SQChgy9b2GM+S0932VqA7TlYNRpM9hfAqd
3jX/NdnYyQHFPh9z4TV0e437A64R0rADDjmHVB6GKy3QGc7/79RDIy5KCWod/qH5
/R3o+8icHSWkMQFNITbx7q8Cjh0lTAkiNuU+Gf315dteUHQRGRHSCfGGbq3CN6oV
a7QAs39hO5AlmCGGQ0C3AXPArQ5q+pf8UJuJAfNDPRmNxXIf10RzlvI10zPiUqHd
IAhA7ufRWdYSsr0wcbsqXrfTWi2jypuBxIw22tY81nn0CwhNj0YQK71HxTGPdH0/
IL5zL/ULSLTDH8pp3urZgo6dv2jX3JZe6dgrPIFyddzyTAksUCGipe8Gc2GKPIuf
uxirVemvDHkBdAcLGPsAwfDkXU05QapB3MFZUJe4ktZi8RA7ah5S2zOCBwdxKrZZ
tZzKWGDv10gPB6R5GlFibiyBwsOMaIVwmn+9XccbVJhhRADXZg2FNj2ng624bFfS
l4JbquMN0AYMsThP6cwapjdDzV0VUwGSfnLHPHGOieDsP1vUBMXXD6yye7TsnVmN
s0Ad4/2PTQiJIu7jpjUk3KNCoXJoANidltUnniBRIVe6Qpn1tDIehQHxurOUKblF
Zu1y2UpSMkjLOq4eqPwQbwCDUftu/hNprcrdh8tgKHP6sYDZDQYYcIS3qMhiuUuj
Q3GQN1/mfsjQa0n9QGHCfRl8RqInHPQpMUgHdu/ptc3I3rMzPpvUY7GuyD87sb0Y
Ei/KrAAEoP7SChka34jVgdeyFSasXGqFW30zMvuR1/pMVeHTu6wEho1Wt2PxXZeb
ea28KC9UPe4S9yG9Z6u/DYXX35CEVYpzzZFC+HB+pMn3cMnjEDGoQvsy2/IdiOcl
bxlyMafenYqgh6d3910BeSKX9FM6rNwZmmeiIhtjTcHo+WRXimne+VJqJ3ok4EuY
nY2FQK5PDM/V8PCVNPej5rrToW8WJFkPVk401YKRkbnzD9GWtnymorXiF9PBNQlO
ZmsP5VAcoE5QeZV1o70RGF0FU5nIvrpWm6XbbR1U5bVUeKciit4HZLi95E9pAKOk
V0RXYTQiruo+kak8PornAV+bPXCNueQCr7z0Hw07JyK7wc4a+L7mzsAAJLe/s2UW
zV9SyHIddMNtOyQStCx14Yz+iFs8qQdOzltkpbqQYgliXlCflVTajU7RxkvC3kHc
NMGxNnxYYiR8l9epTDOid3TqoqlGUcUldoAM3q1w6OvoC8W3AkqyQ751SeDGFlBV
ODKRY1SkUwviw3iStUxrPk109D+4imZ6Ltqz6zYLVlFiIpTJgqy/BD23fQ4MuJHe
p4rCW4AZs5jrgL2lbDgOYwXwPg3xSlcmuH+sA29OEO5vMU6DhXUO0mIFgnoUX5I4
XIo3kf9THMkPZhhBgAur7697wOrSBPyqCkxMwDtcmFeU1b7HNQVsRh1XooTmsGYT
nnql5zx+Wh/mFEzsKLcWxoppGjpDFyV0IsNGSuG+YC/geo3vHeP7MtmU8U13Oy/g
zqE1AUsRdj78HH8XhX6wWN6vNKO8Bb8/KTFdBxmtdsQgrdw72wMbywVwjVZ96DUu
QPxJvziiXhI03M7XeO03LZEplqZNGP2MhqC9NvvNVCFDQ1/YkdeCHBdtvhDOoOFr
H0hKlzKKHE6oXgLdGB9hj5APYmOrv/DLLGx6qBZTIbhvpc1DbRmT0r/BsUbwK3xn
whfc3qFQqi1GqVjTH4QJi+RwStylf0Cfr4YW8opxyk6Sn1kK+X9ftb0NRAi8NIsF
0zeVa70+4iS2F2qdr7dZN4FNJyEg1eXIV4rxLfhHMF023T2I3Bw35AqX50AOdwge
CUE5ASoZLWiGAGnV5lz+Zml+ThDZ99q5xaZm75Il8uKYLItnVwplyQuvr3WDirKI
sbk1b6qkb6MyZXpzuZ0q25hSvozh1w1fNH1nuJBxN0bOKtuAErpdvlApDLO1ItTf
2c1lHhB9rGpp49ZK22oZuRxyNY+12QuKW+0I7ltejrEj+9jGxNUDAxVRM7j/+H4z
CA+/qdr5tXTmJlJskqEN2uxI0hOJ2OK1E8eyDPB0Th+fH5bn2ZKKAaJTf+XV4O6Y
AtfG/Bv/Q9IR2t0zpEDybzDLqI3PzOw4yTlCH98yXM6BzBe8cin2lofhR+77BFG/
0id3y5YYF2Wp2okEYHjT62rXYscXh4bl+qfw2xhUyz4R7Ax47TEby4lNUpqBKfXH
oGtjoppx7OIhuLCYErHXnGLY5tv4URUBWm+Q8pfsx29TZJoF8dPNdED4KbSx5zdr
oiLHZWQD+VKKvBctR4qk2e/8JAWUi45UJkxRImwKX91IlNv+H/2G359vPc+GA/7W
OAq6yjRtIMBdOzilBa1qTOBEt9qHYFxX3RgRSirt7d/slOiazi9UCYGcYZcmZERV
AZBhTcbt/QIHEm/YlbchkYYQQRhgMmEsFsqpEjG/ie034ii0Z5SeJtIOkmcklzc+
bAazdbc/s9BpfMeoVufTIe+B7M1FC6xPdekg+BRMQ5qHzY8E4jL7m1+Ghkl4J6Md
pHa85DVzUOqdYwf9+TELWujyuZfx/NAw2WF++7vk9CZpYJuisCRm6Ba+rHhsu2+G
tilOA0lbXV5krhwMoeE39l2MSc1wA68rPg6luOmVWnyhEA5Up/exVyNWcV4myFzX
H8ow0KN9IDgu8SAbwGmZ4rk7LeLpBPgDXBWJ5vZClFpWoowKfGL/TgVPo3J0rK0d
KuRKdb0wATNPcH73WD/nrjTRYqId/qRyjLwfxc0LnWOO7qT320xy6DXThVHWThB/
NS0vwMzwMs4gpERqUEerMRIm53SyzJEAdS5XbuZDH3GqB8QGX7nDpqXdXjGrrAag
ZcnmUOH7PKFHfMXQQHCt6qebCdI9a3ufrY77StvXRdxe6R+kNC02QvQdgcqi2Ta3
s1HXKd5m86P58NpmMQRhbCFFWjoiEIIZ1Gc5anrjUfy1bpZjDrlWa2udu4QYzBn7
YWx1U7Uz8TD+yw5azRPejgyhfrdC9dE91xkygZAKqU2i1IzWEtzk90KUxU/wnEPh
10XgfHRY17zuh5LgPS9N5i6bj2RKpPDuKqOlxvv7y20d4rSnkL3q+NL0REEnTKdA
tcXH3n1gIEyavHaftp+/j+0FB63jOAA3EOtHkTeX4vDAaRrCW1Q5KMjYbeY28nGd
hA4GN5nor292BN3p5D3jWmvxr9pg13NWA5hgjpevTdMJ8KbVLvRj2qiP8OFJQ9I2
nSFow+rnQAulK7vGjLThswxzRS+6RKx6J71YcDZIY04l/DnBLKWwhYDHDoo9caFU
AAsz7yOjCm6MhEDcYMb55SJlRoOJ3ZkK47T5B++V1X2fGuMCDGPutdR1zQ0HTPPC
1I60+KtjFNgI9yhf5MJ+3vXWYMVowTdI5CvyX58G8a9NDY0nIR0htrpWkbGBrjHw
leS3g9TjL+cytgGdDVeVUL0xn59UvzwgNXEi4xpkheWqadxOEPfU9OPM5WssLtHH
8E+NBRYkIsd3nUY6IF9LSA5viaCy+YQ4rNr2UG/gcdMKUerTRtOISGKP8DmoLZqn
qne/fIUj9DwcbAV+xvsgc60HwvPJrQHGTr9vGIz6DNZcejVcM8ljTl/ZT7AvQtWa
n3eL1aalUboVBcsiUYwIyW5fFUwP+28PMxP53nSBfFRoJWsQwoHHl9vcva0dRVYA
8GYTeM0jSewdt4Dkf/UvlSUp3Xqi1bOxp42+UdoO/Pf2u+HPcIZHUaoszVaJ65PH
5HK63wc3mL9H7e2YBM/wjsrWABM9UkN+WR/ZZx+nOzSADwY5SoNGwlNXKsy8geN6
Au4h8WlH5a9gbiNUTg+dJ61Xfw0/dGSKMMejKByImuCzBAbJCKaE6AA/DT4ccrmr
R3Fi4RCACi2JR8G2VadtBaq5JnI21XEuCbMbTQb4zmy3ucpXmSnhu8BatM8KitNZ
FKIOB8JllD2rVCsUZvdf5JSUU92I8xDzQ89d/qy/HJpZ4U66pmZBko4i4b6vBLY6
IlGgJGb/RY9RoHtLzTCARp25r6w7+1Y4b06jVOfdivQLGS/Vra5MQr3zEHva03cq
+IowqYpJedhwhUsR+0vsOS1FkcXsDXskWQnpn+mfsZODZn0uzyHvdKG+LTJpbk3v
w8rBbYucsIoko0HvEeUB2Uf4M7inXa4I22hJhqQncxvWOAGyCcCGY58Cai57slLg
btB0nhjz2pv3GVkpHhQ1X1sSSZbMZ8FX7eB/16C05V9merlEn+h6iwhKj2ePP1cC
MnxxvXpB1NSiivRDRuIhGNirUP4DUr3B8Gv9Eg32dfnXHBFl5Rpo6yh/ogGHDWOl
8ccaPm8DyToxX8+Lkx3Psq+IUsmd5HaI5A5mgdFvvnPCKREb9+6T78gMAi5iI1XF
VNAF7PJ3LFf6fiVo3AiGI6J8y1qiZiCCrDo2uMAigCGYYGB1ReUOnub+FU5121B7
TQhBwX/iNZDEjZtnMxlFQihymVG0+g01pQWU68wevNsoxlauYFakNJG3dzdrOxv6
gmsG7eDrsZDmWHdiPujfoHKtvvx+LVp1+UL0t+F1M4Gvk6gHyNkASUf7cdolZc0R
nMf10n1h4gmu3RngVMigW7mRk5hyKmOri4B8+7GO65r8+72+ZYvv4HeIzQOc9Job
0slpBGrGT8s9ydtYoIA00tKhdsvFpDRi0hJBOnX6G/ZOY047LxvL3IRZZPfFq+9X
DczM+bfrMMdakLBviYuBXoBbpnFzAxE0g7ypK+k3Q05Gva6nToqSDJEsuAYuapIs
LZRLrO+EODZr6Me8poMbHK1bh7UjR/sD2w6xKUo3I8evp635sCQZAr215kfVYnev
2W2N+1LNAmTHKQeIqmQASJcQLmZn1mXC20PUnzeu9smc+BT/qAEeIalncp6s3LwE
DKYEp8GmKEumLT28CIizYEayHdEvNJXh+V1aAdRiuEAfd1qchjUdKJwmJR7EOJWC
djL362Qnrx2J2DuSE/JB6v5z1IZqn93RbJEcdvrBC06iBnJJsGnwHB8qE5WGaBB+
Mg5OK25xKdpAn3YRDpIzdog3XAaAUbBQgL1LBlWXFVV9iZTRsr00YbgBKTePHjtF
rUfgmM6HXIdgq8K6Fp2UICI8LZkz9hE0R/yRWzBIKN4tHm4KGd8MnlifeA/tEHWP
gu2yq8qHp7KZ1tNegl3Y9PzM6ZeZ4E9yTgdaG1WAavUCWW0WFNn2tDB4IXQaoDjP
T6QSNEnfZ516C9sIfcy+IkL785lKrRD5sYXqud6vHWDxwjzld50ZCTGXTJIgDx85
gWwZwJyXbRDAFHV+gWA22qFHd9mZ8p8GDJ6dPEHA01FVb/x+mhLnOoau3L9quStF
KTraX2zbW3pYVVivfhMEQxLGRFYJ2+p7FsVM3LnBHRjakswv1GyCC0UQ9xUep9OH
bE0ZWSf0uf8P9YLDqO4UVm85OArHEWnhcBeKA7LC95rf4DyJ6KKrML53rcPxeWem
xNj7awB+7P/mSwDfCDGywm11KfWZfssBn8spMQgQZ8UXH4vi0+jXaMOfU4M+2XSk
uz+6bLbIH5NvgR++56bVSHqZwH0Arrv4h74pPDlq0jPSdwYoQjcuasswkSv5VWDG
rrt6sKA1HD887IgEM5lTBkCGNmr2ZjLNqBeI7jXKfIwlD8qnT7NUlTqucvHf8Z5z
VeYeJ6JLS4QvyNJx6aP1Pse2PH9KVE+ZM9I4VYq1FGpCNXUS/m01sHMOHokOkKoO
m5JJh2/ROLTzEOgsrDbd8xEzHa7Nn8DyToCKZMYA2ng9XCT7M6iFmhmabWz4G3Z+
+S4C59G6KoU7sDldgrM7t+iCMXajEES2upISn8n13dXdbfdkcJY9H1uGeiXfcFbo
LKNZYh68HRi1aTwoDe1ut8B9iQWcfC96dTQcplE12E5lnIA6cMs3TqwK0ByZ24wl
NfpJ7jZ3tTeJHEMRVRU1n3OjV2TIhfk5WXYXkIbN6VoYutqNba3LhcHvsjuOICP7
3Mjcf41Ibd2rCO5DwMUflBtUk2xyRF1PMn1+xxlFRug9+BDhslnYfeLTQywcD3Un
bsXoWIXGU7RCo7ZfbXfowDlSwSd/MtMW5G1zQTVJhWcuCAbGVDJEMjT3q6L+v0Yc
Pylr1SKx4OEbdX2YeBqxXjsrFX5JkFX6xRcziOGwOwC8XDeebfdpuXRlyOJJxTHr
I/ZZYf8yr2ySOTSUMARfhx/YJG2+c2HkV0FjAiLZpvSrZ99nFqXcggNbt2iz4WD2
oig1NFJU7ts/uMr4MoH1KBU16j3X44zhC1ifEvfxNsTSQujyQvG7NcuVMKeIlPUf
rBu1bUPKtE6uVG06Bz98JDp8soBezhs2BeTpVwwQrOhptvSwNkMc9hVkQ802TWBP
blsh5H3Fjuh/4oDGRzZNom5J+ni2u28LEkX1tLufi5701GrF78AKTjV5ci/V+Dit
tbhbJrtXV8uOhG6AYZaNKAsqMUcs3lxLzyQifVAgmX3mn9X68vVZqLy/XjQPp4zD
KFegBuaJ+Ep06VEU1JXkFBVfDw999GX5TWHRGwR0w0uI35i2mYC3ayxRTyIgymyG
6MzxSKsfBftvT+lZzwb8Tx9rLDxVxFJRe6ci3zT3Lozp+zYY12MvOT/VdDq1IS3b
uRlbmKsbIK6rEPEVlZaFf9FtBv/jj5M2Xptcz0YJ+XZXixIwFBU7ra+i5j6chGoy
lxzzg74SmKLwX9V6yjyXV4DfcfZeqMOjU30M6mWRGnXMBCbhyvzzG0EopU81whv7
m4Dei0i1T3vP6fOypwHqOeJZn01pUMwlqN4fYPNyIRZH3VObmyRAmGhgpVwuFVej
gBJceTHlNVPBKw3HnANUqpDS71XqYMSfIKwi39r25kVtkg1yziWgvSARq+Ux+1cl
2tj6XL5hERP9tP4ljg9irxr1Y04z0KICMNxTVIZ3ICYycShm5aHFRttHCUTJ1+aL
IbJdV7/zvE0J/vcmo5eYuKFl66Q+YcEeLWLm5SF8m5VqGLTxxrXkjl1D2NLaY4eZ
0QoKqlqVmciwFq2rR0gASK2doQAoMe9p3Wxh41guTJ6VKkxWB7tPkYyv9ip2mOn7
xkvP8yIWtdREelzMsvtV43YI+n/Kk5l4LBpVD7n82CWvCuTOEXeiA9T/F/Hy/xkB
q62DyE2Hh170n5rmmq/S3mHTW3Ut9dGjr0LACskuvH3YUc5GKUp1i9QOxi24xun+
PeOoCJzTR5KeNnaMekdZ0LdnMjIUFgcJqM9WOCkXyB3MCci7smICZbsbHE8p6dI0
gIHZiCbNMD0sCVGvm5AbHPFGMIuTLFnVrstNszxB+OFkscfPlFRlWjaTJwJRQoKS
mQsflrfkw76nWPHUOn04fwY8QVH92dzfIh8IWLkRtTTbdkSuHp3CU1/j2dUBaBQo
xZ7a9bMzWtajK+wC4IT/PuE7W6u0Pc3C05QET8nsaGMRYgqWkA50EVHN9BfwNXxx
dmI0T7+PPPIzG5eluSKFfFu9Sa3GiKQyyaTVdgujLaKFhJAlH5RKuEWPqgfGY7UD
gk45/dCUZrwghk2JNq6igqiQAWV5z6bdPVGjW4budvcPMBVFx0exRUDPE6xmXZjo
d6BwtLNt+UHaIqsdkmfWkYG7dllmNQ6uzCCWJWj2CctX6Eoi0a8qb3pL5As9Q4PB
5dAcnZ2MSSWzKH+i5JFSvWgkdxyFhb0mc59tcyjXhRltNIOZDFXD8o2d+htUe1SX
Jmvg95+mSG9B4E5oQFuOpsaLvO6ojPqbeTssSED2k2MBu6EC2ATr9w1ApnaO108z
W9XlXT8EzhJq1qwHjANH/yOx37GlyAGHFSc+floH/4IqEXeeX4W5Ga6BRswlR98G
QqemUc/z8dbKm3rsXU8CM+57e6jb2AE2XL/tj9OlVMYGeAd7Hmq4ukLP0Lhr50hz
0Ba21Nho+/RF58CcezkSwDH6dlblBx5IYO989xFzTfuZ3UL/TxTb6TR4Jr12Q8PB
hhYtic7Z0kncf7BcS1xRAm6kGyNO+3OCriD3ZlFbWwrcPtNFowJZ15iO/Z9U2y3V
PwEQYrNkT0w8pC+6baHBmD1fkdNrb9rV3sWEd4tRHWXd9odwP+3j2sqRY7gQoCue
szCEblHk+aRzpu7buCit17o1CPhjjdYyI3HtgQ2iSByHdEh2wJ2Z1KB/t1Z8N+ah
5zxqNjq2QJUNDvmllDRF9PuBuetouMUy6qxPb4ERJdlzg1wVkRpAvjNcfE3GDAMm
ni9WSZ3+4xkeJPhu5KrlkG8epavbCJqHDEMuypsvDQX2IO1rhgGRMkdCy8oflkHw
7jP/h9Xz/9oFbDOowC5FkKbMhOcAlTLrVqHwV9l+fCHofSOorA3t+Uv+8fXXuLrO
NQC7cT1S/Udv8h/2d8+vdcpVkqn8fQeV/L88/M+feWN9ARKWsuGMLTCRxqhjUx2K
4sV2x8jQoi9x6jSujQx0VJVAI0gvYAnlcEBauG/yFbtWvE1KxMGixiTV2TmwPz9q
kPR17e36QRX7bg5EyI5BgpmldAHTGd6rD1oe39+XixHgWH7S/LzgE+AYzP1ZsR5J
v1+4lxF/xcvgRnqktWEWHiXHACmByzliZkq8w16abp/8zbCRQnjjaABNPnzBkeSM
q1Xqdd0p+aX0kzZ8GXi6Fj0UZ7/SRqx0WwefE8I15yFWq1LfXQu3Xj2rJfJ2b+SD
GJE9dzRTgmKQpzm0R3pBDcoZn3xD7gW/NVqDeiw38clPnaIlb/MRi+DS820Wrhqn
wUCSqNdnKLZvzwnZ5Zm8mQn/X73xyzmC9UmEvrhzR+2RmAYDN8d2HygS8EYMCJoG
GUm9umblU8fEFvd8rzurI/rt8yBX/b+H+PpgbMTGA/dp689eDLKqMWJvFwI3yCMQ
7MV+H4ZGKUc1g2gAEtwtcNOfpfG3/VxtGiz3wAu7dKhk7TxdwEYJLWSmqjIjVlfE
SEJHeU4/aIMTdD3ZzV61Cw0YRHxeAg7QQYWTiKq5R/pxreURWRQu5u0Frf+zbjEF
hh9QkOHKIJ77NSvR4Lu34gnIpv5P4MoQWb6IPuYli0Vv8oZ5633o9/0BA9oBD1oy
Xe2nzoAF27PpDBfpGouPLZ/BZhJzvFOUwpHV7grmTzwYPpCI2m4MSjcoQNRulZVk
zNhjZDHwHpWpPQ1gbrdfv7vlc7LMJkGM0Gn4OHUETHZybiRgdsO41/JVf63ZMqt9
0tPtpfK7PB1/iCYHlaCvALHOh9z0IZeo8hc2fZO9WwWGY8NhkPHi7lnA+c4LjmNo
Ly5OSXeActlbF9tsY7K/0ifrE5DDZjMykvqQt0dBz+LZzgsPWXlC63gJGQZt41Nu
M2jqGgi4RVUc5IIIMwAsI7VSBU9a0cRqIkCOrHnDGDA4t9psb7zYuqAHBTXBt8w6
OduT2VCgrBoAGVGIirEBrenNxqDvfSFubBTnC/7PA1ZeEH/okpgrG42ei86chTal
R0X4Yy9dKQKf6Seh8HQLcemYFrIAPGw714VPCIK1M6QtPUpqxpUFJhjfF1uBll6Q
WPWISmepjmrP6oDWucPE0f7OdJWrnJZAFEBTVIxfO3IloqGLiWZbcyf4iu5qSWJA
s76Q7+zLBIZq1ewSbGf4LXEnh3y+TXs4p+IvCHNF56pYyrVy5FuMsajfYfkGe92Q
a6mpVy/YcTSA2/EulQiaNa7M3uLhNGKAw6FHrPIFEff6XV3eurBNSci6P5sTZb6F
m0YXlvpMhOlji2WhYSqxTWpZsYFzHBow5mq8Tc/ioP5YH+CrwUBNuzRAQUXffN8a
1D2isjb8i1adSaqV/MNannqgshzNKFmDyg9o2jOFJA7kgY9vUp6kVYPAiF7FI9rv
n5Nv7KU5fVtngySuctJ9uYyb8J632bCnKONp68bO6IijzjSChuiYQq+HBHEfIUhT
XF2e0vw2hbYrqNC14skW3nK6zPYlFY+Fkiyd+cu/5KIkK+ZwQBBf1tVxZhI2vxSA
LaJvVja0m9tZ5fFOuHO8qCtIRSAjSnRo0x1McsiRvKS1rJnoFnc1A8LCf3gSwIOh
n0t0gxmrwlkRuEKLnssiIA4OagsYzFFWaeMKB2OsDUg3FHQ3coY3i+eh0HUFGxY1
fdrNBnxL+2+S82einFv93Lz0IveKH7Ku7/8qLavTP+ErJA7iJ58v7w/fdrysN/98
dY1A/DjN10l1G04ZRUHWj4+/Zie8tGE11rvdac2gNw6AVQHdN8hE6/WTx7/ooFGv
Gw6b3axlz2Ba9rUv/7i3xm+U1L6KVd1KO2XLWXtLqH2rx25uDyf4RszYae8ZYimk
hrVeYX0RC6Ymdn0/RNu6ANXuW7kYZ0yq9vB8ozRngNYQXZO5zVQ2fezG1xdP3IZu
W1po7esUxA2/BJ+YITnR1IeHS4LBryVzS1zWSYLlc8a1GfELtpX+cKkkBt3rMtGI
0iSLiCB0bAI9rjujZ22VNOWxVXqawM58X6R2BOrDyYhQaUDEOFdN6oBa7W8pzRqn
ozWOja5ebnSXgSKF7PvbFHG6VRhjzvfGUElTeR+EQLOp0bwdczCHmeQ2/XaMlwi8
8g+xoDxKpZ23CBFYhwI+f5G/9LMM9LHtZzAPCuAUSmLXipJvogWBcrWWEiBZVL38
+OsTpFNCI4lSQ1HkgNsvjHn/1zGoNjI9EZsFxaauRjVmZS1EVjONiCsZtkBfZMi9
bfdhbm+XGYDXvGBi8qEhBKIwyYJUo0nh586KgatJYCHv5m/u73pR+Y3+iaMjC6g0
AZgHJ4Ovheu5AajATSNcn0OSi1vAKPV2RirG6+k5QU/YXdwgxotCyfkTc/ZSmTeE
6w/npPSxKISad72E+UpN3x30VFjoeMWzYl7UXoGQSwAbfUX0qsmC+N35+kLHUPCh
YOBJHizAbfdNzyFSyfvAa496X7/SAd/MvZn6TeIsbwhfJgwneXA/2gBceicycAHB
EaAyLszWGmyITzc4AnvTKfxeUf6XL01bFDcuV8MuNKhq05SW+rAb2DLflg1J5SGz
EL3GGgAONO9wmbN91baGDS9JTIVjzDIrfU2tJ2bA6egQnNCxgJg/sfimZGKCydvs
XyyiP5FkkTCCkQrJylHCBc3mJYNMps3eAdjFkPs0+Gt4T+PrVyK00g06GQ+Y161C
pmJtGGnVVUP2g1bvlRJKfeVyGHxy3slFtFx6iclYsNFiqORs1pBpMg5KSsVZnDRT
mLnDd83RWdoTgz6L8ZL5VI0uM/Md+0WMlfvcruQNU6U0FQZI6/D0XpHjYa88dmJS
5ia6cWn+c3ULRdk9AwlEYs85pxCEfhEMXne/4Y65X72oIUBAJi+J6ynJe2/XSrVM
a4mHh2kQthcY668FU1s5ImFIPp5kFhW5DuOyw+4cfb04f2sandj9j0iSAScrST4Y
JBP0KPzhdeGc2CeOvZVUOwDG0MbZazAx9YNHtJxLuDi6unUFYqrrmQzxYv5rKh66
PIAX9yacb2vyXQgNqWTXch0gUewov5D5aoND6O8FyaFYoeSckUzgaH/9qLYu4yYL
Jx72dx7yJpQkX3/aN/hDt9j1iJRlYu2mjyuHLI96qvxd6XsnPmOF/qjBNXHo3Epr
CgTpbEDqySHaRTRJ71kJal+HvtxK/4va8Xm6FveHSBx/Q61t0+7AS5POXatE9xl1
uKvZxDs0eJ4EgcG2EoTAdYmdeBrga7BZ1CX/Z3Ti38TFX9EZitoTQgneDXmKoyJo
0guCNTzfOpCHBM9+gBntI6+fR8ViqeJzIMuE89sDzaqkmxMYA6gknTM9+SMdv41k
nTQSkNGhb+a585LYkAwEJKMyrpBWQWX053m0frK8xsqOG77T9mFrQ6HtbgYmbTPZ
UjX3D5PgN+zMTjYUWm/RLmV6NBZRAfX//mumy0fTVNyKE6O42yRGXsryugoty517
XmjJBJFmvVCVZDnjQ0zpKehDN8/9JlvqzE/sWsTFf6WBiBvIrrGzrAw6+8mFYqwz
AowvPk2hecSdYoNYySZBxWLuRe9YNreQf6qG8SAatjHz03UL2o97mFPhuN4qpi+a
RiGv6pIxWaJDtss3XT24cY684hXoo0geIydr2iImJ/qZn+jQPhH+46WmDLBsXx2v
OP1bNXEa+Yxo1tVZfbptJlKWDCoRGbfjIhORIJcBccZXRDwMV2XX38Q+vNXCiciX
22RU7zWIMEbbqRQZzbuk2+FSBZkpWpiysMjiapzNUrElPBod3iHL2vJIXddiXDGT
phsfeY623Ba7mE97E1oMK59hyT+3iBxkMu/Ytp6NRiPFq47zIFVwkhDu+WHqMcDU
zVzQCkBnGghR098GwbEg0dCBqGONiXPsK08lqFuscMjpq8x4/J3Nqjo2SsLnuObA
uR+SZl4SVnZB/cC/H0rqq/Jhh9pzAddmpMVmuJ4oFZX3HmurBvmDyM5LigmbU07T
o52KlZQ8s3a+AosLRCb24o5kqXcJVtyRrkGXpGZntJoJ+D/nlbS+ampE2/P79Hp8
4rm4+1Z6HBF5Lt+b8hrnU9nSS54GnTx26+SCE+XUWJVldu8TnlAXUDaofyj/R08S
VYJBCoeujpXSCIaxGthWusnGG2h3vSCES4O1jrwWhjHlLWfJbur8PeeR+ndETFuv
RpMYMXf1xmsYpZCY/x+gcJUxphRQiuxKOJxSOyBJqDLLGH9Z81CZv18OoTMVPwkL
VlbvHU/0wnbZqg/lDax/iHAhr8zuejPy4IF3kFSO9PHaxTqG5XsGb2dCksSeMVrj
ieiwb6UFGrKk/Aj7fK+Rn0G5PJ/w1WeOADRsNGPwsP+OYlbJb9e/qjLUm1dAuIS8
0qJkOx2p7wj4efCAb/6/O91nTx1QYracCvHJ1hvWCWPY21ZyJ4tU33pYiH0qwbbv
15i7IDTkuQEGLl/vwBKwliSDTCWAe2IVEy7f8IM3XxeNP0Mqdo0bK7FQD/Miqpru
S+c3q/ZNIFv8j+ajVNAxbzwSmBx/ILpfT5mj26bxiE0iMHpz2VAJaUFXqxWnPT0u
sZs9Vv8lrUNvV+7U63rgKilH+b0OxOP0smgMVwHftcpvILNyWfIaho/UswxaPSX/
njuJXhPTZhWdcpY+gw/iL9M4vpr17olo8MnE9rNaGwUu8gp8PwTZ0Sk/La5KHiLL
8M98q/zSwkY3ZPpj0sM/jltBtp9p0jBkCUTGXqfEzyuocc2kkSj13RiMROUefrb4
C65ytr3LZRv5/v3s8No//jf9FPUal3jrEZlOYj1PpXCodYPsdmBohXdcTY6KGPGq
/+ER7zBCaBQ08dQjpeyRUYvlrcEKz7WfRHFi9TGlGfvUHBQubbIL4gDtnlt6Wnqf
Bkn4jcoztUArYHN/i6dwKmR6o/+psZrI7X+feM+2jLg8kBK4HWos0F5q7+hbbZE5
OALgKZTaMYPAGTEACCD68yKE+1Ny3kg3NFCAyW8yOvzpGV/vQawatEyQbqDoq5jX
WOkrQAJQ6ftizut4Vjs0qmfq6ZibFzuR5B7/vheQQRiIz+JjGMbfC9YHdDRkl7u/
JP0Y1hk99BwDZQr5xF1yExHjJ0SJv546bPuQTVcmjoyHxCFU8fe8qskNelU2fa4V
1L1vKlZO1aoARNElM4ex2X2+kOPEXC2WGdNTDuUZKWqJVPACsRA8NsDV/F5WNcc1
qapENK3AYCERA/L7eQLU4zx+WhllTI1f0SJdWdYDtSvMqTT2rqaWM72dtetXXEm0
JqM4pdD7UK4WPOsR2op0rXQ20zj04w/uUlbz5e61Lafyw/UqLhT56NaL4/0Gcj+2
2i/CL/iiyfr5Fbc3s9D5tfnbqloxBR+dVmdgEX2HwJEm4s7vW1xi3lyGurHa6jPp
4AHeGdvzEUTZkJYSVmb75H6/cqASG3ARaTzTofG7+LZpCscLnTUlDjfKehR37BJJ
8QQjQPad8Cj6DdyBBqyHF5noR7y7Nax4GCTVB3SxEJSojMQxgd88BpI4TDFOoXS7
s1ANHSPjn9yP72fkqDakGSBTvy40SKoSRs/VINTPCwH1JygPD4622U0ESnxmgAtx
sLIRiV0FxAqBeL9GbfTM/azP7azLHk6Fd+QZ/e8WEbAQ5lu+W6E7DW2yra1v6xDm
FFTUkJVDXT4CKFDnf9jtYhgJZGUuGSn0tf1/ApC4PpAv1USJxVSueoQkRcj486Fs
JSG+xqCXdZTBO1ZGCtEdHEil72Mek4p4uwRw8anbW28/31scHGsxD7x4b3fSFFtu
RBSB/KUH3VIQVGc+E/o+FHBJim8qVLcbRHg7xVi6mSAnqE9UxKU5Ew3rC+SUIG3W
rc5Kx+937sqWyLB13bA9xXAK9r1ZBW9bguo38uD7S/CVQibA3Wxmjb80kB8wgQvE
oQ6NLiIe4+CGOxfi22B6bSrRy3BzCo4wcNlcitlXvLJXJN43e3QB8dxCPv1oPvTN
MgzaLPXlWD1HjA8mrriDM4ln7iuon5vwBne/qpcSzNoZOsj7w+CagctJ/EzlVm+6
EV8pE0++rh0QsTo9VGSUVKS/RT+wiJShONltntsS8PrQW55xwmulrLHjEr8BPOXS
XSvcHz1/s/4afWZDCnigR8jk6k7jqBSNpqzG+TWUCAuCj7AE9tlUVF8vkp0ffvsy
71DPOgn4KinODYQZNX2Buo5Y4Sll2QYpU9YFv7SH8NmdnopKuxyO1WExrx2umRYu
1d2hMXucrdmYOPzK2+jdHy4M3NbyUCu+/lxPSOlszWkxQRtjCIx40VpH8QhnCxV7
n052lad6zX3afDijxlNuo4/B2h2hIO7XerABKbBj0NxAVkuMQsGyObuOmWnhBiXx
/RdovP5jjw/rPv6FrwRuV5Cu2Mkidn7L1NBXTcutRqu+13loOIuShYbYZUJeLGHk
XiE6s4vwALj06CyklvoRtn8wysLmHUQ25IQ17ftWctASBySup1teYdmm/e/exRkh
h9KeQZXHlTQJD4APRyQ5guuecSKF5SokznG8aw9hMRpWdI4/m88ZTwIfgU3Um3TO
4YAXZxVHz0OciuR3+sLP8pxfXw/NLKQDNihVTJ0dreJskiKZSgdrFA+UJ6PZhlS8
aZ6rWO05UYg1dXIfbr3TUfOdBLqlOyDdih3vxRls/vx3JZ1bOmlrB1KeuKwLy6kQ
HCmwautWGMYk87Uhvty/QtH+u6djKAACw+iRlGHBSCbRVQkHt5AtjDEoeF+MQ9LN
Ww0eVJywyMBQaNz/5eMvcMIMJ8zx/l14BXXKHPE/8wtXWirmq1GxUVewR+5S90Hd
lPK6ofJkAS2K0rV+wa66cTUToHU3ZJGfinCZRWh4VP73FAYSzydMgT7LG1EHw/Fa
nazvOwfZlpHK7ZOvNC682DCe90usYWSuJ16FCeEe7vzUUKd2ftq6fW2HphsdaLF6
3EeOdlNvecpAYWH23bSaV8uiOduEDeXXSSE4wV1FyBOWTxIP3gouDQxh2SeB8fTu
VjVFONgDGDRs4FF7DOH3CeCewWrQsU0ve/5R+9qbItDU48WSrkHnc9kGBTfOwPT+
+kP5hxyyBl6/4gKNuo+TuxQxvhMTfhXys9GcctrieQS47hUQy7lrLos0X56y9qNZ
pRldcxluCtlHhwo5jrZ5+wBYKnxMCKhmGvwk09rAD1CwVuvXfDrK/ZGsRhxd1Fc+
WaYbRNRiTcTRdQ9EhU+MgJYeQC4zumcVtzFQnrlXLjnrYRZsPYbkBUaU2WjyfntI
yIG4XBsdZ8OcWIWUDG2fcOJf/09bl8+Bvfc4xQuRVS+gwO5IoDt2JqfGMgC3XICf
qDG/5IsICkiS3bRBAMifZAQyK0mFIwWtCvWA/S0EH2l4cRqtKbuMg7p5JOj/UPDR
DiAqG2RDoz2KROgPgOyVi9OXCVmYnoZIfUWaEh2xvmRUG7e0/VSEZ+wtZ9UiLVy1
GfH8L6tk82HopYOXlODVBmzJoP+5cs82OrrTHqfDciOnGyiwXMh2l3fV/Cvjz6Ey
zSUVhToNF5yQEYRKXWzou/RdNZa3iCJKPr8p6ULR4+oG57CbYbstdUeBVRkClFeX
ZVCsos3NxKsmO8y3Y1oyy9J7W2l7eE94/xQKGUlNPbXWRJAzw8l5FALSaDNj7iZf
BtEPC+WJRmBpoAylMe2II9RIHBHMPq80YilQwWnRIU3YGfxZO1NgIRAE8hEY+Xzl
iohL6oyNsj8pc8Ukb8XYlnqTlTs+2o23dztfaWuHtuYgXmXJhGwuurNfE9GQ0Xhb
OiG9ZS3pDnX7l7gainMISVbDSOrZDlaQCcaZObnT+IGIypMDEYliwjKfW8yrS2x7
veYY47kgdU/dfrdD647d8GLKuuY+LRXKu+eJaBWVKRZE7Wf4sAtynn7qfgsr+a2b
+07gU/SPQ0zTELaPD5uMzSuN4IUmE9Z1PDtp1L097XzLSiccYgdU3heSYIaD1AGH
1PgDPJrj+BvcSYfZNq24rwWAYtd4XPcI0xWXrHwUa/z2UORO5JwB5OVZnTyC6Erq
ghpMIRbOAocUPIr1YV72Sd5fl5FnXnIWi6Q1ugigcY6NI9uNrIER5G2kM9qXW6rl
MhDGRoWohdBiYoVTz/XpPcpV4P+UxK/bDxVEfDLImb2i8NbMV4g6JfnGO5DJfpGj
HN3QkhgCeQL/ZMykxMZa2HOe3gCIxNX2ubIJ7udYOXNu5Fg8q7Xq46wk7beGkXcu
Xo5JhChPec4oXMFs+CvISpUx2/GNNCgID3V5h8K35e5RGvu8XMqDddFfLwnDjs7x
Qi/rlLWu1yFGZm+AYKOafbDIKjF/wocEyN/iJ5dvY2PaTVpnTgiKZVoP2aSCKxlP
rVrxlkltzM7wMbEff9G7VDw+ciiMLPDssdIh+dunRAiMpzQNjhoeRaw2g5XSxOwd
9bsi/LixfV8gpHVWi773kh20BtwDRxyG3ITR8V01pQGUJYEFLu2n5Qvq/ZpfQEb3
mtGKB8PZscUm7NbE80YocUR8qmeUW1JdvfibcVTxn5h5jgZNxCu/XPAaBMPHdFK7
A+2t10dfX/KY+CIISL5olfDUAgTr+4lsTqd7sKl2tNfargYBq3DFMvaRDubi91UW
TvLIHKzNtqiVW79lJoPY2PwMGkt7+Xe/7Wq/B1EuKDDeh3gQ4b+OYWvNtncRdyTu
G7Bf0AvfAK6lJz4kdxpIrLLLc8V4uPkzWCqJL8bECZkcSGuUX/ICihHgCfUcH1ge
oLWsP7eVkIOcDVnev6yYIwBGie65UqDQ7kYWyuYgbDP4KQXmH/UNnFZqECmCxOS5
TAimYmTE176lHrE/tVViHMwvraPas+VhmTtakJFJ/pJrUdKLdQZEBqK32Ccm251H
yObjCExhVbuJMz+m3DngGR2QY+qGP0IAeUTjmW576PTHNAtmeon+55yNlP8qmYyA
b+hHXW64v9APlNSbKOONyz3/yQa2ZPJNPBkY8LpmATEngrihObovAuci7DaTVjIP
s5sS3+px7Xue1+kUbFOk1UTmLo6K5OZ78Lvbz4r2pwFmtOXL5kDjlUDDp/aAMfqb
OsmvaQd+HGl5PeswADt7LpdE03dl9+64mmpWkbAcu2ERGSa2mFrVatwn4ADnYXzy
lcII1+Bvyfvg0RV4oHfWRYPAijv7oQJAa9Wf4VC2/u4FewwTArFr1Fx2pujJBT9/
9aTDDbqdY8lgiSiAgPPyvEsuSG7flh6lDEABDmolYDv4AqhPBcUi4Lj/CuckI2FG
juC+OJchfdQFU5pwrfxIRJIlMG0m9TjwQuJRRS9LkE+Y9mBPByHJJb3ZiXsxYqwy
InWm7FXPsDDD0Q/3ACEpyjQdml2Y58DQD3rpBClDmkX+Fw3f/ABdUHQqkF6n5tWT
DeXhdyNFxRM2gQIWIUvgstwzwHbb+16tP85KdVOvozCl+ZrYoCYz7/IgwFcSmS0z
tJM1WNRCfyHC+dbx/MvAZ8h8WHNkDzu97qo0pUwSuuq6z7oQPw2A2gnbOOrtktoB
lmvG+qUJkiZgP0ijXNfVvHezID9P5UnrTMP+SZe6D5RaRpuHqbpILxtJq5d5FJfs
1UT+vVH7P5Kmx0DNEdYCOIhs4Ao11pxOhZGs6T+LbBoIo6u+9HQn1IKtezDM8kkT
ZhgdIFQKE3Utuqpz7q128sh9MBCE//xuRDZgodcuoAiYG1551yzw9w3UgkibzpkG
OsDJVNhV7Uk7r+Y5s9VeOe4Vng8RiWdzdgKu9MsK/v0ErsC6Viir+burXfwJ/Biv
7s5Oo3idzseOX7tJSN/t4FlSAzVFyOwiRA1g3x+n79GnrfTiqK1TiHFyRxRuMO1P
Se2XQWusnCtWLf6PuRY/rle9gIkqgxeHK+jZNn8fCg34ubhDUQ2CKECtwyeNXaU0
so3WT50PVWgKcLU+D4WxeWi7t50S9/y6zYQzK8QTIagYVX6sYtFhfwaJKPZVE1Jc
4Dh6xOu/knsxFDIl9YjlUjMsDd3QVce4fP155VBEIC6pqTRG6IUr8mmvTT9YWWHH
Xiib13/L5furq0uC6Faq6NpVSieDP7XtNUr1YL2dzHUaGXBSEVe7fy22QGlP7rF5
rUXzP4OWehWnLxHN1SMKdcRG8aLBLglk8c5ua64RmLY2wtr4KWYfUooxIa1ihapq
s9UXhfGM749Z4abC5p/bpQ6usYqdMIeyTQ1RUWlRX/jECxhcLgV61Mhvo8TCF5Em
vKcXLiRU5o6EtiAteLLWKA54KygrbMOX8SvY/z2WlqWsohr5qwSpAlrV4TjFxt+w
2gJrPIg+ulXEghmqhs7IJe9A/hTsB02CZEVbyJsv36F1F1SLwKXbVKjj3c5qydUR
zojp3C6KieWkUSx1JAZNTtUNODTOuANZaHTnsxo+farBuL4Co76HqFK+7J+YN3u2
kdgrqpBCWL5Lnu9+VsK29GAKCMXudpQHv0i09BHjwKcmcnrTXFyBqV9SKJhixXsi
wfKWMOTtyULtDcZLIVH9UOAlBjWoZUUHYXJUd8TrtDg2zBGwUqmMMkQoEXR9dpiO
6WQiG76ooVw2jQQkf623F2HWmo4roi3MGPtyopXMmRU/jKJ8rzENMVqjqA8DN4Hk
eLnu9ZYnN7vZqTiID7X9UrsHH9/1HfWMSkImBTrMIPI10NCpTsXOBpeegpo+Cn5i
9tRFEons+qCrEbN0DJVf58zD/olkKMGAkCREsVvuqXLuxfbrrRMly1MAUDfOQ0Tu
TZqLm43pG2xdQFmOAnQRErrta+yiDLw4ELml3lU+5YwTN+b7Wb1belA6PpQd04UW
IWmwNPNrcoCuf2UfxGn1Gfh4eG02l8FjEMXGBSIZLshX6cnV9gJsMuyRL7VjtbdO
acPMHvmaF7zfzlbEZ1wQuoA2L9cnTb7hMPuANjkxFaq4MKUvckDxF5Q0njoN8ioI
6/bSCSwk5V/v7j0x45TxI1mSa7feiNL2Zqk2UMgeCK2Mc/jP9/JDduMk1absBPOy
X+TYLiPyTnoVskDj2Wg7mqPv0xFqrjpOkxr0KTmfVAeaXHQIDN/PyAQ9omPmDBLl
yNNoEVbkREcWf3DtE/PoJoWUyNNU70lJNMGwB7c9vMk0xOOPdXbXQj9RaH9F67tQ
XshSfbftfAj3ge9CSm+Ra2Sj+hhTI9bW1iH/8yC7/3ZRAc0GpQRIJ66EPZ1O8sQ7
pYrrEZgv00ItJ2ha55KX4j62XrSHgrqkIlKFpzqOHgfZA6ta+kVBzIVLxc11P0ur
6glQFa2QE5ECLVe8lQU6bchWObuANwmtKjd3irVeUMpF+0IeUZpYkOXPemEPr4Ci
it2De1OKsAvKy8hNxyRMhpWZhADxRfGZYbOM+yNFxFUb33S4x93Pbhwjt1YRa3wo
D3dEv50NuJ2W565DsigMlEP6N2jQupR903KMXI1Qp9DrN0crgGY99EEjhzN3kEsB
7CGnZq+mmB+dLk0dwOHuiwmDu01bEd4pLV53rp6FRV4z+yNtWJqLdeAI+NPkAfJi
YirVaWpv/xQpXZMVhQGRNVkD+uf4/kmMMPf8FiOV06a2qFhlfTxKbtb8YDupKlcJ
om1FOl8o6PImsVFAEqZ+hb+OYfOB5osTyXHWsK8cmWXc1OhU/kXX3jD+vce4fIO3
LNmxy29I+YnZ/T1M3OjMPucHcwFIAhTZ8g3rBXcNrOTFtXvmke8xhLY0+6vxscNI
KPTPN6SzzRe/95qga+o5BsNv3W2mZq8Cf6sS/DxKtiXolBuou3K+KhqqGnS49QAd
yDI3jLf79iZL4TtORFLFlKkKDbVqkhncETTAfSiGwUBqz80X6AGZ6+Y9Rgutv4TU
MuwqoWEhe36GayTSVYHSZ0v8LgARtH8p6KhYknNu3JbWQhk9mUdBQqBxQZyFwK3G
HlV3ofPJqKd4JNpVSrMxlGerXpF4Ztvxs1g6xwztOiF8njBVViAW41F8Hv9M4d1i
zhFLuwQkbXSwF0B0SzdUPd6uu0cyoLh9ZtVLFqj1RYJeHs9VsDR31Y6r8XImQMvy
aU5uiFzR+D0f6nRRf1DwIgGtVlvagSYwWnKEU4+gF5Ile1vsk/pOJj0wbhAielnw
frIYo4CTD4ZV3TkAJZF5lcSvEnrAmWBhnYGrOnHDSxsK6C2PlwKNFjOzd8M0C9Av
JmRdLknszDEzFXAp1uzAUpJ4oGsyC1XtXQTqPB6StWKcZdk8uQ9RcfDnz+HnvYI5
8noWc9pTp5hW6Dw55Xs8yunnshR/nvcvDjWUzcvOE4kEZowOSxi0Bskwf5R08ToM
qD6BzqXzx+aH/xoy8Lqn5sut5HkyzAwg18K36lMNCXy3pJu3P8Xz5ItDV77UwNGD
jVJJm6hq/BE9AACgCmCCOK7SySs2EFgdPNLD4dal62zHwEPt/1k/JEeBSpW0Ek8R
hfvpybndenDPAbPI8JSf7/fZqiUV8YAJsU/LpsvzSCaaf+jpObzVU+7faFqk4H2h
LdGn41IpvAbQJKvc9scUFOYFzMZWjqIC6nKZxNJXi4D39OZ1BZZXPPThIgLjCGaR
yeqUhkaeYKFkHYzBqTnyWqCNbLOD0O/OCbL13UTAeuvB7HS6sh1DUiCXYLj+5nuA
WKj3cozWnlPEAEKDbFTcYeHbr6AxJr0P2TCOf2t5LzA3sm6TACW0v5RkGEjUHoBp
3K0hveZbjL/SzT9stevvP7HWLqcpbY6QXJDfLPby4UtX1xk8qDWyXpcjXuk+q5HQ
dH6JE1a4r8SxMDvqVre1lqLuwpGbE0GpQhL1ePppSmzrqaAsNlCpB0Vk9ON4So5d
UyjHz07n5fpR6doTYa3ftiV6tIWbYY1kejZOksipC2b54KbRP/cpJJpX6Ol5Mt9f
Od5iVbt25qXVOfz6ibZ1ufE8XSrjg2YE9sWxKbru5W01Zi6HvukL2h/DwDr9bpXa
PpEvisVsgfGXWqfBig6C2h9h7PpSKTfA3JuUvn30b2k0AQHkmttTc/5/Y08p6Gew
IWLzNHK3pqL/zkpgUH5HelT0rDQ8NHf0v35aDljDdz222mn+1VRpt9J5AwN8JGIW
uu2J63sfLfAQzHQcqfBZWPJ0lG2GTGp2oFZMLRXvKLL/x98/RC/KKUQZNohlcgtg
9qN+smE3hW8qtJN5ymawouwYXzX5adacRrppP7TvhEo/kl1VH0g6a9LZQ0gdkFyL
Ng1Bn4pAAppEEFRjbhqhOH/zD0xK1U8G4iEKFZGxh4P1uJXvT3vTnBmepDKDlUtJ
vfW6kfK2taocgxie5e4AKgsVh80OtoM8KWluLTkRmS2FQ+u+SjiPi2BmCtLwqOIN
9y/VZMzSFHaoBwvd8QjFN9Bq714e2/EChnLjMsJgYT13D7vQEw/XZ212j5y0GIFd
OwCkU3Emin7JPAQfEB1KWDQa+rjZ46hGBEi9k938+6GbREz769oIxL1W9BNH5QBW
RM+3KyHV5V4Vlmp5Mb5X9Tt6kcw76VKaF1jcgcMc1KZzluP5oTzG1zYIYlDLH2aU
j/0KewhYetG15Sy75MD/HoS59yWh8Iv+kw8eLbrYEVw3qhYl07Fpp4gXFjQmltBG
Ef5Y0QieVBclt6WDrbAWGpAQhdF2iN86pPR4hHFd186kscN5dE60LE7zOypfjdNR
yBKY8/hi8aNm+RgSH8GWi2qn/42TSpk78bSuTUsGXv4aBeJgT6WPOgFEoVD7iq+F
4iOGUguayDbMy2pej6wJN0F4GqDA4vxPCgZedGwPhjDxk+UKZTGs6YFDphdALFZ/
LECd8XPwBkbDe6HvZX/Uou4i6f6cd6BCkUabIlzZdj899+RT+MN8Tm5Ug4AEMiT2
tLbeA+x33LuNzyi5tznQTsjpegVTor/t3VXEkfv4Ad2DzDK++BPFw/GePUUFOI31
gUwp/IdXRwQhlLU/W1BqqKvij9uDhev1El+h7SpkQEJZvzkvnCfyz75WKj6A5Y0W
zGFzIe3yxeknC/4XCVA714g/iPee3H5xxlPhhlWHRoWSaoTih1YCJJD7ooKpFuYQ
oRHLZ122h1j4VNUSImHbJ/FVRdtV7OEZHEwBz76bWxzfRpsxo0hF91MzqKHF8q9K
eOkKuNI6tCr9B8QUxm81QJ9HqmrLlLUYKcqTcc7LJP59Oh0h+wKtDPEc9+b0DSrt
IdRr6iw5xYn43b5y31SeQg8JNFkLKuoZS5aK9dnlcQYZD1YG7ffJ3KgVNqYbc99x
zIfuNZAlIG89S6EX+7wmchVit2pYBozs7T3hQnAnIxrNjX1i9iJh+NAxYu3TtVYh
KuhsI0bp4ftgLS74SpmjpYV8f9GBNK90hHuq9N42dIqAy5QUWhOW8Oib0W+/DQS1
4Qb0tb0h3mbczAwC2v9K0ADlvDkChx1jNZzfdobCAYl4k4zrwRbuUO4e3HcChHbU
IR9u8QbX6NzMwIYMXpNpy0lxzlqrvmV5GkOs47NsS6wFN+1o2ooyd28i6/NqJngg
1kk4zru3IpcJYT6fxi46PWsDOorcsrod334Z0LFQYcNccIp48FrTK3Ie1vg+qHsG
lag/GqJR6WAvomHjwMyakgH10l0gDnWcHcUn8Rxj8l+yyIGfMh8g406u11So7Sr+
x5UUbuMRga5EBBN/pfW6jA2YqM224BF+1oVDE6sksgcNW041QDTilPQNxhrLGZcT
tqLWiDezXyygy10tZnIYdrgH82zqrkWv0pWlj3EBVL8ETjY6V9nMBdy4uMom5xlQ
+8zUpm5/D9Qhrtkr2HMcaDkqAS4W4HmDgw5ferdhjWIUA9MXTjqN6RgnY5AaOQrG
DV1cp4OrcgybCBhp4+r4EhNiFl1F+5FSQittawam1n1jUkkzOcJvCK9Sp3Y/NRQT
mg/DlN4Y7ikQXgqwFFsfXY+6GMCRDhTXNVshEWRjhv7BUVKOtQL7ecODY4VVt1MR
spQeHkTeK5uhNOe9aR9GPVWMvZ0ri3FNs8v44QEkK01xBtWvqTAW+fFdxlS3gC7K
BZNSXa2YyP9md3TvqUhts0I8ewQQQLQmo+GPckwEC6MRew7oNwQDLUmZiTkWU0XW
OUgzqXUJqMbMc6F28Gq4njqrMktf3PY8yNPCBhhSinfA9yZQNUC4rpHYkMHEn0pP
XGftSqhsS1VS4p9uNPdJlwnmlRi8m1+QOkp6XXkPx59TGXsGx4LsvjnSP/87IhRc
iBAVFHYR7qibMrU7CWpg1xVtej8067JL1IKE6eozSgh+KSFnIoBsZzKJBtJ/XTec
FLebqWa+0D0oUYuT4TJzV4YGWAkRmRpQctXZBPYhyHR7hw1MCC4TCP8aJkaY3qeB
snD3UTb6cFPdZW/pikPAHuHw/c10aD7odjNzWd+f+ZSsRZX4mkdYo/J5syfFKU50
Z1UUoGWCNbjMGLujlRs0rgalFcnWr5fLmdYRYBgN8V9tIS57O42mp2cUOFbaF41d
s/vXJB3k9W28ObhQxdXfYx62FUzJpB1Mhbr2V8thiAnxGRmhYThg3XcYfPlb+PuR
exKBYU5t9PwKLtlqTbpS+QIV+EjT6NtgDdNDU4HslLKCib9yswHnjocN5lL767Gx
MGdfEAOY5HVZ7+MBDkxvrPw8xrIDJ3vSrvfsgEAUUDx2jKroOk/MtJpXVvv3g7tL
2zhgRSWSfMP/uavz3vSNKlo8lsUDDWUlSqJml5ATCW4iiE2jQ2OKsV6C6BByXIef
PIpBkeHE5bAAsBUqDKNzLls+1CpQWqyL9pQfSoEQ5YxAB9Rp/Xvh9b77AN9Xn6Ql
UFigb0zUHPHpp685f8hGffjuj3cTh+oJ2fIlWJVydKX+DrlYLWDb/kRL3imLTqcO
hp5VTNXX/rT4vl23+Ot2BiIbFFW2RSGpZ+vRhRghBSQ6qoyQDPAmWv4wAlkEuKB/
QNMjD4wgl/JQg0ElSuxDmmCA8NuZGE5sQkf+Aoy7NYmwRcFgep8QIIVLNVvCGKNR
3g7saiMDYt3odtWpVBgN6hH10ihCvNb/lnZCznX/gjzS0dnKyTEZtx2UC6Rgk1xY
8W/Vg/+R9WIzGGa+OJqi8pFkjoP0VhmyzcEEBGP66quN9o/BMzIQfcPHKuRLNnQy
ypdmGZNkJbldJ+IRmf+aPu3Xv6nxHKyEgeBSbSeRHAgF8JJaUGoXMau4Z4pejqrv
VzRYcrPpHCZCkAjojGVaOPq5pckhfM+Y6u739frDZ+A4sGy0jK5EGofL9CGzjYuQ
dtR77qenc2ixW65cm6oS4EljKMvWeUUXrVReDel3OScmmGIdGu8UG90RD2RcZbL+
8MUXkF80gs3aEwKcfR/dxzacngF5aVJzW87BhOdoH+KhaaZLkpm3YLGy08+t4fhQ
n1C0gVR+S+95Hd/y40GCn1MjZs5UpbrFoXwP1ZsQ4wIufKBMG0lTH1p/3zZcqv9S
LK1jLb88xVR/WMnxB8pT/8EeQt6JZD7jZ3NFi/93so/7uiQGkXxj6/V3ixMBy9xc
G+vzn9kYnW4bBcNTQURkBsNJwGIT6KInp/dqcEp9ICuibAbcyJXl4SPqoMlCfQta
izsnxNFkXUQ9kY1egc6SPVBDgxiEqdSPCsekZH97V/9AihqRCFZ3b/QcoSYJDeyL
RynjF8lWgAx9sik3CzweQ9enT/1BXV2zlW5ipSsYSvixT9pgTOnQ970ke2lzmAu8
THYfF+beJU0KhZgvwHaNgkzbgzm0V3u5IRPt5rH3jiGchJoqpYf3ZykUSP8qHEzj
7y3fZy5m+fFTpFPjfiAY98ivdHgsRDkB9ntt88yqb6pU7vifllIqZde8cEO/r/33
gGQjq/iXd6hCgFjRopi87IPMuejj+I9graaQsoT+cFta5dnTmPMs0xMXqUanI2M/
D8//QwT0e0EVLtJ2aPEIsqxA5OyAhAO+Tr/Ykzn8O1NsaiXvkLGXc8K43QzgxZ+J
vQlVqdJR2kUlBIoKqh/grHDMRhjmP3Ocn2Olxhvm+vyZSZLtoBfTJc24BYHdYEB5
iU8Cbpjk2+YnfxMYrV74uWVK22Tp/xi/AdmCp2Q3pBr93gT1/Bn7+hW5L5uyiZvv
17aA0maBUf4mbPiAH5JEvRQjMW/U+kUyiFcp57r3GhcmPgIZ0w+PXMEXkAQa6MDB
eOVEJ6NPyz3WYokVnkegUsgOSLAIG2+pOOI4kw3/3mLJb3QSofq1CvymzcjEiX7L
r1vx+FRr1KDttQJLRNbiCmu08KN3tZfTlMuOc699u211LDYklnm6VCtoAVfz4Cep
uexZBP2YZmMQV1RLGZSdaqq09H8g8BIxKKnCzXPq+br420EzVKkDD1bPYYRBnivr
F17k395BqXxFcMjx9RA+h8bFVsHRavFEfNmzjj+fYWsWdQx7Fd4OisfYWhhxK0Qy
10LZPRdr36QN24ViO4jVqBGL1TgLc7Adf1S/tPePVsJ0AspxbhVxqTO+Hh44PE77
nFj3vHgH4WoS6S1Z9G5rKO7AQz1pLRxe/YLUHUgav7hasvKrTUgIozr0zxEeEReN
h9cxQfkkkkhYr4kIz3h7o/vF41+OuJXb1jkSvvrqUjVhXrNjJBc7ppbhfhvC7ZNZ
DqN3jdsxhKQenQar2Ip6F6ZwEBsIbAOd99nWSMjAeNpHAHUV4vcw1E3nBqWAp49J
VpVHH1veERkD0ai2abRGs10b6fF3DoLggg2K/cmQhhqHx5PHPOuv02FQtbQK4Ayz
u0R3KkxJOFgMSz1QzF9RCyiLCys4cCo7gIXK84I37MEoO3pXurkNtWXE+LN8FjWZ
/PDVArzquXHmPEjPkM4qsOVAZv6JM2cylMgKwbqrUiTCJj/7QAzYkZLuVAheEaz5
PmM+KOWvIQmexglxTzfrckiQhP/tSwxP6iRWtjUEow6oaoP6bLYggWNfq2U3HizV
0NCm98ViAo8Tk5UrMMan2gsLzZPWSYuL43Ugev4tKa8XqQSrxN9y+MTJSxURNDrp
MlRWB8/mpW+ZCLMvbg1R9zgoh1gEL4J13f8OMFSwDe6gC6SnhopcBIIu3Fte4pS+
KGB68gZ8/jdn4GCf3Y6idtE4eFeROgPxLHzdurdNJtPO2SkQ5icNVXfJFj3Tr7xk
seA/T7oKOcFqXwD2aozsxOObQ3P5+5Q6Z0cYzOTJNnSTzZUjSFKFR6SEGMTB72sC
R1BdVsm1pD5mQ85Q3LdMFuT1AZipld7P5alj02wdtMgfsmtts7Outk9AQlMDOQ42
ViJVUNRf47BA9fBCLKvaTTTfK9jcwqpi7x3EjoOXZVg8iXSkB8JdF0w9CW/4S1VW
huVUQB2aHqkUQ7m5oL/sdyCrAdKU8taKoR1sE7utoP/0yw1JtE10ELsU50RIK5uC
XQHyEAaUuOSvPhbOY7SjS2ny3yeduEnsCPE2CoP1CAgvM/IiQpR9Wiz1rQHhWKvh
I4ehIqrGfb4XVvjbe6rENeOkwenP6RPKGSPOl+CMaePeAcXuwhSxLFxkV9A9QS+g
b8DLSdyDWkUDcCg4qBesuPfk7H3TtsVlQHufc5PlsOb8GbuuzI6V9AHqVysiqg4m
Jbk58lGSB0v+0sa42YcGCB9MkUuIXR1Ugqcd3iUqtguSWWSOO0vHIkCozyh5i+yb
EpAtHMUCi4oL5yk/Cg8jZJ/6Ix/j2Oz7p8qnQ/4iPunFIpuoEy+Vml4YBb3jvfPa
POdzSmuaB/zOOn+Yq8HRi4janW85d1cYNr/5FZIXV6w8zNr6HxN0CcHGB/1BhDdj
j0MK4DxqipaMXX9eGaLWdkyqDQuWMY/boa6v1OBuy58cx6C3kjdqb3tf3iwuB7Yp
DmfEA8TWTHk14gjMJkvtQl/Jo++N9Lverp3gCd3s+47msQ24aTz3YCR6cggtFXCW
W1nZrRlXIZcY3OVGytF7RZOvvu7LoNrRWrBn9z2iFcx3gXXpgO98fuXUgvZGZAyU
9sxAsbIeq78SnDu/ctSWnvskNbS6pO8qXTcZ2dHEecPqmHhHhu83p4L6tNB+OthL
9EO1rUb1mPGyfyEwte/4Qj74ZqVUJcMXZkGiBOn26NN0FwO6s7BzgO8l5TXPgkBp
PktgGlE7KaaxGBhRSYhldKzKdNpqp4XwhvmS/ygxE3INAnHs5ssteLWq3Qooo5bH
YOf2cVOEJoy+yHlguzl7Bd9D9WaX/zipcTjP68xiphF3X2UejdF8x2/TZDZQ0bEC
BbW79wK1T2hYkOAf3/k1QS8plshVheSK+dNqwiJrFF7LZd603Okq0rccl3Vcjs3I
TSJNLGhnT6N3TbFnVr8rKA089zDVK9si51k9IQ+vrsSvtK2KF+NS1GpnXPrKB+Kd
ouLWBiThmea0LW6nUgHhBFPA/lL3WuRrqfsjM/bMkT9e0zywZe6bjRt8+H9AGrBz
BEVNOYp24dgYpX3Uwqz+7dVGpgwR8dV/QWFkBgLg2jrTioa7vtqBK94kz4JILZ2T
iUb1HaCaVdKKd3DgXh6nTF6JbR5JSiXhL43sFSKVuWCls65C9It2dE0gJFDlKxov
FPsmm3ByID34wW3zgPz+igqM5uar/09X/hQfUw3kuAcHtbYfuJ0lhr/PduowoYJk
kmQ59av+Jjqme81J/GvX+Fh6xYlyFOC3gT8jANvQQFGB+3QO8uB26XlYHWGXw56W
hAW8ZEQjssqMjKpMppQI54hkZOiAmhFqXSKICuy2AqiRwGYmrTRzxTv7d576S9Ul
HqIomoHHO8cWA4BXKgZsrcNya1QzHtIdJMGqDfjj0j4+VfIajPJiQ0pt7Jp6cSkY
U8khVGnELGFzusiVKNKCl2t1NZ2bvmogIMgSTDY+rYgY52shDTA29o08LtX+HHgh
st4oX9+5rxsibJPFjzRMGI8+UccFwOIxzpLouBHui42HF3d40vuxJVXQxnUAbqfq
UpBNaxOIxjm3jc4s6WxM96+8SX9YjRYTvbfYgivwWQ7fXMyY86Jgf7KgZ2fYARfg
3Ku0BUSfbx4I9ocfF0so8HsXRrbh019TGtscCbWwFhQY5m7xV/mzpwq/mePYz7gE
PtWBMkeV2k8QSI9d9euFrIlsDKSj8Ou7SBzvb5z+cLE4ShIAaXt5mW92a7FN2fvs
MAle3/2nbINXXBxq5JngfXk1vtyCRE+lfZLihY4v4uFTTu9Lz7o3wza+TSr0D63/
RLk2BiAmO1cQkGooaXePSBCt8saZ2bnjW6hKJSx92JxgIseoEkhFIzWII1NEDxmB
1csCqjJV9MKz2FopJMtJICnJeFzvgvMlPQcHgzi5tnwnqf9X4SSTLo5ucD6RCpaj
3Cgkxx0PPhXCEK9Pl7pRmbG4wUQ3C4JqZUYdcZtnD2POJDI+EBdRqVmAbcD0/B4D
oYqfsw1NXptov3L9HYcWq67uUKkEVpf98d1qhL3UX5c5YQdJuoEYCG39YZ+8jO8B
LSJ74P2GwidgQ2CaliCGBuQjFUE0spmM/cVCojujnCkqTMtIHXtZPbP65vw6YIBL
p4+R7dGh7NbfBjXzeVEGYx++/Zs6iS+AxcU2xDdVGv0g+39HdTyTC9ywU2AWM45N
4pPI6EOoIheoesuRhB4b0JoroXNflGMgDI4VgixRz+L1Gycfw7OHh5EMHSIg934R
aDT6r8ecZjMowSlThAyCD7DqQdD0OQKDfijxUmcZNZZ6N+/KV8jsa+uo/1JqHZfQ
rN4/SOzZUWl6hE4Y878E7UDG7hngCSmEOVagbyoMFSaS52LghnKt5894ohslUAIV
H3qwLGNYj01tlP2bI6hBCxt43zJeL49n7FmUj4uYm3w4MdqOLHlbNFSVRZLytjWt
Cef/CbrSJyNzWG9Rd+cXozU0LfYvAA7JzKII3r0EdDtSCSiaJTkbPzd54/ZemfQk
uB0egR7VZ45PHQvLsxOBbz3ne2tfCAeBTavU9PQ9PipJczeEsaWHTddKmqjcOBfo
BmXssfX55YcZ3rsbJ73abLmsBS9eTEyQu04MBDrxAjDuGGZ6VUar+QdO710Jjdce
2nh/jTZ/RzoQbOPdtcOS9uTtE/OYBZ2exppAOSBXpN3gtN/Qj+l2UW2ZrANwkTSt
PK57f7ZOUce2IbQg3enD7p1S6zucw/oIqso/QU9jXJLlPK2tqMDdpOGoOr6/1Nvn
xvBqADUHkzpP5qu2h+fee/vvj4ts1pg1ydCZRqcfq64bBX217it1yoUCvA1e+MKg
82ynLRl7N3yji+Mxi2OBiCLalOKLWWn2XlHhPx2L4K1L+l6ggKGsvA/JB1/E+B9R
zIwcEX90KNvp7iy6aUmopyWaYdw/FfQXKfeCe8OUmCzZ3iNaRjJPmTIvwMQRT2uy
fARiUnK2HWC03PMp4vxUpBJeFCqfNQK4c80c5dH+XLQPMz21uQ24TlzIRKqjc9kV
9C9MECAT1sNsVjS0U+qF33h27XRmnshcRVSSiG453d23s4dY0aR+PXfdCzF76tgX
BMn7Qx4tgSCWammSi0YFlcx6yrg70mpWuG10iyuhwai8aKSzRpcAXbdxgydp5H1h
zgubClpBMxXEFdlgB+vtzDRbFKx/QhEURlhpmuh+/txY7Mj4LKok9WX3pG0iDebk
S+clVZ0JDhJNryfirJZnQvO7O/uu91IpzoMSNqiASVbnOXSp1QsYouhPoi6jV+Sc
ONaXR9E60sXYfV0WIL/XHENSFCQ32RiWzxMe7W4WmE9eI75QXCBjzOXm2wMyZNd0
gFRXlC+lBKMZLdl5SC/c/tSxnoS8zjqreAlwTpTpQU4j0x1FPwHqqmPnlbUIWqWp
0GabyuoWk/GKSzJlP8LxhhnQrQb3Tlwk20vzQqw1BV7mi0VGmHvlZa+zeg5pfZx6
rH65hPFeSs2aVhsR+g8LhPO37DdZZZvKh9E/3Aq1lQkx4DWsfDI0/d7wUOEf9qmU
NOlot9HA7MrZQQl8XXzwsXmPa7FvhJIImL3GSuS0J7+bBnmGl0sN2kdXcfNS06Lf
d/SjfsmBBteCuznXsqe5DNAwAi5xn/kBjTiYi56x4Y2qygmFEBTxFueiL2vExUVJ
VZ4chB7HwCMFNaCecE7GrMeMAhr6+KlGqEYq8IG/jAFaQWkaCzveB265AD2f1Cod
VNNGHyS1k54TwW7RXL1ObBWrBNWwvVUg2SARmvYKsx9ba096NUdoIrprsi5mYQJ6
5CeV2d4NPlfgBUaWvbLpxe2yZ+EXjQU22EZbUTXw7jehvgU1wPEwmA7ETLlaRCpr
hNJiDEb3IsF16V/T37Sb1ekzs94AoT1KLoL43hAzWf9AQIQOMco6nFPQwpFTOLvH
UuuCY943B2OuLX3jx92EQRO6wnkG5sFEGtybwDHk7IyhgclpQtp+tajmQXj8X2S5
IKwPOiK1rJhZbmoQ7oHmV7sgZORLB1TgpiVyDMuI/XeHGv99t/VssUeSadfwoZBW
4B7f7XS8Uv+z1OmXQQazbpsGvPKZvURxsu1cWeKQoG8Au78yk2KSf7fkTTsDdEHm
XNZiHZghiQ56t+wuueCob/8pK9/Lr1IkKv4WpzXnvaB2VtfQ7TC99/s/d0UMX7LT
cQH7zxvbrar4Hs2rn51KN9clKSDsJAKWwD5Z9p8ynacp2uVrK11jgJuq1qOjtAVo
Q07tGtn3GoWPY0iWJj8IV+UhvxVOxkTwroKUmD35sleZW6mWVe//Wf+6dJJmFQcK
TKxPR6Xm7jsZjPbtdJf6Zgn41zJiV16pVoFMR46aM1O/rkEGOntpOVMcSqEiRnta
mdkt4A+1RpxQFchjK6HeX+CzkS1CSEIgQNtbHVbKk4u6SrvCWEw6kVXRawNEt5PN
EQfOQgAhDGRpRCAhk3h6SUy6B7NjmyEbKWl2KXx+dDyxZsYIAo56YwKnLglCUpYl
OuFbZKktzUji9OCy6ybZc9Yw0HyM1tH4lnm8Sc3kHxLxq7zE498aS1g1Zf1vbvWh
MnZ4h5JDUlux4CuunfZGUh/jx4pKotc6ywfivuHflM8gF3qNzQ85YwZpMwCmyVal
TTDFapEerLK5WtqcmK8aLRUt2Rz3VrnfdJ0+ObHQ9SGbfgyQ7PME2uy7yytMo2Yp
c64sY+l0lU8sVV9JhKMslXwZb10zBQoM4Z1dcyipssHgUNpD54LhceFO1Wb82wVl
9GuQngRmNOq/e8e7cUpfzEiE6rW45l4moo9EefaZY8Rwo9yZ8/u4+rWVmGmmzhgw
iEu6/h0ZR6gmJ8B16wnib8wwAGE/fhZXBoPnipMX8wxBNhyCGsvOxaTLfD0HQcKA
Lh+jNLnsoomK3RRA7X1xB9xL9pYvsUK+0R1SsV2P55lIUMb1PPewfWGiLrHD1aoc
ByT0qvoOwg4LDCNT8tOKkIQs0xEZ6GE0zEgm4yRU++j7IqaTNMwhcd1e11PyEU8Y
kPjnWdh1+GIVJozgsC1RvHkSu9QByyM3rn/0MJGsf1vEO8967n9uk/xZ8ULB/wy9
UxhYj6ivTYrrGep1rZtVeeiI9UbLjBH+1mNul1A1M5hAQSpR7+tayU5NfKP3ihLX
yF6RZ+D0LgbtF4OddllJPAzH152URPBnPb6HuVb5p+91G9zSBwK7P93jqxlQO+Qc
iU/CRecssxga3Ds/hAIsJX8qAx0hW/QHfJq2Jy5Zk1u3aSU2/79kalA7htUU+qL1
g39qVfSgyByEMHkHoCMfj3+Xsrc9Yh9RhnkftpImQWlgrqv6HTS3En3kWsZCNZ57
MxYMytrowfkzsihttNVQWev3Rwu2A39rpIX5OP6qbraUW7dVchXtKf5xrsyvbY0D
H63/RPcJ7YCf+J8PmuWKsl9b4+ct1arayJPIzIcMXUgj1Zf1VUDH6KfA29HYghrZ
+5nfNdFpCldXKfKYAJbiHlFXtn3bP2fqJFRtqk7WzWqrhF93mfq5KptUDQGoZ8Tb
U+Cab9WOgP5P29+iVfrnXihJwtTaOJ/WgyweXUPxDzYfKnvZcF991896SlNGh+hD
D6fNjlsjMA8p/uNs77Fqv5XPBDT1lY7fWBOOAjn/AKU6k+IEXHKtTbnZW+zOgh7l
xFwXJx7fJ1g9VRkzAaa/3rZp/aIxTPjiCZBJz7MLSiz3dGrQMBYc2ST89xYHSm6d
pLMWAxpnRb/avobLx8K4GebkPS6cb4zxJYNBNf/dGbri5okKTAFp9ccsmaAvp9al
P2cxSMRJdSDxHKsp0fqbVMuKflY3LcztOFgS5PzBUPdydQGe4959xtw9D8gbZjOq
wglAYeYR8TP3ANqUj+UqNWkbsDr5qo7/uOuy35VZldCOv/k5T4EbDAgKOvBg6WWT
LrOerZJ8NOC0RB2u1tHTw6DRoKBxvaYSOzKPDsA+JPaxJ1SCqMrjS3xJtpMMj0Mr
zhiVyxEnzO+4n5z0qU34nQIDKXBlIJEI2zfxhF6szSe4uK/qCmDhx8UJxjydtMAL
NSlg23NcQlQAm6ZIzwMqvhS2Skwk8vEdjtUfaNhyG3kSf1F5i0vEpgCLlvUXSFpJ
kKN3MdV6wi2c+dtpIF9uY21MSJHhtRkI/aJVwyKM+c4KeXyMHr26AvKX6wgwMQ+j
qoPt/QIuDs4e2hIEKi+UbAJHphoJQcJYkUsJVCPX4PTRRX1+ObBG7cWo32qtsfLL
VevPxBAFb8OhhwZbTvvDUBj16s0POFDgfjjCnxT9AWO4SCBZlJrSlzz01MVP4NTv
CPUfveUZlJvU4l5J3XecJkxAGbnjMWkOYT1mVrt7j6REcaQQBzn/YSIPGS7UZkln
WPJTT3mGO/4kA4okmNDJwAYvE3jOLgz8KNm6xdsNz8CClW069TQu6/WHcD8GBy8p
isR4VGThX9AjMlXOLg6AZmtOxCig5RdXSiBqknl55V7WCq09sQW3r01UPy+szHwc
Qi/dQPAp9u7DcnH85PAnlKAL9jBZ5Jps0+oSl6vkAmAU8yqUfr9c30zFjPHU8ZW4
WEeoDKamINu6jyn6lnnvxik1asrTX4Zwlf1no+ZLlv/Nepu+PhlHhs/jEGAHq3NV
d2scMXt5zZ35OOoCB5QgVnTklwxFpogAaSn8TnTe/0NumJClwaHhZ/3LIOoCcnmS
hJlvN2HYLwzBssdkHmxflUeo8KCjXHs56CL11w2WMHvr7P+iyO6/aPMyfy8e1XK4
2tPx/Htpg5nQpZT/We39/nSlU9ufAsNazUH4XHShPKn8II+ijHMXHKQXpx4ZIQow
C6BrmU8Jihi9aKcb2qgS4Kx0HjfNp9EV2AoCF6rmlelZ/bnvAsNInupZKO2wSH9v
JYER0s1XEpJSehz/J0R/RZ377vCZCzsW1oIG0I6ExgL810HF7QbedndIfcSX1jkq
/F5w1Rp6Q8/VbiNQUl3LnM3vxKe4vQ76H4dBTleC7EUkOABPFEJckZgz2B7AhN/H
BOIcJLyN2Yj+Xpfu8GeVFVT3lq+DBnLk5EnfCELad9bsbo5RRRQWqIpQV3Mv5T3Y
0tRmq+/6DwhsPsDYc2y5PyJhETz4IyqhIO2ZBKcPBRtJga7C7OLT1KghKJqq6ZCM
TzBJub1hHxQBjRb6vT4ED1Ll1mlrEIm6X7kwK8gSZfCTOXn6NXvgLLYfa/b3iEMG
2Dpqi1apjGB7ekQrWo6u/4maEIi4BMCPfEkYsml9ek2lu2brhwYKUb9MeLfxtmC/
INDkMeSGRONF+aYXaBd2RjVkknru07+BwaLG+GsD3nE4e6tZzcNJ05i+cGKuFU3t
sr40x6rOj49Y/c1Lwvh/zRXNvFuzZqozRxTZ9f22RGeuwaNfbIzgtyIIuAK9LY3r
+UX+mYVaEZT/EsxXgHMddPf6LI6xGkbmIPhXJQMMMGlLdX4DSWonxpRu/3wKO7px
k3yzp918VZ1nkVkMJW293Tn0ioVG44ifHPpbCot7/p9swfzrm7NO2+PPLRVRteP4
2gmg2uugt7FwftbCAfT9RutphdxQKyKvsY2x1la0ooh1JXamsLgR4wLQ1XwDBXUV
RqQEs1Sk4Pic21aQ29oTZLKx3nmzXhkw3y4yhsjteqr1QwbuhMG1f8i00WhBovhk
/vHRdZA/9xPfU8NCPsXEf5XjH1byUWBCtYCCpFLcX4ZLYuVuJSfHdKwuKAZXkOCN
F2wrtq7F4vdKBn2HV79dHaHbEVLqPScz9oDtbNv6F0PwIRNrg8iG6WOZKggs4gLI
NASq/vjrcKn2neh1hcsGGzuHdhBJFra0VFXhx8KfmZT6k/rODN7q40L4STlbf+U6
h5cy5hFF0TB3fd+7w8ZO1y6BDeUyrmzaNm1bt/4dUMlR3WuLwvy4zz3U9/P+Lkxc
yAxMS9FB0Gfp4cBcnYfqIa/0WOr8hUwk+ChQgvnxsRfAp+2tTtFfprykZ0gbgeOu
qp1Kg63U83yAyx20mbR2L5DzZLmE0295roy0lHo/AL7fc17BY5DOzChccr1ntC9z
/FRCkxj42KJraUvVa/kIwNSrR4Mr1+VT75TMCaJmEqajG3Hq+rAvf3dTMXiOrKWD
v9R4pGT1DPEi0vA5Ay0fGs6vqbo1EeApB/K3KPFUoIzb/SCy4kt1zvsPmJ4r8MVX
85EqSXGyGyvrw1DyZNg5aaSHiMLd5Evfi6+3Ix1q0wKvRr396D6JI2pNC1d4rFhf
FFQfvW+rOf+nr3WumDU5+qAhtu7yrOtug33ciSovvnBHSn1OC0ttMAllNI7Mv/MC
8y4y9DHrsxp7kYJCR6kEUndsx54itN1AXj5QSYg8OQxBHtocskfbRG7pd9r1CzB1
6yXaSoTxxot52MHlcZ4016b3GptirSJcADY0DzOsCMv07zz4z6K6zyAv8h1zI9Dv
N3PJ71poD+ejpkFrBDJeKnfppn36M4YR6wfHSygQndK0FtesYG+zPk4FoB7WQbCl
s98FhWmlY+BkpaHgVwk9d6/gq3jnR7uEf6WF/3EQ4sNXcUaLMmmhhmLRU2r78ZOl
Vdk2vGrwOZj9Oo9Vb9LO0lGkD6E8ImL09+T+inZh7FX9ER1v6p7dC5SXPZ3Vroai
PNugLmI6qPqAujuudwO82DFY+lcC/tLFZw0NxGPNN/P71L0DA1VObWhkrBQ1vy+U
Q/F0E7LGHFkCLiQi2WixR0M3LUVuud/nhHMV5EbPchMmKmyaCfS7jRL3DhYU0Ljj
2GUlyb39nvVjmIHU6cUiscUwtiXyVpjftQaZtu4J5cuUjLUkO98mWS3+HRPB2xa1
T6cTTS5FEyWJZvRHQQUrvK66CbTA547T4/0GzEh4op0eevWCdkYKqToEoXZa/mIj
Kg63D9dqeNhn+rwEE/E6onRN/STTycuDd4ateyITxJl0w4fwJg1R6AkwcWaF3DzQ
ZJdKU2lpPHJZ/ZwgdNLEjSXqypg2df5rOB2cu5Amtfa04FT3AL0NhBLqzfvGUnOj
8dVUHD46fON5c7Q242sGvWXytUP+mkDOr4HAEEvwevdmoC3ZI5TU2HFhCc42Apnx
ka9KfU1GMVj1DDTzPxHYWAXgYGzVERIzGxsk104pXoddwYre9r9o0ozZeHrOBtZr
QtrpqG6SlcQYAxcom1xCzlmFpasPFd/Cc5lTUJF6ko1+RE8QfrcNzBBL4996OCeu
q5+snnx+TkLcIXif6s9l+TpN0DR7GS1Uw1Sn6cblaCOY7J/SPG10rtInGiG9NEQ+
kA5yZBQFWBNJXWBwdE5JvQkX3Pj7gpI7IO6pvp7OaFLl7nhhabdG1ekE5VryaqnN
c+wwqa4hkNhBN39CKVKure1aqyzDGWKK0t/f/QBwYlj2O3VwvJav5oJQo6nRw1XH
/LNKMAK5ukC05C56PVap1oC39pfz3VqWO2NGWDtGnGuD3ASeyZHXPYQN6DH80NZG
Q+cvZDzccX5WnLUZ6l3oQioEeHUcOmL9CBp7ywHehzuHQbJt262oKY3H1ANsB4nL
Tra12ACZl4YdSwQVq47B1o4UZrY4VEtljCZgNyq/eAXA4rZL7KwWCmbCQWFhJSZR
m1OghK09cBQ+KyGbjAWDkUzvxh/rWavhGOpVvWyyfqEaa4PwfM0XsqmnzLWnCFLL
L8vDYbevw3CXgmwBA0r25Pt+7L0LmsKE4KLor4MaBx2lN1p9gw1tdOWjrS5Vu5QL
hk3bdjMP7/UhlYrg+8H6KCFHBj9dAINXGNt93p/ClBbN8L0YYb+1yCwNPJwYM9IR
XklgE6FKNKcjfmGh5x9zi32ObdKn5puTGuJAqmpBUoGb5w3I2e5Tafi0beKIP0EX
1tb1rqIEaOqHm3SmM/Nqm46fchbapobyNBXEp1EttbIKIrIKN56bWb6e6ae0J0sa
zVFjY/If+PO01nfaxlJWMjdK43clGPNOeudxSZeqlKyMWAmXySVD5bYT1pUBc+MB
py3pEnScKcsnYlaWHEP83kTWurNkaubGiA9QpBRZga+xDTlVsaATZTnCDasBe5aR
6vYrS2mRyupIn7gO+hPEAwZftXsNnypi2LjGiETKxAVGAm6BzfGGlJYwflYL7qWk
df9S2Zy7hvA/l+i57b/RhzYrVIqTTm4f0DHU5goW2PqqRrMP2qKGFt1dve/Ob+GB
uOVuVRUwmpC/77Yniq6D+WDCHBvexHpMUHWX9Vl55twH81luzoDbz5Vn+8tlCowy
W8Ki9S9XPJblqGMUTohvtFgdxmHIbnBYyBSZsXDOp3ThUtywxOFQXSAiQBRsVPy9
iub30sW996yW/78GSerHCCoqfsV/xxhbiOpwA0/xSwBL35GvE9L5Uc/rJAA9n+ma
NXv1dtqOOBjonD01iz+eH3dX8qAYSVxRzjKhXfJ6E3AXZhVNWJYQHXeHCW1z9RXN
08B5rQrxD+7qzzOYMf9fXaGXCvtCPsadYemJmy+pa/Bgq+/0p8Vy2cGzIUlfZ8A0
QRvVOE72Lvv8ydMY5lRjLxSHCYf0FIpzgBrX2vyfXC9FHM/6SC8u3xQCT30b0zwl
pPUBpvfp0JMzwuJqBjtZSq13353Ex9ykh6YixL11N10vElyGOii+j6yslZUA/16o
H0qVND1lJl7VHWzgLM+GBsPHZLxjg4DTvzxj28A4mQni9oFRIQiJVv920SC3anfI
hX1LtduRyGNRAXyO1HLEzH2yqcdXXpZRIiFg5ClMef+dNcHVQUts06UOPiR4WU/o
feDJ5V8EfAk0V2Av3icYVdexCwpz8u0Kcf82aB9zqPhItBR7kVrnLH6VWoSAy8bu
uWb6NHWDIMPAHiX6DckArhydhXmhsl2HSTkysOIROiJ4yrGKnYwEvD89GjT0bWmA
6zO6DfhwWMntapgGqp9WxGRDpHEPI7SsOG8FESRQt+wTwVbLPIBAXY7K4CToe5Zw
1QOZUBHuf6N3w3YXKM4RAdxcULfhfN3c+P4VYH5YFBBNqwGC0/LrNBJcXmQsQYQ+
Te4G9ntcAfUnYwniVJELUDoSfh9LNxCnGGXZv6AIWGEt4iLdxbm+1QIcOCSzxUkw
EnKADftYahqM4xodeSN6W5/GfDsu8dMGxGEocQaoL9AdoHot1nIDPKtuPdezng46
R+1YX1o6kAHRO6j6fAFVkHUi7AnejjjH+Usquf9nhiLnFeKSZBMfSrtTu+FN8IvX
E0FYkL7eSZG4VGWfzdztdvWufsFI8/H9RBzXpwnwIHIMb1NDSkAK55JPtk/ZWkLg
VePFaG4557v15bhO9kGIty88OBBL2Ys6KocpiPZhzTj1CKiQOuk1lFINTo5yBikN
ymjmwtQLBITF9HV3ck3EhwK4gxkTpHQjYMxbGQKUyrkPAWqJmeQU+jKhgqY6499g
Pxt3S5/v4McJSPN3HuphjSIvRKmg0lwo1/CAXS+PABF3pVRB9fPTtwGp3t3DWSZR
R9xfQ8RoGbujd7lVz7lrIVnC/Alo+UtCSeiCIT/jD7XUFktBmZXMah9vFzpwz3Vk
Omf0KdiI97W0up1GiNNdWpqjy9gCvyye3H3UT3dgzSAfFiXzpkFjZByEUpy25n8o
vlSfXROljs2UxYLbcwXfjz+AHM2DyZydrou9sy1N36ItctvCBHdGlgtnHQYKpAq/
uwRAvmc0AKfEkXM2A3koeeiHgwfILDy+NsHE/mVujfmonWQwm7RXBrAESXbJ+Ahb
Rhjuzo4a4EcdwQt+FNcwLiGic8i3OXP1COPQLCPFjadOOSblJuNfgQNu6HtGv8Lg
UTUzgF6z3iZDI4SEhl01m5M034SmmFbB9NPF3uwp2Qm8NyroSKnjqst5+6IWgO49
SENATyjQfCxNx45BISeHeHXIiT1uE091sYZFJ93309bx7iRd3+ViwUILNxJBSvv+
szDArUs7sz5iWIEVN64b112TySrRBoR4QUI95CoO9J6qp5BBZTqWSI+5rNRXQ2Bg
nRWEXTwdcgwiPcuc+j2hiEX4i4Y+ZP0ts+kffAr/2chgfBkUJntZaA/9GemLrT5U
J0alVzgSYLtXUjjacmpTLD/NBVt27/IyhcCzBcHNRv/ln0omOltQtCxeibX/t1qf
vQtpQo7fhlAz9H/5FhnSU5q1xxInDmokb0jNtoIeiY4zoFYU16b/mJL5eRKcdFTy
3OMCwhCsKDRujSdQkQfNXnPqacRd2KCB7X0oFaswbETOY0wEFtzzq5ksPeTjOWgG
XZtqTP68ueZN4LhpFTcLHyr+nsvSrINqvegEYAZ/6Z2gbSKPVnIS0J1hAcV2pods
TqlJbFgQR44/nCHIggMkSuCTQJ4SHqPjnjcxS1Tj9YFHTdJYGZxS0loAonV7MZx6
V18jNxsp4R8oHpvCqezvoaTTkkbZxMCJBSwq8iCtaqlg3Xp/P+vZgMFffaXJ/mnI
FWqipTjrFckEGjo7EW8fVNqM0JzrFmOqSFqGuc4T0Tj42x8V/07itC1LQW7HWGwC
Gz4hkImToAT0uJYOIyBZj5E6zKG+gH4ht3JQjEQ0OArt5mw6+muAVJGBVMapSkrd
rvUoMjFJG/xYkqni+lakBd+gYfW55AsKVP2A6HcGRDOgJwAM6IR6r3ZdDiM1wssi
C39lvJSpV3Gg3rPyTsDgkuaZffHQsqJS8Z2tStZx1XMChQKlTlUfMng68sQiTonE
zOkKRU1V5kJK94UgkmBpz3yRrAw2av7zpZOChpQvjbyGqaZfwPFBnzuC7FoZWgp8
U63GvhN8+sIc+YT0NFY49MviIzPI4pNDubJkol/sL36pl4Ymt7vJZ/uxTrKhXW7x
GSxwWapbL2oI6qxQIqqnlUx9Q4/LG4jmMhtRNkji1iuyoN+6WInqIUqKqso3NUHj
0Tf/9AQPU4EKN5XWPkBFqxOpehGti/Y9NDihHRVWDTqL+f7ykD4du0+lmSnRzNqC
2kCpxk0yxfkxb4OfasH14NqPqIiRdb/5w7wfAi9+VKsNvIoA4ujSMdNs3bYe6dS/
jkBVpbgIzgitF6fA1O/jYguuTqtEf1ObdH0fdXC/WBwYpro2xvGmAIkyGpvjEmUD
eQhzeLU/3D/65+igLMdx6+fQ1kStY+wbvF5FhJPdN5tItFU9MFbGpOqZxXR7oofv
A6Mp4jYo0Xvp1GNa8kYbWWljj1PAybFwSDjp66OK53ecwORdaHy/7DYRU7wFFTz8
n+tv57OpF/to4LIE+DCS6rbLq7K8v7Pe9K9nidBmLiHKMbVcf1BrmKEwGq4tF3fi
zUZDf+U23dySd9YFNTRNQNCGBL1K/JRg1+OqnvkPiogj0XtB6+fiieM2ZLc3kWMQ
HT1Qkfx/0Q4sE6EdL6ZukJpzYdivm98N8teYhRjjNBzHtJpPgHJe7vI9Ijqzxmez
FFvtrB9Sxpx7D0LQ4kWQkwFMBHeXsvmwn7PenuI5RbLRiYdza4rQDQjABtMF+Nnh
pKPgHymQUdtR2OcqSWHiWRBPuzr0io262E8pbZJHMvJzfYG9KjxBrZ1wCfkq8e3d
GHZOKodeSSpN6NyvLdUFGlz5TDw63t0TEFBz4T1u//NG8arMkqDpOYqYhilCVJYM
pKHofhqKIZ0fqDyZ6DexGPuHojlJFbSfFzAtc6F8o1SuvFH/V8xMskFWps5TOkBN
LfQDeLjgqjcbOb5NZMSFOFE4wsvfw/Y2Lg9nL7LCefSYQrt3cn8l8RXtQ0CRcOsD
y0GMrBQgFm1fqHCoAPRIKv5RqGH+eC2mZ4rFjcLn9UZKPAJhQT5bHxfPWPGgysZc
2UZegToDTXWNjwwKjk7+d8jvSAWZB3jrysASVwHJED8Ece0z9n89rGUwZZh2cL52
GbbH5K/fMniandpb8hVvGar0q4MR+bXj3PZlHgqtG09RDzkvVvkIq6npQ/VwJEZh
JCRYE6HPTuVdRH94qszzxThbcRjAceIikQnZp74/++HApH6YXOAWb/uzW+NuwpBk
vv9MAtMa3a1R0XQAxabbjjIJ8zm3cc+R5t2HriN8GYHi8g7o1xKdUyQx8oTdwMgH
npzShwl4E789l821J0J157iAUtVuKRHrilA/vnMa1dtWHgURO4tujSW9/Kbb2DwR
TrbXUcLXQnJGXU8e6fltCCsj1QmsHzcDVusMLzuh9lb2rjmlxWE9gwIAFZWFoQZG
MzfEFW7lxSDk6+AEXSzTJtkGaa4P4bRTM/srG/Op70gsPR1Q/0MPp5pqTn5o04qd
6+ghZR0EKmkiW+zumzfPQN71Fn7Yu4LEJTlE8HX7VcHTGB8/1PzVcdj+p6+UOCia
X6dspHjuaRRkZgaMtqBapHNHIzaWnkf695v/29GfR9WfjA9A96GYuybyZdxoAvqi
oLsPVeQGN5FukzxSi+pLKuclSH04hhCR9AMwrXX9iia4HpHMcRBJDbjlWCwfhkU/
vk7lli3WuBQ4zzjQYVjSORSiqO85pQHeQWkAlH0oZicDxWetWx0z4N1gJNSBJ9W3
75yaBTqHtjXHKKY1tHS08kh5EM3hsreFdohu9n1ri64hA/5i/5GmHUOqoaUTrxcb
R7hiBjdNl4wCVx4wEPpflPNKL4gJIIeWt1+Y58Q02wt4WCf9ATjSpVLACRFy4NWW
loHMzyju3hqDKWeyEOdKub9DKsY88DvFwLzK1SZEeV15oF+dDtWgPa1dODYIuiGk
gVscvr/w/RxRkpPWIHLLuYazwFTptiUzJNjmfC2Ivqz39B6gyyOkA9DPcIaPCTA1
lCraz/dgIIepYhVyGukUxbZ4m3a3sX9MffR77lC1cPbDw74K3Xf+jTpIZUnzriey
JmcuNohEZbhmaKTgm2bxiExTfURunD1uRvWeoONTQ0BZGj+iopVg66wQ85/SJ97G
zl1pXKt7/qetbpZubNfkMVRwlnS/XAYLpOT61aMRqfCAffbllafayg666zR+zq6W
5FHqQ0flIpwogiPNb1TKtfn8c0Av6Iw4fjkWOKJw/necHF7hJKYtDDOkz54tD+2P
dQg+YUfvcFwhcuEv9Dvl3Ysvoh/91WNK/riLEg2aoIrCg81fBSs+40cpMrBIaUXf
pSCbhRKn78N5FVe1ZCdMSbguJynz3eqK9LzSXpFhbZccIX+ZPEchKEP4KYkyjwI8
j9qeyCEgjVMdpoHOASPEah7k+TPikSqB8KwtT2J7Pum2S8Go/k+i5Fo30NAF2wMr
gqhcJAVtxfT2QxuwqfTyssAYZ33ETkAhqx1iK/PuWby1YCZ9AYEeI6LDhZT+qxRx
cQjsFigU2am+HH6LORFGKiQOcQWsQPx4z0XR0+Z/3Q4gAY/N1P0DQqSRreWfNJ7d
XThXUkb1HfsqGNzC/vEt0eTtSgUVQSZ7p/xmMl7ftWlNJUNBs35Kr1ggVQu7rF1p
4YXmxj2siqYXspT2XHU/6akvsCH5Sgzkgs8oJBPm2Z+WQuxhaeNwH7fXxM7c0TBu
8iCjQuO4feqMbHlgVdRZpCkGoPgk0hcs5u/jA6aXqC+/IWOm/yHtA8CX6ncZxUUg
0DCNsGG1cG3nvK5WEV2IDpKbO3vF7Es4fBCtc5gqm9ztYq7E0KObse0a7ezPaQSl
oIXOB2rASUqPFfhQYgPF6Fy3ugsyrd1JBc/sARMvucH1+EJrwSpMoX5nItAehx8R
6fwTK6D9FocGEUMfb4VcXXcBGV4oM09r7uCiTdS38MbhBIyrkziPM6MmN1DE+6ea
DIIk6guhwcgGKi6H3AMqQ4/3iSqY1XJxIX4cEn3VwuG+c6UKZKlycZDaAmAyNCeM
hPuAmxE7ZS8I/PFqlIdexY7i/XzTgE/jfz3HnV/FE7l7gV1VLma0COEw2OhKyww7
7dCA0mz++NtALoWawIt9VLx8jHTjpEMdjguupEDeSfx1vSknvRgoINJQHTOyH8kA
xlWlVFK0kEimOH0w4f1xI6rBCzT1IBiwdObfKo2Egh9VX4ZnA/pgubGLTZ4bkyPJ
JE3ywW1L/WtdHjNljhNWHJzapWjC2uUPpijmuT5mS0s/R1I+KhVLklB6zOJ9xRKD
RZ/mnBotZXMnft0kXMc/XcL0czM2lhyDYIdcxacXwxhi1SXeOLAUirH9b1h31aVX
5eHeClg+qAd9skCSD8z/9vxyrOP+tP1V5lD0PPaBOMWAxIa0WfTjZ2zeEnWtvA9z
r3c+5AT0ZUdhVAlJmCmixpTPTgzbFxQx57kwGqMkzOiT0qvLXf6hj+d4KnwotxZW
kzVb53eP8fDK7sX7n+poAMG/EAYOis9gNtw9wlvn8z6y9eHLkzxBPdF582FSsUtC
f6Um6x1TUYyrIfg21cH5Z7mwN5MZIOyH7v3zmLCWxrqzxYTUG+NNdqizC1qoCslo
mYmMOKxJ81kW3v36MCUiCt9lAq9xI7fJs4UAJrj8zlYPUTbMwAp74lOfal7U6bp+
CBmVM1zFCR8kjm1xt3FJWimN4RYlpA44A5u0YjpSE+R7NzvoOecse/zpcl0gn1NU
prGsFgbMtRLANGKS++qSTXOFtV/H8i0sOo8JRd6LaH7pkQ7KP7fhLsG+sGChgdW7
Hw1jhO4+y1YshWjpIBPA+zFoLkD1wm3NSbaRWAPQgzraCKUCvKL2EJ6wzu2mwTtz
ezuWmUEaN/dQnIl3fmb3DXqKcVjJQl+96HnDhW3L/B/QwQpPmehaIQ9xMOny7NBv
rsR0yWP5FqF2g88DNGJE2th8PHBdO0vVz3mMiWwWeyPB1hEG9xDans5rxKa2WEKs
1U4fckV+mjAsuLmECZ2Kn5KspP7/2WLN9QUMPLpFdnhV22U9tKVGm/msF3BmHJJn
o+pYtkqyCz28yHUDsyPAYRPAbkfQg3+FiRoiKBJMOLfO216U3U5ZsGRR51Lt+yzz
SgJOoh9cbKAcnZpqf8YhTtyTf7ERACu/6a9N9FYDvtfT9XtT6/ggfgips6baJYmp
32eIdKsanRhmGsdA6kYCbT34lup5RjagTRDwxZITwZIGpPUfeBxIH4MR2dq0/JTN
13n7EwK/L6yohx1VOv2WWbqT8hA0q9IlI7fVONzqG/Jg4jmp6+UVw/mZR/xLFuET
imoh1hWCfQ9yIrcMCtU7Lisj3cc/iKVQRL3VLmMqZTzOP5CSYWE8pMpQpFkqD5yO
wufErRwsyIGXZUduLukcSaPfE3YyWh7+wJfJuEK6u3notYChLMsCkuDuRT6GCKdf
SE2yXcT5063Ltjz5GW2hC9b0/O6rL92qBhUiVArGOxts9yJqXZswUAl7L+m/Jj0r
R456CEkHFU+mdf21Pe0pZjx988/UMAx+lm2fxIDBPsmuxUyXzfnIPDSUa9WXci3e
rBW3hPoIOIRJRchccHI14GruRru3+VqkASAWX82TfEnfg8j9ZMy1qMjEDem8xh6O
P/rhH5NRVRxzimNZsBmWa6B89U2yQ9qhUfIDWBGU1E2BzjeJZsbTBlibGTKMvqsl
KyqU+niQXCkhO1rkb9Lb4IiSmcVKrVQN2IhWREdEgQNiXRjaRnrY2aUEKU6XrflS
sInlHYRM3uNQNKR64VqmohhQpTOzjukWdCKrGBjXwsTno95lpbeT+g9NPOQQGS+Q
pRyL0vHTBfWhpDyllAKMUl2JS74K9/gO4MN8LUfu+0aa9Ibyi+kTeWCXo9GpXo08
Pg/1v6mEeLYB3zr7puNltU9jPVR+vnFhNfkFN+yE3kxxc+SN26MWFFM+3AUMz4TW
J6bKTXpjI307l9mQeNl8j0rLLBnv34ZpVeonGszRZv/wgJAHctUYOROh5TfqPQPB
aQpqjvryc3dlgQdU5XCUsHL2HD57+59jTQN8yiPad/TMjd/d92Id03Pm/e/l3Eib
Smm0yScUTHDxM0a2j2dT4llHrsfk+JsdAFiva4vO68blF0JZVDHV2GAD7kYxP/lh
ITG+2biY65I+Q9aA7iiBFzNSKdaXNZlIXSfI8YutZ852cLlO3nzXrnPOq5mkFnkr
FjusGA9v64obT/IHPfJXW96e7zwkHGnzG8hqbqHdLhAjf2i+ejQtixaDel5TyXqS
aa/OM4b5X0nUJHiGi+LvfIAxxJjfobvWYf9NES4XHXQ53hDSSnQWoW6ZetCnRYyc
o6AE5UyxZ/MgO0dix2VRfw7Bz18YUl/o8FKbRnUGUbZonug5Q9OZzXbpMc0DRRjF
wOmVmPsWhuf/tSkxiVqZspq65tAk/N4AFV65aDqKP+hus/Q9ia4r2y31q1OKppGR
G2soYiNYpzJVBq39qFb2CtN+hVzx7H12x4M9YK08WX9CdvIoVqTAat+wc88GPPxl
f0q9T/VjQVkvi3TdNETTA0KdJ9z0Q4mK5ekn6uojTSrl65lanlmjUtZiCOk605g7
iSfNuCOvFqZ36+q6H1YL07l3LLuIUxwB3s3Wq7TD5kdgU6KwlJpUEGfmZ9RxzUKR
s+vEMN+lE8PexCiCyrKerpkd8h542mzvTZvrBwNywFM0zuygmjfLRFwAWUYhuZ7k
3fCYP2gFLrojdGbBi0v4O1VJT22TmelLHnV8mmnVXF5xSipNSCeFuSti0Wd5V2rN
LmqQlhiqJZCs4jDtzwtAC8TUCOjSk3kUpsjtkEBbtcytQg04vmw6k4dg1V920KYf
O/LT6YLMSnsNcNswQOn/diRzohvF/Du2pMpDOFUO0jayizgSr+WmAENUvJ8cJKwZ
c4FIz1PkU6q/bKPMb/4V38NWszgKrW/RzJvxd4uqupfiehzaSmO9vsn3jTCbTCgf
XKpcGeQnuuTUj6gzKQ8VHohEOolp2oez9NzOzo+RVyDvCu2pUnWsjWGdV38pSVZc
NU7nhq07/GaeBKjXG9R7F0RHj1uPjQtezLcS89GA7ExLNb/h383kQ2sKfXXK3g4c
Zt4Yn9nXGzsgIOn+yKHGxZAdITnagmNWe+4oD8zpqchvb4/ckE13Mx1DwzKZa5Qe
IlU9sqG7sa6FdQ0g2al+57ayJd5X6sY5YtMeCKH4VXu+7ZyprgOt9I9f33Qd2jrU
Y9tMfHxCGR0xmLeDWgpu0Z6FujWd+/NDZWgSHc+VLPqKzXjFrbJdKXLl3GthSpQZ
Nx/UxS88K1TStuzcJaw2akRxocSLqPSBzLP1aD1a4ZG9tNRzt5q18apd8TDIsbHW
amACOeL3bTVyTWFhlUH928Wz8Nkr1eoam9qBthe7JXfdPY0OMFbSrdEy5brn6Lza
QxPu0N95GYihFDm2Yg6xuu1YoOAL1cUJuh6P5yvWkUDXA5LadS4IrDP9hhkle9Bk
hInOxgyd5ISzX4WEYO4ICb/rwJDv5YGZAV7eKu/hjfbMlWIPH5FRvZOTIlIvgA4t
VEMDZBJ647wV9Bn9ch48kTZWafd91YAuc2BzW+/7rxAXqmNeSHEkuUPn8SQwoGHk
ylLf6VbGZlvBO0mJoqmGxefMXDthigs920K4p9mJ5ozB8dRKmltMbbadXh9B3GEj
8XentAuikbpC4Fjl8eeM+Oi+QZZBKjZ8bZG09ZvvNSjC6umNLuBuKn6OfquTlz6L
X6Zc3qNORp61+5OTGmJbMkubKom+gy96r4IKNR46LGDWN2YkUx9YXRzHtO4hk5Yw
N0mkDHZouvQ3JfCmJ3YLTIJPxc0BO8esw8QYnrNmndUMxta/8IE3kax2zv+4mt4h
g1KnSo67Wr4aSu55yCM/Vo0RICWv87OhAmpBO6tMPNSfYR/4yjUHKsWReUR4tevq
g7fbgT+gOCSEnz5Wzw9te39+5OLkVcx9NPJNrzLshSnXHydKXsO0t7ElXVmeVD+9
icKkeDQpxI02Cai7tpApVgxdfoEfK7afW2BJeeoBQSYrUI07KmTfy01jZBQhY50G
AJ6eFEJbFgYT6r8YjJgH97yIH7nm22Fy/ACk3vkDg9Z2DCt/kirN6bp+kjzxMe3Z
uTV/QZvSpjmLS6poPTROOwHeF5lKYVYgvxkT5/WW1nW8gGOMGnUw7U2N/SXCbvp0
+rSSfBpEceysgK4RIKm8Mgg3JNEMGxL/T+e1pNh1PhZOrAcqhVE6bcE3DZZ87w7O
lEHHCjR4XwhVb7Hz6tQcLeTKKP2uY2wWyvvVYxIL1I47MIYVX/PnNlwAx352OPH0
cM6ymlmltJRmDRU/i2TwO7olN64rTTU5b4LHahcpMeFNEG4RbCiAYZY8pgLX/rvT
g0U7RKdVaSsoHQY0iY2y5WVjlvCTwXhx38M2/tRMoC9VGt3/Lj+xLZC7dkP6zrbY
sunYGgnMaA45UH1eDBd+G1NvQ6EqIVeZhOY9L3g+tsJ3U2omvXbPzs938oil9nm3
M7H1gbBaboby/SjhaMAHaG7D9pZvLdPoMNl9Hp4ELGC/X9NqpCbphGnVaCRVnvuy
7Kxdn61DVDazuYeS8+hlX8LMkHr9XqVd0dLybZrGCzZ3psFl27cpvwUxAcaJntU1
id6LzWItfty+ZcxBkRK5KwilRPDptzbegyJXx6pIafxwWMp9Cvy6EPowFS4lk9F9
7oR65vJE8N+1l5XPVDy4nq9B0UFW9mBprRMuq1IYWhuZ0j+aGNH3CDeVtlO3YTDG
Ue68MqrdYkARWT4aYqV4etGYerNgjDK8twn8PPPaIm61YgGdoe8Y7/FSp/liaCEP
5Xc5Ag7zzSktaUSjUp/pZAfR+SKKktRFsq3a7kA/skmat2OFailEXwPX5FGTfw9h
fBzpRWq4gV3yIy8joVS79domcNlgnN2QisYpDMAuCdeTtDf5gUkvbKcSXqKfnFeF
vGwNv5p3whF3qpCMnYJiXNHUiYzPL9b1/8bPlSK3vZf7lARiUgRWdaAyrHrDXffP
wILJqW6uaO49asP+ZeLeK5ue/YKGKXUkKAQeh1aKhUEHyZhKcHuv/XsLfQlATaSi
uHnY6FlQFm31bLCKY/Fs8orUaP+2h9Vh8Hfa/7qlFAUB3Hvg7JWwbnohADoNjoNW
RumIQn26ooT7wVPxPL4KD1jYeJHa43ZkoRJQS4n/skRZRP4DqIn9k7HPaoJ4/bte
q4woHZVkZe7lTfjHkttwhB2JzanlZzXVQVwVtLZGVq9/EATv6Fkpp0KQHJ7mPnso
xhEkWfB/wr8ZmkqyDn/0es/JX7i5iUFFnKwT+yhEsz1pQSUQ/EuAaMrOxyUqwqib
xgtngDwoe2NUbXxew0f8B9O3MaUcKXIOgDXKrthjOoulQdvujmiqUXGTdp0tzp3g
9WdhEmtu+K/coqoSWHCNes0GFFsTWTNehHmSjoFAMEIYzxVFyoiPdrwNUi/jURuU
ZilQGCRj6bU4FnDl46FpD5ranhE4knnGJQIpmYWM7Yz/3jjpgnTAt9XpEWp5S2SG
9+XrbmHP1iJ/jqHsmS7rddCY7QfZ89Qt5789UsvxBWiwKvBQp59U8zGAFRLApBYp
3aWt0T0ScM2AQnftQPtSwX9GaE5Mu/huNT1242yIlmf2MrHO3ny7wtobPRalwQtu
alciwrZge5JdQKzKfdld22kiF0LRQo3qp2S1dbPDRK4GfW8pQ26DVzileLexbyQS
FYZf3PAc5Z2aG+fAGxY7TZBuLQ6YZMbam+iTU1+ixFvzvQxlI82Yfbv0FaIgO0TK
72UyTVhbj8lTh4FMTq8+PnIqQFJgv88XUpVsE8vBrWvVDfrvjTijdHyVOta3vyyo
o0L3kiJ6+8g5Ej6FIVnplvMyDxntams0/TTe+Xs1DJnSySp/GP2YGB8c+9uayRs7
wB9XIwPz2j7mRprJeS+WNx+V9TKHkea2PRKiXgKMdZYtqRKadOMuQzHuV7U2SrbY
x+fMHWL/V/kViO6cMUG3BXClD7Ce5m4YKwTgAApSSZ/V6rKS0ZVHRBLUm4MaAYAo
+NwwOZpkQ/xM+35ZCkD/Pvz8mepPbqbNna0bMQ66O78CvnJo6UdXSQSDEfEw+H/W
NqzcNS0tYnAwapEYWy+QXM3XOJViQG6RHxf8pad/TcF06/N1tMKxoN3U3TgcPCpU
PSdLUgBJ+szkqLlllivC4FbeisBym3Ajm6lWIZt6UF2npJZiw/Yg7jdroqBFHRPj
5VtVREzowQvNrQaBSmj0OBX2sMXVwv7auvr4DwiA629AYlEwPeBHrz7a9XCzuZQu
K1hDm/chzSCC9iaAtxT4Xxdp9CtxssixJBXctYAlWTOaZSAvd6vZ8VaAH6gtvcJq
8IVj5FyWXWGUVwUM4MS1Kr1wlFpWZSpu+PoAs5DaDz17At2BDU3T3N/FCIqM+3+B
6nYk6i65HTVW9gkaa9Sn5RgyU0wpxNao76pb2pxsSwTs9KNpyHz1z5DqwzWW0MS8
pRd+ilHRBr7rcqLG34MNMhf3NFdqxkXxBLwXea4Lqf4/2nx3qTtCY/y61oASMgsT
KIAmxaQ467X9gpfPM7ckoR+zgnoyZ1n0NuQkAFTcKeMfOO5BYSZgL4j/9LuwnP3c
RuUrO61fOEji3nbYn3MdW6rJ4AmeGJA6L06Rsh9MvyDo4bfRr6mZS54dT2q5CNt+
/91W9cRkgpTo8HgN6Ot01GV1itYJc0fdOzqGGyZz01Z8qfRlhxke1sWe9fHMt+wq
C32mnNshKdmeZ62OX7jImCfbT/ll+j4P+Kc2wPYSmfRwTPki8AfrWsZbScAaOz2R
Em3drRLdYHj0lTgO/9hN8Qt3tLrQSbwIkI1/vUiGUIS/Lb9MoCBZgAOC5/9xxSjE
BmzlQpRZnX05HegOqKOYCpnt4yh+sM45Gzx3Z0cco8ge7a6HLToLCTFFzBCD+2D1
P1GFgXBASwMS5uHH/7/Ax92q0jYf0EAvOdJz3/SOn06hEwRCxtKBoPD9sDrH+8R6
7oDwlHI+1QjosnbyNCtSzpy8cJmnaiszGO4qfjEEMn5jRao24Ri1V/mgt+tLlp4r
3gLGrYbbfjxqIBgBsxWCJC3rnveqtd46tLEspsO1CeIuv+nLrOxAhNHG8fesl7ah
qEb/l+mNWecAd119VTxPcFGCskqh4EaKwRrifOzoHECGmChRkS5AzM24TyuJgoXr
An+lzQDPAo8X0CCY7pftGbUE2CRDYlGFvnNr5B/ZinGDsjdz5RKLsHjCzBceRCdu
bD0hmGYzLfykM7e3Z6ni2IvlgcshBIGQjtFfF+djh8EOKkz5svfPhzjlc255ecAg
y98Tsromtyw+Q72phOOFpEJz0WJO9iS7jTGtW2KzjvAEhdXmJYrMIvb7wpjILjzx
YJKFo2EZgPBC4tByeW0NA8I6FONg6WpXZ6mAWvChNCRAPL56d94Dpi9o3Ro9o1ro
V1eTssNIjjI/cTwWqCc1zsSD/Mzzr6svDm6KwF/5z5v6SOTx1qx/zdFYpZaa0jQI
jT2nG5xAyPBNkgPhxgbXauM+jhasx36HEAlpZa7BnbqwZ3DcLVzFn8gslRXnjVuU
Gh9Hzjfjc6eUO9whfJvVqUyNypl3t93o0eQl1Ao7pCfDe8WScofkvqFTGdZPkonB
GH8sOYzuK0bfAOmJ/evSUJV4Qm2WrXQ3nNtTod/KcQLu0X5DmJN7RCqSTY2ysq1b
0tQLniFwfqiaWrT24CLChHfQ/hJObtt2k3PyKG3ESYDdoCzOKqNSpmCLjaoNdcTX
5IpoxiXuYBHiGorKKa3REBaNyJuehuQMqt+AnewzAHpefoZRkJ1v9roS4Hlww56V
+N8Y8mdhgRaB4qhQlhPndHPKXWg8BzD7V9mEXWlLH+evzN5p54ozSrvbx3M9syuz
k48JnN6UWyjNg/igR/LKRBVES/XLXHdGV/YQdMHtwEeZAPzThTtJbD15IW086t9g
Hc1oByTHRJzD1N8DGbO7tVSnTdNnoAl137yJIbKDVEuGGn36QEisboipOD88hpqo
bO6Gyhwj1trVuHldIfMDq6I1ZY6uOuJQYUDN0tscSmj3h/MtQvddXX6+AjB2tSlQ
QHmlLeitpQvB89B0IID6HNURglJ+tXPjFZTILklOdWieO+qtLiV9354utGDjrrK4
ML1dUC5pfjawyZsB/n8WbQ/XWqQ4uYTMrLBaF6hN2lKoIyXR099CdwrW0FR4Lg2v
DM23QqI8Rld9TzaRS8fnop5HyuFJUepoONO3Wa9rP8fWFEr3gH8CddOU+F+oNPCI
3/txxFtxu0Ai8ueHZIWow1gHJlBNKju3YCpZex/d+6NdFOmAnGCpPYd5xRCcYz2b
5o10LOs4qDJdw8m9YVibnmDen4/cDJpfV6i2GnCpCos6WUVQtyt2sy2QiekKQlJh
6N7r/fKi/x2sN+8z9+FfZxpSoQrpE2M66bfmKtHqPxqPgxT9RoALB2CzLhLeayPj
yXA1xC/urSS9Ea/sOzSk1d9Zf1gIuGsl/JIuhhdRaS/xnLKFgV5+qErcot+WHRCO
9lOibvXwPSteSar3eBg8Nfe3/6OfUWpgVy9yxmtCmY2jGk/fsetJZJzdjaEtqqhK
14qZ3SgBLEjnY98zFfgjrfiE/gtvQMMPI8Qjod9DUgkpVTRD1U6SgT9LNiViAq/j
NQ1bE5xQWL8mgRwK8ua/rsj4nrSsN3FMIcmzF4YQHX5KIbCVKC/K5va9jTAtKnc6
rXShR3jJMrqusRSpcDvx+n7qXkYPyXhUOWWjpaKifGdiw+RWAet5j+hO7G/Fghkf
TDdGmyvduTqKBDpTeGcJFKWtgW3e3VZ4r3hppY1JOzncCP0Bu3gyUnapP3CVEFCB
byE7WjFvTDstFTY3VhHrd8KjR8H1sPjdH55uSqb6Tz7vYReIzZAC1QGZu70+hAoY
v9x0cZEye6VL3o0166uPxc8r056NI2hx9jy6B7tZ0g1oXx+ssh1hWxJf7Lcle3Xw
IuTK60TmTIxbXrcSH3bqarPXfCvwwFUTVwmGlcG/g3LGWd/OckTlW+Ac9ZAgHNGO
WXKWwaw7LyhQRSKfsHF/4DnScz7uqf36Ixosy6Tnd4Xm2djMwSMYQrqBuq+rgnf0
UfyzhmuOT9bX40mUnltX7J6s4bCIDbH7Mms/mB18CFBZ01v50cpdxAEmS8eNJOYs
v81R1ug1fy1syXJGLgrVC4ENN+NQJqpqzxYRn2OlSF2ByvoS49wfFNh6OWXbULIp
WJrIr8dHC2repZYW+YNPkW3wwvLapclr0t8wtNSeGThAjhvAD2+R3atO6iCnMgbF
Ozap6El3XTWdtfjzK/dQV3QM5PZQfy2z1kbfazSqbDCQmHRwDC8NIfFRyV802BnT
GURgjv5L3jVeNaaKhQJRyIjyZnfhAjaPfqUomZWT8oJpJZ9xpQC0pvNTPz5UsyO0
3W0t/U2HevTMuGu/JShvSStq/HvAaHRZtVzl8OAJ2dX7/cEqlrJqsTjaDt3oETZg
ngYy/ND05MZoVkPkhgJYrLttiP8TpoT3USdSYQCB58C5aPdh7GJuJfoGrNqwb0A5
xKLvZOfEwfGs1OkPXOj9xzQ+ZV3xA3QGh7suQCI5uBvmh9vKTUm1rY4hEWGhQKLr
QpS3JRrHQIHHKWvbQXfShC/Gkz9y8dWqA3mEzTpSfJdFLX9Iyh1FGr7+uGn+lFvU
eqI76Z/oKd1tcNMo/YL0h1cXcrOrSG3p5WNPlrFmT4/+nPxkEzSdzOA6irJyAprq
AB4Y84Cv0JOlYAK0UCmt82hl0boc1oNBp7rK4VbJEDCEbIusudwAEsJYtBsmKBho
xFArT8k6choOnNzGCQqIIiiPcYwhAba1NPI9M71zZJizxT65ID4ZnzTc5aNR28vw
f8bYiKbGxTPUzwDDRGpOCyq3IwVG2epKbDvaU1ay3ODFdwMaipFcP1rBi0W6HewA
yU7U0pwSK8kQVKn5QlOyWSkkPxZVAHY4Ta7AH723R/q+T8iSHngAtwzKodnM8eEu
KCV3kwvrZ/9i5o7tPQ+FQnFmNJisZgUwkx48JRtH8t4v8yeir7qCKk8PhCvJ8qtS
3IiXonXkY+ZJZYpJNBFS0/ChIY7LM+43j4W3T9n9psUPPAZ0rZ+qK0TioAZEA/WQ
c9K6uUR2qj43uqEFd9+uR95iB22n6igfEHuSMAbMPqEfhTVefdFHXLGniwuIaXUl
iZW0Br+KHu32VgloWzDjCJcpC63rCD3hzcwMSteSkYFE5HDfl7zgnq1wbyh586ia
sWTk/rKHbRgsK5NpZmJYx2dX9JwO/5wgxnqVhKayGdkTbhlMGocxJTFpT5ec2wtA
H7zN2WLn8AZ65nTSkYx83ou7f+HXlzdHYeoHXknnHl6076ydBih+r55Icugv5f+F
Ki5x8zBH4OqmUfsQKCvzU0t80vnIRWHWkwXx1EbP2QemN4XZIGiyPPaJZ7Ulwb6g
SWCPoHuWz62d4xIDPmV8wOK6Hj79AkN/ZtbGenH8PBg6gbcpuKPQnuUwp4I0ImF6
d9W8nqpGZrwN0D+2Uk2OoJZxRy1gdHMYSOiiG6kcy0lNqEsjZMsfJPvL/kj/sDp6
EAwgX9Jqc41SMSKoWj6G3+Lud501DzgUZIukK7ghKRIG73l6i/NCFZyXuLpVIYRK
PylzXZQ1SY43nF2bPwG9cu/9Fo+BRJ4mBqU6p0+InjsC+e/gm9V5j8mlFCdUzoiI
IWaRHfRtrIxzpG9QvI63OYQ/HycFSrKI6ytr5lug4ZiD2U8mvSC3JRm8RirL7lxX
/BLOuthYzgjR5ObPTMIYAABvvgYJrISz2ZisMOWmIv04JfxlKmXizKLfhz+hNcIj
tf8weg3+foYYduo/NCVKg0842wa0OrXx38oYW2oXHPb+xsnWuEalId2CguOy9yqD
bzYbuwh88rcrs0jH0RNoi3xX4C+rmfuk8G/uNbMzxXuW0dewRBz2Ks73n/HkW+3c
8W2GbB/fh1S7CEogHkHOr2fd4mxHWTXN0pj89hANkpr+HRtt2USWjDtQ0gR/tn9+
lIeS4LgDTQgU6GZEO5LM7iTGCCSMtAWKmcd+nBMARdT7p7SoB1LxepmpEOEk12vK
e0BVSui/5C+15kjmWb922QAR6qM1gYxZ+Y52GliCdOEz/oaVjNyZIC48YJVAq3Rq
z4x8prk6QKfLou4wPvvrN13y1tsrzmEO+HhWa+2+EZMX1keqybFYDhdndU5ZthOK
S4XZfRKLFY8OCnGdz8QI0P2DObXijvbpy7snF8KP+KG/bdkEMZuYbX3kXupnj6WJ
xWSSw5SX0cudqKZczUfUEtiFbEsUZ85sw49+snerDVUUSpvboRgyoyW+eEo5TlFZ
G110jAMkSk+8A/TfmfXDMsqIHf4NeLqrrP9DCx17sVnpl9/JSfm2DuczJMvJOMzm
MpwewpMaTa0uiM1EbbcIUSLNTIfz8bfvTF9qxSPxUaJMXe/MJFpjRUHsVcj+mRbH
zKW7ZswQuGPQiL3QOWMgNh5Q6g5XveGfBIw+yTEHRgwtuaGzDWxJcA4MbJTBFeOT
TZrZ3chfCYpG1ZvMuvi/JPW2POR4gZGlbCbYr94L29E7tb2qIX1fdh4G9C9jSYpV
G4oA55gRJFWgvsPKjwiazaRCkgpsSLOd02Lhf2mxexC2hyLNqhT5vgjg4q9JMDT0
Z9cXKKBdtOHylPmkMUBRJNpaFK7hCLd3phAWjHyPFkC66vu8jeBpeBV/rddLwCMb
A2Z4ywJSMKwpCw2Cj3aoh+dZ95IPIG1/Rf89bmpsYSNgWmTLMsSEQlCy972uG11D
e8GaXY0lwQDtHSDAqvml1M2h35HQXbi5gsCAiB+6VuO5P/Z7MBZ8EyEawp7TJTLc
485kQrkuqxRl3RNOyxkKzcyZjUAFJnBQ7NCr57CrcUBJoC316YmemjuGBjkrgqiW
2P8c7VZ7wT1XAPJP7e1bZjCPDPHYtJf9RaPoB+ZqMpojAZXVL0AaY4v49tHF1dTk
+H21OvoEBmSe8tGAHJL+d/F366rhAGcnR2LrDmg1KE5xWXHXrsoik/nMmNPXG+Xv
DstGVeuXXEmOwM/vgRSFF8TG96vWkWNN+jzjNzEwWhVZW44WcHvdZenMGAynPEOU
uAAxEHpo3l3C3ZqqlgE/enVgrcAuJIxcWhjxRGKhP6X7GpzN/Ft3uD9D5BCeMhR3
pnitM9lUszEMDKsNmglKvZ232o/VqBdMS8Y4G+PKn8vJ34JZZZWmhdi9wXqE1Mhz
D3/35Syl927/X+sQzVjkYI4mfUsS3CZOQl+2A4ThPL4ZRZpHQ7Vzu2kzG2W6EdDd
hR+fURuRJUZ7i0q2EByPC5buVVyF5cCdXc5RaOsM4/r4xUrk/ISNSuyfw1jpx+yq
ycBx+lVJu3kJ0me65LaFcTVslRs9oId4ZNYbEY6ChsrVJVgUVNFGjrjo6Q6yvQjU
b4pbhd0e2d871/vuP2pLVB7VsVjjjrBPUeSHFUhAi9/WhXxQNAgFNKtwLeGlLbuZ
55eGTfMzx9w28Gf9n0jcY/UDLfWCs2/CGnZAlnN8Q1o7xdpXWeH8DZTxbeW5VUR6
pXEf/5V/ru6Rfx98HpAAQ8leL5bxUvK0yhhmmtmaGUk=
`pragma protect end_protected
