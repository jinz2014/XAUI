// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PaeoAg23in0DJmnSoPH4K8ZTHmb8bqiqza3+eILTPViYvPkxjOsBXRPAjghBQ0dK
54a6K0EISAxoERJuI5hCJPRi68qzhnrHBGu0x8YUiU9f2ibWkyxflAfXm/HkWJgz
MI9gbnIKDadb6C60Zwo4L6ZQrpDB+dZKjJIiq1pf2G8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6464)
q+mayU58LidJCi/cCFXptfsUi8T107PJfE/cVLcznDbc5MUAco+U6cLVUyJdvunw
I/WCX/B3JhcWkb25BjGvz6mFBZvz4ylp8D0qohRsDqieua/xxw/ImcALpSuAlRsK
tvAWU/gImZPsCdddRZvDP4DiF5nqutYxRJ5a3JVozZLTYU7pbMjRBogYu0+MP1ax
vdyr0B/qGn+Kz+VtN5lS3porPOyz57FUTF4iGWC+CR4+RMpEYictv0sqMi0YjHgp
tylLbfNlfuWlWtf8TedbMyyKkkBC7ixXKzjDKL2lVxoc9kwrOm/rIoU7FzXS2vmj
ZGkVkRB17zIHd2+agMkz7xKp1jEqYWd3sHuX1i0IyLRkSwV8uv+6EnFS9R1ctWfO
R7E2+CEEkplknoIVTn8RoErgMGFOFcBnibPjHVvyu35phKG1Hy+wyqI4DOTljLUu
I+PEJ9cuge5ESpb+FvUzC4t9Vb9FdVkiyYOJ41kE+FK3BkDYScoykPZnBpsqBRrm
07YGctZAdklwWkSU6ImoXcYj9g84YCLoLX6rdT/KM+Wcrre1w0dui6P4Gsxacvk/
Xym4Be/qSGR/bOSccDmdBQdaxmuqMI/XIPEnynkBfFixpqx4xsAhT+ZcuuD/4BeZ
xGAX2Um1jXFp+nGq5qSjUbwnkld1pQrqmkanNL/d7z6/6WcXXoOUSGKCDjP98hvg
GnZs+Fp08EPA0z+3+lNBPfM1fMj1G8vtOuysfP2SYBiv7evUsmrTEqfszoS+S06p
nMS22ysKSqMiSUcrnylsEeXiw1oNIfID/dCIQrRNqmYtoSNqG/rxbkzOSluj61eC
7hpMfSWasXroegULmor0PFvWnHHCrxZ9xU1setRrGyFwweVgWVNs2gxLlTi/mGp0
fxRazq4hyD/zIq7hBPX33Bm9zVVxYRCrTUHu8ZLpWbip+IxYLb8KS/r+uQb5RYId
/81FLVOHmkt4lrm1O/h8bgVkMCxQgpW8DkIFRWFoPXE7tSv4z4+Vskqcm3Cm8TYQ
WqiXc937dJQu8URtZII2F8xeIqFTtf86G/KZb9KO8cnJA7We0fKdi57uLeEBlarM
hWtV/zsb9je08akJRJqKEfeIWejCaZFtSvfKAWcIpHkGbkg0qFIx6UiZqasUN6JV
KCaNcV/5E+o/j6wT9kiqxpyab8DHSU0Ph1QLjC6RTluJp0md2MmjoM2X4yTfMj3T
ad3Sex4KZuJmbGEMKZsrOk2E5EyCZHl7EhICVM3JrLVx89nPS50vMoMJ4B00lUTU
Sq6qtWjSy0jAUEu2gh+7iWwJKAY9vw0AX+k+NCiU263rHUkqsgTomRDWxF/juPlQ
nPFJ306qE7pyBPyUwJVqQaCsj57YCwrspBeZztxbVi47N3UPhO54e4owc0CufKaI
oMmFjHUxRqiockAPKROhClTdVns1kVCDDXmi4ndYSezOW6i5wvaX6p65es4UcOIV
6uy4P1YqrzW17NSgYxVbCBhKB3Evzau/gPYcY30QOvf0V17HZZP/THA+nN8+4GPI
4j5fgOyVAfa+WApAo2LLfbVuwn7PAsMAW+dW0f5W5wILFBMqeJTzE0p+0MjyRrnZ
oJiv2JnKcrtbfgZxkMjwzyTdIprldhyqjn7wQMDXYQLxzgNipvYn9uGX9pgvbNPy
WAxi/gj6V2WH3i9VAJ4rTMuAwdPaM3/A8BxcOUEPjMzdbZOzrxJ+rvWFrFYnj7/f
znDOmZPXUjCVWHUekz/RjUSg03t+WoVquJ0YgffcJ+SmVVp+qmzomX6WdyF+EMB0
XB4y2XdZrD69wxE8VZEZc6KdrqGI25/vD0d1sKNdFOBpDDEbTwpFJ925lvBDr1aS
0+b+ukuhr7daz4nQraPpLc+3fcT2FAETNNdSXKS1yVcOj68g2EwqZlx6YyQAhINA
rruxWf++C/xGw6HsnrOZESNryt2zD5uHOjbEn2W8iKKswGIskyG7KgMkM8YFEmfb
5MAb+tXT1AaYH2W1ttF3IB8PjtsybQwlHGCPpW4mXN3MVXUChQTF8EGaa7lVOgAI
mBcksBgrBPT99mNICchchxoLQyIMeo+BrrEBW0LlIJ0mnRbiPHCq/J/vDGJQ7cMr
pw9xvCL0G8syPeT8vFv1/DxLyfEaC2TwEgLzxDIMGxLYJXxme2BBtTZi+aVGLNgs
TL2sC5g+uAsa4Osq60M0Xb55faauFKZ+0lg8XwD2wn856f7MO4pPtj72ycsy0zld
qTvYyEdFZnUCYtj3Nb/IWv1WkxDyKCrQfxtdEZ2PypEvqJk1molIugBWXiBgY7+0
chHkOE/WHJqAZTpHz/RUoSYiy0KmjIURdWtQJqmuz/YvaLQrZIUQndwOgVUsgC4r
ZQljjG+S0R8ychqDHHvtZFjlPoJViVw0KV1icdexIiSe/6jD/1EkSGHDfwgPh6T8
bmaMPC+i8FxqYiZ0uvMB+0pALkjUWdMEYR8m34XY94cW2LTM/DyHvPHSSlGkhzDH
uGNHts2+gWeVfNQYc6VmcttnPJ68nnSGypONIukCYuLWRU/fm4KMucODmVkHy2j5
fdxmjjD9i/awdugyFtHhTtgokt1mkvFa75+nrgRm9GYygUityu3zD9TfJ6QCqIFf
4wWn58q25pRk7HaLnjWEbgFvabd54xkDHpshXfvnsN5gPe2+J8fJ8r34l5OjCwbZ
ijRDlsBrJ7edmV59ybfY95836SpF5s83mbW1RQarpuT+InVkeGV08GXNaocasYRp
miEhVmQ3Q6QamDDvvcdgdKFyMQ+WiN8NIkv1J+Nnd2b97bFHiD5YvRx4m/MGnGSv
tRzQazsJ7YkSQb2aKawBYO8vApMIjb4tUYczUlYa8dokx+t1iy+/NX9JbHbgxUYg
fIxObgE5/S3d7HV2KDqwGLHXb16nskS/3GCe8d2cPw+UJeLJKZrKtGlZ0ldPZ5ub
fNr5fGvzxyRWuISaDOeB9iAE+nJKeeSZXuiuAAi+fzL0DKQcC20RIYPtuLttscXL
cNWltLsXRqRkjKfOJtfe3ap0Vdy2C73TaTY+HiqJ53HPd73TXssWoPkGb4xCei0Y
LitYRYgg8GtJ4iqlXUHHq5ZFVZV+rVo0r+9zyblvjl5TLvKTUbF6vYERxmPxDkNr
R66kSmIyhvmteejgJefsZadpKV5tbXnIeo5KyfnmyjW3h1V7Jgp9TNUuYp9vaWSi
ipLrVMPnbdev/Zx/ZIjd4s6usk1Q9zeSro4ZvSgmg1SxQr4YToETXtgCcYz/tLgs
798DwvwoiLyvVT6pwN3JK77+Qzax7UUErnH7QLxWGO7Qeiuhfj1+uvvzKQ1JYmuw
AdasZ+ypon7TSIB+01g2ha4JsWd7GxGSHg+ESo2oG8Hxm6+l7K5fo2u34bZnox/B
f4/m65k+h62cIJY0jOhFEOjSoBh69GIoIcnovai/xwXumzFT+RrQsvPH+FJQQ+H4
IFcwRsg7rxcxYpA7uZjlfby6IIW8FZXzUImnASGeN9Da7qPeM12ouBtll5H2zVgF
4Ts2+YurFqa5yakSsk6WttN9VtxUQaJBniWRMjEZbWEx1NOUPqWJsz8NSp4o99Bo
b+ZZIwDgeVepzZWPpgBmpz/OaEbXaExed/qh7ENudKcOyuqeN9cuwWxEosaR4Hc9
5qhsnY4UPUoI28r0N9WaD3Jrx0QjAtkYZfAr3uC9feCBc1hYLz8hq62Kbf1OY8Ig
2CUgHLgOar+mIthyKCnzml9f35iM7UX77Wbs8yVvjhX9S700W1Xy2J4VpbFpSDtW
LTBuJyxtOHPrxIn3BLTJ6pL7j2wOyrWBBgWilamRBqoB1zBYJ4IzoEdMvldN4sss
OQQATfyAlKlXp40pQek7Cc8KWay0AnKrriJSpIWqjAoumueZ6LLRql7wPiRjVjbo
jMdRLV+p7xee52QZRf6JaWOLskTadaPIMP09Z0CWsqN2Kf6MIKhRArYtqHY7woAe
rwc4qSgbGWKwui9e28O3MDyCp9RjHd/FiUNyC7lWMBO1UfW52EZziWlIYjO5ObbQ
niyXY+6lm80gMS13ywdvCuOynMA1f2Xd9hbBcT4ivGnIZT0COqVXNmfvd4szSxqZ
C80j6A8DvSeeYaxkBrCp4INZ5ButwItnzxgfjOQyQtMpl/mOsCC6HFyoZ/VVukqh
sILMgjw/9L5orN01xtTnbPIBm83tsybwQ9FBV57mc14cHTf6vqAiU4hR646lS0Eg
EKiZ5O1p/iVBmqXJEDJCyvxoKR2IJF/qnNvUpolZGm+eWO+JdZLBjX0kOF6WW6Ul
kxshV4nVW/NUzAynv8yBtXcFqkOFQJde+1v/2BXCufp6IljMqe6EC0HMRl2cqRaK
83KNImD0igXqJKiKV25gGke8RJsrtS5B1SvrYh8md0uBDXPMhYtvQuQzlMpnndbM
Ep8jyVm84NxgMLWIlw1kmureM9KX/uYKfkDo8qAebCvevnhWETajyrezFRQ8Qg83
iC3GkCfs1YEjYMbHNy3KgY9aGM1MkkI7lBmxHoGIm3PccqEQ7WKpwL7+WO9WSBKq
V97tDnj5ri9YsbkKovmlWKhX0COEmK/eiDrwYKxI1+7Cpe6LcAWOgFNep6cysxcN
GWCl5jzcaT38zeWo5P+M15JTND8W3eGcM45pXDrL1GdtAj2ZZQsrnYvCYpNbR06j
QejHVTL46IH0cVVJYjXhkf02HCHZLXY5q5rw3rUbNbzJXSLbs9cDiklW0RHo2l/G
yAG3RJGhOGwoSozNntuCUyc1ymqjz/OEn3Bc4ueTLhy6g1sXYBx43Gm08RiI52TA
j0KrJdgBEu5LZ5hL+J3eovhnq9Abj6hixiKcGjEwMwd/mr3GvH7A47zfn+U29O8l
D5AQDSvKW4OweKSwVS2gx7WzHhj88kKAMR69wC65SuRkC0vr/ImhatpQgt/Pdp6+
H1E6kFwXJppLu4f2AY9L/A8nBia63s+7t1S/K783lU1emLcL+TXJaaJ9xEVxswqN
6aOaqk8RCRrxkeTh1lwai2YJahPFQukEgbH5z6V7Fx42MwKESUkRdikJ+9p40PuU
RSRFxRVZVwCQr4tb5bedU+lJJmvu37+eCuBSxnhatNodDdxfpRAzQu0Wor2hAGV0
8UCKk/p1lOzN97iN04wV3oVCrk8UnvBykIrpxClbFbeg4WjtkGXgDTKjY0Yjh/eb
ge8eoUgECCmulczfugjpnzPADD3zrt3ZciHUElNt7S5mc4phTiX1HZ3QywrXvHRu
zprWdXWbY94NWRwdLFn2kAHAMvM1l8gXDabkc0cW7Y7/sDA9ZeJEPW7i/lg/DWJP
iv5gMIe1Yrjk+mBkxoHzJqUVoKQMlOkcImwxH43onnPFR9H016PZOLKhGwRi6q7V
2NHHrC9Yo4/7cLOy7M+8KWQU4aK17GxYYigVaL9pV7ClI7K/FwsqkA4rRO29QXrz
rTt3qz/JUP1QOlkBmzmEs0bJC57FT2djB3oXPqQ3pgT+JslRNXk5ZHha1IcNzZ/B
rqVtWqiqCoIJkxWxqDuaN2sjWc/6gsYpWfL75CjLmof9a30S52TTis/UfeyPuI+2
DvJPmfJJHW5L3exuCGwccXZPHTlpl2DzW9W915bZhQ8spFXLxinag+l2C8pKh0G+
942XejdsjshF8iGwrZHTK8HUkCqD93uWmZCQhAdDgyfR+ikHF/hEzZVLQwGqTHP5
9f6EIkNW5uOSgwumkgyyisqbS5zstL6SiPc89dJOQGM8H6z2L9ANCW4RAkPu2luF
iUCGY6fomlK6YJvImtrS9RxoQyIbRPEahjMcGV4mzamuId09sxgY5DDNeSxM2KsN
+uNyoA528ty4zxhsEPlppCtiex2W5W2+JoJqBRTF7Av9LGYyx3hy/7E/ix9SUIu9
rh2rfGLnAkXXoh7KtJM5QUD2oOePnuNQ3CA5wxGJV2hfefhH/l5RyL/04vfWR6L2
yWs5gtqNU0Kh8qQ3b6NRxu/4KUuYyrJl6sm3KDekcR5Pl7/YkZUKLyx967T6Uv66
bDnmJe7mvjItV3DBgSeqpsR0qMFPmeT13p2YpsjCwicnn8iTjOKMnMU69n+NWL10
uN+yJTuq1gPhUGaH8eeMghCjOyklssgBy8lITEhrNvglTHKtnBi+ss0aZewBWqKU
wIBW6rhhHoBnSwWikyJYxP7+HhZu1sV7E5l9JHXWMg2bQU+QVN7MMal6DdJAapem
YCQxpwLV6TbP0yI2lA0E1DOsb3rKtakgRz7GOUk/4hildfu1DCQc/8miKTOFc2K4
7fAS+tilhc+vVJ2l378xLHYoxm6BLMy9lW4IW83qENFM2XLLim6mO+aa5o+Ps/iw
bfuWybNZl72U6Ll+cEODf6UDk8J2xfqDPnoJ7mU2fG/BMKgn1vi3Gx12mXlfyqKZ
c7HaPaM5Loo/KMNHJTuq8ch8RuPnwb6k3HL1WXePG6cIVE3VqUem+2PzTMqfVRzP
/yi0WvbFhg91V1ce1o61ciFd0JArFisqgwGQaX9NSuZtZqG7RenQyEN4lGMbNqdm
K5wJnH0hywDKU3yHEm1bgnNBfiTiiKE7jvXY2EoLbUqwRW1a7RWbkgrVotS1pIOn
q/t5Eu0sq+lqEkpEDKAAtwPJmiqCrxJrOPGBWNhEHWnhVHWVd8wmGEGFsVZq/6oU
j+8zXe9qJkLJDBxrigSfNhXRI7E2Vf4PUdzfOfnQhX+lnAsM5DvIwCCAbmKCQ+5D
PySl0p6U0BhmfWqjAfKgUHjE6gRtSirv7Z1q7LtbAEmDrME/Mr8k83LimwpYmLJP
LVeb7pDo8K+uWeLxpGtB0MG9NqkWvdd00sLkx0z0yf/g87Exo+8i3/hvnM4DB59+
+fkrlHkPEjDdRJ0ulDPJbNuer1E4eyrBq2d91zBB1HB8aLujyFzGqEMSZFRyTWY1
ILI0TRHG5aCeGx+jzn93E8wvqOg2tAJ4humEnWcl2rJ1WETp9SkxVQeAF05GpG0Q
ypl+WmHkip4dPviuuLM2jk3GHUjsp/q0jSj7vQgRhhyVTpU1tCQ+d+b9otvPbcvd
gId9O2U9zhZuhk/6c4mIfuotywuul8VopQGSQaoCD1J9JBoZbvp6DI0zwfAp/aE8
el5v/+lmqL50sgTU8wTmTxEomngsYr+9J6uhIwgmynH520+3fW4nx7Tum8/njV7c
nch7gWV8HjMTTHZ/IOI6ubJF6jixdQeeDd6R1RdjCEjZsUBj/FpAzYQL9NNBsuCT
a7gOidDtAb4kmF3T9av7xdazII3/Mkbk1Ad/rpSVSI70Mmk/r+nvoqJVp2lTxA/M
7YFwVF0YVGS6Z2g9gXctcnvqDo9Gu3wEOZHDCPjTMGUgPNsOeEZAAAhiUKHIalW0
/MTuMGx1jnsL63uJWUJo4gZdMJTY2gsRZbGBge6sNnWrNWob7UHJnESQZiLkbOCZ
eEqLYk1cbRr7LAmGlf6uq/BeNtpuO5nzEtoaLsnmPzuZztt6fJQz9xM8O3HV6Omi
hgc7xAQDbeLSTKnHOnSGKQ/90ZtRYE2O9G/r/6hSIFHOr16+GoKsgG8L30NPslNT
my1r/d02jCEqBlP3lpLouqNg900YpIcr+Yzix02Vx6QrIFScXK/JHrQrjye1tGA/
m899VZpMafWBzMx0PkcxMyFf43gjabybw/F9gtdOdaT0GZ97cGmHvN1rDjWV7IMf
UlPKw2qyI0j4+9W5Mn8cMn61mCvaMDbv0891eIWKECs+jHPWbTBnkM0wKwmJdf9M
y1z//h4b+DeJAIkMmaDsk2fpPJKGtjsS++Nbk1TTub1zRqY2FjsOhW8cMtG/SLRx
xmfl6Pb6VNhVAkvuLWEkVK22UX4SvanrPEPVBRImccmQDaNJV4CJo791ZNgQ7f6d
YgHMZ3h7euGo1bmFoc0mbjzpIhVoAM5eEBl6DC1P5VylWVcB8O7KevU6atjtluEz
bbk6xmfTYKytGxUQoAIFNVQtBgse6rigaJ9axuLU+4K2qrEZOYgqjn2PvcgqG4L/
hpn0uSoU/OD5BakXeS8pzUDedCIcEVKFjFhfA0+G1cU4x6lx8KJvzlSdISq0dni2
n+VsP2fmcCx+vVMz1MF6FlsLmc1FsQ5n6c2F23fym89VFH+i65BvWLHXr5fDdTt0
WGjTjf63g59H7CbzIpvqHrBFVg71jDJmOYQg9VTLy8b0LM0TS8qk2UUgOqqQ9m9j
aEqNz1Wi3w8nphr7Bf08pGFNy2mQMc6rWMXe+2DSrAqY78JW0UOgUMs2CR9KOTFu
+cHIzNdZfnnjsDY1yzXi29uDwtGVoStE8G2Pm4hlYt1PqIXlj/bkpppBWCR6Li60
e4aDQm856sovPDHwChEwJFewg0zwYnyisqWvpTfrvadw4zbhrwwtZBLAv3Wg97Tz
6Xhz0wZ73ofuvC0vlfs6gm1cOGCD89gw9+Grxnfz7XkQIWNizilWb9kZTkqDF68f
vOUNai2bWXX8B9FePveGAjH/1pYmQCjLs4npWU/GuCYcmE8AhH6b6d7nLVHeqlPW
uF9IvdUVre/EGPuwt5ftKsQNtueAyRePAeWPgXoMBYPMgvKJIH6sQMQc/pWUYA47
UoeNUdxV2tlE16wMpKhX2/Ec+QvHZqFKF5d2KU8TPbs=
`pragma protect end_protected
