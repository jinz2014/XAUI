// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rXmmkwFPjgOrImWQCit8i6WOnq8LJTqAf8mB5wbZZyE023FE1okLCvp/QIYKp2GC
H7BHQoGFDm21xyNH33/OdL+RPMVGZ22wLB2YEyycdkHzPKHnP0xynYai8EBaIhki
fyY1uCd0ilW8WYwOzZ+zgXMFxlchkmeYJ47SioPrEVE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16656)
dXUSZ90ppYqJk1p0mi7n9XYH4BXnF1xnNuFsmRtCPLVtTjR2ITeAE8yrMPp2TIqc
XxAwMqROqXVCh5IFk+klyLSeBTZ8av9kEhDvz+tSAAGLBANKlk+DBhfZuFNifj9W
ogQiD51QBszsv1q6rni4eoEpOzlhPt0bK3E4ssPsNQu5D0d1Sy7eatNE/zmat1bV
KoiV4dTBQ/Y62EZATIRVmKVlXUKWhyoJbQjw4aO0XIj/YI4y6YLdXu90oDlckw3D
bqpwA+6MCLbOWF3TEMg1yyn1B0/dnQtixoVQOP/++kAon5BR7MXK4pSBvwszSrqr
R8UGcFUXh9RQeAj0D0XgTfROIMeh9ucfv0YxlGX+9itU1n4iw1kmEOaFXB22/aBC
uhLTHlBUNb86MPX7LbJbp1TIfVBrXZLfGZzM52WtD7k227LiqIcaYS1zFDJX1wDO
/pBX7j1qhVyYLzrjQ+1hn56pxeqyoJAtrPBhhWQX4GkX7JSm52tJxn9Fqb0eDaV4
c+0u2JH2TzFSpSFMq6Cp2HZqCjFLt+KQnOvA8CTFXmwFA3EjsVe/QV7xchP2b0ta
XORpHsxRDODfiLZKupS/NeYwty3dgbHLEtjqm1x/4M/SVYd21QrwrLeF5fGe8LgO
ZZdoeFZGwmcrr85/DZ2zRHfQ4YuplnIY8NlhxRsDc/yAj85Z1ikF2mEmtep/4Uk4
HrPQWnP1gJ3+yvOudJqy9ZlfuH1rHrM5vGvWVhpeEDVfuXRVyHstUXvIr+Zj8t5e
Em+6jmb1CI9JjP2o+4z6CbxaI29R3pAP/yixKzkkc5VGgSPyPw+HzCf84sP3vl4E
UNe8rmWA2fsBo4GRTLIrDVhHzyMepTS/YKrrnUqFoafQrRfDzXbr6lwMxcEeXLiQ
xXmWCPApWyt/DgP+F1Mh41Pfiwv0Xxv8midp8G6rwjF53inRDmdLnk/FFBc2Nxn6
CAohQLZ6Ujy/cK2WXuFCXgFB0inBtQfKXMGeOHIF8ytBq0qMU/DQuO+vqNMWxJvh
RKQ2cQ9mosmsrjVYyCkhY3bUrHg9sML9eaj5k2At7+gn2qp7LzUrsiw0+OzRhulB
+HhOK5EyqiRaM9EopfuBtXL23SKnx9yNVIRb+Lf9JofFDHCUFLbIDnJ7Xwa98L8E
nLb5nS0ZDleQfNKzf6df0kWbnC+m4sWjg8sAE9DTiyj9v3Kynl8L8e3oIwivX9l6
X/6j71siYi7FaB01GXt91y7ru/UIOCrRaSnP2waHzwYdoT+xT1kIE+mGotFdxKbx
u7R+2ZAkcF3zmqFqfspbWEupKttdGfgnHfnjdysSFye2ABZFQvzwaxgUm/zKpVPb
s0qdmQPZ0ZYocATFCu3j5ax3kbV5kLG8K3To/HV9+KoFzTepr1E40s40/6xRHKvB
oy7gLBOwOKAamkWQTMRqeWB5xKAKt0Y2qvrLOPXxNkoG2QVzbB/wpkGgIUbX3XTQ
7EaBQhKd5lAK7+K1/wbGno6dTOUw2Af4PYWdejyG9FIxrVJ116uQvBhxBGN1YlbA
wn1pIgATuRh+wlSVDFJyC7n4fPgPkYnvLUupsWpiEse0ZS1Jl4/kYf2pIZUkyMpF
d/XHL4vkuJqCxKbCyT1Dcu8KKvRb8rOaNbc5NEjXPNP2tMDbqDV5yj+z7U5zjOB9
e4wqrkvnQjXNk6THxk3dLTgZtseQQfezUkF0SpLLZ9QsK1TjGm+JbTp7tYr0wMMs
sUItpY0MTb2fGkw6Ev2e9jt/rsFTb6qBIpvN1qUVoeUgmhBXz7Ckzos4cre2qjIf
55AWJlTv4LHS/Bamd01c+/kHZ8ZsC/hlVNb4AzrsWyGYjU3codPHvLbWK1NHPuw9
FA4SAE5C18+sAdzZF9T6lg0Z+0BJCnWDdEeOuykwIebqQ7Vq6WIaiwH/X0Dydedh
CzgQXMdXHGzgc7KqTa5B/1KIGtPeYL1GQVmVvK3N+ebR34kOgfqB5bjONPSH5WjC
hQv8+XpNg29b5eT+jWHbeiMrHV7dxgi1NafXC/9XOA09NQUw9xk3aZhXKg7ypm8z
4Mi0bXxr+pcGJK36GIpf43Qh4DARyJyWqjPe8XwrtxdoNWLlvUj3nVfrgZQ9S4Tb
MQX8/gGkiPC76BnVHqmIgyTaPFH8+bd0f/+8nFjaPzmC49bXIQ2/F9paivAKmOjd
5EsrIDajA5NOVMLQV9lLtHkQWARSYz04ca2UaO62OUPg6x0/Voxh2HnsEGa1KonN
AAvpR4xPJvsHCrAerDcfukX9H1rfUKQwAHEOm2HKkE0hOF68hXlRLiTzCzTu/fdZ
Jh29RM5VyWVG+aaKFARfij/RDuNreYcrP+lu0MRyME+GwTNGz7BxoQ5qudNoNvrt
mYDv5eFLlF9iyabqgi+AQf75fuGf6Patdw3XZnq0su/3M7kvtU5+d8ktOgPp+13+
zUEnwyXD9Zi8WUZuEdwo9bpwqxIQ5Rj9lzNBNYpqkZdciJAv1VfqMAgj9OpcBXTO
dx/Ek9dQH4H8LCHU2X24n6RyHEtkNiH3NVN3OaXqTaTdjYcnd0/BEXUz1hR6Mo8H
LO28WPquHvt+d9Z1vXBmkBdcW0dvShTKAC5I7JDt0JZrXnCur51tiUKdHptULf7E
kRAnkHdC1zZ1IQ2c/l+63FgdpUUZ/qnCAGn5IRUmDdvAhLZIFUU/EccsTPtPdh5A
Mhi2DzCYTYPcG1pAipiG32hl92xK+9l0H4Cnasok3AbOHVrZn+GRTi0nHHp5MbpH
EhJ2ZabX+1F1tofQ5ov28YaA+uWfR+E3qXKeJC4qdhkS7VPkgMlqyVN7vKQahjCC
HPYmW2E2De6/ZpAeEVhQa9iwAuqNqJ5TTwG0f7iJ+hF45TqQBRUeCVRU8EjNCeLi
Im5Gj5rHqM8tVNWptjPRkzNP1vm0fyqvAgQYM+TVb0gdJlFqR6tIq0dbGDdRb0GV
2GPa4F8+oKImcOfs+uzcxQGeW44Vhw3+sVXWbNgh+Np7X/dAwLsVX9neJ0dX/2iG
fUk3Jlvp8cKdNSvJC9vqlKpQnlLxV/RE57GoUp9xa58GgRo47GO91uDrYQeIWx5b
T6k0YjPW3BdgXlEJ5Nsqz8W5u0dxdZnsATeGKVkIHZlNxNve5mzob8RsDbDwtCkd
mD154Rk8P6GFccInkbNe8FNxv71yJrRMH20JKZvBnYTKaQu3f4ghVGhKrZqyK+xZ
H4ooA6O9cEzY5q+CHtqoFTPik5wW2/KHu63tKpEMk4VpJxKu5UUkzWVqAHLGWM48
gWcFQbRJqFaMTPFhIEsv3KVw6S0tiV5ngCc7Jvq5PDwkeHjtvPhhAhxgYo0VIIuZ
bdYgPICyzUeQSdBU5LeyfSFtOz5TJaOXL02YGeR+dfQ6232SVcaXOVZ2llV9WIcP
TfAhhwrw4KFz7gHzra2N4A4IyO0is8ECTaxrbRNsZPfI2yxxOq0YaKoc9w68aflB
QX6cfI8VRW+2/+7wdtLZCz1+VQcp5US1PRk5ulNgZnQU+UHAlwh6vwp222/NFFSL
G59aTfF0Au7LKh5Sksyir6+C864dKlYupi/tj9RVGC71H+/HIm1ZXZFX9yxljCsi
fMzArqxUGaWyo1njiLDZ8OoUQ0tYFFAbc+6HwygBnyGOIHARuFVYk5BmIDnFcMGd
HvrUH5mPCcVZz3iAun+GTA9xCqppetBDgI4NOBMJeRMRqshj9M2XERBjSQYET+3f
cFR4bb2uZHxzcydruMcjvHI+n2Q2CWNPRyFpA5oiH518Ao/EjtlM01YG8NJX7imz
jXY8yy73c2I4yhNRmWZNdNgFYHbIUV9bu2Mq4O+2HGBY9c7+0ePBRlkwISuy15nx
SV9oqb0TGYLOhv49TIYqUTgyq34u0cA5jChQ1XhpWBtrMM401/c48vh5I4elufQd
PnmyrBdrYxCTATnfQJ/TR1zYSEwgjr9gpqQp/algKJzWt68tPAdNXNA83hk9JPX5
TWdN/WOgYp2vPAO25lOYpaGtNoLma/1Dzs5mGjYjQ+uv4uXhmldVv8B0kke1C9kW
HAf8wSCjPKgtSM+iwEMZxkUH3C7LvIu11njF742IMMcQiOlZnb2UFo31gUIRkZ4k
93ulzecvmi3bAY42j8I/tBZSOFucwQgyc6AOz9OeKT9MOP8H6zddtCt4/VXrQy8a
Wkb5yoh95oW5s8MnePNTHVIW3wSQ+hLCEm+3nSQlXD1eBwjXWOA0bwwLJap6SQB6
vUbvbFRGgWcH5Ss5b9R9qyGPOVK9XHR9SZc+2gIwx+qBN81xrrxfia/fnk8M0vbG
oWWgQ0eRdNgEHV6zVcb8HVvfe98va/MhTRDQBTUhDKzwbbIhYUQvSqLDlQfD2V6l
QO4fQvvw8u2c2B+5Ku5JYJrG9P4swdlg0gcQ4F5VEMF75Pcs4pbRTLbisyzbZ45Z
2Hw1xZteDg8Ca4mTeZnudD7W5abUtnK7lLZamZQErrVbtFwqWaC7xhEkEZO96vvD
qkKQZBSd4AZUXoEjADy9s9nzq5kg6r6gwKhiKJqjvy2630Pcj/xPrgB2OE4Gup8J
9jlEeXSaEgAO5xmbrs/qrAgOC3GwKXKbDPrIibcvqgxzoSzaqD0fQtbLcGQncANz
TYfFZ1boT0TSrkEjXXNVkefczcCIndzZxBXetSw4qX1x0tJf8ZsZpjoHd8AUhqf3
AM5kMkdZ4Xpcj/ZEUT1ViCXzYPnsbfsvMnHXKNs/zuzJbnHlt2Q+jwPASp/SB7SF
w0SGDDPvjlLhT55lIyIvrqodJKEwNXIQ0EsA+cETQfF+qTwmI4/umvzoljKnKvzn
hbKhZKCkRx3muOHHW9MuYFAtpUPg/W+FvfEdCphTbIRRgsGIyAMwITp4gsdphO9Q
WfBBS0OKh/6qF+i2TEBekfKWcvI+rS/CGhoOJqfoimQLHIupYKYwFPOaHUL9eH7d
Dgd8SRqYdTdtcfwd+0M1OGu2GhWhNjaCm9bhD9b4YB6FgDzzEv7RpsH31op/+mPJ
BAwsqcMzMnrQmmjVGNaeI86c/fJIu3W/rFNldV8ryi/77erlbLTXlkURWAdWTiZb
cjVo8Y2dRnazlziq3BI4OcXDe3haAKvFdtQtSOn2gnwRsoQxX3MX3BSKY9OtKmJw
dWUNgOuHfKYkB3uGAlQq8T9QyRCSTy/0+cct+9RkJknc+nTg60wwzkDaGLl2t6vT
TsWguNH5N++e5N/HB9OBqplPBH8Q3AFgzRtRDplpBknascDPKlU3XQkUl7ASDTip
iz3A5fWugML4tDNT9tPrqpzF1apleUofqs+IpgMkwcoVgCviJrp2joYlZYotOtHc
w4SEwXL9SNe8aUrf8HG9DP3nOeeESu9f40lc7T2PZqpl6CQxGAszxwY//wb0+9mt
ewozHli+IARMxVVDtf82XS/YK+88YG385BgzoPt+4gxmHlzbiPr3eC+BPtMHj3Qk
cDD3kZny6Yt87+fgA9/iL6JRZkXCRdWe6KMVB1AVkVQNgkdYuZrBmUEF/DPYkR/G
BjHgqWyRvoejo/ugbU/BBPmlkWiYXYsRoqc7YXseD7sYaXFxROADtR0aEUpRNfjv
hnx4QPRaWEBT3gi11mIeS+ER3axw5izUG71wK/RLm9hfhKzaHSvFRxXVYGjI9/Jt
89rlWnlc3mHl1O/IMfgmHtaZMJp9IMFhiayEcDltngyImzZdMl8fNuNkL6tAiDek
bAGXRRiuSbXZEKqxxuNkElJvV9cqyNkd2xoQ6ETUjArpXB/hSArq5PImcKHoCu+N
RFp1y1Hf/wjEdKSYA6N3b2gSXSzduPP4DIjQBL4JmwKkkuICiu0SPsQbHfwkITrY
/LIDyFe+RJTDEGCwcnTj69lyrfSkk40OG6vdHpMHuwyop86ZXN0SGLRSTdkhefxM
my2npmydbXJOFX77gW5aZhrFOk24hRn8z9VLyRotcrg9/dodQwgWEAzHnNTyf6nn
jYbAOnj1xlJ/va50TGydAzUriDjIerp50zZqA1hlWwSQKbwGCX5Q2rhlMPUd0/Z7
HmKvOk2PwI+6rpiYpVdmSoqvyhup07HNN0m2lXTCkQaBRmtd9HvnmuEeYX/HKcKz
LonmLLm/V5y/N4ERDHSC7Tskr2tykD6SwGWbg++GTF5hIQyrlte+RHUnhBfLE/rb
wjKrSIcBKxPJxgMzm+30XkYA66geSRP11luXqAyg/deMTZHJvQNeyHgdUQZ12EBm
Us4oL3l+BO1yOPe3aYnIF6wXXkFTXXDsT9cUce4S6ZmF4ClknklpzF8oAA5cVp84
kjIom/qUZlU5ApvHfJQ48yX8Y+PH2YrLfAZGzM3THcCw0fymp6TtIYgUzOlTED0O
0Sp1XY7aZG1KAt0FBr0aeQG2p3HdyJjHfazQbBQvXVGJc8zR/LHxgeNKd+iMzg8g
Q7GS1qT3ivmgokxg6Uay9ZUFq6pX9/NP6JsyKqFcDenGq7ILYm1btMTzgW5D3hDR
ig9MmOiJTJrPdqFb9yRYWtLzPcGEumHRRHO7PRvuekf7U8gVKXkjPNEqdENUNQVT
Fo53G11KiTBq3Iy1CPw27IuexIM0Y58NJ1hoLt+ub8R3GiUq7XWqfdOdhqyxNTdf
Crite3a1gCefqG4X9XWYiUEcgo8ZXlYstMheMMvIsb0EjAgZiNcOxyOw43j9LpW3
bjYwAp45K7IaTIjMD8TRhsmCJsn+wbVE4URacHUyKNhVy45rZyP21vI1YeCexpMD
c0bGUKF4852q2YKVDeIF7oiDc59+wDQhMjEA/zaS9TdVTy2nnT8ldpGLk4qSmRYM
pnrxjhA21mc72dEOY2fRNoTgxUWnIGTls9uIuREMMCGrH5mLCM13KS/Kr0wAuWqN
Hq/+8UojwMs4PQi9LVKh+HURYHA77vT8ud+MhKOgUqvxy8Uxbqwhl5CqESk49A64
8glZRTT702oEcgMS7Ccs/Ln4BNsGK5EUDTYhBCdtMXgdqiwddbxAIRLnZitWyi/w
BLD0Qxhwb2oU8BgwMaW+pK0ih10G3VD+Py0psXUq3+PNgTu4Xb/DZ/AqUIR9k6vr
rOkKJogHrJudztDNYjVzzi+LN4tkOPille5PzCgdobzCeW+SkNEIsctckwxwAHtZ
7m5AJ5SorT25vs8AQHBJPHn00HFIFudBXzByhMyIndioE0dweuEp+inQ/uUCBTqp
cSboi59z8i2mWpre6YUyHcf3qFTarfgW1ddBC2a+1pMEPbT7wy4vSt/tnLZQlGrN
qP0SmKtLr4FRXveNB7o6EBGqPLTh+hbLtQpQMIFJ6oGKcSPSG+tqZ99gFXFJcY1N
IAtuACnR4g2ieoI8GLB5YYduP8pIeQFCe0DI3984NjbrPD+p5HpdWBcO0269K7EH
95cTvCbBezsM8s8SBdzP2jYMCQIWxb7y+/2SxDlcLQPkfu85pVFIwWcqZZ6318zy
QZAlFxaZ4jFRfyIJiAryJwZnx3VwXpJmCyUFKkIJ2TH92JWTkOC+sOSuC9wcLu9Y
fXIoUx2zQvTFRGo6J++3PdJpynaRrpgW6nFT3/pT4EitF+JPZIpNGAFXfk0pZpWT
spX6qNy4NYqYMLG+KX1xFi9OQS2mLpFe+4yuFIpqIGdgjhM7GoPOFskUE3GS2/ju
bCkz434cmW//v5n25bc8GHAmSrFiJ3gUUV6e9w71y7nuTRbHXv507YbG1oMSf8yq
6hYyZ1I1Pq5h5La2LK362VVYc3EyveYECFrXGX3xjMWsCxyfE4dZOp53RI6ff9h6
7IdU31Y2f7YHIDj92tqMrlP0KArvLeaG5x1M6fFwDZ7zhrtkjqwmZ+fh8SAvDJvW
syU5QD9u1uQRNM1eWiGyfiFVw6AChlFwGDot106j2sSkqkeDZNkNZEoRdsJiAxm9
zebaAzTON4HnBGC4sGvPBZyL221caxlD/+4I3KONRPZCMPdvMTpzCysgoFa7QtGo
7rjKblyMW9IMEqsgyG8YouHLRDM3UtyL93QhiIK66ICoEJKc/ax83gt86R0xDo8U
QrW7iJrbDAqtMa4byAy+YOlF9WRpvCLFyhg31o1luEt18i9BA2IYg8VCB5+S9pL4
+dB5jzmtOymL5FCkvMgkYKJISgydBMmX5o29JUjZkcjBz919ltbpw1DaskMJNT9T
brqfOLNWN3g7bdu4IFCguV/kfXPB0NE4mAy4oEgsHo5pQYPRHrtxEZLnL6BcWIFf
WkGIUvcXkF82g03SGWmzXutiS1y1Q7ZvKRhGOOlOYMIPCIPs5xX9aOJ75ScJnIQp
MENicBcFrAxlprJh3/D6svJG9eKC3C4LEcAlcTGvp78Ps27kllkeyq10tZgajhbj
W1F3Rauyar22Mbr/qc+mS4MDHU5LJko6r00ixlGKOte+gu3l0PRg9FNf6MXgy+2I
uThzg7x25285Id3exsUs9cG2RINqpA8kEYxuZHbOU4dIxHyEt2mpq0jZwpdKqGU1
vxRuH35wIlc11NeCapDKApV+ojvlUVNzehv0FfWdaWX4xcZvhYtw1AqY7CHSnflM
Sf40pzI6EcXsG5klkycDc3q/wyd0huYjfqjpy2O23ZOONf09vRQgZZeN7SBiT3R6
rdWn06PkZK2OC7v+X9j+63Xh5zSMWUsR+10vO1n9tRjX5z1C8Ah9ADJ1W1ZLHjid
Be69KfnH89es3K9uPv3Whk3ALFcCN8e759gAYPyOx2e04ho6aHjvH1e6oQqx3aa3
iI7d8L1rBZvjI8wiZY+xGej46uPmSOdErs/99Fzz4E7Xixty9CqSY9TB3sRUvqdr
3IOS5KnQpAYholr3qyJybwp646GFu/mzlsScKjwSBVXe1rKcXiN5oSEYKLajdlII
DYHXo4fXDoIxjbcK3HiBAHApqucEhjQCQUiM20/GM5iI0GxAaeaPikxOeoQw0ML8
v9iO+ughgVnxJNtzdwn8CdWs6NTeRJw4pk0+6p2TBsZ/RmQEMn/wwrwVJylezAL1
JkRi2PXcP+pkEJv0yzEB3Pgybgl2iR1s9FSAcm3ET1YqekmzVk8I3y4uRvvcEage
7rT8UWamuAZLPbGhLW7+CxoLnJmIyw7ij3z53B7bvHfqIatry71l8g8lDzI1Bhcf
85LWuQGw87UIKu+vm1EKV/iebidRq8Z5vqTUKT+Ys/zUTjacPRfE2hzeQACMeoo6
jlnZLwBhVOybdkFpSO4Y+UK/f7lZac3OTPfpaWpACCkB492xIc/ooY5E75TSxTzq
b/LfrTEkrYZoHjmq/+uQslYzUWJ8otWYHFmg2wkgAffXQLNBce8Tu9TWztPQUI+E
usZXgFkIFVq9UJOFpJ0QkHB8ASH930/fSqJoHpE6SnBxqPunrp44UV6c8tRKDnnS
SEFGH1vXhG+ZQ/BMGuX6AxzXFWX656E4CjqD7KKFs6BqNf6Wkr1YPte547SQz44v
lXvG+hL1P1EJgEQRwes3sloe6bhD2YNez4Ykhn2UMA/xJ5/aTFygmLB4MZq3fCIz
usX0J4ceTWSUtUsruwXKsOiqyTZPRvJ6z5hcN0PUTbi6bL7VRxC2VeyGGxJB+oCd
ftgMoqHvF4O9WZ6mMPr81xI/hwpXKn70PPE8+CNPTLsPcn7ERcYKNBKMXf6X1zXD
BJzuPBye9PxGUTcsQZlNxw1vh37Mh5+wzjPzXvmO2qRqPkAf+j5NI7NWBbsc/8wG
uYOndykNoE71SmihW078Dq8SYBLjB1EZ5bWEAslaXP3CJzrFNzUcKEYSfWJrntyT
sAdUhzW3GwVUOx59FHriIATeqERmqrokT96bpkm86xVFehk2sQCedPcKwPQrVIrr
FRo0gEzbKsiLIIAOENUKESu+SXUEYLaDnlQheFlM6CiBsNIdhbtPZQN2okwbsUd4
xfSRCfHf0G2d3CNGENk9nItngmlYf5M3FaVLaLRCHeCTlMO91D26L3qG6Ez6jIY7
OCA+BZz6eMQ3LCDHgBxewdRGA/eB3+uBSnHWubNH5muNXnKAuvhRN7lSKOcBwoQt
BBObPOZW7/eDI8ZNzwqV4FbegR62/fKv3HoUwHrC+MhdkrzwCsf4qcAZYVzWCy8u
3UgJ+YtwR6y0yjbfTRGU54Jf2xbBh9LOWR1ynMzlHORZDYCf5EApN5ywvE7JK+58
km0TXHha5CGnqPN80/Frn57ofZNTO/WxI2jx38SOqBhhUhwOMTuy+jsjP8UL3jsO
KJiF+rpwyT6uI5rNJicAJNEGDA4j4NrabcI9UcroTzvACt6yz/EBOPty6Q14XxMN
DOrJtRZQ7sI007LtO0ypK3zJB4hrCCFeK++Gn+3y1muRjT1/wwWUNn6SkgsvPaV2
B9cDWRfFx4jxqdzQAOK2g7j+cObUJxDyYuMTYBsgopCWJ1X6KfNuMfdIlq6skXlO
Dj1CZl2ES1uAThrLpLDwXDu6PNFarpb98flY9EpsvxvswO+P5SzooeZReaSBhW4u
wsic9cLMUz0z2wGuShrWezXeslZshc1qO0INWAjYPJP2OQDD1ts98CMjYS5sk2Hc
4EWbfQIq8QrS5GG5rf9q2okzvVGrYwtf0PEnXcUYSRvHBy5U1zBbN2VrbzkpbYSG
KyaGOPdbXSakXHqKkgbKI5DkqN0XaaN1BbynLk023L4Ar+Joq1ORm11HyEqcqNrm
CbzgyKiWHEuwsxih5tJ+NurrEX5m8HQxOwmVLcSH5h6+yPYC4xQ8aSEhh4B1oAvR
Rd+Pl+glG08JhCZQYE5eQiMULYhJuDr4mOD+xMlBLPFogEJSIvcDT3cMfnA6J/PP
56SdiZyv4C49CNH3f38zzke3R/LUcDSsmgmnuHc9DXQTyeDE0uc4iGoxoe44gvUB
DcnTJ4bhd3+y1rJHOangt4ghKg0V3+89+6RZP9dbcy//JICAiuFCzuDfLJkEQFP+
NGYnDHqq7Gq/9+MDljNDI+xxIG4FXehTI/cQ5+Ss1iD+x5Mx7nEXRQLGWNqmZHIa
HpYUTpXvVr2ijM+/fXfUpDrdolzcmOTSuVd3z147a7i7Pt3q7l7Cq/3Bgzn12J9N
Px2WSOOzt9o0UbsSu2IswQaah2Y1vr45xjam00YqsExHpxbjGBCbcaLt8W5ad59L
xm0eSMytQQD+X/A/TfYVRkokOYbBOkQ5996utEWfODGN0a1zFBu+XYsffg4oMtKv
yXl1McUDeM1IWYBcQ8zHqW6xAkDhRGy0dNHv3TgmgwIqD0AJJQeMaab0gu5M4Wk3
3EW0iF0M8jwga11jyiPc4QRKyXSi4Cq0PkSeR/X1emdFFre7+4qoDhFNPDUKXTpI
OtezdJXLBctKCpvYuKMUoC6w405wi56jhd1FQ0DC4rjPXC7JdIrSTgRuyGVCVLS3
sUDTeNE+y0GYR1qX7Iv4/BWuM9pFx42zs5LCcA+orFP86qh2gmN3WDIXgmNBx8Kk
r1S/5jXEXsDU4ILA1q0c/O4hcpdGsZMFFVtfS2Bo7iD95NrIX8L5TnO6CJQ+E04U
AxXAYSDP9AHKb0Z99LRoMjEKsVZ02ZIgUg7v190ZRijpCnpYg7ApvJVIDkh/Kjhp
d3BGiXMTAB+/kq7B9iGOdHWNne+V2XIqprSf3lZscJsx45+B9Omd4v9WDa31YnII
rSh2KXIjeVwhvvTMR0W2/Hxpzhs3d4B/3QJI+Xmz+DoB9CYWsUw9ZLplMaBpw4Cn
gUkwz4e40rb18FHJ63VqLkbqBUFcbMH1BPBbHJdDk6jTiDYekDXUWTVnkPep/u9A
VMUkV6MZJeoeBS2ZSF9E1pOwmKk3WxWZ5CrM8xk8IvKGwLHn/BTTNxgLVLMS770j
aoPZbIjdxGh93cYCxrVjMJgkebf1qpF6up3aGufXep3TbroMssYolNaSWSuWNHP2
6U6FtN9aj5qan515EWFNq56NkuH1sRQH6U7T8eZpWxvXCXmPOpWrPGSwdMUPZY4n
3FQGyiB4YP9yswOiSU2P0pcdp5VQFJluClgGvBQ71dcRRbd5whk0cYZiQDilkjmY
Xv5H8z6YfonzU+IbjGQ/MvLHLSe8w6ozDfaane/qFQweKnzpd3BKYwxp8mArnLSF
HKPdlmDZ4zacrBG6/Hzuz0NC86GT6Jm3YFb8t0up1Fq2bVFp6SOkGlGfS+3FuJas
fzRlH/mjVNWxnjLvH+0BWufI6Y6rvXDpjd7Mr18yBey/mV/CpEa3kzuG5dhEOyvb
VWZHrdhlshchM/uziZc/LHNJSTlnFR+MdqGFBEmUPzRWiRMsch9IZSLl9fIDSxgX
kRPNxMcpNiyWReXpilTjVy2k5zAZ87Xqk1FxPZihZy3Td9CvDhD0H9UWchVeA+22
vaMVXLrClueVFslz6PL1mzEoJrivuDp+wjX53qPUPuOw88GJ2xh48potXB1F/hMo
/T9wVsNmz7uOQ/NF23RWARvbaxgfeYLnrdzxvvFSfZSehuIoLudHM5nrrwcrp16/
Yop3zLRNfEGP84JQyoGWpYXW6LWHQOYbOuvAQKX67r3XciovSEPlm59aWc4i1/Ln
uSPidtphkimxpyKNhrQixhlNCVS2Qr61AaBRJSi1TNBh17lGHOeiE35Txr3nQfwd
WUoneIQVXOpiyFsG0vlUmJ6ja1Ed4Hh3xGeX37XtdTXCH58X3IybvxnBIPY3wbxY
Cv47Z0EdhYumDv7jdFc8UAONWqYb66kkrkjoTyDpDwifZPBMgl/5PUQQHHkQ0Qng
FkDoscGVDOWxvDo6QGNvDe5JbIp0XWzdCHsFisdDjE3rQt5olTN4rMm3as30eb2e
Th5/8FfY+PeyDVS38SDU6p6ds+GBFs1EW+FHk+BadR852tDirtVOmfiiLDaw8TyP
GFCJ/rQmm8aOSbT3z8aEJrnS9yJzu3r7SNWzu++GAG45ESnh9vVsrc8twu8wz/bG
ogjV8i+ZC3Zp9/0OAEGQiYOniDHuA/W5zvLbyK9ApLbmZxc40dWJSYaP+1oyZHYw
x2QXca6C8Fg7BtFhetOmk89QJQNF9sqGLG6kvXGlkY8nb7Oa1dGJdxE/9pyCiW7K
/xEUGQQOJ7s2QgPMOkcfBFBZB+IKNpFcqat+zDBWkz47at5swHPqYK4y8PzVJsZO
zzIGx0jLVM+95B7wsHfcdyg+Zjwl6luBDrXppJKgLt5jmxFrxLv/WiZwbKtrxKmK
cJAjynf1MbAPpeh1xMoRUzWvfSu6CD+m/RqLNUPedWsHTVwQ7Li63MfDJyiKSwRZ
UEl5ccwW/xIBmEj1dMtFjYZGpYPa+q9NVC/dpOFiAUpg1CPDANAzxXlyaqybTyzG
X1lUWGm/LDvgjpmNe5z8kw3x29Utkz8GdyvWSoX0KUVGVDOsFHFki2v9AoprHKSz
aSDEyozFwJOqLrwrBrgDsuts/qhjMPMQDP3qSaZSPGWPXAFGDBHpmU1V9FfJ4ASW
BAQPBuoLQBxXJ9vJm3dBnfvYu6Zf5jSPr27I/nvJ0+UsEWIM11YSiiGdoCwB/FHB
qi9SeRe22sAdT4aUvZ/h+BTFTInt/8Od6epWFRRu3+kcpBht4uaQAC/U31nZJJGD
VZFk4sQM9ezOyilvvUv+bzkiR3p8o/gGSxwzg1N8cRNNjHAFuYwxuUR/woJaI8vw
Zz4Vil/5GSaTUmx2mrVpbjJk7Or2FyMqRn34sbjuiL4jxrws9lleCFZ/kIIoXIT/
IuRJAq/M5xfvNFTS6uuVJk2jnxlecVmd36+WJQ96cG+yBqz+asfM6ycFAhw/XIAx
wqsHxd2RPCJ5MSBb++GANcyRsVTeNfketFzf2ys8lnzRywvdHWkYmhNKzWhUhxp2
Z+QjdtlUO0kFP0hmaSGrsgWtgUui+dzc4xTfglRUJSEsy80kJH/xy7VljvWsJJCV
WaXIafX40Z17i9CdeF/985nXWe2nnmogrIQcTB/+aPm++5MkJJjWgYQbV8AOxst0
xb7P95HaSyshovjFF04eXS8DKuTRjcmQvAwhXnndSfvqN6Fe0ayOzbXe4rJ8b67u
2dchXbZ0o4oMt0w4U6EWVtmqy8dV7md/vVyh8L/+5wFndQJipt+LTFhF0Wg+KWq+
xmitmaXKqqTUHrRknWNwLBFD40wSG8aMzE1dWNGU2gnV1y94IXM+8EoTIMf2JCYj
KWZDSeerv9r6XGxp6X0l57w6mJEToBfPdIARIXPpiM3sDhXOyelsoYMBdV1w9d4t
OXj9T5iYD1S4j8/2qxcT3XoZZelnh/lS8dF6w+TZ9NEh3h7ih3WR/4uf9e6Ss+xX
/EFcu8liIhJawgnxPR/IhDHmRxBHA4Opu2JRweLzh+R0xArs/V8M5SkY5YpM+BCy
TJGPYn8I471YWB65qkvFqVcETbfKAyhjs75++yZvNEPLb1CxOZ0VG11Zhbrpw+Ob
Rv2SIn6Tp0nVI2Xs4eIXLd3BZh0S8yTsUpyLVFB8jc7ulYsmBXbGDISRGZefPskZ
8b5KiAfsIyCjeDneOGwn/rbViMSWaMnVDr3PqahAK5fGid6Td7FlxvgQz4OH8yTr
kIXrfCsSfOM2kLf6rqpD8NoVPnt7Z/5TiYPD7iInvta+AL1G/Q6eXSvLYcZhwNQB
oZzNrdIyrJS68R3cp3V9ZuSe/ES+5g6dKQbwbnBUC3W7XLgDQHqZmucNPzmgF5V3
P5uSoJ0W+zIkhZCzAqaodF5x73lcxdplm9Vu4RbCnecO5aSqzqrphCJX0bRznB2D
iCkgfAD0KHf+3iRkEvkcTf3XVggrQuj9ZmtLrFYUcSHVfFGDnxE+lFKmmsK6L0WD
iA98fpny4OPVy3XoYQrM1rCBKHmPqKXBrSTDtKyOdiQlwssGoW7dS16V2xmhTtZk
6i+02WzbEZE/smqVb2dml4V1XDGHngnVWJxvMYloU6FNtSvDY5tr7vPoSEMXteX6
N2vpnxqkjr8YqzIU4w7+GIPdoQvDS7ibSPbrjUrZ7IY/s6GfgV15Od/IRGdDLs6y
JDXmtkyEzKa4DR8r9v5rTyudZJS0RGanKVLkJIBJe7mE1obxuMumHP4FZpxxTHTz
ABcu/wPkK0woE8JZ7AknFeYSwj3oH+I6/v2SbFfHqtxN+YT/xMPsX/ggBV/tHVHy
25XX+99Oiy9fscYTlJbRamJiJWWiI3H/V1ze1/xS4QxLgnVWSgAfmeXLWdfY8TPX
lC6sITA5BtTinP/AsBIS8SYNvdoIV5F/pfFa1ZXY1VjRTdKqDQJgc7iQGTZPDDhK
Xr42ZF8WOEKS/zhr1tDfvV8kW8YNO/YoeZzUSRk2tb2kXPTXHoo+hoXf6VkBkj91
bSZnl4X8Uz/EWp/pv9cIo48R4tOyvog54NHJe0IUai+RQO04bw10tpzIdE8+iqni
WkDC2Xn2i7mJAV6l0sT3syce19GJWa1qsMD2sLtkZ+E0i+socuHX1wpp3Yer2dex
nkPQSJCJID6JlFPgEqIPvqY8BaDwDHF81HmZvtsq53rv+Lg2wOmRt2JhuAM5RR3B
uMmZdnFx2JMvyy/d1LiBMCEpg2aApK/yJICLtFRJij/vxLghX+SYANyN4w4Q0Yyr
CmmfBW64DHk8SRcjDyOj5NC+RDlTXDzXD6sJfwDOOkqRG+rN7Kb+KkP+s4UqnVDP
p2Y2Zksc0ixmnpd2miT/vC8CBqnz44g6dFBB259duik70iiVtYXX8cZP4OXXmHlZ
vpQWWYx+m+9bUZIIHPE4lrPBUJnZ1CaEvDGy70Phynbfth44FCvhQsNHRTM1FfGc
YfzMgaM76bqb1+EGUtHx8qB0OVa0Xxwt5qBUFQzblB0USIAYTf/1vURtRftiY6X3
ANHl/rRaEN7UrxR5TteAA6gLOr3cJ6x5v2/9zplu98zjmRWm4yrPkyc0TYBMVHRX
gRalzbQsgQoU+RwNIW6PK8RyYJt+5lmgO5kvyQQsoPVn73ceS8sMKred4ydeDiYf
v8xVcTiBb8Ve1Ugu1Vnv2YpGU++5IaN7Ks/hw620hle3qFVW3LHRqTV8YNppT2x9
Kino5zlV38sJFATxNrS0TjZ5gcUaBZRQVxLQEsRfim5ChhuBNBzMp31sVfn9UIj/
2uicElI5K+ibKtQYVN7N7Ot54oXN+iedwEpWxfeTnUhVwAPWeH3Pwk2Al5wbVyxv
LHVUBtyBxhDiiEfA+aQQ4xE7yneWk6dk9I/qHT1JGdN0VuoVl7zXU0YrjXsAURUT
2c7say837c+EiW883yRegDOtzlPaYp5Ql4gYekMZQb5qlSOPrKCzTYjaDrIgCVi3
+1JzWisUKtxbGsNCwTc65/48xrmMi1W7IIu/x7uhKaWKfBaysBAzzapG10dsXbGS
acEZSqUG0NwrCu4YjImpU40hv84Nss2Rb7Gnn1XnhHabLBrTuNniZf867vHwqA4a
CxqXMzo1c/wUtaYhe4kqpE8JSoTEpAoUmp8KZxi2rrPZcgETZC/gU/+96ErPbdZo
bRvtylnkxu1rT//YouI3dVgMqdx74m4+rX7tnlduqDdXmERew3Iidr3QGB6tqSti
PP/3mhsmpkp3qjFDdHKPKE3sihA18rIsuG9CtTF+Fs0zEycQTw+xlL6qaUi2Nzhr
+7JxEYd4bidNjEzsfGJNmkVDklSNRiD26aWr1Zw9rKPotWoE3qdvIMjPsCfbo6kt
m2dHjyU5y1SwctK7oCNedAuYE2G+3rPa0yX5+33wTs+w78t4pzMYi7jn+/0Al2h2
DV9D9ZI07iKcXX2XI1oQD9U6pSv7ygZlNtuxwgDaIZoiT5iC6HHRdVNuYEpkTnof
Jyx8hsI2yKRYUztGVAki1UnOmElaIMoh7EdQWhRIbLBAjBrqgwDJoOz8eUJVs1dS
QcubC7I61I43TJrWRjUV5hvtATwyF5ddrnc7/zubHoq1WEzUS1HTagIvCYhIWpj9
X+eZavDXZw/z3wUV89ZIhakyxz1urZFrqpJyn1J6/v1j/y0wyqpz6W7WbjdFnTMm
5a3TuyV7t7ZzMlgp36oZL7L8z2EGcfAj6mFBG3Ri8MlRO2Ami4gf688kFPv22vbx
fW9mMsI/nT4kzBgK5/42D4wMLzn4gE7G7GHXSmRKL1UoXZnHmhhoOa+v64VS/3Cj
umOW9TScI0Xm3clQqqBlFI/SYVTrWH0vLb/eJJtGctdwmix4jH96+kL/iuACXmKE
yEYyZC+fp4WRcbsYsSC3WmNqsaup+DEri9heCE0A0AlLx84FmZ7T1wiJA0Y5P5mI
WX1gzN+uoU0Vgy2M61B22K3L7dQxfZUXXgcfvDBH7XiXE5gYAE41aiq9NLWsslFy
fz6eBW+nmbvze9k854Xxr+xSd0Pt7x9Ky8r+cdoS8++lJknqIG8e3esFKfd5aX3e
111EvDfS64u0VDbhjZYsNzyzklwBcVEA5EihZxeGxlV4RAQTW0v9nDUedaEKpfTs
i3D11agKwT3qprlnPxWFWbpj2HMtS8rEIT1zCa6DUcAyzyr3LTfZLRq/0AHnZuqd
aJEyz8MyZNn9x3qOYqEdk0VsKKCWGBgTxVqndCfyJyplRGDzbrUg7Qwbqz6wDZ0S
KROcAiOh4yrkzMrGTLlJKDxmq0Fw6XLq1DdG9OC+zX4KqUAwhtWeNG7vx/OXxpe6
/uDflcsw7xU0mLCCMxGimOEF5l2mHLB7XO0gapuivDsnqCJJA+B6TZAgiUzH5M66
0zQdd9DYMGWb8L5rJ1SmYkTyFH0oRgtvMhm995jy8ohAbiJ32KV/6ajKGOoUyKvY
s4BsRlTxM/3rRUDtsoxzhfAHFfnqn4B5buO5fopBD5kEdHSGxgNdF8xm96auPllR
0tL6WaQTvstZetUrnuQsZj7Kdl0vqyqJ9vWg+xoDjtfeOFF9Mc/lKyOmjACkRzAh
HNyI0eY/jHJvWlRPIk8OfXnIz+7BaS7XrWRIdcvZvcPov8KjnWbXw+SK9TmvdVqo
F+BRXiEXTieKICB7CSR6EhKW8oPOZiQpsUZl9YpzDIXL9nr5qGB+/cU64daK0OJ6
V61p/jMwfbJGy+ApHV7sm8wr1Q+lf1HUWA/9DAPHopWcYhO8B9dxtm7YnGTNlOZN
eCy7BHjNqYXdULIhaV7N5mdKTWlzWQ9R8OrqeiumCtQlIdqejN37fjXfB6N5f5sl
6NyUKGBU+e9A2bsZx0Y+Doz110adCXklwCP0w/AwbExbNm9MdUOD9ekmjJBgiSYB
pFR2SVl+G4Ihd5+4CTESRkWIkquiDHqfweKUkNenvwpFBAyiJpojWtP8uPp2A+RC
ahducFSYN/X83htcj+fSPLfNbPmZjZKipEIIVn6z7H/V46ahlHQIhS15vu9t2J8l
eA3/zdg0UaxqB3+aAOryZNAkpjXYVMeSynmAYcbXMy3hxBkxLiZVzQnJxZ3jR/IM
iMczJgl4qdX5WNvTG3KSgYvUExtmlxa/u3Ju3pXFy9GNAqC36elzEbDL0wi1Xpx2
scxblcCwqmKxmJhnIK32hEU/xOGiPwuAEjh7ZkGJloi5bprA0EtZv7/U7im9KL9Z
5i0TyilmNVIyE100R+dBypTGVFPmO5lyfExlZIPOJu+zrqRTEnI08tAiytZGZYeS
46nzJyn3b+7cTGYUWwi/IKz8sKzcTo04fP7VAUi7MWvmaC9hK4cgjO3kFluJJ4rR
orV6/6hxhNdBLge9Drx9x5oktlBv6bo+uYyS9JfUDZ7/h/Zlh2GLLE4Y68lXizKY
fN9qmNIH8vTf8FqFxoG9f7OFOgHUH6vxDAh5MiJDZK5PY+U1gLBiw2xn6vbW6ur4
pNUw5Z6s+8xx/OwXPXuwAV/w0bar/jbpS0SJzOBFOL7711UwzghRlSKnLivyi1L0
LNKPT+1fkxAGr+Jo3ADF/IgKTlBNnMtRbakzNHj1OBtNHR1+q/lFdwErqGyn4uHu
ck5K+NucQehTFwSULZsuRWMQXKWoEzPXHfbk1IiABJfXAxXp7iT6I1Zk/IvMt6Gj
Nl5IQy1kltNOeP7PPcPldl5KwEpfJ77i1CGeU+qCyQTmLtgkpFkVH7qFpvZ0FXwu
Q59KXTrwl3wjgZnigglyJwULOz79ETJjUaRnYlB6PB399IP3rW+k6z7EHO3kMEqA
751+Ox+tLC5qOWg5jq9urq0M613GamNnub3afp64ZCuKfOu4jNcFY5vgfPbJMUy4
xn6gjNK4gpvbpwifyhSwZry2JRxc2APecemV/ksnVuYE9eCk9czoGtlu1mz0hN7Z
x3VnfsjNW/4YCfuFkN8QTILoDpOq+iEXgokVmNugxr18k2bHdwgdCKPQrbfIrGxG
6U3JyF+RMOoEhYoUA/pJLvmu/0NsKw2xnwBDj1x6X8OojmyeGDKzOcZ0h1rLcFCn
GJkUzxlsTSemFoHLn0pfkw3KpBY9OTMalIKXocYofk4YIdKvTDcrsED4WEZJpIH4
/jOUM3jzjFkGQFuZkxuvHDvssV7iVdh2AGNKzTwj0nWBzr9/ToKoSoNuM//nHgGF
dv+uXCz8tuSC0aTHT8KcA9/c0vNFCnPthXA0deqmq7DwoXGrRT2i0jsKGSPtwL6r
r+AijgWsMspzIUu1T7CPYcq/GNdSdKPFZ82P0dEl4p3kIF6nqyim4s+UfbZBmcKy
Ptzu2Xdyeo1zjkvTFT46T5ivUoCJnsz3uAlRAAmmlcwud6/7mB33NsSsYVWc5Irv
k7JWXIh7R0kCGl+gTBgLqfO8/qG0grzsqG7sJAIwF2bB7NahYxQDNBwmNUTPaeK/
pAE9QsHaSz7dO5eD1uPKdjR1WBax85touHEE2H30mTNdMQmwqOSN/ylhRbyxA/Dn
2wH1zap4tKRdAp69sV/zPYBtzFbceOFM6K0QJdgPPVOCmipbgBDyrYFIH3hDfumH
2N8XZCuB5FKhPrxmUtqSSCw5eO48X6jV2D7O78DXbVnaw2N12NwgyxxjkdzVpkZn
b7dGJsmjmW97JCye+FzbBFBdds7EP12RQ8LfP2z/SHjQb5svelng9YiohAkf5xx6
8ZzHiTwW1GVCDPQVl3zcP0e4fImLDXeImDvzvVRbRUIVgoOpSKEG0o+v7Zfyn5cP
zVj1cE2Bk6FOlBLP/lQ6CQWrIIwi8AVpyRZAHn+bq7Y0mp/PMOJkWejaJrNL+1pS
q7IAgPVDoFGXlAGW7pN2ppT5ZAoMxl2VaLsl0s7HV54LEeJlqTcEsXKPCJeHl75Y
mf+3M8C1aj7nohxhJJiEgDoaRGaN+87VphmUYrDXVueGS9OMxceyGwFk2wHHw57g
tkR4e3cp4s5CBFPftjmqKxBuzvHZzZBGBUD6GWPcij6fIKnhaqToCxl5k3/2naIx
iHq6dOP8l5roArZk/LtZ+rvQQgsGNpXbakla98LuUt64XNYLz0rlzUrTQ3BSn68Q
HkHRUBSSHv4J9FPdP1NVvNxRSiFXpcpqH++JjX1/tFHC7g0lQ+t0j6anexFtxcv0
YiXZmkpW4UEjXHrdjstSSS2EVd5J8Ksa4GejK8cQFGHKBZExvu/4dwFkAaHyXg8j
L4bwnqtPFK/sBs9FOl8/mJB8eBFlMK9FzryvkK1xsqdz3BOiAiVcLhzz0GOWS1kr
AYiQLyT8YaGnINQ9no1/yNcOgwrXCK3bsQpJi2dmZIjnMJPVTkrxhIBQPf+ch8lV
8+jbXOyOQqsHpZPNdfyWnSWN1WUCuiGYTjiNbryLZq+bHVT86KEGXFqpNG9vk6HE
IIbLDq2YJ4io/c0Tl9aTM/tCwyj+S73JrPdxgyLNQNkBIpUtB4VuINlh0VWZZHtk
EUvFFBrsFUmnaKgaz2MPj/FCxZYDNczHAas+eUKlmfLeXijCECymoI5H9aXeSRoO
GxdDl7O5NJX7q791Ztnv2l9UkZnNfx8WBsFBPo2eSO2w15mdvI0JTNTNw+6dtHXe
nudQrpfq9S12inycJnJfCQUxQ4XdeVbXFo+mu4DYwtbBYuzUIjnstf18BZer9l+p
JibxPCelZ69dps3JgkuSpsF/VV+W8CM9wxXZj1UACDyKAsHWEqDH0NnWEY22l6G8
cO9MIvezSMIZe5yvXr6wkH3cOgK/v9ZFyg5Wp4hiC1SME5DJqDoATJKB/J8EyKUr
d4/P7sghDtGGUlHhnPKrrXO0XsuX+/lhiR+HNJj/ZaI/VZ/SqdU2ZTDRjxYQ3RvE
s5ThhHtF+VmOc5eyBptDmXDIv3Jbj8oy9NyXAfrL6ERsy9vEJEr3/WwOTYvIumx9
p0JjjkdL9alEU+V5cmX7+6ENfVdtS3pdtHFvHlujo+ET69Psc22czBGo7mYg9prm
vVf2nc3EKVV4IsiO9HlNNw3/HMF27QI4UDERUjlRCohbfbfOX6amo2McCJbtryf4
iYh0whXmAnVPucMCoCxFWcGu2Ie3Ugc43yE4Nfq5cRNUugVxWiDfPIujZtND9FvO
4mF/QNV77+72UkIOAS6y5wq75qwc/gQvhxrgPHkxDmILCaXHPqSsk7/HSdkb+MS4
MYHSDwKI8/fYkF1midzlWduiDQrYQAG0iWNQ9Y6CbkaJUcBLb0+/tzBbLI3thCBv
IaJQFG+YurTh8ZbCMFM/NTrc8DpPAqEWtu5tPY16Nai4U3x8jSmCTpliugwLwM2b
qZWPnGSQNG3qEqk4sxPeRALZKMNjqP2pyMRkVTbs0wHmvN0LdOqJp0ccy4fk490J
+yGYwOqHsOgGDsVUW70pUKi+58cKwp7eOeNbCzFubFfWjp4uxwFxojKsE6wy8qYG
vGlng1Pz0mw8XaFyY0Vicf1sTS/UK8pEJphDZd9TFFwtEjlSJl7wYDXIUHnUHo0K
qOAexv6GGWaBircK3WI6Iq3+hjLs8hpsVeUwZ5I67vOI2jIol9J8eD3juCWgEvZT
GtVKStEbJ3x6WOzao1cs1sRSZQQZQrPFRLVk5I4b3PBjPv9MdeuvIqh1OGQEGCzE
0f0CpkgWmlPOMDniC9Kfrbzg7auDGZET7UCqLI7GhmAsxUYRFsF1niYzhgBzkjh5
/1iEg/d8NI+syDVHXzytX8WSWDl04Fd0gmZHC/uLtWQ2UITrh7BbBXShANhqpEMw
S1VuqL4+nnS7eUhswT2kDgSJOlhGpNrSv96SW1baerbss8PzRhkyzpu+JObfCGYK
F6KpFmiybXuszurbnqFboNW9cb2OSpZQwNUvTmDJRHlNVKunVvxDs9eqlXiOQtcN
+Vg4ecMQdFSnKIz3skcXjAbb8B6irgv1ZlDpUsait7dcKsFbhqierMptCRIv9kTY
NVGRPrABSpDHuxUwIQRgIM4lCmBSgMaMSIy5HIgfwl+CHiroK0PYgx6Xn2FH0vRl
`pragma protect end_protected
