// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cd85dbUDJQ098Qpc5T5f5lBIAax21SXjMRiSlXT6926j14gur2mL7Ul1HQb7mMHl
YpesRDv4TAIJCuGNkj2CnbZLE8WiN4c2BfoWElfZ3uWJEYw/RWRbtvgewz3RCLav
R1GjGN+EsccYz/5AsqVDFYxJXk9gxUjrCvWBTeauTWM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29360)
7D3l/bO5ZXb8b9owT9C3q6BQ23enLWXDG4ND6Ljc/Zzj19D1uKbzkYSlgbLcp78F
+7kiqv6lfeuAlOi65Wl0PAl70I4AFS67fFqPAYX8ZyRZd7llg9bkhcK3RYMQueI1
P6VPHIOt737L5deC0igBcVIM/hFu3ZJbfK8A0UoQ13VSb89oFZ05gTzIsePX46RS
P614B2zQpDUj7m6KAyjMWYjS1MdYslCBqi/dhbVrqSH7UGSPJnJbRXqPT8UXimLj
rw8AOkiAd9B1BywHGkm2+9zoNy3aYiCx+OAhSRa4e/md1E6SO3ZWHho1kV07Iy5m
PgBjEfXqAEUpK5WBc+A1E9db3m12DE2BMBCi+jAMfoBvYpgYMiNafu8kDTPMREHG
p5q+omUEUyIZWAhuWfLRHcePHtHIfBp2G2ax3dGD4lPr2qVFPyXUpynYWyUEk2CS
rbpKmIKb+Jw3d9sMNur9yKh+ap+on3HmM4SAXEE8e2DdY1zUGF1KAyiKWT/ulfhP
Z4QzOWjAC+UVq31ZQ4AoEGcRItO2dMmS1/v5g0IYr5IVaClfJj5p1MmsZGdoNZjA
U3YQhNfXNdwm99amOWDo8WHGMX+c3owEA8fExZfnjCitSDCe86DGnGWWATEVdbx1
CxfrvRMEuqrUq/cGdxNCPUZxlWCcu+VMlmKjrpfb2TPG7Gvb6967NiOg4zMQluaW
Ep0arbYaMiN8jBfMBxG2NQHDxuuLxW3ixKY/mBLFmK6Tdnh+/rW0pKuExz41cDqu
mi9PH7JdRkNsEpPCiI90yxDeWiRSDUbRPC77k/2WKksEPTzEOjfe5lezUnnKRPzG
M+sRpDvoqaCNMAUHx9+8JkfS2L1CU3w17RsYEFTWVqukTN+AfySmDo+n4dQMF+/t
/fwANK9pFnjQLztGLv8QX8kqdk1JpdIakoXM+Q+c1IB0jN1P6QDcv+qA8ifklF9z
vUbqHWwTcBMUTm2OS6rGfU2AhqsZCL1/P8B1YoZIkEaHoJ5RLvmx2/wd/cTeuwvR
fhZRXr7kP7clNlKdU9EokinhhvW6ypkByOgLIu0NgZCfWmMklwT6FllKkCPlSlTB
7I8sROJVNHtmsl09KD+dhTvnF/EsMH6zOYA2tFn07UWn2aGWPrCrP2OE91XVMvvz
ftH381mGXhrHA/7QaG8p1557aB17jB7iAvI8bYouryaVrAlBN6BCCzpVATNN0tYN
Zvq4K/mr8AcsghZSyjQDPaS0G2rHn2xCdjPRgkUZrlFaBkkbx6KShpyyTcI3zhLa
TPe3hwblnhE/cA5Ys5OSS1t2KWYrgU8OQKKnozQbgAut4dc1UsB71b8ICYDza9em
UpE0GpVURB+6LrZWGEX32+L7RD21LHiYy9hTuv43ndyZAejNqczR8zPO5oknDi1z
5Z93eikwS5qKqK/ZZnfIFE+wAnhn8QyGA+rkaCYT4OEzULkIvTQ93hboDHqpFgCo
v0CubQINlx7LAOZ2fhh1+Q/pMIDHO7syShemjZkbsaraOgmGKwpFRDGe/R5eAyzH
BiZGSBjU3Ybf0AzCG8Xm0Anml8qzPdHgN6Md/+DAOjFizOeYO6ac0cBoLsO78fdQ
L0gcSw3SPuM8XxYFWVsHpwHqr2jk3KZ70hE6jnEPlziSCBD/yFobIthvhImlbBgp
qDIxoQLaN7mprJzqzTUCv+pXqoB12VQz0162Gh6/zMugNkco3X+59rA2jDZDogGE
kiTJTESCwiTRZbYIQmFU7ZTkOXYXPllF4VmwHqSBohnWV6cWBTXcb0mbPhbdDA+S
+DU2UQmIggri/H7mh/IP06MeyBaVlK4o1/piXUrXY14HcTO2qQldQ7QfHh6Wtva/
wXp7nf8aL8PGuaS1uQM6cBeeGTmlABj4om+/L+xJQOcjJX6xTFDnR0RilxH4io1t
S4rUJHgTw5AXbxcTsOtP9RDi8qqldBA8hxk6wyIuvva0siPMoT28DKIh55ZgZvOb
bbCZ4KuQO28VDB9+0eKb/Xl1+dyVWH0T7JIQjdT+Sf9ifKxZowYIXxnTlb3Itl/f
zAEcpvru5WhW/O6ydv0y4/aCyxPQECmWtzfRRNWuOiCGGeTzXYyiQSmkFC4wam1M
6ZYO6phCCS5bUploohaJMZ12CV9JJUijDLZdPbdUYy5kxnJQ0/koT4oPVvWAoGDB
XNDFaR8bYdBVrKX5b8mDGm3nRmKnJT8ndl5ionQ93E4dj40NT2qPN6R/Ur+GGVG2
R7d9TSjo0vtOYYvZmTfaHkKfA0r763kATcab4/Z1v8sK34uI1Avr12dmVpXNWb6z
IKO84iYZXplu+O2lsPouqypTSsrAhtkZPCp3jfaxXvq1tUEC4JuSBs3lTKsmjB1/
Y/hN39BVVPBCWeZCVwbAL52MdacYA5jFc7VeKpo8dcvskqloHU+e/PjunXr8m531
+LuopGJs0aVP3YgrIhbPdDh6S96EVid4FikFQkiMKIYBQ3Sczy+ztvwKqip/ap1W
O3R2zxZliZ+QHUYy4LkuovJ7UBKv1lblzTwJ9i81zvxscVT0VXwUF+FFBm05oR3E
N2FKyTEkq8MDV6VKqQnyNz1v5yx4S+f1y1HlZOi82+clN5mlUcPHlWT/iCgWcclV
WEESR0hHWprCAPI1phDfBHhrV2mivl4h8HLDQ1g6q7SHdUutW9a6Caf10scaS6fS
i+9DFRY06RrR1CvYYhmY+KmaqBmpG3mZsZfquSDyhkNfOap625vkQbVkwBpUJoBw
SKfkGeHbcyetlbSaT0BXCMBMMVpDj0L88nGfclDbNUy51Y0hkLC5HSsK1tnHP5O5
VQYlMw0uIx8yg0M3MmW4DJYgSu/1sjt+aKCssbXa8OaRNE9CEQxgqq1RBUUudi4p
M5NvYL7h7SanWN1AYJe7iFN9JwivJ3/0t3sEeZUZFkT0FDDazG0JWtxeB74/Mw2h
OZvS8K3mtEH90uRMDCwfVb2EoGFLmG6T0bHq0PzVLXLm2mj01xY59MicJXReXB7I
KAEd8y8vH54uTVzcukX2ufP83dXAJH1fK8Xi/TGuAczyubKdQ1du7sLfc7SIMnfL
R11tU7hHv9NGo4OHOPSqu4xh9AXDoq601WR7LUT2Hj8pdB2jmBdHxW+L2E+yBE0s
qeI+QrvGChUiz6iXR/5AP++6fGSqoaAkTsrJkz8g6XevxnBs2uRZzZ5FjYk9Dm+a
l7IJa/nKXcKuqmwsdEAuY+yxybEwPU7hiel8MpEfqDq05KgzuS8VLnXJddqkl/Io
HIt+hbHVcKb7ymSEsyHHACtpjAjKBd7jh5AgXVQhqn5O08TeTqXdScpz0K836Bif
lD0Orh1wQBUccPd/xxPt3X8nfak59gHDrWkiu8uPHIRNp+bJFMUm0tPsNUvPiZVY
RziGgmiuvvdTQEhQYnirCR7QblWANcZf3q+fiwpBBBpUYBSmsYahPe6DTP0UdEEc
cVk3uaY28jFigRyjkJ2Tm2UN1AqhXVP5gFrVxq0dpTGSBxgJMW2VfR+xzpq1V0dS
XTySfsNmyYEC0qRcZAlEo8lqTqjR7M+O912ELx5fZTC8XfbIAllwRFeaIg/3juWX
Oa2JmndilvaLtZizlw2Jk3WVPyTWgCcStatne819VPhh4nQIq5FlMEM11vc83kWx
ph9MjKDPclIWPXEp05RDADxhpcmb08fcW7KuNxEPXr+/qJ8g8PlBnHxh+xoQCNk0
4N4y7AUoQZ6P+HGaYopRQI1mbr8hxUemVlQ2BN2aamxsIHdx36VN+TflLrDAyoPm
odCJgghR+50q3JADViJ6eLahLptb12CnNIErQ+/MXorSZDjNcEpgR4+ZH/cC4g1D
xjXf4F7uOUe+5nIQQyiDW/FTzLC+uKLnTjhLgbSvm06S3prFsC2yVQY+Y9qAkbYr
Uz2wNf3gGePzf9UPHEPqf2vr2sCCLM8Fr2B52sGWWutCnZdDttF7repHFpvo45A/
NqUJ3deQ6veBLEajykbu0uk/sSLXNE7jOZcoL84MPnQEh/9Rat5+3etrKdN12hZU
s6aspossWGsiShWEKVwfjvZ3/0aVr08SsYXZJiNYUnL8mVVXJZqQYIOvVI3DZLVW
IPRP5gJ0U+oGEfw8xOOKbivp5MsIp4/bsgiiq+3Napx1R26yiSiWlsyZVuez5N0K
0mU7HTXgqxAy8/O1zQVJPTjz0NU+BOP/ZMdJIpZjZnKsu2K1ry1YMvojYw3qBYy9
NUyhyHBhhQ+bDggAklvs/s47RIUIZ9+TDlPpzgJ40m2VdpDjD92Ks3nRZw9mvf5s
Pp+2AxvmCgBp5Jm5V70W5EteSHeMS0DHxbHSVJG6pdluOcEhsaFpnhdfetN30EQA
g8wtLTjbQdy4HtVsHZ1c0CYBdcfky9WnQYWQ66V4K34voE9ek6IzBm/GL2imEZTM
x2NGSkFl28Z9blrinZjn9mSXbE/aWBsp0Bko2d3D/uNdnXSjP0cNEv/hYE1v1eMX
467w/8afSbXHTz6VabrSiN53bBDIdqF++qvd4OD7/Pqu0SZ+q30v2lrxT52iDthz
zU1ssefsUBv3suZVv/xFn/ojAAsiqB0BzqpYlvC7lBh+Q9fX3bXjWDcUfB7g6j8Y
WTLbBuEWwU4wrZxf4PZb3y+MykDryL4vjhOVFrxI/Ho5WJQ0uRP0Y9/H94Ufzb9J
E0VkscUEZ4qp6MBvsDX0KSFVdRJStj2YFH52RKZ5IsNV8qESDwbhTY9yfzJL0Wac
9882Ip94IkisxkPm/ls2rFHbvrrdi0u2eHiQvipaOesaxRv35wIBS1r9UdBmd75Q
dqtcWc+NZU5nTS5bWWhW/t36mhXFFo+cShdPP/urJyojonvpzQFr9VTmVc+zeOc7
6VVluHz/tQq3FKa8dgcJkvKyKLyjU2rpiw2YFflxNsTp6SvzP5kmdxXh+bF1Ei3B
2Fac3waarBeOcDPmJFro1S2RvIg+LaFGJnBFkTsndkV19W9E5XU1m7dkxi30Po91
LMw5eVejSC7JNABz1o9krIqAdNAWsjiHjKH1jAdwIBljAyAleqs30N+D21TR60pp
nnmI4BRBtYSIKimXvuWBVNfaqaiQXPOQL7HhLni529MseMkzYFHLsKyJ1Ff3T2gk
46s5DwIgpGrB9V7lfspJIrJOajc9dgTUSi69wE7W3jkW31gFZiB7fvjsHwe7Ts2W
WYB96+X/0tb9Zyds/qDUxp61JEvtrrnWzmltrCmYWGLuFhEAesKL3+6kwhhRPM9G
r63j7mIvjkX8veQPz4dW29dCemPcRB5B1BNLhxWkAz7P0YKBsOhtcSrtUVYbymUy
ePnNLfRBljAcjCaKZ0/cyFcs8F292kx4ETilVltVmRn2gm/n1oBPqnGAmDFrwrmE
EqzKWR4Pq3nn7LFk1ZW6YGsxK72otlPIlOZZQgszvsl4zoP62TDm+r2QftGJbtYr
FNGPClEeGC/zR4GOWmkhejLzjetcwS67U61xsgm7fvVMEKQdEKz9j4R6UPceB8O1
bw7sWugLzUQOFZyAlGIHYCLKokS1ZRE0c/7RAGopRLnxzVhVjETWEnZncB5B23sW
y+HLkF77Ue4uECm0STDz7RXPRg/PQZha2AT+BvSUZboSahrHw1pj7NLVfNX+psPF
fKaB3rI9PsKOIyJSj7ustQRREkcUPa5uQc1ymV2g3gCmPXa46H5Je6Hici7avM2A
cjxfoUrafLLueGWSPqbMlLPMTZU3JHm/cLEcSw3voM4hhtimN2K2DCxNRolOtVL0
AYXgSaA53xwubaSJIX9Ddk2G8OgvP4vnyghSKXnJkRF9/SF+ujravNX0v67ffzhp
+v4weVbDDyp/TJm1pWg9WWkqJcYAzhprxlobyBR3j9VFztbsbXP5kwPE2Hopl0qw
w5imULYpJULBgT+pnGRI84CiuF2HXAjxu4vLM0Umy3b7Y7N+0/FNtncs/bVqs1mU
hKn7R8+k+CkPvr/QFNWDOz5F08eUx89ENvGeHnfIOhwS948fayIT7Wg8c+2/dRn8
u49n2L1tUPpuvgP82SPly6qnnX6t/aBh5Le76XJi7H6t5ddHd7ACx8q3hIro1r1c
bh/ksGhD1vz41QEnzIZ3aiexn8kuiF+qcHpuGU5OiWMOZ+WScxSQBgBEX98N5Vu7
DRmkrLkqY9VXIdkNrjxm7J+45L19Oj/yswkiJgvE+6aH/YAzGw2ePgLltWgCqhaU
eKS0aVJTvQqjLYPiz3mr7TXQj6AuBtZPzwH1+RVzXBLTKKhgfuew9BCF+4GIhoSG
tE6Hx6XKxJkKfIcSGfm+q9QjsiLmfc0xQEidWaYtTnfLQkZsaPriOcdWWwrpPOEX
E3T2PWzmwA35GdIfAQI1EVVhaHPMX83egZZQsw5rdSbmVA9unyLO3B87Hot9UmoG
TUAO7drcSw0WS+TNUwkAgm4leywdupfuwO3h4BIlwpzwZgujkBsr4GHl0ZwDYeje
V+rKapCcG4Xy2PRmqIDTg94Gcl2EUlq61+vhr55JuDZ/m8yiE3dgP3+ga1dmBHj6
2ePuS/1KSMONt3u3k7bmSYRc7w2RkmfDUjgotuk1iP97R6t0mk4baXIuoRQvZD++
xKQGJgRADq14iLdyQvVmQICS47VwVwuE2xTabKOXt+3nzm5ki+oLZ3GINgtImEJU
TarZpDc5J3gBIkVuyHfTkGNwHDEQF3bSYqiNuFIDpvYjKmVx4gnH5Kz4KhOuXkL7
snW4FSG8LR7TD8RnHHfDSLIBptcHJOrOgL6HRTFMSXAVvsN312gfAIQFHs8/1Enh
vwXya6xMYdAMZ/InMisvbARwcCmdAh2AENzeJDbeU+ViYzRnX9Dw8h4KFUdsYYUi
hWi0u6zF/ad+GGOUUDX4reQe7CNhEuvuxmmH8CROcd9uj2dYlwR9XF2UTdVVb5E3
0qhLz2MttPj6izl+9eYvJ35scWtrcgtaD1jYSpBfNzKydIJJ8FlHj0f31mjHWGLP
kpFrMi7uklLGt/Rl2bq0rLhDh9T0CDu5MspCU7UDTMcbWnP65AL/WGkSIs0PcUpn
hwYVtBDibREODfum+VXygis8inLlZsUjUxCoLdurXVyWgf7rFTof8ejgraV3Xhcz
99raPtNFEXU8KVHY5QARRoynDeg4HBZTTn20iiemq75gcgfk765v2nqwhker2xys
raNEglF3bEhtzKMHTGpxk7Wctf65qfocE+9rVHM0YSSezZtFZXHHJlLtpqwHICz6
kUUnuP6vXS03UEda1c4uLjtqe+8T78kUF9OWDipJ4i/iVReklR+EcTpod6NDMZN+
tK44JFYFInsDmKlpCuDU9aTf9V53k3cb9mrQ9DbWTnO2Trp38Hw6imycAMqPigD/
PK1BuV1MBEXIgGKv043IjvaTusTZVKezGCLH/AuTJXV0/KdN3Nmx43F2JKleOrNk
Pco/Gimm6haEn1uRfVhJKjPvRs1LU17W+CvJMj8xYObjg7zvS0ydqU1jPhBytyoq
CeQwgsGrckf4ccczfg3aO/JMQJDrshyPO4hMhTXKKxhbcrV+xzeHCfgb84mRCDdK
whl3CPjB+SDtzzY70ONcNfmgEUZEI6a9hL3MgpeLGLcOFMOLXytHVjmY5M40quD9
r2dd82bm7rdqgHHCx3A+K3lAVPjiHaljLYTHmNgAwCR4p8Ojne+eKZhbDFZWJWcQ
kX4D2J0wJqwqrg4HEvDdSFVqlg2bhP8AQFoy33gs+q5bzbx7x2FX2/R+zDa2g328
G3r3BVI0bgJMq19qjybuwAENBp76bm7t+ataowx5KK0m8jpSRBIM5q+3xyTVsw8b
iHGhX4kG0fovtYJNnqbrCBikQZjVvOoU0Ywo4dDZjjwx/lULddyLziLn9J8Yxxsn
Xb0uTVC3PhAnLS//T2YW3Ck94jzgJo59ywauLMcT+rXnnd+MGGV93SvajjixEBrl
cRVehCrGaaX/CluOeXlOqEErv+YN0sb5JvmGbfchFAQIW9jwnPOcztIOTo2UcM4d
Rz1EkipRqPLKcLXk7MVGnIiCiyHxUqU7fRIXrfyAwr2VJGz28E4howxlnMw7gqpE
RPkzJ7p2dM1WsROkhAOS5ANGdfhts9cdK3PtZYKMdpwOgtfwL2OLYGI9AaaKHbYT
N/48tT4pvWMRrpAdIp0cXDJ+q65C+4Noi66rUF5DtiKwp2cSdfmbixyy2uTSF7HM
/DQbnFzx8r0DdLaB/wK9iG8Mtm+Sja1xGDqf3mBxKRn0qjQASPqGDumUufLTPzyb
BmR95hqK9gj5WApXFjemwMM0zLuWuNcH6n8YtAh/016KDPbtmzbRBZDrFbpzCB/c
vPeFpaEaWp7yEYQdYnjR2CmEJsmXAWEJtmIYPvT+cXjYAriBp7XJpt4OX8IOojqL
+7I+HzBK/1+zwRczrXjN3Umsnwau4y/ZfZkXdAtedmEhP4p+0yabPRCprapZ5bDH
UT25uAtXCEoEcLyyAWko85CzgHVXlN53f5KczvQWAs6CJxkLsQwioIFcmX4EWOrC
XkHN8T0QCmslNr0uDTQGokobA0EsnJfUoGCakBhRjNE5GJCjd63zXRKeJy1U2u1t
HWVKNFjW5o2gUJPKcrX26gxe9fjMYUmJXsKPLPtJ2fmNxGQE0i/jM4+ECNhWayCE
Em4XOkw7DKe01kkdPnaCMUNcrO3lSp8tLDZv123eX12f00u+REfUHJRfAGl027iK
LAPZhBgi2nBfyd2QQnD3cU9VVa3H4cfCdsmVtIvZCy4YBziKlWxFs2mjQLEe9rPh
vMFTK0Eiw8ruLF/kii83nOcm4yWnciRXOIJe0JKJepcAnUm3+G94wdfH62YSKNhc
dLrEj000vV7H+WFz3yK79hpIb148xhIwFdQoH1PlWBR2pSAYZoMRK43xPY7EcUxD
39nqLkMi0qBGDjHJe+iIhgDDKX09fpGr9JRK8EdSEXE5qaI+20kjls7RyxmoZgzd
CZot1TKLjVgOHEaapGaN4RAHHxLL6oAPzfB9TSsl48CrvDsdlAv2j9SKdzQxxwCn
8X1PaQGS9XfmXLfBOsR/567TeU774nplk2eK8YSI8zA7NW6SZ1+u0BVDGwTVTtTG
kkIhvBkSTQIB0KOnzpXrW7K7xRoR4/DmRvA2RWBzKuyIjYXRipuoLBHGTGuRFqo3
AMFLc8Jn5SxnEd63jKnCP/Fm6RkHCk+2SIu1K9bHtBvQDYuEzUfOcDHRAPIuiYx1
S7Bh4u8mC1HYbapcjbTVduOZ1hVrMr73d81qBnEjclEGPKrpJOnsa2+I+QNxosoq
IxzBNae5DfVcNIJIotwwjDV4WLjvmfrzK7nMpDOWxJ7KsuULU8A7fX9UjfoXr2U8
gzPjFt6NLVZXKXqr4gnVVWd229feDRnOGByXsVIfmRQh/L4LbwKQufLcXH/QLuNF
FkZvCvCNR7REymWOyiB+F4ByKTIyCyrQK8qI5VA2dl4l2z6LKLvMojc3U9YTWNLQ
mIMHiTaO0PND56ovufCfr0Drt828vB482Il3itLuxXpsO6nGVuwoXJky/R8AL5vg
vKFFXr9nkI6+cnSOPzMg+FcGnhVBJLbjH5U6QGLgtvfVt16VDy7JL1ZU7HHHJDOP
BGGL8h3MbkTC0EMNy0lyUkyI1I4htr6ow9blWkpgVJyAIZVXpjQoFnHTB85MNNGZ
Ih5xc6apktBz46ZwEtXkqQ+LgDLLwLjQWfGfcldZU/wh680Es/czXdFNNRWOIccq
w4Ej9nN2HzMnXJH+tKwVNrcJCOoVkt5L25a4fRnNb4W88zx32OV4UYz3d+0DHZ+f
AjHJ/y8TUPNcUEQd2gPWiVe2Kg89m3CjoC1TJQrNd1DOtmPuArVx7YeoZpmHp7T7
bhogIy0iqYcfuQ0f6A3oC+U3tPKBDdfNSTIfJZioQCXZglDoNxWQaVarZFkXfQls
N8tAjKnprvqy5hzWAsr0NSFs38kGpuhGLz1ZHPO1C5KWM8fLAcY3V+d1j7Ykq6/1
l4A4OGqB6JbZhhjXdwJACXE12yyNzD354ssg3z9vX8Kc2yoyD6lSEYVnSoSEZaUb
8iOVKxbx/tYGUTRw4oo+6TYvRd2kth7DsLzTSfANmZ/X/Mngr/vpBQG3kYTfECDl
VYhbItXZ0JdPbRZGhwz5BM/8OTZEUfeu16Qrp4KNvvdNFGbEBIf736mOnIgvKvSR
Bj3PxiMNL/aETYOo8kJcVhiAcpfUS0oCGE1z5YSxpLp/bZK+/mGVB+/VVcnVuq23
h3ueQT1pOd9/H+QeZsenDN9X0NqdnCJZzZagtbJXbiR+rth9FoN/jQXuuk7Qvz53
yUtMjwWhDSL9IZF9hS1Y09HkTd/q7d0XoPIpw0fUl3hMsrN0BwQgZ6Z8Fitt3i7c
WX2+MfmqfSlwejOK4Jjv8dyYW292LFbyhESQRtlN7xVvNLf7evEc3HFQdWvRYVDV
mb/563vtYFFCuYclmhN1paYpyGOU2Qw6GKVoJZPxD6i+2NSxnxB61qJLVi2I/zLd
sMOsyb9EfdckENtvuO26KEDawtKrkcUSvjnljmu95YsVfWNNLakkRnI9r7JeeBXv
cJv5LA+0xJBWcd8B+QhUiMN4L1ZO+Z3FZqBaAPNaXJSHO2/1v+4jrrA/2NAd008L
VEHQ0PfHPKe5B5SFJolJYzU2Ah3d3+1gkSbLGbiZk4lIT9L1FbSlxXDJMwvZzx4h
+9wCyHRQjMjRtBUvavTLprH+6YGApseRcv3E5IHnX4KBIi+YEk6ZyLmjc/EQwKRf
y9zPAzsMMs/+l/YxmIBnXMO6ho3yDbK0JYplxFNRGiQ2qQzqg+PYbXHS7ILds9js
wyS8FtIwg7C9wojPIqW+3UjcxJKdvnr1zG4T5ttS4AwfgGZPE0IWDjD7j71E+zOY
OMwC19vBsfKwiI5THl+QMx+hD0lcO/ymuy1VWWrEOGVprcbpRZhi1jLfMGrvSbvr
AcQJEdFWrgaP++tu8g21PpJePVR3MZ72vOSpHF7UzzhJzAGgfokXshjf2px5ABU/
9b08b0Ksd7vwMpQ4/PhWj1Ywj1OJPyhrQQotGCCD13DWiQ3l5HmV9FE2r4VGktOv
J0MjLoWRhlfujAI/9idzrdcLI8cVTLhPbHh4vSKU23OVJ58nipLMX6IpAqq4Nyk8
alJ5aF2ofiH4aQX5p4+F2VttHQhx1GEBDnjS98Mo8q3xsg/1rfm0MZKvPxJa1cVf
LhKdBCIwfgLv8Wo2GS2MZhTiGbw9FctGq1rwQxwnC8U3qc75mqTtH93TnfQdJ/4l
eDA7VD8QF/1CN6d0TrdHgTkfhwMKEHM0KlB0qr0AW3TcUq1U+eFyI9hLW1O72ex4
CvbZxHl18FPYUFEuBigXJjyvIgcx4AOipri3IuibtliWVg02TS84zBXcoiL7MOMl
KdRZKIPYViYehvvgxrgVuWVCvhqc1LUuBEgDQ/o8R9lMcoyz/zrvOUDPX/yw5KvF
ew0Dae2b2wKOwv/bOWefzzVlVFY51t72W8x3KSJYXGif4k2WprsEOV+8wHFZusN2
o9ZNJpykHuJMh9LQ0j2jY+lYxtF++j1GR9gLjrD4SRzAldDTM5yW/8AlFMhm6jWd
TOX6XB9zK9VR9mIW+z7NgavPN+3l8sp+CNdyRZCrFYV6u/n9AuupCRPNfLAiSgHH
6R+tehRFN9BFVK3UgTPsK320UuSJIbqG5Lc2tkw50q0/8ERveUHy+ofSvP7imXkb
VCMa8YlfDcM7EY3Tt+9rKcesJOUsxMKNYodEi9LLhY0XffRHDETXlDgY+3x31aiA
yKA7NAbfOKpJR/ECv1D6baflT1UbZQdARRKqzUBE5hGqkT8ZRuFjzQ9cneWYWz3I
0QpgztNAzy600/1vfOEQvBo47wflG//PcZyLpqh/cgoWU2eD2LcdhBpQ+PoI82Iv
yyc2B5G6wK8/zWg/C/QJuTpnyDFd/0cOjdVfXZ8c3OR3acRXqfROsQOmtYkwsfE9
lVvRFmxVJFJ17bJcpBbSL5bZiJ0NHM5Q8ckyzgNbOSUZ2m5vIj0rqabWZjmiCDN6
v1opTchLOyC2JRER60jV7ewuc9lJkIX3H6NOKqpNV7HuyPBHhp1fzB3TktB0pNDQ
sReRRsIujJ8LskfcBZHhAHJH+JPZfijg08RsK8BWByNMGr2TJP0NyhajfJvnKgog
tOSI/PLs85G6w3r/2C3YqxP1IahICRrgjRUy/2M7I/H15lyboQgwmQUwJW8J8GVZ
SjgEpqUmT3w9MyShYZu8RY+Na116VxAfW0jtnmYRKab78FAHj5jfsK9i5bWXalHr
Sc8/Hw9QbN3L37ebpCsjP64YkgVi7pHkNxz84I4jR4SRUouBbUIInV5TQcPbLLA6
b0h0oSoKZbR7AFu1i2vsCPlIKOaPsQ+LMwLsyX0adGr5+wKom136HE8mR5D+6k5f
ETSrul8bg4uN2mCfB8W9mo5mo5lVyyhusS9E8V/jGpqFmVwn3RgRLIcECfFLEFoL
AOC20frcDQq/DWmmNOg9++bBTP8tarSaUCEyYKm8GwfLDeA0fPpB4S63LOCNImis
lp4Z3JKqE3SmI/lOyaCUc8PcPIdUcE4Ix/rczAgp1tABvSIDE17G8j0HV9CimAYP
wkLCY7v13lS+MPsaZqvhlNBv2IzfbNys09Igt/I5QXbtQgZtusH4ODueMuEknamY
KJAc7tEZsq5zwpcVNU201NasoCdMS6MOpDNqQrMLRRkbpYGLikBw8uAqiGkdmNiQ
8Q1TkvBRTu6GASr1Wj5bCFH8/0DzWNetSH+xjQGryrfWm6UvVkTvX0yzWEkxzzAa
LJ/z9UJ2rnL+kfZf6PnohDO3vUHSoIciCjKrHJWmBa7f1nueAkXy026dgB1YjtmC
ryHmApo0HlRgTyf9IUybsfqPDPbdOq8nVc13Sry/ze3yNGkwKWjpo9cOb0AMVl6g
CPy2Z7XJw39TwIUNh7xmjo334+HMLBfeW7wBuKQThmc5pMY8ui0AragyJbWAuz9d
nzSadxx5XDz3d2BPegPHn3PgCV7KRvDZIUFEIGhNBchoiDPDH9HjL14Ebla2tIW2
XTA1tzU7wEuJhsz+4Dqt0q/0LS7SMrrf2HB/XTFEt/sXK8Gn/vkXCvZIc4g9HuUz
1jlkWf15CLD4Om4YrrzJtXfFtnEQ+XNAFGH7OvJSExdXDyzAFakVe42xq4d5EoR1
bcOFQr6yk87AsHHnRrqaHz0FvINHE9weCrWRdhkqc7Tg8J07psYIRcSNm7oVwUm/
Oh2hsRWP/l40k7t/oK6ht9EVspCe8NL4DOmobcX/DHgcdVJcbxYk10LRwZOP8JUr
aQKRzq98GC9NWTl3IfO7nDCXAEXwvqqPZwKBmEUBUMnW+UsUHL9SRX4yPxTuUJKZ
VPdxnMx8Tts2KaUaTG4FWR+5cQrY6U9TQEJ9RwH8QCjmfc7cTZ+TgCXVfAVAyb9e
t1J+1BSOTlXSYGmDokSl9qnL7nE+2mBGk6n3Ue593iq5Ef+3bJQAHy/SW8zETC9V
LLGImHw9P9/m5k2J+3nonvXaAvhYr7MKqcf3e7jYcZ4+ZmgySf+1dWXR7Yrc+83Y
Xxrycn350y/mSLAf/8bCi5QauYrogtelDikC9Wt/hK8vlUN3HVI4tgoBjHnsnWUp
pVq4NWyAeffXfoGHa/y/a/edaxJTvHb1IA+hCm2+k68kNL7Hjnsql5yb6xfQiTuY
Ze1qlfXUPbqKFtfhOmqfEseoN44f+URGBvzp8UA0ybya6MZpxh58UnC3+0UconAf
KzymZFsG+AieDxmihlJVy7+SbRsp+X49rDNdeMn1VVi5W9YQGJ7JGs+hwamn2v5e
1O4KDzVXWpWNigN8ryDRX+y2bC0nn9mPdjaiQLR3T841Oly2mm7uoxzRDSn/uYoB
OdN2krH1Y8yhspvxANdefMGsObdnXg8Y/X3uTpE9NXRSFHsfW8EZaVtDk8nwR9P2
r6L66ioxYfAE7ynGiwpu8H0RNiz1NzaYshm7P7x1ZR1cCKo+uT/TRlgIPIQjuOEN
m/zZ5JyZ72zoTvzbMwqUfWaoNNTgMqujO6BKdrmvY3T3RRorV8mxBnWiYMsw60s9
VDcyrrVuRNx7ZKkBa7NHkHM/bbEc/fW5LHOrUiL1dSRq3ZsIMMGK7awkFriW/rUr
x+f3QzT/IhJfidPXDowMGxK4Pe82wNHx83HcXlwOwR9hFkNoSawSocmf/UNMuwSH
+4LvE8qq+pkv+5/M5F7dGkUwunkh/BSreuolemesdilzJ7YgOk+EiyJ3Kf1/Fb9R
NmLcYu4B7b3NVRsiPKS8FJ/Gsyo1C1G68FFfslDnHgjoc1ErWaytzslsPwolMEYL
s+vrjTVFX0M3SUz0SBFtf6DB6P31gKU64/gtxFjmsdhy4YKexbgMF8u6Yyl5MhNT
x4I2+yBN4QBIZtSE23sn++EIC1paTLysoFbbzMhFIBdu31RnEEZxz7QLBG0+xYR5
bu0vqFiVx/Y3aJ6NRJe1NE1ZHcRTl8FsTgac+fYyOLjLED4CchKsN2YKQUH/D8Z1
sLbKQrnjtifKObviKW6ui7H6JI/0ZEfmyncftDFyDZbqGkm0x+gMnrFoh5dHxs6l
R28gQvwp4NPNbHAvhk3gZbEMp24wrsEyCLswhzklvBM5JCKvkTHeoTiJe3LyefN+
wMjax+FKYkMQmxQ80fy5evN/YezeYNL4nqTOnHqDBq1k4CXuk4j9/lVXP8JdiYAR
g78fPhSeRuaDCR5xIdh8lSrT5SaW75n1SGYTSgtLKcN4V2rdAOZdZlAi2RtTkpas
XWsHaHXxlA0ioPWRRpLtSsaQFnsCXJZSiKr9wcO46/SxOJ6gDO++qvHCT+tiuyOA
FabP4HfjBFFoZlDT+ZEnbKfJF7jYqHyWR+3gLFwFqchiB82IeCTSYMzHmoQ+G1o8
edKssra5mFuJxV4b7rIyZaumSGUN+js0N5Z+3wFLfLEI2ctHLamtTiooL9zv9gNp
jnLe/DaPKjVXmRxsKgBpVIauFP2NnLCruzlZ/5G/hUVwUV5X37n2gpaj12WXqevB
vYkZvy8VmW4zlS/PCmp+o7XSnqhD1s75A6r+QC+RCO+0Ux6m5ymNz2tq3qfFuSwW
0o0ClghviyZwznKAxBH6XHLWIbn52u0GrXC9mvfrSYlqxgeb/7N5qGM4a/MTdtyK
rPkmqSruENQfkzUsS/OqETBm0pjSNWMbP6i2jdPm23vFUl38ZKLBXCegPj48eveA
GytY1gBqI4owz9sdWDmZyoELuRMudDEsHREdTJ4zEltBAw53zv/R4n2Mnhp7IxBD
cZrDONwWVgXhmHpIWL9lRtvxy8jonnRihbg+nKwk9SY2omtpoOlCcdOYZge0HFUZ
WDVD3Ybmc84o2HlCo0mH1cdnhUulXt/9RFDygDDw25K5qCsWYDpFEekO1VweYMlm
4qi4HqwLS0v+XLMJ9n0gMYfue0vtNVLoXuU2evK5W5lpwiwI4a9Stb0NhBXqjoMm
zFny6MpU2jhp42SkSnNagIYxFpt8Tp7KDyQdlDTm9zbLo4nABy+BsTn9NZt0f4oF
GAG7pWAFxnpi64QJYTfmZ9+1lv1dmFOdob55NN4lGHZKXodyJIJNsriVwejcNnlL
H7asNLJ/CA1fUKOq0Sa+LZgQ3+OCEddI27OxR9iHdsvUv9109hy24C4fVnqHX9PB
d5cSAk4qD86zM1O0tnK0QJ4X/+PDe+6KRpp3Q2+Na645FTKQQB3FosERoGbMWE2E
e+ED7fjGkw08TNv8No4bxigfj9s4NV6fbE85BBfOzDINpuw/xYcrPR42sjJgDmHy
D/LPCB8LrSReApLdocqbObTUqwwG8V00AZ6Id6qy4fSTe+NJ4ZgyjdRosgb1FNOz
OGRPTmu6XzljSJUnZZqFNvQkKaxbIaCPr29yjfnBuECHhooPtnEM5KdA+I4gnXgK
n0AVrABnXJ3gKcsO4gBYtQSI15wyIJqUGjwH4A7/hf1WhB8zJaEJKPh0EgTh3os6
EBxqOBDlyXBUDf0e5xkKwGn0JW+U9aoWxxw0lLZEmr8k+Wqq5VnJ8jg6hh+o6o15
R7dfHdZdasQrxHgq4fHnmwfhDSZNaBFy2W0Dj72lE6VzL5BCEjYJ7HWc6QWWn4sP
Tb1ZLC0jLO/YLCfKaq1Dmf8evecRd3TqehrWBbrpvRSxoCMXkROyp3/xXbYb/fX7
0MHdvWlwO8d7ibuoNTNXFijF7qLqZo6zqf8Dkr7sgqTjtg0AFKuhoGx53+apyp4j
HUOBGseUe7VG4Bv0l4BAt2GaMG7QUyYDErT6Gp2QX8cX4ho/V61fETonRLCrmL2L
vPRh9netYwrBgs/EqtmTIudxNdL34EaJND1MYwLdilUFVFbxZTnTYofd9FdTgtwG
hADU+wI+eyX2b8dAOK53SJB2qJjp53Ukl7y8YPPzQ+aJEvd72D75ytf0MXzikT9r
J/+7f8dlj5+DF50pL54tIdTTCLS2avAn+kIlZVfzMJpaaDhEiX7aIgap4SblUIh3
YH1Tvtc43ea5tydOkczeSEI33OULnuokPKKG1JvQ/cwyxR4QpKjwVFcfZBeP5ifj
z9VVbioLSgilgy6yCPQB/OGd3S8VOSrkLXy2tcTrMdX+8jxXsBLkrMvPWiPZs3+7
jZl30Qtgui52jjdgnDQPSLkTLRAvWh6EC1k3a+5ML2qA5/IjqfU6dfpYbvhQm0Fo
+z8doM/wDiwkwXNlWqaO2EF61kGCmLMvZ0cmxio+tkAa+Qytzeb4Ci5zPM/lQyJw
4rYr2FRr2KI7EZ+hmD6+oyZIjrIZKeBJHsjXd9cq8HkSVk1lR42o2etco3IejSjf
16Iy2VRMof+K8KULKi1zr+SDGWTvHNrKNxpdYzPu/7vNwzpg0oQMO/a+epjzycnd
a6NlphvJqXniL/MerNkUVRgEni3As51rVtSdEmcdrMqyicoPPogwSFPXA2No0A8A
onYZ1eNCsnHs+Hk+mxZ8iJwSFdTWr+4aF5Kl/ZN81BFAgR/vdJocf999CY9jhmyi
XIThDmECDO8Bdpcpp6IrXgCZ2EWyldHpD0a+mllFKAE5TWo5AIGoa5bQH1wxXLFr
49fmKYTnocoNKu/IBemftYUpkcrsJveUnZzPO6WSnKVTKMq6S/FKHzxz3JUWFvjz
vldIT0YBxqi06F7P0ybNgA7qiWgJJILaQxwO6IZN1tdlLUWUjLminFvN3LZ6sx1S
QwQg4kmohIF1O/+RXsCsApGoLUI1IZMJ2l/DZWPAJHsyA/erx67Edeua9gvxx+6s
/SxbFrVRAu6DZDLfsO1En2qwVti9hPEZFHWbD2J4Gexo/kysrmicB/iCj5Jyev35
/itMAccarO5y1rErqTGWKVsv2szme3Z1cV5fZtQxN95xAyiTBKqmScPG1JhvqL3t
F9zlhTNi2pLEbxJUxSDEflOTH076irbgOgfzBzJrbPZIq6FH1tcAbek8PYeL7tcZ
XuWM9+KIU4PTIXWRQ1RMlPQVEiVq6r1ac6n4DnOdxyTd/LY6LpXsrNGItx2v5T7g
t79KLgQO1RH/Mx28cEU/enVtSJhbObITiObgI90np0Wo07fYdxBFnlnxtWeT3YAc
ZKq0HI7YnrGDn84VhkwIYhbvUYgkb5jZG9c824ILs3BEb7oHabfwDrJrQ+lolAGC
SVuUC1joLEMD0Wy+vZEPxUGxmbTKIh9xCoE8lWnLqWx8N2Ac8nI1s0RXWA9RUxGE
6S+75OZ0uBzlOyQIFwanoov8eGz4QPn5u1VToRnHb02+sb80eEBY67zMcE2J2qwx
ZCVPzLAO9o4KoWkyt3wJBE6BhDws2hYShCh4GACM+agrLoXaPaSoWmSzpK9KZWP4
gvHZzM6fHH8YjHd2SifmSKSyGu9S+nCmOYt1N5k4b68fQBo3tCubLzELP+pqCzNW
Pd2sz8P1+ZN3ztJpOCNpyF0UjgHTFleSuSrS+WQ4/BSOmreTG/pcGKdYgB/OFBtc
dVfAudWalW0cy8dNnnoJHyq1VAqWhUdZkC2b96U/gWq876TvSQDVuIjaVfLeKKYk
JheUGUD3+EV0Zi0P0UxbX0t9kC7S5K/i0Oa89raaPHvZ4sUwYJRJskLTmoLAPMXo
ElSFVVQU9RB+QaeliZcEv2pvpSGjsT1ROxLLuhyxP+lcLYqCNPAS+iTpsTSe4tFW
zSbsJJIAwGudqN4LEiLxL6tX9S1BPkC1x385OvYuc3qqr56Llx87JGwQprNDIM6M
WAPut5tbArfQf2EtP63gAptsoTcSWm1VqL0kGV+ypfUP923rYIs/dFbndQLmnwNZ
uAn33Xnl7ry+3Sqzmxzv+NesmjQ2RJzT6/l3Rdhg0MmW/XxtEL1IGI/mNLtA6JaW
vBRa9IDHHRXVccsbcz8f0ipUmXex1H/A7JI1TYDLHEHpvSPg0VuBYOqAmhZ2gALX
2YGg7eFWgHkKdmOR5L2owPW3itK/l9qHKf03kOEfZ89AcKHeGgAq41ISpx8XkgXg
gTmEEQe0WAUuoGUquwD89UIQa/eSFFycGhIWsUd9+4sc175nZ+Le5aNbstBHoe00
gT3Iig5ARjeKTDDfuhYdm4BnQOV2XegN+5eX2L5XAMw0LxNMEwxdX7vSaO9SMd0X
TvYCtPeO76U+Q6LkBuLaJu683A+YJQcAJxxmQJy70D8dyoVxtYZdePlYeSb8rA87
DWZ43p5X1McjwOWF7/1sLmnFeaxaSWLSO8OXl9j5KZAw5nJUptwJgrg6+y/avx1P
aBmNPhHym1w0lob0QWkgU3bHRjTH1RtRoxvHoKAodMbUwVdTlROwB9PRKTLchWst
j1uy7TNg3cQKjZtoY3mnD05lBvdmP5XXtdUI29IehFLsTS4PorWGdEOZrae3XqRP
u2T6vva42ioyVAwMNiz1v04Gtwf9v8ugS1AeC7cHanGTMov9ZGTMMucB/Yd/aJwf
B/BXRWOlU/BEd/P738dpy/iN4ILzEY4ns4xR+0WQpj7fZvEG98dVPnSGO+Pt0H5V
onNPnxsHZSHdJCSeq8bJ9lcN8o5MztvxIfSStgK/e6Zi18kyxUJyew9EqHNfNnip
zKeSnEnyzOq5zuabIoYIiYb+mTGnq8l9RfkQ+Swb9uBh4fGCU1fMxmLnxkr9BGcU
IkHIPQw1KNwzdLOEj3DiGX4zm4/aIqX4QNEtdVRUEYHRm0rA9W2Fv+xbWzUSmiG+
qsqDC8w7YNvAaVEvOLEGP11UJvCv1/ov7EWo4d1gwBKktUq2Dvphql/qbNLSG65b
xFcnVvqR6uIf+zf8dTjm2qm13jYt85AdzbtBN1ufD9AfU2NOxG2Byhv7w8PLJIG+
+ctBcUxZNxjvWplPhYyQHJq73rN5yXglT9SkXMUgD5cfm/Ltzxce51nTDTTW4Obx
MP3UHRhHJz9rSlJ8CyZDMyo9RJ/syuInc92e70i8XpZ8hmAQ3vJA3u1Ii3/jogbE
8kRhCD0angO+ruwK2wyKa8qTX4NpmtWcrHa6/ieolKyteLMZ6IXCx56I2UqXZeWv
XtIkjRiI6CSu42ds6Dh1MSlXdrnNxA96kd7Qwkt4ghSjWKkYJ+83akGGfU0NTJxr
qZD2b9zP9rEzSQo9bL2Nxdf+Vr+C23UkcGP89Kl64I4NJwxVGGuCC/GH+Eyr0V8w
ARgl5zsUXkgQUYgQK8mSTq83yRaj4Uy92zdVuI3BW9I7QExCvbudLBqvW91BHm6R
X8zqEt3yD4I6hF1ZBonx8XDEvB1ZeCWWfKdlXhhoTzu7BKVyACwSvJREm+yDVgZH
iTq6k6WFAmyHmH0+c816JsmCnx2MnK8U8gDZfV47Oo6XbT8vanQm9K1GMwIGcTel
W061H7iOUsbA63yglh8KtB5V/X+9n5GTxKYUAI31oqOiDjqk9KQ0tfW4GNjttJoq
YCUBNhA4siqSEqhV+lxu3QyTA0wwGz5Kwd10cyS+y0iZmjgRqI3FaBJK+O6+xc/Q
ec3DUOpmFKEMf/bUDSWwZNpBqKnYfMmjid9QcT9N8pjJNHVCCfsgob+bwNFdtszb
K4JdZ77xhrrwZXueQcPHz9CfcY/7tpYZKSF7LoiHBQK0rrFxh5f1eau1HfiVMD72
2KUnve12g2gzLF38VO563SC9486SWrOpD/NqpIK65zr19WMHp18jREOtAyKzrSDd
hpT1MmWv9sdSyT0huz95WNRtKfg9o1zRF5xpdS8sKFbIvHvZYQyUQkLIHoYwTWXe
g6MwVJus9RFRh9Xj51FkPC5Hw+4eDdFfBow+R+UgfHXjY0w+JqmJ+MDPAziegtvH
EUvYvDMpCH3S4EKw/9LJ3AX6M/zW7L8UmZyoF6pDiichlua8MJoG+Mrj/HBOEcZ0
nJWJ1AyDFyUD+aB7HRN8GUtXoqUTV8cghDp0EsmEPUHTWFs1S0AS7joW6pmK/NhJ
LSeQlbx+VYXlDs0IvBn1GHbJ4nuu6O6hdB9osFKYgmj6OI5iEtmBG2qX+vYH1CNM
OKpd/BJ92d/38nEBbN2tyZ/zCqy7x/vgrvFA4Fs/NeUu8xyFLl14qPBAkq4ugzZm
zY/u6hGZZ4uxzx2YnK0vu3TaiJzymuTkd3A3Jalo2qNeHX9p5OiwLmylxDAKvLQ6
jZsJXw9FlG57LUcjRYmA5KEymeCDrd21F1CGqjT+veq/1gSWblNu+cSjnr1olvUd
wsyCWRQW2NDgwmuDeaHtBwv/4lO9BoLbUByxPUUOIeNHNqxY31I09VVXhsZvK6aM
l1gqyrT8Ihux2jX5ZOKKFTwGWgI5sN5p9fZsXmwmwkumzHXKF80KwzT7mlEWP9W4
p5zyOVMkRZ5oAyzGTApGWEUde5D2fayBD6BWLupGmtSpa8+2ioWjfK2SBW5sGw3d
gGy+Y8IMTIa+AEH0dawbM4RaO5t0SoIoQcvloyA0KP/a/OVf9tQc9BRArtw//WjW
DHDkZlfLSoMmrgbB+PQE03PVUINK5ZAz90MVCYBP7Nm8DEloiApLOouV4INcbSPk
rqQn9TojrsvW8zajWAV8dhpHru61bG6vjCRg8MZv3DLBO0SDyZEWsa+KLiCXjBYT
6DC5kQCxC7LFoC/ekM6EKGe9nUn8zrP7BqNRm2LokHgETtsv62q3jtOL8v+CFBLq
SvMItn0tC8XpPzalAjSjr2W+c7RijkFn3OZjAu21pIU7abSjwvAh1k3u2IYCdu1h
Uc3JEbkTzgepsavNaxKGIw/JqrYgHA/uR60tYgk2tUjstT1jU156OeHowT9vRqE+
75F2EJDeTfWB8qZ/WzwxV8MhW05p+mqAKiY1gN3DWPKcjdPN2+ft/nAimetq3bDn
wiysUzxht4sQN2SwvKhQZGfqN0if1c/DYX9XupV8xJ7ndmLkWbRPgD5RRE9Y8Oli
V2vArYOqFJ1HblR5xztgkyOqTAW3PBKGLUzP9RcAF97r8H/BZpTfGsI2ZC+fhi2k
zY5DPUKKFQYBIr+wHFUmV+tdhrZIazJlaOy9K9+ns4xzeAgGkOcPviIko4jk5YOc
5Y2TIxcakolOHqwoKOZk19Gil/WB0pf395fl/+pEwaQtpZ2InCStx1Dsmio/A/7w
Jcj2M2FgQPk9WnwY+wA4dUTmNcmN4kekSVAjvG5+1aeUkYgcPDazKb9hcT9pE0w0
p2LtXzxd3ms7RgNkDg1EzCU56cxGcsKneeB+Ow5syb87XCeL+H84ikcPOSTHxUs+
GDKGvEtIi7jHdkLQwydsde+zdx8Es5sUDCR+8A5o2Hi8Z3K7xLlfi3VXyVDu5b9o
1JiTDRJXpnlL3cLb83cZO6gSRa518zY3oIpY4k9uYvPBNXwhCGSiAvHBvDic99k4
Fr/nPcKCXBeRfrnvdLU7b6vI8/dsMVZve50OytsLVrNb2fsaI5ztu8bYtX0iCcub
fNNgMhW0nSmB87ieMWa74g5Ynt/RCaXQIVeRVPOP6kPfQeb9QXFHxx9MHdud5sXp
9w8mYHrNZPP1daBGsun5tO6Gffq505kh40T/coV0bavscH0oCzDTCtf0jnUGzhXx
UDuzZJK6bRB6ZeENooh7ykk0ignnuz1+IpHJyQjx0Yt6860hATuU0+jqjsztOGae
hn9BsvCm2mcxIUvcQdMm5jP21gSWR5kzwBteJrSQ19hDELx2XZnBMh31POvY/9qj
AMUZ7hsS7AOLskr+RWA5xU6kri8YKzGsgyvoE+HF/65wVEY9OZhyL9HuMcl7kUa6
/y7NDcRs2uDjwrVtETOTcKa5WlRoV9xoxupT8ipeJgJzSnCxyVG2DG9kdBw4psoq
7YVSZ2PhPVfvjCktAT5Dci2pgMbHQ2FBXR8oLln5myFuwUDb3jXeRcf/+EArvBoE
kHYm6z/U6QNQ3C/BH8beDBs/6bbDkAuPT52NtHTojnt6VAFDcbzDUFyV/Ue1JW2B
16/pf34yBxwI7ORLgTbVBrR8DVdOZFySOVwuFzIYDR9relOM4NctOEK2OKFxnN7O
+ZgzYPE9e48e8FBA1tdWQoeakVvTYvDaIfQYI1QRP+2LkbFdPGHoZVf1h4r+GIwC
T+bU1ZFGieFB659SOsOi+RSSHCa7smqLwYWQtzb0ED60nT0lIFtrm2RSEbha0F9V
6+epWONrXhHu0X/0MuNGDWFL8yIPcEnN0SULdRmMD28zCHkcSqa3Kukm6EHErUwM
B/HxVHPXxMLPZu1xxEquW6iTcqy/mNcNmbM7YpULSxkYO00ZWuEQIlyGs7cElDhd
sQ2QjhVrSOSf1L7uBB22ZlTRT6Y2yGRvrdVAt3yENiC0CVU/9IPU/B0xhiBTsBOt
hlGmCSTd6TAJVlqzUBbgDYkKSvxOBwcVtJmRYrnTueomyer37qqFa1OA0gTuLKxR
gVbEAqMDcKhuAnS9BM69NtARGd05WTlrKO+DhyR3SOKDLfp6dC9i+J1s1xLvnXjB
ycPFKCZ3kfruy1T7o5Do+LLHAXDx94s0wSF3cz6j0VtcbqZ2psVMFBjUI6SCPEDY
zYpRVil7kB4GeuDR8jgvN/dPOnBu4w72xieu8c0cwy69i2a3vT6lrJTJG3fPaubp
ZgM33cY8n2nce8nzNTzgVDFB5/h9FMvJmCWw28SsICKKb/90214vdMOE0i1dNVrb
qirG414JECWrcXX3EwE5HwCscTf/Y8oWDP1BpNdr3BO6oomUGR3qUoc1eKYX3g45
7dQTV/ddihF+0CXvvWccYAUetdlplvmhp0yQyIxEg9TauozytGgYQy/p6Lp0dHHw
4de18a0iT2fVHb6ChmQauXBo62RFq6vaI000G9OUSOK77I8OqkHaPAQndmTX9aMF
umcdIEh2ebTOEW82MK6mrgmi/J12HDu8HUZFNxlNxPKzLy5oS+zVXgCVeFoYjhJD
vgUBaYD96CeVFPeKvCHjjx4/6xTQ92Aq9upSWMVEqPtQv+nQzSP2DZq9rIbZIHP7
3uvch484hZA34XgOLkQTCbyaEDmwwQqlYOFSW3idUDBzFR/G9oeS/Hdn31rDBhky
73+gOV+GcmDZDiHi9CPrZPXtFAobj08kO+2qHNwqVjBvbE/tuSKvv7sNRb7mgPq/
InFPU5zWFwykCNUcBWgs9ldnAgr0NM4nL7C4+7s0odl4kippQOFMoaP2+hqocpy6
aFzLY5etdgvCoDQSajlV2HyyP4/ApvX3WmAgbGSbr0859X3Sn/nDrLS/wMn3Kw/V
yF7I6++9rx4Go702yZr+MxRoQY9xgX62KBQlphVekVakUK9vy0f7CQu8q83cKDOV
i14ZMdBaAYWRox5/5otHA5RcTOeotzpqFNgf5pobBu4neBAWojc5tlaNPx5fvCR/
2rdRSOGAFeRvms9E9tDBRKw25WwGPU294VatrmJKixJqWAF95pbjNO5xwpUkeg2w
Xx6KA51/XhiGwU70A/v69+iTG8iY1iGyV/w8x9h4hxkiq3JCFKxJw1n4vB883G2/
DZhrDead4AO/5EysnjvUStN7j8d8Tdi6/Et9MvbKHFl+1mqV3dTTCNrzjbcKxk8D
W71c17xs4qJsAKF2U9bE1x3jJjDfb7uleP1hDVty9hVakL2L7+QPPoHsgOfMJdNO
NmEHyNzhefebCXBWQEriuU0s/i0FxSDNcWB52ypO7z0jUeFqSgvm4eFKSSQfK+6F
+On34KQWuKvM9Oht/8hRpBDMBP+hoCZixhHOaDLwScK2pX6BLvqsSBYDdG+oSIko
XBjrCn2BU9Bw0kpfSs7gt+H45slygnOnmCMtPIx132JhmuhC/8R9Zv59/ycNqGwf
Y50jWid2MJZH+3a8q+wbKN/hAwpEeZvnI+R+C27lsLH/P1LDxDEu9RsDWdJ4iMMy
dwmWr8gFj1QYxSkM2rFHxKyQgpX3S/mlgZyYuG62I9Fzql1bzMR2GTMBAUW4Xvwq
JVivlyOgvVb3hIm8ixUhK2hOixYMvSov9cf2b2QwEve6bru+vHSBxMZ/yIlbbGLZ
icNbiVeUIBMAeY5LGV0pIMA5xsPJiggHXq1nkeTVqJCNsIrOxcaKwpdXWb0YqwKv
i1FCUEiO9lOlu6IS11NO/8QSQ+cIWr1Rj+A6sIsTGYJtrUghoCZ2hrhQ8/Cm9o3i
mdKQQiqhAsBUsmLBS0Gh3X9OC/ckMUymvCTAefe3OoVpxokhFAINaT2Z9Pv6sStU
C2VWlmVSmlx/wW/SPgzjxSZZ84euW5FNSuaY3pdBkfNtspScdhJxW30WkJEXloQb
6qZ1HL4YQBv4natXBNhWlh8O2Z31ctVOEh89mSzJCe5Let7tQvOk3lERpJ/zrVXD
1c9FA0SqP+f/n8f6oEE9BCMqOVh6U284qcEoLNPWgCo/TixZP0V08Lb4WIM0CXg0
tXnSbfOA/c368sE0r2go8J4BYb+8GtRZW3SGEFblFKcJ14Wv4owB/Cz4suhldxDb
ZyXdlRJchQaB/RNiWUyNV9e1kI0yLy4PZQZTJbrAweJwDcaEoZKUdZBRXrSxMs7g
ZCrn67AqJOALhLvrdm76wMXNn7eOdXryoLmWsT2Dv/6B+M6DmantmyMIsRjceG4E
sDBXy/KBvBJ1sCY+mdJZXJ29Y37O5Clvm+Cakj/v7EGq61f0rUDR7XYPHoR0/hjh
JOO7Qlugwma+4K7YGDFvbqLJ/R0JjWrcurpGwg3gHMmmajAGlzaSWegc+50gINi0
7s1HjQznxg2S98Qw8LjVO5NvLn0gl3xxzolVIzik+R+OMXqg6y63yzxeVVoOKtGj
0E5KfyLjHAwU/IQpN6ifFGx3cIQcajfSRTFloCx8ipG7yWgmIyX8xpwS3x+73I44
xnTHC0fvL4LQOzykR9dm0fNQKkBuJwIpg7ZBK4yCjK8ZvC41gGyJsnW1MwVSIZIw
C7NB3pjfRbGG98n4TtPzgxWIfZAFnta0gFgcR+XiqUBWfmEzpD0Aqy4WqDijfOvU
C35bz3C5ynoMgFIzL/fqh+IiH2ROzKBtgVTkxPuTJ4W7QwTGxVFxzIMmtBnUs3qa
jAH6bmg8dAyu8t4lLYEd6Uu5APz7ETpjCAdJWy18wuadJ0GHTiUOMZD6JQP7KYvw
6+tBSNT82u6pI3xG+9JL21xyiS2qWjygMDn0It/clKR1z7690ZvMd7pzVX7FY/TQ
Didly3T1sSN1iVRoQuHtMngRUXP6efQzztF+vERumO1ScSA/61mvxdf4JRFl/MEJ
G+KpBpDXXGS1jk47QamM98EP9Zug9BKH7pfHCbCCsjgpseP48JTfIIJ54BcRJur/
grR5lDUieTvFTsR4yPmteCllBN4LbHZzz7br3TQ/g7a9t0wxfh0tAxEJgydUooZq
EhvFBTqIHfrylDmIu4bAVrHf4AqYCgm0M8M5NANHUlO4dn6x5BbhSl4nbiPegwTA
0n+y5VD4mNcwBp3Xmrersd2XOfPVCtMAL9xFNFPMVlMKgZ0VHcKJfmgSoMH4x3Uh
nwNcNJ11GWZBH2NNaDV3I19Wt7j53+pQH7WXsA4czgpBV2BlNs+y3MsQLcvcg6vR
oZVx09YjX7+n4Gsg0K7fSESIFceTbSb+P8i/CNkoRmgQa0pYZ06aQ612Vts7YVaX
oJCCQJcvFaehx4TTPxpYj1uBpibqdr73F9aCmWD0k/icLxDYkvko+uqv6fNNUHA5
LsFVC65Ca+RmBjDWSFUSLLJ7wF9SDZsNrUBQkQWDWXyhPmjMG8EOMnsN9M4nucRC
h/+dXDE8TTksHeqdROe88EpZGQF2Xllxqi4wiXQh/8/HnORDvb3fKVFTjqaVF1Ut
905SeOhB049TGnCBfreJOdrI8YbG7KOHif/6MkKEsydtP4SVtOpD5LYMBss2hbnA
lRixRpLTx1prb0LhC/sEIZyE6/UdlIc04OpOechBlItm/Mna7vvzdOcz1Fg8BVnq
KynxIah/thzD4cilPW08WCJQn64KVWq0kRvi3+Xx2I36BbOaFNoA7mtHaZgrpOOq
Set2rbOfn/n+9/pOEFE46AoP2wkM4dD8KBU0rSgFNmnpQeo10qIQgjuZgcBSsJzj
MduoKeMlkyBvUOQkiURyCw6Tcgz/K61V7kWv1gbuJp17h5XreCwBVlLA8ryNtFk8
eyxJQYWykXgIk00CinAC6QqiYkQe0y+JQGvp1qCWmxI6CTztVzLwI7F/bvCOxae3
n3rWCUEcHepL3CB5RlmjOS/56xc7GltAvM1O8DFefE6bL6M/oayrZ+yf59n/wMwB
WDNTz2ltZXWI267kMfI5XAgGLFRxBsDtWQRuoiHEVaC6t1EySyu2VLupGB04PsmW
0ggS6W48V1X+RTA4JpU7JlvECrx1Es0TWGqrIs2MWqdWgg2UL4pfBy1gxDtgkV7Z
qQK/i/pRWl0SlUvGBD/BLn3npetxCMh81NWTogI3KE5aWTVnTcJHGG83lGsP3TYy
bgEXb/SAsNcjIljGVfvf8cjTKIw1T/lcXdwaHuyV0FUptQnnIUL/VwGhq5FCc7al
3hh6qsrzpYMItF/Qpt2fuo/tN5IVFVvRIUA3NHKYeqDrsWeFGk7dqkxx1KnxOPNU
tslNf+KtiMAUJisL2RsVTK3/jyl3MAKMbUPWfndmiYrbp0lULhr8kEvdtPv55yPY
SUPOixBNi6OW15KDYfpxN56qH5VJUh8ylRyjQjhpASv3kwZrdnVtLrJnTHSART7K
Cf9YQNHvGLENFR42jWm7nOo8UZQqf+NPFR5CJ/sgiLMJqosi2j2HTZrc0MWdzFJR
mHAextvai33GdNI1mPnaOcjRe+XfpwJXTacf1J9bLNCcjiDjpzc2tJ3O/mhwp0O8
6ADlheSk9mySN8tK6/ESWLTkrGsKjlyRDA2/Euoo8U8kUf0JSjxCOyhnM1ZN9Xo3
plmkluZpu/Dx1iVR4+ZHcTDXXtkb2xuTqvfI1Z2XubtgsFIT0N0hqH8WrwirrORg
sR0pTe6UFc+ItqE2Ess3LGB8JFFP88rewAOFDeSY7NoG4eXOf8fCX8GOExB6wmMu
hYfMShjLzz2/uZ2rpe/HePK/2/Qaxv8+XdSAjozwLVG1lryy6UxkbG6Gni1eFp6J
7m6FMqftvWBTqnnxzvtXOuhfm+AJScHQZmWzJx6xYrsInB4V2B+eCCo9ZCgS6FTf
iH2RyhCD9vwiTEBdABo4o1G9AudsJb209cjZEylZk7M9xQiYwqtF+AGWI8tJnF7D
PKtMM8yaq4Qucnc4ypQV8tCa+dBW11V/vQdN7kphbkUyL1iSB2GIBa/qQzNdettW
hTkm+ZjdxJMDLlZiK8Ce91UXWr/jjMQSfKALHyyXOaIHK+UKEeRB+UA//cZ35zgy
gDx39IG1EwkKBy81frXQ46t8HyuFDIGqifMgo1MxQRL7s/s+sCC1klPRH57uN+xt
zowEJytfPYZNwxWwnDi2v3JsjQ8274auAsdN4VGsij18e7pKs1nF2/4sT5Tn8uM9
7Bok7JC/kcDaBXI2ekG/ZmT593PGZUM0wsuUfpPSj/7HWDuXg28e3p/bPas9uFk7
V0rbVd8WzT899W92XlDHEOm6wCTVAmJzSTe78UnUOpx9aVf1BB6FoyxfrZh56i46
JHj2Ruo1/kSpXKzCu9ZWr+gjCH7W7xBmtI2ldf2UmJ7Krutn4Txx3N12LS2KJO2I
tSmYyIvurE7QZI1bNW9ts/qQxNvlFVAd1D1xx+hhhoyS+JYHu50AlDg/HPO8ct1X
8SDiggBX6RnxgEosfIZ4KmzlqeVYMwU3/U5ukcljc/Ag5G0V1CaydupIrjD/qN5x
M17ta8JghZV2FJbUY3V2XKVnVrLtKKEp/333vi+B1FDleRSgzJOu1C/I7jHM1/+1
LBgJ5Mm9moH4HUBY2SLoYE8Vl6Drw2RtyynFcasXVEngB3jRFi3g80raxMOAt/v5
c2/5fsVoyZwb07I5tV0caBiNv/Yr8z0uVCuJBsMZbj+jvKmqoiSnHpHtYvJBLokw
r0CyZith67y7Xd1zZHMPiJqGO2sN6Cy1heMYzt9qJID4hO9QsPrFrvgYE0CnM9SE
dl16yZFEeFY8f+0XzOoJYjAqRLQ0SomCbg0qrOaAI+8l/V+WwPI/jd6aCnLt/jHM
Oo6IjuZvjz6BK6ReraeEyRUD9/8L72iJBU+QDM6sVeWyx86h/wasx5g3YEiouMIC
ElQUUcj7CpWUiOt7AZCom36cczieC7ATeAm/ui0GaH5XxEly5GPjxDtDdwfuYRKC
YWHqd11qT9f7sH0o0n1ecOHl8nq5XPccEOWRnuJ6duhLYVpKInMAnj8Xrmqo+2Er
8bQmI32dgpXJCNfBi25DGgEOqsps+SaHMEvhdGklSCZnEWQc/DLEBzwwy9G4ScvU
kqkffnoZrOIJ8vrmthapoYkn041dqwXkCz/nlEKr0YZkFS38joBh8VxnDc7YkOEf
8GYHD7AhXWpR5PajBNiZlwAO9aOIYM/ScbgIFPifZ8FFU1aJRmGFq8aH24Sm9Vn3
JlkDfrmepx9s0mL87qhd6ionQIlRblT7GSdpKEiKu989L28etkWt3bBYcgEcFT3T
6fVk4lZ1D+S0mZiKGELe9T1VAvN6U54J1BeABS5YT3m43QHZ5f5pGyQUjKq8J47b
6q1maPi59a21yi0Fky0hRakKbkyMDHO79dEikh6LmoIDZKlma9P/Bhs7I0SeS2PS
oekRyR6xImhGVg+RuMqgRf590ujigWMUQ2REJ/p51JBDN8X6yo9qGFRBoOeaFYos
AcLYjnvmF24SkyuzGXnZd+AE8/42Wrv747zOEt8clygEDPjYpf30Bq6CCU5ufsod
G+Z+wVX440NNv6vMGLZiGvWos6mYIXhlZcoFYgEO1W5qgB7ZDM2tuV2B9pekpN+n
TYK4/549gTdNETGL2mdRBCyFvQ9eLWNw3+JaB2Mr6mQVQkHB5tQRl/l0aPH2oRtt
ZTUGlwS4qH5+/QuZrQjiGwsJXKqTEuur5Bxto+22kPQvtJRZ867JCg3/s6uHrFLg
rxBtLCX5/tM1v7FDzjfROVlXcAosr6bC7Kc++yQSFc4GL6YzmxSuE2nd4SurhlsB
2xdnNcZWIALObL7Z0cVR9MJO/cD+oXrTmABZHwvVxAR+v1SIBDjw9HV+T0WbuFwC
WKj4/zIvu8lj2US8cspwo6ulOPLo+2cSKUe/DCn/X9fdbbFpL6SEcyVJkHv+bClQ
OuhCvD+qaOl2l+Ntxlmbd7n0FdYtCtR20pNQLVsoihjCoZLX11JHgnwqB5PAZrd1
AfpiQFAxW46XO+UxwIB9e5zqZG8p3WJB9aDrc+iG1arIZ1U6Nm6+Hwg44+seU4Ju
EKFp9OHN5/Ul3EIpXB9PhY13/dC+DYiuEcZXv0xV5Oq3kHTJjWIdn3peraiGnGr8
xDS1UNRlIn78/zvo6R0E/mrjT7wMbNQk+Kt3KcFnXkm04LECqbGb5iUHQWfe3HTW
aQCNzFXxM0Q46tp8TTvBwJNFZ5tM0tu/XZpTytHxyr4wl6krWCbnj1uA14m0IPdy
71F5jaYbk6m5SF5TkP2f4p0/SdFRn1ZvvAsw9XOjWaBvmc6H5X6KTVNecQCft48a
OTmxTuHlYegdjlr+kJC8LElU5kvtk4kqOB69aHewTCAAekLabPrDGBsn7CB+OU3Q
hKbIICvwLaeRj4Un4JF9IAJ7VXY/hrMRj2Ij66MaRCvbIIUnZU0BiU0s7HXqGlw8
LcfkNdWaGsZOf4qx6SAvSWbF+vgu97rlO0NzctFcDcR/eRBbE1/XqNXBHyGctnim
S2uAP/9DB9tvawwL0Oyt58ddgAOccR13stVagIjbdV0iI7mOY7IH8egm6NFL/2V4
NnQHt6pNj01qGqi2rd53LgKhHOD0uvY/WH8mcqY/goZS9eICm8AIwQ1PaeObcFGi
RDpDDIBEBhupLIz2yxsQFEN0dIhqnux9dfuz5PChrL8dnFjHEjBlPju4bWzyimWt
vFCkZR6pltHciipVQGcEOf7Cpz+nn/upV80OoobLxdVibufzq3emaxJUhDB39SNK
MjDLZWLxujrqFMu+9k9upwSN2URRJ1LfcO3dcgi2CYD0OgQoWiTX3CPeuyoI+ZOC
jaUbExTS9n1B4vvlQdnUT15zoNqYPtnlAXOSONJI47guxj41ZL/BXuisfyknJajr
E345SrsEwG49ZNnUeBCFCQ3tFS7ZP1cItHGJHAAcd/yFrYdF69sW874rX1vh9ro+
4RN9MuK/gj3Z07Ko0cdAIDz5Y3cDWk80uPabv8gylAiarjK1CqHgreWA19+buuX5
f+X7sf0WAjTUfz4aF8LsXq7yPhEdODTfqA5Gbd7fz0l2XUqZ+O73PWCgZqYzouUi
coQfdD9QIkuy4Sso53B4lz0cnagBAeC5wHEyFifGWje46RlkGRzMnKtyIE1TnJpe
6YauhxJppwS7/+W2NTuAz17DKELCNWri8dWOTFmvRXsD4yVA+EwmUe9HV9WbbWB7
04JQhJ/QcPDIyhkvH+E05B0sbLEnnv/SDhgBuQXphGwNQbUeGCdkjJzm7KhqiBYo
C/L+1uRLnHopGF5mFbVzzGkZ7liIj/+14+cZruGPrwSCk5w0s2KYZy9z2Adgu0ha
ApqeiLadHwY61GrbMB97Y539kvQ5kw4FEmWTOgJbhcSwgihVygJdAHl13qvVoSco
qg25LTNHTPQJOA+Q+UfsA0Zc8NyuhXmLsmv6KbOrNzoD+XJkVqAwAfV+5lzU6YTM
QDkmtQnizudnIGxAOWkiGL1muhsh9wLmbsRkP0aFxzQo13Pp33kKFfza3xsukobB
cz+6j+V4j3Ln+OWACd2b8Q2jLeiMF4lpZb6pbLHTRQYt6K1KI0yOFQdrjzIWErTh
mb5K21csiC6zVr+LItRUB+avjP2DmvwcIok0ZuiE5fCySHgLgYQ+AGTJAg4OUF9I
bmkizwT23VTA1pMU0L3I8BO0zi4kB4hlLxdbg6Qoh8rKo5+fiiL3rJDRNPxI7FV/
h/vAUxAOaDtqbZiJZXGPQ0lxMUJW0UsWvF5YinIQmz3ToxJfS9oICw23/9Tpgy9Q
jI8b3oH9c0T/Et5Rtie3cuxMKN/GLj7c8fXvftbsLrm0Yy8I/4a2Vu53Sv26uTDi
I3vrQrbq2B8qyi51MVWin+S7aE40QIrgwaOjlsmYeQxMx9Gsz4upJZvQDosiq1Ho
UyNZR6gYo3tyDI3WmW5qxhJrgURnp6QanKceEhQiDnHD47iGkjzrHNhWbf9A7gzy
2Gh2neR6hOi4XJATTC9WMyireBWfvPKZRNIEEKZxH7QU+MAb/APjUWDGEsvLqJBb
Pjto067VtntrtBwgI9X/0iB1DwlAaHe17RhDa22ii10/16DPMlTIq7RVpANc8bh4
3iS2IiDyBG5EQqXVVqnU3iZzNFKGGUBx04ZBTBQ8IouGAVZjhX4zpkkeDQtS0Kg9
GRy5zviMiZmQFs8rSNAdaW/7d4udQMc69We0GkPDO8woIjihgd1GrsB9pcCyBnln
w4wnkB9ahKz2/2++1sXwouShyK7d3gJjw9Q2cMMbN80a0NAnKFZhu3KORcGQP9d8
dntDVoPB/ku7DXw2qU+v7UkIwDT5bwVf+2ZJLww9capdITmpapDY27yfCJNdVODA
WKLj4tVYxAfb3ZMjJRQG+eXSOUy7DvibV+tE6jXhjHkIiDN2xFHa3JFEiMTjfNq9
eezQXEkCHNn9NMYjtinfPNxLUJNaO/OvDyE7Pjj583ytBPTvPh6zCv/AjUSjaJqs
hGJOVyklvigKbvEl1m5oZy3TGx+8JQw+7qhQrSy2Or2UuitEXpWdS5EaFpRpX9OA
e93k6P7aZZvj16lPC1dF7Isq0h0SlUtJb0BrUsc71ieca/FAfvmqhfczLBeV4nQC
Cff/krDbOb3EuG2SHLXC3gyZh8FCn8K6WlaERVdjk9h3pQOkBkn9yVpoiPiLz3rU
OYps4eeyvH4qBr+qfZEi6fFxBC39y6CmxM9s9oTmoDndfRv/dvNmqOkg8Tv7iZrI
sn3vLOmLNtFp6fKp/EMvlwD58I9IsWP35Ap7RpSZLOJWva/nziIZrP4c8hRvWXRk
Aq+bi36MjAZ2u9W9CuWEDKoi6hTTYSAt5cEBIx4ytoDw9FdTEMH+n+TBg2bb+K7B
a2boy5CBOMel/tiwCZjRQHA3GT+RnB3I491T/YrwxeQpNTPcvBN+lzp/x9dZl3El
eRm+jcqPfOib4WtOjwxTkxCE/LnxNmn4o4zWYLkxgpJP9cvP/RzqU1dAPSeSr0oN
4nUBcDcwatJXty+Ufh5+Lrp8247d+HXEINSQx8G1ybbS0u4//6+7QuwlGJ99N88g
9s3Rj0/fnFYQ9hJz12jfjUQIkkLC3spCqhXupQiGJtE8vs3z5b/2iVzV2mHgpqG/
9YJW7q46V3m5ATiGP4FAkHbrOoxvfpopqzlLqWJ0V4/h492+cpuEGBv9CMn7EVOm
4Mq0EMALBfyMJl5XrvaX3ushLEJbOMoqerdAT+9QW56JSMXkm8uhAkFwAE8zc+9y
F74/l9CbVXMvgaqI2D6QV2et0uVo78+QJ5Cv+KaPT4XueAK3ZSr/Tp7hJkKqXLJd
JqQCUfl+EjWfdSVq3L5fdA8vz7nnv0x0yIFuUJ9sRNAGTQSlKmHN9sVWd7ggQSbj
wVmGRkWhH3TmSKJNhPOFG9FkUiGsWBoAbrNUlWZE3Xm5oACm6WPVnyXGlAKVoZR7
WxPF7SHQvcPcmnWKbAYACCn8pgHfOcDpYFQ4Ea7YfBCpLUgAc8MD7sRWBa+rbfZ7
d0BvPEXl1pCDHz0CcSQgUJG0GncJAGroiarIY+ycLLS5E1RAid6TojlWox3ZY+eZ
Kp3MVqfDbVZkxUmYq6YRCnC02MaRtzdY5Qw4oBPepb+gJdG2P3PJuirY4R2zF+iE
KzDrzSkQDnfiheWzRMBBzb3hUZaUpou/96mqM9tD3OZJNGtR9FbAVTwuCFK3rRht
XyamXVJkqJkJpHRN4n5DeGoWvr6LNMZNUoW/aAjGFKra5ATsaTCpZ2qYLFBvZKLL
1K4rhrizEP5QoVccFmqIhs33qEk8FYdvSeCSwnl0TWYFpnkptgvvTZj3KoOYd/d1
E280hEwjLZthvmJg/DOeVpVw9cosG21NFiqaCrDGXOPThkEHBVNkFNVTPZIrkAg7
MifToAb6Zu2W7HPnrbmHIipUc3k34DzWQDl+dSc7l88ZuXggDPyXVTmrEI4IVMCZ
XyZzKRMLThtJLrlPRJyG3UZ0s4fHX4HK/4NSSbl9Fot3YylI66t1+BbXn4xCOQiQ
0BU5Y8+xEz06s/QGY3acilZFJWqJcOD9Sb7TPrbWER8pcXTvFEM0fW6UkpEOOuF2
VfVN/e1NeLmCbDnwWwSSqI7PpiKmgUL0iOEBFfiruDgs42WcsqRw2AHXXamjcVBu
iRUJwjP5uB64/iTTMNk0rtPaxy4U79uwmL8sF+DbTUz8C/EVDn+tE/lyrlA9vG3y
biH4C27pRx0ncOE0rFAGN2CBe3s3Wkdbgqov/LyOa8pQLx474vjyff7aTXrgZxJA
E9KHqZp/FdvW6MBRyKX2+YgA0iLQ/quc2l3SfqsHY9sh+ye8/l119oynoA+Jrz94
OtZNB327t2NE5vXNDPHiK8pKXZlm38Oool8np6olXh6W1aYmiHsD4mr3cOoWNxbM
rIwfSRgTiwXOlmj81QcxQRVgPJazVfWdAa+QLDUIplgSirCYfB5qkDGfiPuZQoeh
WJPEYNPkSriIC3B1S7P/GdOofOAIt2VqAnQGYVHY+wjPtqG0J0B7OipudE2fb3eM
ez4MfMNKArqMrX/AxINIYKi+9WkwCqC4hMNwBNSp9wlmC0cSDW1xkn4WTtXy0iIc
uKg5u8I6b3QECZD6zmD7JNmDXTShD0Tg+ySGbmrNH1m/RZq+1CWGWECaSAzqoQdT
3djgPkRJCra3TcbEiOy4ZQjjobNt+443P9eWHuidXwHr3sqNncCqklrmblGZCgbu
cKxF1TdMV0aSVW+04+1MV0/E9nItPE9dXwO21woltIa8b9SDir+nhbXp3z9FXmlE
WmlVoOLnEY+V7X46L85Il2YqAEESx83IpPY30J/RFxKJZGAVMGdhIl7Pe2WIwRVX
jdfVeafLGPyVvZLmQ55jPAV8oPdywrnveY7Lml0NdTqUtzabb6OfDfLDKiRYAJYH
+UpDNCGDFex/rRf6Dop1OWew2sRYqGqBNrpxBJ8zleQPNHJxgJLRjdSHLC0eVV15
beKHByUEESUJa+Jef6dm9KLWB/yK9bXgJVYDPaRdgVL6565to6v9emGQ/2Ny3w5s
RHNmfUAwagGd8oBL52uXJysN8WxFIffKk9VnMoMcI1A6MXRg+EETpXMZk60oTNN0
1LndP3jBeW85G1IoZ8tMt88STN3QXO/aOw4+4CZcZeLc405NalMgBCgkPerMdxSN
ZJR+PLv2Aoh0V3wSzHLZn1Ea3sK3ns93N/OOjpNC5BdLC56J6pe73tgHcE0fL/UQ
/yUSe/GS1MoWRXExJC7Q4YeLPV01wDdE4eIIv8r7OBvPSiKGEgYQoUwKdc7Za4hf
ElW8cotTM5GsV2YpVkQDqXZruPUskcJFc0CAKNF7fDpYNn+9gWvZPq7dJUZacs5/
kVbtDSBuWYIUSCsAT9crBZIy1El2ASvvyZ4Yl6bYkL6FicLbTGIjA80+bIfwM8DQ
bgnrorPNU7H9DS2MQz7Axa7X51nUKFZ3My2lXdImhcADRZcSkjb1Wbnl0kAJB5JV
SI5ilqXyQD4L8jHVOtb2+N61Yzo0kl9uxuycgdv5B+kHRHKUCZhs30phQ+zTEaKw
dTQwhWGGDohBBUa7vb6hb7P5a6k2pD1ioKyK6nwwS0hqpTOQuk3hQAxfj6UzguVX
zksYmcsIpVk3+/GPNl6pw1d2ezfmymneMmpXgqwuwI2Su7ettPwCellS0OpRa2rA
vjlNgbNBClUy+Dslm0yEEe23HVRXtWF102E6L+gsUR2O2JEtghWwFbxwU23T0zlp
jdLrTDFhiFJzEe+37BQwiWeXZvauVVBzSAc5gk82AseSdbQS9wC81r+PVzMc5zm1
OgdGWMzd9gEucps6eRcoWVGs/NNZu9sd035XAPJR47Cp/gykatiWqYkb6gbATaxv
mT5HM10INXBudN9sL/Z+7tbxA75yT8x9FO+zkVUeZX6Klc+QZb788NgzFSIK/+5w
RsRpGxtyXPiEMc+vmywlZSCytQHco4CffpNblqNDujGAxzu73NgcGsyojWasXE04
A0pGLWQmycbEFbk1PBeGyIc2VGgz6DbeE2SquyPBj5h/D1wog3X7tKb/c3jrlY6k
DhUuTKU5EBraEjjzRUd5l8m67eSntklr2iCr1yzg1vI6WvB+TgKaKd8eT1mEdUXn
9nHw1nIIwCYiBM+OCBfdhy8BHdKyMMbPYUWpGHW1RtDUK0+AaFf4loxWmuQ1G0lJ
IYthC4Z4ZLSUIZ6ZDtHA61+idCSuUEhm34RQnXMzzXfoNU0lTpVYCJdfyM6kjrw6
pm+74xNfrGj89YVVg1kR9tjxc0/xhirNWbTgUYTttNeFN5k1PhKUDVve3OKMmQLC
po/OOTRbxYdkq+yj/FNoPQyItCFAepLM23y+vr5abUvaQtMSIlazy/b/dajKWmF0
sAw3GSMUeUGOmPPNClempPYKdq/piAamp8r6h2hRvEfdP1AbDwusqfxNaANznZ/O
UWwZImtSaQYU59LwKinILi8eC3gJb5P415yVJGAphbN1aad1s5fRRwbjxZaX/KkZ
Qko661qxJHpfa7gEylayklq/xN4N3VBv2EtJIYtmv5Q50+mttgHgHkQRBnN0emrg
5naBDI83Q/TZZlp5ZgQ+VTitDHRMTskm7CYBUOqMZhwkC5q+0sOYEkuBQM2rQu+1
jBpxRqGOYCVXfdtHM9mdZNememobxx6HPfXP1n3h2YJ5z33F0+uFtmYxuq1GAi2C
Z4Lmu2rqnoZFCAQJW/nsW0oFM5cPQU62aOXz7VunXWmTQEoascH8VLNVBYBFxtdo
7AdolASsYXFGNvbSMtYuGw5iNNjxu4NGQhpxRVflcM6ysI0x3oSNkEKOP+UiwCXn
DtUSRUZLD/1nk0e7+uHMETa++TOp4jf39+bcqinwOoOY8pb8sdlVGLJI6XMDR0Bu
6gR77ysxI1jmM7Pz0KH3evNohJGN0HaKF3p1w+cmurzZQ3fklZNEicyKTofrCkX2
zpG4BUqCvPAXaxofyyAOAMb/y49iMDVOKjCakeWy3zRaWjCjihywknkIaK2mVg2e
RudsIPsBbHgi2EakFC86c2j4oktpGpRCOVkTRnK8TvbfNw23Z+aWbzK5fRrCF2hr
PGYndY2Y56DE0xovjnf8V50BocExjADBs86ohIgX7PfkHp7vsMId7rVjopXQFaQX
i49NY+RnrvG1xYEIwf1CWO63IXep3dLk1COOz1NFU+qJQ/r9YwEwezzLnowdOSzy
Wj2u889KzFh8v6rnSLJsI5vRQWWNQ69LQ2kcD+e3AcYt408dxK9caeHNOkZMtYsX
/zepr0Cxmhg/Vt+E2jAl88tESxnxLTOuh1DeaVwhuO8R54asz+2YS9mxfXA3hLzt
K4DgxDJ4MqMkn76O83OkLdHBKhHX8DIzv089y0+dTa9khcX6TsZpsFscQE3VOR/v
o9DwLAut954LossFtB2Ok2t+nvI5t3sqVbapz5O1V0uDdeAPFUljiZX2yEkqYLP5
ms91avQjpCqWPqe8nNfv5qS8PtJqzqbxFoYKxKCcPMrgDzWo0Nl+OuZUlaWTUq/l
iG1aNZMr4T+g3B3PT7ZJjJDqdDBKK0CQxCjlw3tWIafnDBfXGCrXFlVy1klbBPZG
czut0cpisa4cO4+V96ZnKQSNgL7uj4YiM9hsUAcBBSlhN37Do6tiffWGR8ZulAvS
pls1qWWjisBq4TJ+Qhwl0aGmgBeyHz+3PKy3cLsyMYSl/seVMhstrpQ6Wq/Rvcv9
LD8vETM1Q1/vLpcE2yHgwqJdX5QJ3+FBn+mMMPUJoc4+OSl9rMJKPymyEt09jnuY
4jR5AgtJo4b8QibNWvY6VnrRCEScZ459ASo7tUEdxi/1EP9zkevfvUKROnnZv+ou
tKknL2gxDd9W1FM5A1uQXV2zy8s8quhMNOgt9H75/DzOyMyXYY+4wjtvUYM+LNHP
9UuyEgbsqbB5DiAsyR3ibdbwJvgQP767TYLoXC6ZMLfcf5M3Yb5on2Vk8RO0VPPN
76rSEwtQVIY+bkrQXg3/uapyIyVAtDnlxeFkMHkBQcFhZUtRd1b2iWm5wD8wMCiC
/kzCXpeDJDAL06L/9z+yx/puxfXoUvteMuh8iSj2XwVWwAaAzEwyjzEEoaijMfwC
fA4dR9K/qIqxAqo3fatcyjWiLAe6Rnx+eca3a+dCIW67dwk6aqgdnqMtGD4aB396
6CtdecdeZ1duxeh1t/zeklA3Wto5IyPfmjC3OpAnP1zQ8LB8tdPEfDCs5ihOx7hb
Min5EPyR4IeOULT0XCxh+7Oy5KnMHWYi8xeCaGz/xbyq17OPhusXi4e2Ga2m9RTw
qxaciPAUScgP4pGQzYMa2713NIIpTFIUJwk2denh8QfReaggxlAg0hmS8uPeXHa/
Dy8z6F8F2HVV9+lGMBJYNgV5nwl/VttWYK6K8paCoat508xOrfG2qXGEtvoKnYDG
PbFseuryClZJceUyi/RsrYpYxjiKDf2KikV4ATV0CjjNwLdS4/9yizyYPqk9NJ6m
ApZfl9cCURcDk80lqQb0EeGDMajbNZfeqKBS8pLh4O5JWR0vzANKKZ/waylwxPFP
F+KJZZZpOMuB2dIZOp5mlDorVQcCYPpsL1MMQkDTzVCxl5qIJUv+4rJMjfdsM3DM
8G/0+Asv+Z7BcdkfUAuHK4eOam5QXhqyOgw6yMcDeWkC0uzrR4gkNyC7C2HW3o4V
qxmYqMxCfww7Z2gT+JZlVqN3g9q6AloAknZieylXZaDw5edVpo/UHcyNXU1VLejj
89FEWz6ckHuODMzPmEkoIowvBsU4qNLvzYxkCiNq4iBVDJc/+RaPME3v8K5vDElz
pFPkB8Kyab/I6HH4S2uh/1l1E52jV/I2AjvsKluCWv2uzpdd+QyoPItnFQkxYjeo
eT6mb52E5ch1kg3iGJUT6gjZG4sfrplSNP/gM6NwUbethBwlz6/RnYRmBUp+MWNV
tAuC9PCxhK3BGeZb60KFap1/ERLlZHiFnL43qWp84OGB91frnyztziNR0RT/SRYK
a26cCcmh3IUnRy3V1OM7UFp+9z2ceLUeILV3NbNC5riLfeLJAPQk8WSSnvb4J4VB
2Nr5V5vUgMvJjwO0mo5/4bCls859o1E4EYeZ61rsffQJ1D7S5abXvo2aqL9p5vDI
AzGLtYlhIgTCS+mBxY4va414AAzO1iePcAZWbnbq/GCfxYTfcR9ImFT4TNJEJ9i5
DMUbjEnACNTA0MQsynIB3kVUejUgaHhQdpL0krzfuBfP8yFf7rmxTSbV55jCTVVb
pHmCcV+aWmQYRlG9B2EQQYo5wDrZPICGFxYC5fva0UWpt8IlqH9iiL7xEzFPsFlp
J1/bp3gZY2vZv+EZBQJfAL/pIbvyAb3Q39ZQHABt7Y1EaURmpkobAZAU4L9UhkyY
kE+vRnIZ7B1ttEREmyMcG1NNqatxJsOaKaSzvbjK3cg=
`pragma protect end_protected
