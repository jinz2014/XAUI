// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dlX5OwrnnQ35aJIoR6u0nANJUE3ajrW0/Jpp0efWzl2c5+KemWsma42A2b9tT2xS
i1XFd9kK5Q1BQqzEHH+CqSpCq976kqJOJSddo/gCEHOeePPcc6ObbhbKQZvmjYa5
Z6rCmkdEbt/JNDEis8tOAJEjlXOdayUSgR9Kt5nWRHc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11456)
qyHt9pqr7fUsHwT0xq6Khyx6NBXftg9nnK3ZaKRNZd1udr+ADx8jVtVKnNiSm0N0
2P75/erJ827cQLGLuTnl9M5pEPJGWN8nBcIpEZ2QJK48xZhcxdLux86sBIIhI2rC
/rYUn13nn4eXQtk8vDbPI61LfkeRz/5naX97hd1Je67Tizg143vq+CGwFCjBZM+F
pkkJo9bsiIJGUqAokU2dQGnnme1nQfBISnJL1OnuuAiX6K/IQspO+T/2uFxXEKie
8h2oQgBhyBXw2HZlY3AKDHdIjXRX+i+c0zMu40vBD0+UyfU9JoNINhzxKGUP1wjW
kbsYM2CWY3P1lrmBmdaer7t2+W3XCbLj4UFGwbZvCmWHx0q007p+jZzhbFWZ4cl4
3MoDflnBuVsz3IQAS9rBx/I/l7z3Z2v8BrF/ks44tKNj6zxpw+n9o0lNqJse0MxD
TdsfUQg/kVT2EjxL5umuWjSxd/BArDn7Oq9xShd0zYAC2hgDVEUehwuas87XLC3A
7tvTculRWkdpr9aKT4NPaaUOfMNECOXVuD51CpTaFz5FOfd9KRb7QjiwAwzbv53E
siFPBXKHtdv4DCeYiDK5j+6+r+CW9NQ/Zf0r5Bq2keco7beqWHqz/cNOA4AE1AgU
KnWaMOk86f99qEMb+tj4L+36SViiKPxwMMlyrN8dtxDvLEYiBd3ZzQcS+B5rFEYR
wy/OKIRTyY3hL76/VLfSQXPlktETjeyznvHI5rb615SbmJe2DXR2qm92HWqtkXPL
W1yFAt9pshmmrgLOwvIFLAtCdc/2+7ppXq5cEr0ICimpkH+4ohnsCG4DFcEqfG+A
cscBl4kx6Y6NT+9lfYLD/oY4fXt0DLROvOcjz0m+fgoGfFJx6ZWIZv8umMntBHn6
po0OyQeDDdap4YIC63VkNb32BGX+qNz/7iXHAqA1x3rg8+6MwaTOoABRoEmKhn7K
agQdJHLoi6v+8BINaX2B9DdI28tb+yMYjSCVpLH+9hmaVSXixvKTRJoL/y6Ugeno
4qdhm84eUdYQPUB7o6E6T+eJAskZvmw67dpwIwwzBrJQ4vV7f40Ns1oy3W22w4Lr
8YOrHNwtsJq74KY/doV3i+zxG0UssviYfmRhDdA2rU/N5uYRyq3yRmabITDfs6c8
lguW43l+x87I3YHiTu/tzL4VKui63gC1MgZ8EwJr0vYf1geCEhyZApIyrT049rXQ
OCAO0cSzXMTmKi1s4nSknD5FfgByUCjuj+mgriTpxv0GoVq9wGR3PitbQRcUED0Z
p6sUvzQDAyVV2Rbb7deeOLDNVXGdwpoQ2Mj0MxDIIFaVm5457/tWNqTByolmTTJT
Po3aq8pNDPzLQB7MCQxrKNAYZskiLLBWwhD7VT92+I7rDRmRS1+zVL9UdRKyKZzH
jk+o4oXVHReB9Kwy7hHFXg3JKZVgD+yLYIGm8gxyd5RfEmziQrXYVe/oGdXpec62
33Ce8TopV2SC2ert3z/9cYbnQjwZ6wwCxcrEyit3iH3k5sHaravyo8DRc0/GF6J7
YCI26ImieWdXLoa/UTD2gGqj5Qq19Y0teq1cVe+UVG2tsLET5q3UCv5izlS9Xnr+
eQMEfnkxjviiSzmJYsO58JrLp+lxr+rv82U5yD3KBjNa2Ofw4HEeL3EIrUtaP2+7
u6pjOpuDqGAE79bc7EDkerpJ2lN2WxiRdH0IxffiXx3lLWUAs82jXrDlrfWkeG3S
tF5DtMvsDXyKxna1V58ncAZcwLkXNhCx+OkkzCi9yDNC3CjaU7VRrEMTAF53EnEN
0wh8cEfB1MtJSa1KBcU73cVpVaxQk0o4th2yDZC1f4whsI17Cyno51bg40O2r1K1
GlqtjSr8D60Pi4/JEulzzMxlzwDkVTc0HC7tkptxD7R6tTs4kAqySDqa0QsCzkCB
Cmng5o1/4dzWm2y2eLQtVfINtrFTDcEjz1GRxMRCHDxg1Jh9I4SSYxDF2CnilrK4
9D6dAWdadsTIGI0OQ+HauYyJY90YeD90z0D+uaamFTz/zOmbm0cXe9sWidKhFIap
jv9QDd5jm4S6PflFG9VbSz0940OjAj1QgYq+Vg1C+spnjkRcXNZATMRqCcRyKzt3
aJT/JkXYI84gk+k6VaJ9cbmdTqu/5sZ7J1IpBwCgFtnFJppb+xqdDQjPcBY+/ud2
QLYTeppsJ51zM8V1rlXRdY0q1vWx+GIqHfnxeZKpCyIYLOC0XpokY7CGRDzInTch
u9PIe+8EUB9ozh7yzzxVakXyWN/5p3hJpzwWQb0BBgQcMtUjwZTPmE/78GaLpzBf
dxsSFmz9VoLSq/rqF4oNRNUYVSXHqEcNsKhClvXsPJu/fZmRb+rS2X2DhnmfPDay
mW4Hn7ogSU9FM0fJb00dORLW0i1i7xUfY27wB7ohiuTmA7pJRpKTnTtp3x13HAjK
J0p6a+JtO7gVgu1IK4Y7drfRZxsDlytn29leIkYXu+DiaLFEehNs6Mtmqiyzw0sz
AUAkZIP7bHneAzgSCFC3/ZzLLxSNxXiYoIIuEKIDzWUwQ4Buikyu2D3O8WGp5LI+
NN6dJHXgrydCTomly1y1A2gOYwWgqlO+y8m/Ja0XFxVtzt0H3TABbDcEUoFUzfVm
ZUCxeVulpag92rja6upFtymMlHI+oF5VU8OFynd0Hr6JaTBNkmbJmIhTe78zSs/i
3SrqYD7AqubHlw7z1796z9nq45dSkgoOTsvz7r/sY8sGnOf6IBSKEmAVUHGmkYXE
jYXmE9RAeIin0ewVFgLPOf76FoI4GdQn0zUKTwE8GvxTqfURdJXUplUEU4WaY/yP
jhioXQo1VTvhdDNv4kcpE8KH2Li5c6Ru7BbeSOC0BHeZO/x7dVwtyGKvCunr83g2
QNw3+Azb5Z8ojUJSvGW64dHLu5Q2PErv8v9eSP56mYKlEo4cKpnO1fVWN4itMvDU
DqjYpJdq55L1fU28HzrK7Y25rMToEHOHJqN9kWQYxa/TlAKiyPXrDTOPDIlUnPdw
16RvrxRz6zg2mWgxjh8dhj9WsqSroaOd2/qkt84Nz2baO8ox+nHPLf9NHZoV6JZI
oPY+4hjtZYz7pj5Mopl8cigsvuqmqUx4EOdbdu84oixAUhIEPZwd7Gzl/W0Jar+q
m95d//juJwzw1V6qiL11bP30F4vrww/bLhWtOftEETmdBBtR1fuJxlEjC8D37l8M
vmYYeVNF3K/w3YtLSMx3048wwdeW1iBLs/nQkySt1uvvN5CeetDUu4TOAPQPGatf
cZHdYiVnCcCfR2WszUMrci/z2rafC9+ZiFh6jbWN5+ZOStMsNnN9baCO2qa1WdID
9IaH6qwaeVJKoa+0VvQAJDyPEsaeh3KZ37NC6JMDjAHib7URdvqf9pF+DbeTFyXA
03Dsq6s87CSaximdTKe4bjBKgg5Y8Yng/pAO0fepOXCVkA+V0TvcjW0qrqqj/Aeh
9P88I7+RUw96HPzVFG6vZhPvdi25pso+d+R10qRK+QLvkItKgITUGIyKydwZeEck
vqLTd+y9FvYAu/eMvw4QPqi6HUha/xlKsjEDHKPn4JOeHHfAGrANCVT+NwynRzbw
D0kbBzdP7LdRle0rnY6ihH2HnPRzUrD5szdBQ/iJJKfcnxxnOL1OTDRmJ2PrWPpp
iGcz3jhx7FTeD0Ws6ZhOGNAxTTGjJsW0mz6RS9jXB4UDRpmdRl2hbLsYCgVRLRrc
d+soEeLTi/m76uqkVlron3CpRutI1PbmKeHE8dfx6/M3z/hprXhLeHglg9dbYSVD
JAB93EKNol2ERlMWIT9vsca4dZvXBpoKli/5TXeSd+ib3dS5f/Qf/bcyrlPo2DCC
Iy4OflJ8NikTD0e7AD44xK1CY+lUSvcZPCLEe3VT8UM7IsI3i7b6rbNgTn1uX3vB
sAFF897tnJfq5kuuEeKSkuSW51kS+EkEV1ZjJ1u8L2M+B/jlpN2ww1zoldI6FV/Q
akPSsi4ApqxfOfgcVZ3Vwr8j+LSZLaMcvJhn+ESaB8Pheu7XvtaEqT9UtGF3FB87
4W4o2DABp16xhG2I81T4ywYsKuxnzm7GzoekpVvdtRxfhvodKauWGvwPfiAT/uYB
TPLn2Vl+trq+J36S/aRzAi9BkwRpC3d+rBfW4F5+eHOaQwPIxpCMjL1OV0gYXxeE
5IqfZVrMs5UJOf8bRUbjgUCZNBPTgCoKk5BN3KXrwvbbe00OLXhI+hEMYhT8K185
4u94opviD2z/Kk6PYThCXJI9Wolv0ITUwZQsce1lDW4CLInTg/OaZ1Ho5pxdawbv
B6gOEOR0LYnShqOkK9lquuudisjk4iWRqMKOG4z1pPorT2StGhWIJQXmA687D3Yl
d6bMGIbNoNp2RVNVy0eBit1zgXVdn9LI8wanSjbKbZBtqrBMBzKp7dyADX8KfpXy
sx5HUpDaOec7J47YPXisWgXBK9QtAAiX1Wh8tGvunxIF0yFe/T2vC/tWdbawbj9Z
rZcQ4VTEyKNGhpKVVxDdS5boovXUFc5jLSXMEjmU5dfJzJv/BeBOeV/qtnAIpLjJ
dwubdveR1+10m7NGYepoThMh9ZSEIVQGj+MZNWvTl3jjoiL3tucGD1DSDlUquG31
GEH46bpiSnLAvlhI3cUqspUFUBytL0dxn0TIglaXLTgRgTAZQwUpM7lJ9ESpeqec
1RXSSPl62pwrOkQXi6jyP79qxBrpiu99Duet4tofBY2pAUmH8SSYNDh4CGw78BCC
cSy2Y6gjx4N/LW/6Q1AtiK6UJOt8gtt7elDSd/ozX/TZd0LpoCcVscnnN/b8wUio
telUqxXMFmvJnPrOsV7hYJxR/PPIEOhhH7HQy4zq1Vhw5fJu5BAu0WGc08rnslDg
kUJ/mM2P1Y4HMBMDoNyawYsgC479fTxkSg9frBj7/LSTkXWY3scTSi+tV9Oaq53F
47qncr4l567Ndy9gIKvKs0dHmpDAi2rRlBqqO9MVRYrVWnLnt9zkmjtor1LpItgQ
jvysBIyXpNiojKRylY92pXqWnEFl8LjqzPIaYjNF9ejojGIFD2r8OzoAX/XZ+vHb
cuTWpQ9ZVJNMcsRpJ9Yr26j6WRqKAo06llXrcOBmyN5UVItXzdcQcM1Bl0G0y1Cv
icMcC08r2qPlXLhxCWlLuyiow+Md+Oy1O/HnPCsJBuTXPqfxJiPI5vbzO7CzjN2Y
CPlkGz5AGBsg/er8X8TQNy45aciGaDlsTB4DSctJOtfCWcId/ZXRCpiGclnV0PBM
pQY0erDCTIX2VJsUF10MhxdooX8ZHFRZl3xg1L02g8o8kqwjA+Ucd3G0NsPtttw5
Se/0WDEX73xmNybf8JmIg1Ui+/RStOIPqSjzwA+WEocAgyVmy/V8FfLlaM9Imm0j
nyjlHZgiQAriD1wxUTqKQFVWbNIPr4o0mXJcG8H6/UhnkIz9YTNMo/C8yRoJeIEI
QbtPueoQFvQCGfoOqjJ0t0lmNl3iaJPI+hquhdeplqEnm220RZiTMp0s8zm3C+5f
g3DK3RbWP1bvYm+4m2Y3aWjYB2H55iQ6nRFJF58QWOoTQtSVC66NWklSscS94LWf
T5TD6qxLhtVhK4mUoIAqeDrwnt+1LjNT5cCeY6Y6lDVYB63J+5hm7cNaTzNmxubA
e9cyFOjedTjJ+4U+S0P9GF+S3gP2Ed7AiPIivxcKc3nXKwJEL+4bqOIzXn46YeWH
Kp3BT7L1SRY8wWFo94S87HpMIeemRJB7MfCrXjoQpaEq4DB5D369mZRkKfl4drD/
69EdV0siI9u89ftuDklEiAFqB0mP3VVVs36RyWoLXetaTNgnIIMnV+XhPqmkftoR
jAtsEfN1UKZ5cMc48AjOm8RGqHDBy3bk1siOO6pz0rFS260UKYOkaHEm9KnWq+IV
qWcFtarL14k/MC7D724fyBBeURAv4hRuTD1WBGsrkXxnY6hjZrsJp5ZJA1by4oog
ivJBW9AC9KmMyyA0YOhjly0bH/oNDbuCtHSol0LWlvmqV3uwiptEDOPYJLQnM/91
9jAkrdwGZi1sHqkJnbSWBHz45YVrtVtigIc9yV6T+GAOXGz88NXFUyJVdXlNrViM
pt0de3h4wzGDMspwqhVVHyjvaZdyfEjPiNvzP6JZymdMN+Oh9Fu0DHcaNWexSw1R
DlqBS+WT2Iw4qX+YW+xUdnFKzRPSH+2PsTIjCgt+X7wHV/0vrdn2tVJ2B7Se4Xla
3ovWBzenKnhFeWnlg3oxy5mIlL6FQfpH6VWOPG+EdAle3NVS2+jnLVzdylfZM0Yt
wVfe8VcRos0euiY4SC50BZPbN+JGvM5MOZG5r3JPc1CAW9+iqQSBuC1rD98XHnaE
torcRwqzTnjoH/D0mG7yH5ENQr3D733QcPjbKv6djZbdiKrnzqwnJYM8sKIcFm/d
OJrbaNg2qt5+9Nku3Jh7Yh3Rr7doV9R7u2u0rnUWuMCe9Nxgw548aiQEYfkmMvOR
PSGjAJTNVSF1FCMVpiQr8qnNLGY/Jo5XRg7GkDuLnTKBCvxvOMmHMwAiTL5fFYZY
xfjczCvMMbEhM3JnoKwGWLCRV8CVXDSA7ds2Zi1hmvHOreRGEf9bHZuUeygvwSsH
qWiOlszR8aROJGaUltIQCs9DvWDryLBqpgMu/oulhb4VLHgMDzWWf3GhsqwrQmTC
G1JQPVsSUtt/QoYkHTpefwgybqcEs1/dNu56T47t3g5138L4KaWiIoH+l4TXe5gn
p0j8o9OoiaRtzRwbwLDaEunrvWyd5Csd95wxJZ1GCTnJSzprtw54YpkIqSkfziBV
GENeRQJA1pl/Yvb2LsuTMN6sodO8PzhMR6PnGujDCTGMBmXgNbwSmqlH076gtxpL
IFncYbEP8Hp+7jZ7g/qhthj2ddSBpx5LCQ5QGoi9eZmm5gV8oYfCCX5foGZ8rSFc
Bpf7VnNx736Wh35yI2/kKRU02RvJw8W4+UkblDmD3rzI4utjhdd1u/+Vzn12OGu1
l13SSPOE6isIIfqdD+8aZW57PwdHA3A0yVou5HeQEqGHOPLi23J/xIG8H1oXmwYu
Hq49ENAaozZhZFDnLb+sgg1zFPZnUeUvnLjo8bnTcaHk0iOyrdgtSob04XlJ9zsj
T4aiHHLTs07+8dr6w6aCQbJw/L7K5oiwxJUkVqa10z9kjoeDU7UTtsW6dj+V9vKc
V0qnUecKp1JS9pedNrhEAr5d/Q1EDC9k6h6WDBtTULOceoNVoKXrXhZeQMCbN2Sn
FBc00wlPFU0Dg7ya3RCvE/97U5oPzw7Du15SJiXbMYuelqXaw/BEG5LMUTyHr/Ja
yqonj3dzyQqn6RSXWQwUqmw+iDuLsaFkXqVw93ja39tS2QiuEu5O0Zz4ES4gvqx2
mmqpxotrbupdha95n4MMtqDpTkm+/t30M3UtAXX8CsZZg3j+J4NVcQiCm+tQflic
YjNLN7RRBrnIWIJ4s/50MD9a4T9aRUqcI+OB1re05dMvamc5zr83GWzpcmAiCawf
CxO2QXGCpp0JclbOrlYJkge1I5i+WNRSN6OySHg9Ou/7M0O/F0b6awHIHkkcQ2SQ
FedIJfVYDMmB/BFlu7KgBQsH+Q00E9J2OS+QlvxsRscOUUTzGUN7wSVtnU3L52Q7
x4WNsDEvx9hGPJLy4EFrxLGBcnqaqMVEPqkuwFpqNUePjAs6lQDFvHEJ1XZ4+8qI
LwhcmhxdM2UjJkrlG7n5CrFQIJDK419U62SvaEin1UyOIw39AXFRaOXrm5KyCXTs
QBHbcxr9X/7s91ylDt372fUJYPzl8Cvh794sW77yUPg1Pm6sm+i6dTW0lwiO5pbC
mbPxevO3OA6fRgfRgpkwZxFYX3F9GcsmH5JN9srZiF8FzYHo6bpnPq7WvCZOE7lJ
+tKCJban9pGNT4BE0zL+aAhaJLOqMZxeKMttvLK/jIZ5xFrYh47F6/kc7Mqq6ihl
VDF8ypf0qVSV1gVF/LqPczUcSw/4Mc351XvKKooODnG9Yi+cwGDtf3PrIYtMyma7
bvG3grZ385qxs6G9DwUG8OU1+w7lUxKxauLmt9e07ySN3SIjRce0v/zoPfqOaZPi
tXG1PCC3jjln7Tq1sogVBc+13KpRzHE8e3oPDHgwSHXR8nQcfPKb166yvaqHuSuF
pNgxRpof9dBnDsU+nZchprSWCd0GIl2MYi8mCOEg/lR+pIvYn97FVEdyOxktpMo3
YSUu5XhIEZxXhlheDD8CjetGTo0UVXqcZkBdHV35BVhZst7FhKFggDXrCXgWTdpL
4YIlYFMOusfsAg8TOKaD751tjYA10uONHT9kAI4roR5jjkNwuq6+C7dJZs5xLLT5
sPMs3pPLf7I4sp1nR5dJ7CEYr7ek4UzNRqSvBN3Y9glM4GprPt3HgHkN9PzlpIq7
B3ygCnu2w3w9VeQ44jHoSAN2DsnB6VV3yPjmdxc179vzjS5y9+oJyTDV/yXCg3SP
PET1q73RJQdhW2J1UIelgpdIXFL8wcEKhARlU2FJVSEPWB1MCuHisQOTHgy61kqD
a0JC8g59lRbWvBuZJI5xyibHiN5XtuYg9RPmd71i+LIa2qU8d5/WCZSTOIVrqVSS
Dh69G327ckwP1kpQxDgX46sltnS56/KqfbHI3Jt9t02mvuJVlRUrCRdj6eRST/Bs
C78hveL7QRr/rK5pZ0hrtVsLVB8V4fC6Gu8xG3Eikdi0kb2WtuKoqCB9nNBzFlSf
dEjvlg2okcx957wA54B/iH8hHZQvsq/k2hc7sQzRyRFXpE7i+eci2u+YJxlKvFDp
cpBtw0Z4+/Dpqs/hlzry/oEM7/8U3zFTbMUPVsxDtCnV+IbtWwP2wMFSENL7Pj3p
Me861yZgQ7xDgU9GzT4vIYXwpJ15b1CheQYBM1IMZ7r0YBe4oXFWRJDDOIUeN8H2
r1UG2Sh8V+geZI84mzvtVmbIyFU2LTVRZkfBdvNn0ltY5sLNDx50a/c1GasQY+eh
rgXVPYsx3jo/WVuMwyirOWwgEBy/EuHccIruo1Lt7tRyck5qgtFFI0/SM2Lg5P+q
r+3zdNzt2E50eVhrLfjPd6xjP3soE12CduSxzYmMRglt/pSK0tBZ1p0LQVNyUPpI
Kte22CHSEy+4gecdU+GL/wSmJNFz6yAc0ce/Qd0n98goM4m2GtKmKvMl6fMqxqWf
CeHhjpWo230G0OVp5y2vBR5Zf6c+UnA42vakJ5zxNdBDdUPDrxufIoHmgrWOjjoW
MeNKFR0A8Oflpxlal35rtFcy14hNZ12OuYptIeuc4HEB+vboMDcfUnC+e854XZMO
zjBuNMA1+5uBVr1kSSfLt5NzD2IKZhVryJ4zZRWa3HsypEbezfPN+8YLgLXdeNXF
AV6BdbzrvI6YCZX3kWk2d1nBD5BV9xOGGG3yOm01vNKJoigZDRVYYXO6nVvFxVm4
nxDhvaLEwp4ibhkvkCkjRcoKICn51Ay0JNvToUTYQjiN3EYTldYWXojTnoug2ryi
BKi5zogF6b18cxDTLyYvOi1za9T9ks+0r7KRVYZ+JhTL/DSAg+E4r1HpgWftS6JR
tIOiOI102HXKs7doVUDO1hvXnHlaQ8X/w6NjAE1jSDDgcdzZLRWNEaWmBv8Oh2ZD
JJXMO4Qg6qyR5ClCALUP/b0D05J2rIdv/XFW8r3UhPZMbKPYumW4a7AU8MCEbzyx
Oalsc6Iks0fE5ZHfQe/lipWsywLmDG5TTvPGMhpC1fb/dfUwwPJXMLlOovug2xi3
MQeciUPvTi4EFEv2JYB3rRdHkAci6iEqPlo1jm7VeKoGfepdh0Kd65yhGn5DgLC5
w+L9IW7ZfxkqH9UoLayas8a1yZIwsixFAwpoiAILZG42HoeP2H0nxAACfNNWlgaO
QZVU1N0xj9INkxc76vZgFkc0FuX2ZZ57iJBHfEEbJbprQjTuX88UMe11K1gHcOXM
sAPNdxPinROo/x48I6s3WQ0+QHLxhZSLqyB9eVU7Y6pddMI0Oqzc1ToaISdDSH9H
/l7497GtbULq5yeyJC2231M5I9gNCJIBbQg48Cac1jx/QH6s5H1ie9Mp115am4hF
WJjrQSvIIiFkNtEhWPhm7TRFusnY/obL3/EkLELuqPmVMuwsaklRgoPyPxKnXIbU
Zg1uV8OsPBBisy80VW2JEZvUUM7ynAaB7Rl0OlPc15SNyKhKtvZyE0ScnlsUGGwR
iWno9Y3xkhA8hd21cJMG+2NegAB+AYohkovhFF/WFhUDDTWzDtabn0RiHcKvjLF7
/ZS4tnJJ+Vh4U8qZ4PyuPgG2vbjn11mdmNC9dq4MBS7cxwUPGmyi10kJxZwcVPGq
QJ8lt154E+jj8IUd2Rojw7WNHgbk9MeEbsPu5Kdv+6N+jqIDiSy6L4rmsXdIlpBz
Skyz1BIjxvr+vwm7Cmiay1hFiXhigrldu9XTrMtkf0lu3vka1fSH6RQmN7E3E+Ji
FHL56/FBizxvENnVQAuBExFxbiyp2/VRd6tE/kKE3ZfqoBSlmKHAEtFExCSp3MMX
VNPsfCyQMADHFoi10f2NmLbsZOtCCrG5gP5s7mUXwGDw3huoZ4FFCfu3oOnTp+wQ
oC47jY5YD9Tqhripi+R+Wfe0cRESgIms22ziqfyP3JS5QHiuUhhoaivyT2wCxXad
66uXN/d2N9jLgj6W+xoo7mFDRX84boi8MrEP3Fnqq2Gd2/pUPYqU7nddpassLiaz
93kz4JO4I0VuuxHfKlh/AdpKbBMRZfLx8n9fIjvuyGzxXSUySpIK2gXqw3DeWpyK
76oNruwPpPPHVIgPl0hPrxZW1Ysol76shim0uWosmaGOl+a7FCBedwiN6yYzItPa
9Hz+hemKvnh/X223o+X2BdJvn8lZ3jinW+PgJkV98LaUwiTZa/5UsCxBf+aMGFUt
wnaDXao7ZUqTahMAkLwK64AVcwH9ycozHeEdhkEFJrrQ3tD09t4pP+xO9FYGnzQt
0bpqvZ4pxvT06XUGnqd4GNs6i0JdmzRcOBPSpXpEn3UvNEFvsgmNYer6TlAEdWKP
RSNlZJg3Z9+UoymfX5QF5btioDFXwdgcR9A45w8NFyfNBwtYF4TZjSAKA10GG0AA
rST93fVZarZvMkt383CNRiImR4BwEbNPOc0Vh6UYN0nmTYu4rw/L3zkZ0Awzoye9
8u2FEbcKrhOrpkG3XWQxAN3OFTm351q+Vun1xsBPXX//E7yldr/L4jfHWTvP8wA5
JB5qpN+wzM/i9VpGy36R6qdVozfKy6ov6YHsrHWLSnBGKJ+wA8fZ+eVwPj8PwguF
JTIoSlSwkqa9fuYQSrLyz3wFMeTKlb1sAhAB3BzUrMZA/fgDvyqvV+SwsU/vJU7q
KDuELKn+cLRMpdl68Ggg16HJE/TJOK5PQGOPBmpaHcaKY69z4SiWxhs4kW1ETufC
zCMrYYoChpkv0zsICWR1gF9PHl82DwY+HgZuvevpJp/atlXzVdjHxxUP5ysWtg64
eZ1s5qC8Myjf6+WKV2ixVY00/ODvywyfD56WiVpLtthg/KdJDU+LbAoFk6tynJl0
gk1qYp6+OO5/v/Cp2VPTlv3xp65b7l+q7LKiwHuH336CO43MwWu+YAal1cLgTS/B
WQVFA5OE9vSps/wvxEqfzAXJ3t+Vdpd4kMzg0fGArp3XpRFix0Pp9ybnm5btegdR
cTvZL4bZKO9EiyH2WokihSFSwXfiVl0JcmXPgP713R7muDZJIpVQVGQ5Gcad+gyF
nRGcSOmF6C8EUXa9Q4r/IB5w6MViZ58HpMTqr9m1bNk0xqQqVi+2TopUPH7/Mg7h
BQ7Yh6ZAKHYSQOW5nIFgReSv0tM9qFPD9JpKxK1Pre34PNhYHC2pec2xMRS74dPx
YLW3PVTc+YQYGWX3IT0DFL9iTLQGOKc2oZUYfvIkyH5qJuGtKKcDojdUoF2CuPVk
2vzMVKz/LZg8HNx5dHqw8SdpGmp573hh12UagS3XfSkFV9/RggD/Ncj8L5BU6vrc
fexypXvOR8L2JkxZ4PFax1j/cOl8CTUKXLuGWlr2vmOkAOR1fUdlarXjmZRAWg+w
Z7SWxLp3TZY52Pj9v8KVk97lgYS2iugXz6KcE1Ln7CmKBVa2TqI2WX94sBICCOZm
qnFEjp53h0iSZktp7kFREzqU6yGkBEAQtXfqYe9B7kTNIZ3B+/uYP1YWnRMPlyDB
ceSvJhngj9jrxEi266kIR6ICfmWBsJkC5NcJwxde9oLe18xVUQxicFIDad1CzF5W
vLLYdYiLAwRi5I7AHYflfSNtQOFQH9zLdgcdCQA5EUsrBMAMeRofFiddsjcMHQ2v
CxUwFkEPmyUCT7xH843VSJO1Sh3KdK2sA+MSuoHbLxhMTwQYC2Fi2xLLktyI0r+H
Cqh/ra92VQKqpH4ceQFt2dZrhLItnzdiM/2oNEaZdBQT7bwtZx7ex90HyXSqd3WI
z7rkbguXn7nRhXLcpoHH2cv7jOQH2j2wsoiePpdrQJlEamVurCKgfc1rp+8SYmgy
PswRj3iyXdzSKVELrWiT+f0cvOXqwBBZ1XOchc6VgzStG5F8JCEdJDDBEBSMMyB3
SRpDzfhBfpJ6XlKLTVy1QNVGnHYlis08LdWbKAYEjVfVnRSH3GgLjhSxw5NSg+CQ
bABNPd3XElxheHLtxewIHuUpXiZbgUmThoEOABChlT4V43pYEZHzlAkhMgDYZ4Vq
eU/hB5juebF3siL1jPqFTwDOB3Qy3+7hsWf8lx161Aey4t8uexVrH0pw8VMHX2U8
7vOX7V1+eEMpdginy8H3beqlKmnzQy0hSNV9O8XXfSaUGTmljVmpCfswK/tVM4PA
DOfZr8kIb+YgcyFYGDj3oRgAVSstomdU9JJaoeM4ErUC9km0yaEJidFQmdLlHj5z
g4aTdGDfW0/KWQvzo5PTMhIbjci2jJubMfrZsRw/aVJKvAKMVnQVlvCH1DIiEDRO
FxbHhMUNwO4BsaQBiShSDw7Jep9oCGBG7Aycdd0odJ/WgXxTIesL0Y7xArDrlzWS
NPlNdCAgSdZO6quRx817UQsuE7hwpvqQVMkE6JH8ZDA179GZOJ6L7/Y/JpyllA84
zzbkSd9NhqMjR1or5wgl6V0eToXvICZbpyxEBmSKIc66uAcSBBZvp4EB5EBtVSjj
3iOn3l4CYwxJqbXcoPST3gfXH/ax8IirPpu+SwlRrF0NDZgfZjBR1dTQdGiLsl2y
hLXNnEsuuSkmRlL/kkIyh8fCNMx2R8+EaKaBMAxkGIzE3Q++knJOLmJ98VqdhjPZ
5tXYYHO+ITJZy1voG/bQRIr5al8/XWIV7Y7DeyZxd8jtkjHbXA9s8R9ktvaRdfCQ
Ix2OffHmhvgdCfPaWjLtV9vWCnFPx22ICjqN1gnS/9/PyAlsOSrDFgFf+0I3Y3/Y
BqYPpboriB5Hcn/aQ1Xl8zrLU+FUZRICoAbay2bOeZw5rFfWc+8FMaFpM4oF3HgL
+lvZV6HQls56fbFyoeEXoeQ5dV/mRe2DrsyEGLeVFFbq+yIGtsQgF215aHzm0GQn
ti5zarFE+WtbdlehYRbyrZrUgc1+uxHKIOrPR6sc5cV2qPaVwCSQ8K8Bm2Ia9X72
o6KJMLlRLFwSg/OO4z3JpBlYgS/pq8TxjhX5w3K0pc91L5oG/F235OlbDKbwwy5V
bYR570QJmR9KI47GP9M25ePHW4M+k2+FxwWwePEQ5buKmVLQnkMz7ziiQoIyokMd
f1azZ+eF/uedaYHHuGdXE2TsZgg4/V+EmxWm9GcDUE2zfjrflfJKprC8bsn9tVXo
I7m5E3QiFzx9kbgU6nT2tttNOKHqe78GTPZQrcuUr/4cJp/qJgWpms9R/DQuUT63
6V7RwwYXp3uk+pP6MNNWG/Ler1rzpRbQ56qx1BtTxB97bvQmd1/ZdmTnYzin+MKm
1bpQqYH7VpgYaGmDbpAB7M8nRjwdCVLG0xcObA5eN4RF2gt7Oy/q6X39a4D3sR0y
742Bzxcke1XMI6PryLAerrUdClVlSpm1Ww+69GV02vI53oQVHo17mK5PPz//14gC
cPtIuNDJv11rXQ0hLendqEUNlTA4dfLVq4NisclgHhuGM/id+cQBzs97Gsr3vI0H
B8oXFFHAGiJvI27oe7hBTmibrpOyxp/F0PGHCx6M6tvqQZfOAEwNYhu3bQ0AcJQ7
iDderS1af6Cc0jJsg1AaCqOK9VZsiNoQkbhoW7pSTDlE6uJKCtK0CqCW2IlbVz/p
goj3IVCxgCwV/p5hdD+NlrtkYMOcxvEgWK7pNx0YbNSbMDgL7KQKuRDUlqHrP3Vj
sqWrVWeZ+9D8w4J1hQZU+IE5LWAmjmIBa9bB7+znOI2JdAca+m8whFgjk0S1OQu+
UPVnixisK7kz/+Jxse3n2Y81NKWmjrjV/x5tk+QpLvmSMdcBPCxx5iA+Ef5OXaiX
2cGqasipMl9forV9Ux72tPBrVXonWThwWLZKmozcv0fBMfthYr6m95MpyqHCWid3
rfJZiVucGMiQ8VF1sNvPCpkGaZp8XfQ0J7wJ6TqqewFkOivNjI7WLjkHiWA4QqpN
eDAsLr8izBq0Rx95U6BK/rNUSTkGzpjz5woS5GahCjkJ92sxfzE0p+cMS4KAfjdV
HhwNw1YbnLW2otSW/pe47l8Lj6UKcjB8TD5xf9ryXZazk06kYIgCKHH0vvj77LFt
VBAeavKa9tWkt5AlYysrTH2UKI/VjLVdIBUOshXp2UzVLvyz2VQZKd6QW7pe6WFq
Pa/wDRhxSuBQYjXxikun+DRAw6x6hpc5kEd0iPe2KtHAWUpnoY0J/3RRINxwGQrd
8zA0NAa+WoR0M37Jr8MPbNz3U4WF7K/d2rOpRJ/zi5oTAvNKYBM7N4PrsPNpGEir
0Yrg/iZI+JWCsweY+3aspPTBBgPSyjJEVu9jcg3KliqGpk6WUTIayqGx2TRWDTXp
1LmgTqeFKs9sHFFApk4tAuWgbCuxp4SM6TmgFB9+uKskZWRq64Bc7Yoav6tIbJZU
p98l5uh6QQP/XIIVrWjbAoptKNKKunZpj2el7tJ0y1lqzH4ny2cmS9Sbmkh/d8ZU
plgWDFZVWrvLacqSUybckVyFuhI09xwM4yMmzy3dwZKQ0A+UBESeflSpa8zubnG9
3Pf0ZDB4SU9SWVzb5GRm86/f0/H0zk0ingnSklzjDEjZe8ZQcl8HFNHTUCULgJN/
1iKNhSknItxCL5zCXAK/7kne7PLtFhG0pXKLg72Nl0MRvicJeTSsM5JOb5jua1aI
o41LlH57irxHE+UsVjrvu6Nh2yxbwLCXtks39Ft+mjY=
`pragma protect end_protected
