// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YRRsX8q0q1DZ4iMmi+FZZlDHQWwupicvtxVldpDzQOKnohXFGyuXmpOi5qHQVYaE
2kc5HGwQ2C2Etvh7j4SPANVdnTs8/HeiXcp9FgGEMl/Qwt58NICCPhv9FQQEy5FL
DOLPvPb5LoowfBM+Gaqqbm8mqKvRX3i2jCByVFccpLw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16336)
gGpFIy8aqjK2/jFgauMXYa7Aq1qFKl7/GU3oJGLFrnlB5Pg68SJC95zCbaMNQz2a
6olZDZ93XYX71C+UTTlZvcW/xUHr+PLLHrqojk8bo86Hqm72jQUr8UDf/L+o7Yt5
icZ/XqeR0c7suIsIKz6G6uY4Qb2Cg9aD+hLuLxbR+8G8WUJvJd1c+ZfnRupVKoLu
L21W6RdmmB4ZES3+CK3K7wa7RtPKTfwMFOXGaoeGZx+S0CG/9jEvek4qKtAsT9Rk
cFI4/ms9WW3tlETxiDmx1zSCfuoauSJvEEyDRq9avvRGncKvITAjyCcJkO5KIz82
SsSu3ldQX4iBtoR2ogIpmma/FqwgNfP6wSnAwWnONMXygKgeaG3pxo054DbT38HS
UQ+KWkZyvAEC0FMCac+Ang3PikOZL6YI4McfYTxskxahdsy9sbkHATZks3VmIV6C
vFdUGZ4q+hba1ZLfrdbfv5/OIt/PsWloiiUDrX5OLDDZTk7DkP8O2TRblPLtLPdt
IBqyfbMqIhekYAq0VTvnmnep+jndtIqphIxt0T5E/eMnk0//GIIeGPQjVMdh2B4U
p28WAPcZwAb9gBrV7Nsn0n1MjfaQqE5gHJ5Vnxu1QPKRZ4EWfD8+y3HczMlwMyyE
5GKLWtR8MQ9R0q0xJHslAGcgS8getgrzJd2WyHJ376LSiO6Wc0PpvzWoe0zc4PA6
t+fDijs4szUvH2Qct3rkvZBKLIY3lo84OBWi1KQLgkAD2wS+cqIbSmC3zdrYr0Yz
ILscvwh/qgmBJK/4nEtHK/Flbnyb91lhUaDlOLGLW5J6VEWzjSQY0RaVJ+UbsjqN
yrthGMuxb6BWjdB9V+PbBqPG7Hmc3UdmOJku9sk0OP1jilnAODBxGrP1dIqvu3Lz
rApFi8cuCZV4aF1puzfxeu1bMVxlAYDvYxItxoiblLUixgWiNbxmpY3zHC6/tPgz
F17BnOiZeYGU9PhhnZazICp4/DKg6rIXTKabUi03Sa8n3w87uNCTPuuRvFgsYY7I
pkMR77bUZEhMtWXF4c+zSdMLs7tHfQnyi7uUXy1DJRld19sE4ZS16DftK6MEbwo/
2hNALnKCeA3Jw3SCu+cHl/3xo/HhzGK/weeb/z/zuaPFsswVdNNhx+ahSuJg5lCY
KT7/ZoNkoqPH5gi7BlVyGWWGS07iFsWIPw6fdTEZNxSCJ6JBOFVmbEu7ZSKyEy4m
p6SdnXC+RxWCfm9RYWSXHkVYJ0ECj4u4XhdLJMwQx/ZfaoTLukSQy00zujN2KybL
nYoWeLmqMmox+EURleqjsnAHSAGRCHrLns4cbfjBnWGhesedXqkEeeZEzmdqkcIc
ujxBhuuzrZpr5bzmBxbpzFbcWFcFZ096SLcsq7pvhzZEYt8Cp8b+fDeB0QN/2Hhk
BNHqMfb0cEgqTuomyclBAO3utMJRR7aVIIB/7RMt3Q8S3ev04Uzj2iuEwz+xcZt5
hpLKBNfqRf+/Y8LAD+wGspZ2nh+1WlshV/5rk+I/PSJPHRHMTnFvumMxYZJelNPK
Ykv3bhFXgoAFx7eGR59uHR41SepH1m2Os5OWpaLzuir8dLkrFFFqmK6BRc8inZ7O
Yk+FkiLOCmM3n3YmoQ6Xm6JEYylMO/Ym3Zg/LOQ/u99J6aoOqNpIWBjqK9eQaCuo
Vu1wdD3QTod3uYqAbSafRCqtS3R2uWtkMxsWkLLg5n59ph+8vWqPA4ZC1e9YPZ+G
4TyrlyjcRzOna39BEaZH1rACmyvx5pz5uoIrYZZLLpi47CF1utMoKsyRRTAxuV3C
wiByOkhAbH0dtCDH7tNBkA/ejuoEi0eGzGeXYiSdIJIXQx8kliikPe2hIy+EPnUl
qQzOJ6fd+R3Q8rWpYoUlhfGThKLbusYjpMSpHrX46OMVfMk/iBGK+/ITDY3+fCLZ
BkO9uNRuQsqnOO0KJYhIFwKB2BWBlgMF0vVDPsxPjYplKfcScycrOTs48xElwoOp
ddC9NlrRAp2baGQyhPWxPh7kMTxwDBiRVrhy4WqQbRqFRYEtOVnYlGN1O/vvQbeW
RvKW2PkKJA3mgC/cRoc/xOuSxq5KadHWYm5bPlqUq4IBcLsidmdqEjbRwhdlAKWv
OT8xhvubhMI1KZ55sqGWLByKvHcVfu32kLe87KUqwVPa3Um4XOaI6MY4KrJy+Szn
KCZwLkNvvdxIy+QpzR8nZZvNFCNAz8y2jSx+uccGwl27oOMH8F+bvAbMcVUompS7
cg+8CBJ9TW/TdAenav/P5QJ90hzdBfSuDHD84TTPrD+td8TrpEenxXJl/kvAJwaE
MchX4fovR3OPRn8ZorZWvcTkgAPqKLdPsb86xhb9V1D6PIB1Pf28CRhn2evtqg8n
SobJuEWbPGXtTSyogJSw2OO3y71UtBkxS+xs2P3wJgsdIAsyUItknuXKAbolNRXk
IcnSWQQeqnzqPoTpdY2LXeXEuP5UVPLbf8W0x0CxjO30qxo+GkNu/yKxUfUFpxsm
VV4jEe6QSM7IjkMKBKawVit86k7Jm0omRnS0RbyJEgxUVq0X9jU3XQVQSSxQio1A
Czy+JgiZxzS0CFKa8ZXx5WiavdKASIUvgeywHIeC3CZS/7KKD0BKCOqSVT64EXsQ
xX0bfAJ4hPW9lSw25PaDniqB9ESCNjFFohrWd6w7UwDQVye7Q8mTs8Knvgmx2jck
LVjf6wIDYY6yCW65XS7Af2ymWv3N08aHTfZjx8QW2nrvBwLWs0MHPU0eEk95Q/6n
QmKPzfXHuprbTavHQmbnySO2AI0S0iIU9O15agq4LN08gqnrVBBe2o87bFCTDjct
c3xwpCYMVKy9RUnKQRc4/LCznNnJvTNzepc1sXd0l2GaFKgMaLN/0aVACMjpG5Mj
bEv0EgJiPiGwQjfUjdBXtVKsBI4hVJSQ0mCRYHCTt833Bz3pRyWniTJQviYPx7yd
GR4YTP9OiiQemlo8SuxZwiSkVugb3/QsgteICPVB6PJCed6xTt0IOuOhx6cBn64g
CF8vYCOvamJRO1f9vlA6kB1dGll6hH9y8a400ihdwOfhwdlQtrZTnUVNskd/RLBY
+VtyKN/Wtth9pNyySLiYiAUxMxYJKjk5iiX0N2ZCK27j/0Ow7x+BcORYK1yaNRe0
gbOyLBhnngQ6DECdwt+X+nNC7Ryscmex0RjSVrnNgs8pxNWXF238LDc6ckH697CV
6EkOlC7MGMkgRR1hXv5iT6l7KMa55qM5jzgOLlD27qOKLg/RHIrXg3QJa4SGwSIX
7yrT5x16YzjKI6lsq2LqWbBEWafH+t8kJozhTE7pGzFzSCKK1gLuPdb4sVHaSEue
+mHPzXQFf1za9nSoZJ0WqtND6cl7G5C5KA+XMjIiE0U65G3A2o44kSQDf8YqeBys
PwfimmIPPTUTTyCMUBMmD5UqUY/ikm53yGbizZNZuJW6CF3SMVGSjBLxyoPnplA8
FWenkoa1mlw9UFIYwgbq7TwHeHykoXIubAiXMrHdcjvShz9PR5RUWJxvD0sDR7lS
GJiXtZHesUEFcvgrqK4Y0LcwviUllUu1AdKS/NKfNQimZvjy5t7dppDVKAJCzAbQ
4CBC0ecLV3dga0Yx/RGF4uKkw71RNXwh2vxrPSbp5ULSDye2hU8deFI1Ofj7MdN0
ufuDf+bxnkCDwnWcaFLWnjuh1RIk5Rut1ELy4DXTz5gQ0w0gP9lJc0bw5wVXBF2d
cVmKA9C8xLpw9YCpz52D++CgoXn7Hw4F8jKh3+s7SWcnG3MO5Q+GHWy/qV9ABdZc
/nX4egywbYVCsCkgZxbibW9btp8U9EBbW6JlnliKtyPSQkO2DO0xdTOMbERLgCLz
86cQksoHgdtrGYNFMdvNQcW2oKtFgsBhNLoZw1tYwtLCHQafg5WPg8aJi58c/dX7
kIad+U6Sou6i2Xqg60kxA4RfSNVHbYoR3NWDUww9m1cF56YwPQPpuumbRAjrzKAY
XZtJ3wq8Z7vHz3rnK3Z4iJqJDJPGNMsYx9Ie2xo9RcLbpM5mPu7im0VGbJ3Eo1Ar
+9Ns/bcAoYe/wSobkHh2vq3ZBf2j9WZiKyYJPmvK8F8MPsnboMOVjRDbck2ahNs/
2RwydMbi7dlry3Wqx7SqYxJarzUzQXETaLxKvbKXgI5Mx4lGshbtFudbGtgkrQg3
UpjV5dn7RgBY+X3h2c6RaMwy+H1YpVjrMJp0tugnmXeUmpL4wkKgb+R/UfuRUP75
GT8YWmrU6aaujz3KW958hfSIthJlk7SA4h/Bsuq0eIF0S2YzLJCiBPELDmJ5KTS0
z70pr9M4p+IvUlKPUnRYz6I8XENptE5cHik0c3mfsuxj0YWqvvuOwKeyst0BmK8u
AC6lMYhJnLJ4mtmDHfEJh8+IrRDx9Rhb27HH8LnL+1hYEzcYqI3gNEMgSICectmQ
nFrevDItbsluQla2OSmLy/ZXS1aC5cM2McjHau/eLdN1b4FRQZ1y6ejiwfvAD4Kc
OHk2Qdv3AHiXzL3fqfURGQL/dXxFV6DejH4w0KG9ya6gBt3a9IHQxBcBP6snJYoQ
wJgtN/ucsaqSbEFwn2fF2yBloqxcKI0tKg2iwa/P71c+zdADtr3Mtj4fEr4vyw5c
BVeiWjErB5qaM+atmRD1HpYV/ydUnVENNMctQEn7fnriTQ3zR8BSFSATBMW+pRXO
K/SSStVnpyA/XACVnWTWPBvV03q7vUo181W5wuE2uLA6F1UHiVZsRw/9YYodl/JN
UAjlnsWqsq4EpoFHAeTQF1/JjHO/1S9DUpXkFyUow+AB/LrRoMZgEL8uW6AKZW2i
qduk9/DREm4sOm8E0FriCSaGJGXszNe8DSLqRufjRWak+WheRUHRC+1vZSBbqYtz
+/YpDCTuXIGP+jMQ54OJ2z5wFYIz5j9f4eu2/hIlF+3BNAiqSTykWo98KOvdwcna
E7BApZxxz8yIz6XMyJb1MSAqdzOWcJqgukWGfezLUvRFf8mgTRNKPhfYV+CGglwB
7m9a71PnI3GXIw7MPgqCBMyFCShIB656noizrzgYSwvCEjeFLH47gob9nkuPQOBc
Yp1w2+dHJqp/g5etbTXZFlR5QTBF15H6kcAYS5nSVZf0XgWX7i+ZM1GyGhefbauw
PtTuHMQdDjNccmAh2tATwcsHW4TdYUAo1fLdxRnv7sukV8ARQ+sN6OCJMAlaSgRm
pEOnrRNhBM7v6oD+v7Ig4QUGDjW76NcbdCTvP7w9fn/TG+Ye9pqFV8YWgAtX56kC
Nux2/n/R+AxgldmsCFlmMVSoefyZxG6kuirmwwx45K/QJVUml4jGeedIk/NOr6Mo
OnYibW8f13QAv4O8tm9T4v0u3o2L0GsofKaOZ85NB7sEb/SRLyo/DJZzOh1/5rIn
XltQ59WtnhJXuVw8AB5k6AL3BPqW/+qe+OALD6IvEcvaoVgnnQGuN/DELq2FDml0
Egn0954z+SJNDeoCtEVmLKwHNYCliK/CjwsLZBdALJznfBszTa3PEmOEfjGmTlu6
zT7NCSfVWLfFrhl7B8DpQ3hqlUdaaZbiGOAi4g5OprKPScmy2JkAdrXpfBhlQwzr
tsSf5k4ZGZt0aiSdFkzQj+HeqLL8h6vRz2hQ/YdypA+bUdncSidKNZIdil0DzjUn
jlCYZfrgjfq7gw73ve8GhNrI6wkp10pdcLF/t6ZJRLW51oin4JEufbLo0l8Yzb2H
4mEkP7CATOUfrD0yS7sKQ5OmQhGFd7P4Fw6h68tcScc5uWu98oLOaVxBfRFKjCWp
eoFIYIbWh5tLWUZLBNND/Dv3UzO1bJMtoYYTeQEVhhdzDvZjJ45rCYr1DeGbRE8+
n0pmOZBEPgidd3d0/6i74PWqG9vrIxjmRz+YJBLehmoonEGpMVEeMdDsb/r8g9hs
+tkaeo/fA1KKpUJC8jdtGyWqYf1ooc0wdFyaa46Nv2nYmg3ETaPbvwk32PMxuglR
BNGgY1tN185+G5gSqMlQGxWWBCyGgKqsnGVfq70LmqydRTf4oKyFOaQobx0wYQKu
ak9aMMAZRrscdHjTIZpwpwmRyHPOdeGKKptz+eu3tnMIKPIGx0PrwuH5xWPfXsSv
QC4TX020eFV2rTVkhnVymc+yJq9RO71H1/K/qYrGGkMOboTI7cOxmJG1YrtxKn5S
RyMb66iSIlqOfVB2w33yj4kF0LwE5AYe90dNjqTGfbkB4f/5CDFdV44zdzcextoJ
Lif3HfKaqzYiCcvbytbEtWH5HIyWYLkya77JtlAp6aYWTZj/aKjhjTkGHXce3/Rb
qioJlTp6yshsBDYN+oZTNp668f0fd0rhRbDwJlSgM3rRSFkyUQbWbp5pmQdPcXeL
GLZRrXqsm7ydtB8b43KBGPDyAu/LIT8ahIye7JHi8Ec6op9CIWDz4oe4XTfkxfF6
jc+CJQJT3RbFq2N8mHwFnj866LSIbi6Gv3EirU3goAKo9mK/nziFUwfJE4F5yr6P
Dbw3S9N7McEeKIGSFhAY+/FBXaAX3Yt+iZpgNYthcihWjq4JtYVVxGuQXE9gagxr
EXiWqZS7zRhhLmb3MXjFFXi9XzRxaferOftxlr9wga40aXx9P/nAlatLZc/FxQ+I
6TOoCJisVxCH753AOdOFJORedzEY2gVFsQvV2f2fmx16xKtW9FjAIb4RKDF09VVc
IN4Cg4YGa8Xj3SPoAyG7xj75A0pLpbN5WDXdCjBUIfKUVxhFUO3NBDgL+2UR6t3E
z8991+GeDjk9T7olDjF/0tj2UrTbjgka0RfiIFysQ22ST7fKgNpUyjqxmmno0boD
evBjydFYAra8T1JBqLJ6A29GCaedY/cYGohBmbkEm3VB2loaobpRqROwOVVmHbVX
jeOk8n4EMSlpz+VnMgDZGVD0cL45BmJ9O8ITwwi/X3CdKFzi5ORfXd9OymipTGo/
/ARXIfCxQe0oPHsnpr81N7Rpt74ahKfMw45L8ZjuwfHMHRrjNKAvdKhnTd3zKunc
dhGpmVdkWqyUd0gYOSyhPlOznAnuBHGwL1B1OjOEVAkg7TdUC8rNeORX5eOkWSp/
7WdvDLCUGWf0jLgZcrh48hyJOkWBBXNxMj4Yjw4w04zlN0aH+Qq5Irgj79CCMN0g
8CXJgE52UC0qMJPrHelPBNQmCR5aybzMLRH5bj/XX86A1mkTD2/BPMsL9zt9s+O8
qP5Lxp3pNd/F+YX2WNrLABu7XvadkJ/tik4PVPyIyro2JiAC6GEie3dOThhNefV1
qm1jDc5GwxbisQ4wNIhvcz/dVsiIuCXK5O8iXbcIN/4Z7VilT2/MqmdCVDKVNpH9
YHgsQO3XbZnRyv3DqDuldlJMLv9yJ96T743/u3v9OluKDR84OZIR4uiUCiG9C7BA
bOEwI3lXJaeL2gHVKRMXr/xwKyWVjcFhl+PcSBnv/pUdcYgB4EqM+iL9N4lKhx39
OJtJV5/t4ttkZm/XHA/PynkeArqoe7QZ+z2SHJsp3FqcJ9R3rIk93vn8PURd+op0
uE1WZuN+/JNK5HIIMnBM+Vtdmor4QE7P7HHP5+9nt0Im8q9xIm3Z4EjySuHnAfRx
NwnSjL3avLKoqhviM+tDCQKjxmzgGdwF69PAHrpqbJJ4uxjYin+YkJzVKbhcjXOD
WWT997xcU8brK4ZJE2FWDKT4K7AqgRSPA7Ne+0Zo9pdxi7ESOrSpazQpNSqS9uJz
8ssJdkY35LIaqk1DssidBGRLfMBMjQJ0hglk0y9BzodaERIv9xNZyaefzWEFMChZ
8grADqexIEHBdskNQCblMUS0mCbE+CTKwjBzsWlOzWgPSZlOZjdS6/soSMi2+b1f
U9xaecT+I5fhNjDjr9/6ZfbilJ9wKeVP2kppvWFXDsTvNKjrQ8zqhn3ZSrK3bfzL
CDPmGOksi1X+CroXlQ26lnmw1TQYdh+t6PZa7p/rgEnV0PytK8X8r9n9otDYU1d4
DSBxThOzIXHio0W4KwfUi6G3EYshgRMPGGDBxoDTK0jbrsT/Dle1P+SdHTjpHZpx
ij71XzrBCHmqeYzXyY+uGOfiOQBwxbz/FU+8dex3E7+8KCuFJ8CbBbRWXtVItNOr
NTH0d2nWgdGZLKo6FQ52+GK7k7xuuY6dRjPfszueyq2RUWq3IIewKSp1VxdIYH08
HVZezCAOD7B/PA4UTOiFCYTsdoFg4rbyR6HzbPnBGqa1eRlRki8zBOwhd7zusw0W
8+pccNf4ddGcseTSbcVF4Mros7XoQdiJZRNIUDS2CI9LJymFYp6LoBala02Rv+8P
SaDVGkwwGEqirBwnsyzLsaOdWdo2hm96H+XfiWF9B3ceYiohbCEGjIyrUXElkZGD
jkKfv7iS8S4qN535JBlMSIPqcrSKJwIhwADNfD79oeSNpI8Gdffbkzlz8znEzCfZ
jN+xUQ0ozQhqTHVKBnzPWsbJdnXcwlqCdlhYDCsbQOK6wfXdHvytn49BpqyKyjhj
UgvNX4eIEUvvHn4AkkAPriC5UsezIsFiUHAoZ3ltZ+9dR2DCjY8YTylKClxE9RIH
F4XEQsJDf8Mwbfkl9A2Yq5i/zQVqKIF5qX6kS+/QGP5jIbtg6+E9kbiRY7qKzl0u
kJ1udn2j+LVfsD9m89B/mHLOIMLdDchd5nwnlutzIUxVFPbh6u4SqG7Q1PK68OgB
vJX+G9VhcjYBOWKAhJsHOdJBP9kBXYCr144srZindOTdo8JrVMbNEkX4OoP8NGdW
FkvJzrs9pr2fKZ5pUUNDf+zupYACRVfMnATNYxLRXNkM2bix9zGYvO6Hu/5O7K0D
BXJ9FxvmjcBSHHUYB2Hgne5HGT7R7vgVPVlGiWwIalAxgYnRbG/Dsj0Wwjwf8qGK
AAIe5U3/j6HIbibu+EbelNFI39QKZnQ/G86KBA0XVpCWtLHho49dE/kkHdSu1YR8
Bk7TgEhQrJNXhz2yrkvf2yoStbEkH1yN0T/xpxxn/gvB/3eNIU3CW5ewbvlXUvKP
nuzbsLdKz2XXiYHXWTuyy0cdOUfKacLh8gwm7Xj6aOoHFfrfs0QSDgm6oyqqRR3C
ttZrxM0ms53znmxznvoWPdqC4UoU8EQKrODYJeG1nV3JKxrRRQQvPWJW48YeFXMg
e9wi+Q6aYDv0txlDEChIkC/ZIlhqwS4fHD4Im3wnWBwwSqSS21vYkCgfBPQvYdXz
7qq5oCbwGzYvZPYwBQERH/SiDhIH3HJbqOD2i3JUvMVnbF9aJxFKmBCz38csOGoj
GpfNcPuJL+YLx34vUPHpTGg4P07DiKZ5O78Tm+llYVwdIL2cySgNjy6KuvWm87IE
9WUDN+8CNtI8xOX27fCN7rGjQ8e+928k/xA2JnVyZQ6wnBvgU1Tmh98sPDMMzem/
JZpSKwsCgtMbNuna4BmdXS7ZlHEH5pEutR5KRsxUk9C3sDzUmit3LUnsT/E5ShgI
XhZHb0VfvRTG8/g0K/zH1ayo1futWH88zJ+qY8Z/6LTO4U2y39FXCCtPuqU+lSKn
hQ2Cs+rlVgcegdRl3y5wfLNbLO6Qz8uqRr/l+Xnq48rffGN8Fq7FA/t6D/MG+ce3
88cVh9ZrVxLgiGvlUEp8ZcQkMzg/3y3b+zqXlCSHk7BhxJ9w4ns2zJNY5qOwm3cY
EuWuASNy5fHYXbIfniyfunou/HfUo+l2ALgRJ7Ec814nFQrotVN8lb8wPhXNZNfa
NGrMwzjN00OwAoge2hOr/9zmsWadjZxYvKdVpXYLbeiTTfI75EUS8O0Fdv6arLtp
y2BO7GQOfr/V1jIV4NHpaaoEFPJKzSMP8ep68paFoNchEIJ6Lq0nVOkUqtrl08Oh
uoVAsPCVpyLSjb/vrpBXCxkUFT53TrD4ScSqSwNZMox2ZKKN1fmhlBf4WBCUNOQY
LdMfQBDhKzPUsi9CTY6O9OeDOhWgM+2CyuJVHsZfwtJ/tIMOSrbDxvaafLyFoTYC
iFGG74jXCVfKzAcbIUD65Rme/EmoZH09Zl9stU/JNda0hAPHP61V8gL7Itp2IR7k
OY/ZBx2+xUC9E8iqlmsufzrYKnfYuXyZ9tVwVLRBESTXqJvlYc01QVWEFz9kHHiw
+9yVYbQsKiUCWgsPaqRp3NVS7Hk7CP1ye6wWX4O8O1Uv0toPrIJMZzt/ySzUu84h
9EqJaY+bP0MwEjZjMruZSs60bLgx7bjv5Wn3xKR95aSWADdOUwxHSfWpf733KxK5
UZpFiYu7e65lTaRQf9YDcqHi26wffYDoKcTc3DkyFMhkrvmzQiAw+6DnIHdBrvgP
ijArLawlA82p8aUhwAUmqH5AKHhZPHRdVbfeIN8SwS4eabkFBPZq3vLV+mcAgjsF
RGbw6mL6hcOnWp99Whn/1yn7MyO9m2OSjfOMwT3mzz82ojNCm5nHG6gltdVxXNSH
CfXARHu3Wz53/mSrImf6YsQGNbhmAtwiHRZiD6Iy59JmwYISvFxJWam8fb18FZcx
E/irdeZHqImRxKngEvUichGbkC1Wd86J8atWuMOI6tIOhKW6M6yvh9y58paHvPKN
BkCg0UjcVbuCEyjxVvOW2670vGGdciW18P7E9q8d5hzF6zxQuEtQsqBI7RMpcwln
HhjuFYdJnc9OTyXFhEXTEfqcJ+xkrBHHoueYfOd3gqECUFEufR3eVER+KcxQW+jD
TRroPiDn0UkIzwrqn0uV2eiTCJVJC5p2QcZ68NfMMbF/iQtMal+ZQ4qBhq9OOeb4
BL4fQuwkXgnudDoWjrCO9hqaLhnLgWY8QFyu+/iwNENZwYTAxbGV8oFeeBaVpx/f
e+14oqPOrC574oyU6l7kVXc9n4U3m7j7E/ku2hqTbHmdcZ3L0BukrA4IUpXIBpK7
CrsDJyxt1TdjHr5FxDJFMou6QMWvtaSooN7T2hRTRV2vaVMYssq0hvzX3b00rQsO
7P0u2sletGmAJa5+ZIiS/1uT6fXV2iPjR1O+vnHEONcx9t+biY9n1dow3FyMSRc3
JMWmJRTIVl0gGMaajM01f72E5ytVh4wXxJ8plcg7/ciZ39cgwaPMZZTvk5IwAGgp
26cqntCVwbJHpp4M4Dc9oCSfukTZC969c+tX7xyc5CnHCg/SJXJc2IivNC9C6xQn
LktAGEDfvLkiRrml1E8ZLQ41fxxWcVv9D1fU37aJxG14qNay7b3/9s17MAz25RQY
TNRYwaTbzkmeu4kgHuQ70UyhGl5+GqRbHncWH9NKeF6ezOruUdTXfxYYOjtE/Vn7
0HuOnkCrInasdgPpIdIaJDf24wkMXB3BG1oJ+H3l2TyRkeC3Zi/TeitMB5oxoODg
9iQhcqQeb9q59uMblLlIPkc+jflLb8oCJvnKyFYHR4MB+HMyPxxUCHjoh9WmpVhf
h2V6VmsUkP+LwfXRlYDsFwKCSyYBf/6baX2lGmOcSIH+01hA/aRG3K8N/HL7dgmP
FALQu+s68sSJtsupfqUGD6HQJlrb2ynwo4MiNFZbZz6jLyxUKHtEGGC2Eg+8EEZb
PM7XnRQqTDWhhM+gAmilGJrlz/66f8dNdHj++C4gRQ983eC/qp7zUQkrOeO92CC7
R0c9dg54RWxGvxBoIA3lg9xHFZwAFWZve9L8CMd4LQmtDE8WYMgue5Ku5t+G3GZY
kb8bv2ope99j399fYH64hGVVrCB4G2FeQVWQPNP8oVyS1aGgIjOC+abgkqIp0/66
GLLRV0wFwAxgye+ycL+4BlT67eApCcWc0khLdMp0gXTm/Vq1LCqOrGb0JQx4d9ZA
FPyWbCIb1bd1GaeZwiOvN150HWb0ssfOvS4kluCQRBEqUpQD0NlcWMQL7zRLrUQn
1352U7LZMuQ/YWXiGZlZn0M3KJp0tQIa4aj6VfeXKPwpnz+4Um477gubPznXA54g
xsBBnuvo0Hbc1vd7TutqVDh6KxUHc/QPUWCiYMLSSKsc3+jTQWhqOMUNsE5+lg1P
Lu8QRXBvJybQUS2SbFi7MP9WHafGCvgMkgvEqvZQ4HCj6LQQTnW6qtUVfXAK4TQx
oXkS0sFnfkYFqcj42OsC0HnKUzwQh2raQyI/s5mvTDIeM0RetRHB4pdi3TxVaI1o
Ns/wNYNbcQzmhRGewOldcAztPv5+X3ZayywhCevO4r+vnPq4ij2XRlppm9qlkxQ3
abqZHm1sgo9m2k/qUAuZGM4ulEHDzSzQbVNoS+oQayvlzRPS+ByzGNvD6UAcabMF
ohBzEd1YYsEMhVWEtMbCe4mcFTgLVIMupiHdJu4FCZMyCiOeRKSWamp84qCXg60/
n4UXgJedUBdY68iqkqEwqjcZFCLQidRF0uoBPvGl2BQh6CYvNNOx0681okOzbLRL
hYlQCf9v0AgIb/iCR+6YkqDcIaAr4tlN+E6IE8KJdA5rg00ttUzhB6i43yU2fIyK
FudO6JdSmZ/Kxhgn6xL/w+GPZlI9pnbtErz3g0cuWGtTbYJ8Y7SJXS0sw+G5HCtw
u39o0puW9G7XwII9ZYnINNdXn1X/evQPN6fatUCqrMkeibk9h8PcywcYX97nHG42
6psH5LQHW0k1JCgCyNpxlalQqCrbsX0b0/72TMDwmsYg+5OT3dt5ysvouX1aff0z
qp41gHnKODxgWhu0Gg4HmibgreoEPCRes0EeiJl5xs1jLr9PXSosiSZQ3NNJc8BJ
uJJpRalTKAqeDEAWaePyQTX+jMxdCnDcdccZ5n1vMvEMcxXdZjb3hElHW1mEQ+vj
YMF8i42G5NygTfQCj8VzAufB6MS22LHNbott/PAPWtufHKxEpkdcKbmLsWqrasXD
wtaStgcJoUJE/BHSoScnVS4iKgUvh9iGnh6EZE7zdFSBbogX/i6QzNIuwUwSKC4N
rWR3ML+N813ZY8vF/c8LGXSfznmYPSUD6GdnAFpaHazuW5AEvyok8O/SAHwlkmsJ
fgYMJfQs1R0cyL6/aU1uxy4NFmvJvPGcEcaSokTfgZ2uv9bC9/Moo8P0rCHjvamS
xT1cU0pyJsYEBl9Scgb7OKsebDZfzg7lzlY6rnB8XN3GvgZEHNLanAiyJUWCd5e3
3lAIs+yg9dCY4LhkC90v1Ypm5Hf5NYYZd9XYzOAC3bo0ZS5+//h053pHEnzGBiQ3
ci3SHoYPXbQGZpGNUUKyUTrxZW+e8N2eIrF14CmnBPcAu143R7J/LQrcE6K5xKrw
0Q3X0slJR61I7kCc5lpwPpf7D98w2t7Eai6/s1LW+q4T64y1lG3q2BkBlLlcJVr6
rls8mJDPrcYu13LS5asYl+pk/1qjoA34MhSsAvtNcD2x494qpnIFAJU2+4zy4Qtg
8xA2aWEGQttuxm4TBOlrYEZMqmgXi8yUqMwR1NPe+mdGKQIgq7CjaCPN82rWvOzw
H/rIDcZHd9n9AA36YTc2No1w+OOH/1C1DH2AJTFRGeq/ISh4ejhfpHc7Y9t+j/Cq
ipGZkDfLhYdG0anXQ6pWLbX2J8H3En4GMHCk4zzRLXZOQbB0JW6ftVJXNfwtORFG
vMt8W87Ccgjx6T2G8m9k8nI3aYDggjMKYtdnKiAp+F9sb8sWXdurLL06sMOUop8c
XmB/jKWkL4CohVdpKuP+UxQQzrgnAazVzAmiXzaghKppV8Btq53KWvT8q/YbwAzf
OdrsOE72tc3mwL8T7PwL/PWTvq3yilp+cObf6qZF5XTyjRS3NQV9XScAIODIHlqH
CP9OcLPjHC9JlsSpWp5AhMpnmGgaeYZ08c44aVtFD1tOQFPAuSjpi2taDstVDkVg
IvngZ06LIpDHkTX6svoxt5hR+5B+3u8pTlGtEgPWVT4WsLjOXvsEgW7PCRZFwSsQ
az8bGj8dS12OsoF3OK8/xaDN4LRvNll/PM5kHwGOoRKGfaD014if5gEjo+3ka9b+
jZvZLTAm03ctARMIT2PLLa0hf4A9q0vK44PorvejP6iFNUvJNTeEGXx499UQxnlY
KR1mzy6K6hgJygzJfVe8u6V/f/u6P3c7w/8NY7QlFIa0/I58THuAd8n2fr2uOTAF
ke1MymYmj8gMzXOjKs+HzWogDm105ngZHxxNwOAhBnCNBpS4H8ZEUYxVlvwjG80T
0ZArNjJfd78+626caR5SZmOVbbKXhBQ/tCMCtKxWZFIOkdbghpAQa2vhbCqOinve
JGJz9Bud3nOnu4we1uX8016QYnjbeOork2GEIrc1zoBluaMT6ouHILINf8MnFdmq
YMlc5tEyYNQr23gmKMuAtCjt9RGaSE2vD/CMYCr1t43iUV829EAc+FR4z4tjmlSi
9pS3YnTz9SDTdaG6y771RIOWha9pc9LFB004RILaZrJ8I0Q4vtajP7i3zoYRQX1S
12eeKbTrprrwQLjW9ikwRS4PUWwjT9jY/C1CZePjx5A/cOFhQJlVqURwkwejCONp
LD49WF0tKjaXyKGoIj+6NNULWQs1aHfiYgt53URFz8rOSTHWNO5ix0pwQRXjzIQK
dUJlRpfGpxDZB4IkeNIvcsenXb1Ea4Rssa+bL73BssD5QBM8B0tGDJ3FOeHbRnci
ji3IbeSiaoXSfM5b/hAemR6E5TIUKS/UbeCUsfzzHVuvgdCyR++QvNO/qC/2SFxP
5SzrbVmoJ4QDxMHxa37O0LQ3zZdqnH6mhQFFXXfUHe9YSOqDaDgyk1UIq4Wue1Wd
p82+uZp4djoOHhQjVJ2K6rjniUUhxvaBl7WCNmaUPNYIpuXS/v22b4cnkpmYnVj7
m6KvxCe6cNBh/etV0FJqO1vwyzKSPW9LSCUlvSa7DurL4pRcTYthZNYUJW9uWaMO
wjtoVOAdKtI6/ybP7nMqG1zVxNwlQehx6AuocaVjfWjsajsBu9pkQo+2SHGUWXZ1
g8ytkPtiS/ISA4eDT6Uruall5fR0IL9eBeK4esV9lfHZRN67R13/+6jwJUKitjkB
NhFZvbUJAhctiLENfolXqlU7iVTwfX0V2ZMQGYkAf0gG0R1DW49R8tRS/oV701N6
gS9UYmQbgZ/rOvvm3imXFlFExwR5kH0KXetuttt+DeT0PbzX/YGuqjA0tl/ElckG
jxOjK4TIXsDTPaeeKSYGf3RW4PK5JJU3PuglIyeLVGuAVkVlAk6lqopaqz0LeCst
YMZL3di4KLvdxGz+3tEW9V1O/qL37bn8FwixihxP71aPAFfHL8DCZUX4bIaLkLpz
R9N2jDbf/0noRwTC09l7oxX54goWjENrj8wD3hM+iLHqKzptBi7cEScDRJhZmrdm
CwWZouFOqMgHmpM4zDdCCb0Pw6TSkkQ7rCDJnB5R9JTTZfBNJ90LgGcnwunDb9XE
yDJp+D4lOnOVm9myjXawwx3dgKcIvOElTM7F45cgrpzt+8D6ZL/FZb3D3FWBhEaf
+UY43ftoaJFghslu09LkZtjm7NEbq8ZafPOWjKJCPsGOnspj25pm5YdUJIS6qUQH
dJ/7DXWPxX4vYtdiYJCz/s5TX4n/9Zoz2Tyb44zAW7z2+WeeNUA4QTjuVc+eLsL1
+pi5RNGipURN0Rdg4lW10W3fWhaGmNcI2qE/smtZ/ZxTzDC9z8zj4mr/ZYLOhvAh
N4IMc8EDi6JMlA4YlTspN/UWYTlfcT5OQtvbd+bNPMeict3HPQUTND/J9cKOGOwW
UWOxbC7pgNrbHWTgI8dxPLmbNcv4dnhAXV10QLFmwXQ1M0F3D3AmAVeEzdAoXQKE
iddYcK4YmFf8XAsmR5D4yt22SYY57DBnbCK1cE22oB1kkgg7LBSQRnoul6dgif8f
XxEWB4oc5PMchcVz+eSIcBoNSa1i5w3JsTrxR/vimravEl8Q/4zGXMlgzofnWF5K
4x2j5aDYgyIfvSIyLFq3OzlKh6ArC3c2m/0LsexL8lSrxPux99cHgxxzhuuYE50W
GFlfxMM9qmicPVgWiBnGs6+7TnB/gGU5w1XKADLFcvagGCd94Qc43jeyuVgf4EUq
VvqYx7qNW45Tg9OSLU/jNjndSL4lrIvD18ZCOyiybpDGyVe7xs+w5Jjfv2/HO3n/
FjJNhvmSTFIM34wJgrd5rQrQLH1TruEafU48xwO02VWT+Q59iu++SVRTn+XatSaA
9ySADW1qHIuFqrf03u4ApxGtB+Z5HY5vqbwKymA4uSfOjDke2Ybwd4Aj/x0x7xrN
ethjgyMq8hRCMeAqbUMwdE8o0k3YRezC9bsMrhXe6o7B+sf+siAUqhHFa1esbrLU
RgWBtEA9sVKcBoBDW/E0ByOpH6dZxe46wxd4BpxjywbjwTALZSEDFRpHeO+d3LEJ
5RtCPRia8MwwiDchFCXPuE2SL0aySxrO689+yMJpsXlkNirrtx1PwkgNSZZ22J1o
/jX2NCy8e165E2UjjqGfjd9SOjoYueiYlbzTJnaSIPeX0kk+aOTN7kR7KkLGEDJD
QOZtr31aoJiu0o8l7Es0jTUezllQqTflCtezlz8YN2OAuL/fR5c56+MBdJjk5bUU
SEAx7bZvP0v5W6Wk3jW//uQwCDWt9ey/iRUvh+csTbr2F8omoOnOWB7Itc7AHA7m
vFCazNhOOI2Lp+VQ6+7j4vl2lSooLp1tgGs6tf4m6KN73FKjXWIOfKM3vdHuUu7G
jrqHnrnPTka4qENVaCJn8dUQDU0ApUpdB9LZJ+Yf61aOZoffVO4+cGeTBQSRbZ1R
64gpVda34FAwjJsSdWvL+4tcbdQU1kqjzfUx90z/bShtkXK28XVxDoge3WWAAn/Z
zp0GdA13lJaQv073USa9FMZjr4yWQUOwc20F6UgONOn484pGk4ft3vSDhmezok/S
LKsbMFTdGWlJJo2lBX9aQYK0ORZKmLRfmGLle6C5IX8kE7Jruxq0zbkIUzwhJU7e
3953py43J8JBNM/Ej14wPSWN78GmPzrTPtCMgLyzICKPxI9fYRMprQClOZ4ddEG8
4TvxDaYm8a/UHXg1WA+KvjSLkBIZzns/rGuwDmXVPUt1132q73y/v3YqN6Pk9+4+
awn8C9zJop4eyowdB1Up1MXtQAGJ8sYEdWmjf/aALpq8qDkfzRT6jfTK93VqIM4U
YiLKAwOwYejoO8rdiUklbhcGiC81FpdhsgMPnomsHzDLGBKDrYUTqDsbajTtG0Q2
Kx+ycv/jhTChMelwDxaeGu+rKlMPjHfE4ckZkze4zjplGMVYt4mG+NF8QQXY8QWu
xm/AkamgkABKvwBff7sSIMx5wmu8R7abq7vAquuB7Fe1ui01mvFhly/CL8UujYvt
VN3mfkol69QiS1UJ1htDl1XeKmsazMRMH9Eizq6Dy+dxlz1zzJN1vHUgfKG1sDo6
oDvwINNtZeHfSreoHzI+Fafx8Y/IYs/bgjvxQymr/bJBrfpVPh8yLuC4SJOJNRqf
mWglRZn29Snb92eP34CVuK3FgFOufZDmOIILSyjcD5Eup4zpHwwoVwqF2g9Gf2qF
fFrwZ7oFdgdyUKKRRFV/tKQHbk7AOHKMYmK/QTJEu3XoepOikl3yT4S8y3WihgCO
r15BB8VdH5CUszInVhtvl6ozxS/LQeLibFTRyshHFnrbLq7CWCt/al4U55Het4Ve
A+1avSMYSa8LvkLZYtbG1Y9962vFYCTPYy/t1qM9e+MS3Gc8nhUmaILparf5KLDo
fuH6JbhwmYL0o3ZvHy1mp+9/ww5C48Ov2hkjgmkgWrEIUHrWJf9hEki4v8SP2v0D
aOJsxe2ZD8LZUX5DKY1q202xxmtUzBj9rDL8SRa9l9bqaOwdqFNiWiJIbgM6HBht
dRQHCARAlgs3gq4zSjYe25qRiWd13SWbfcjhFXywhkjkxSb0R6I1U+Q14JEPAVRc
8I49ycufCUBreKyUyvoZ/cHjGxI2xVOdK5Fl68IYRtGhyqrk6VpCjVlYdOAishMF
QmAY375ZUTNsfLJc8IorkiGo3BEEEqLnovJU9Ap1sWu9bsWQQgc7HOLoyx0khx6k
3K0rdyhPYskyzODE/3ZAK+MO0C1mpsI/RsOGE7ty0cfdbv22R2jsHl+b4OzdZhhH
ndu+iTcJLmFCkSxH2wWPNc/rwrpQpMO25CTI/qNq3lsyYC77WySZ8pKar1c39bIz
2pdLVecUl7X6DkOmVfJgL2xjN57CP5PomFY/4+wG93wdBYHpbHevdtZMDTIWHdgO
Op3SZzA5jdzuf029Gg5IPGz8k75cNp7YEPvTF1rqzcXxVtl5Tdimud1c9lLvzNAL
63PEEgjGzYC6LUw+YXT4P1yrM1tz3Uq2VrkfsAsAlPM5P6XYgk5vYChspOIPa+Wd
+DLcwyRCD6+E61Ve685fwuTVWI1RCkM1moSelUMrDd9hJydIzxo62T3fKliRY1gx
2zQAzfNVHmXEcQjF0E9GK+BngvqfgqJX05MlFyGyAu2Ciexjp+Sr8aXWD+hc5VNq
M8wl5VPkLg2IAv7lfIK7ned+MHaAkB/tixp8zvtk0+9165reHvK/Y1tWOSKf6fwc
HjVQVbDTaLhYzZK1dhD4lg70jSW/D4zSi3F5pdDaKIJdaMFtcyQ81KW4Da3F0Rfa
ZUshxG5NWbV3tr0NaJTx78sOxMa4he6VHm43RV8ivkrSZnQaIgNM2QVE2NpPGvnw
2DkmPH92qsiaOIgaR9CiSe8/m7na1w7EnjfdNZT7S31gIHEWLTwQBRXYf0bEZYL4
sD/uw5j3T3K4rlByZHQQ/WiCq/ktymcDn3vliowcJJjqh9NGftphKG19+1BzCTlr
ICNVuG/hq2ktt+/YA5EzrSZVCXDRqz3hkDlvPmwAuTTn0nzusIDwEjA/RNaYSg3+
45TNhQeXDCe0yVHFagERe+HAcVafZcE1wEdq+Hwo/HFqFM22MZGBxOnKbwK+jOgD
ZxiNiYE6rpNZMvwTXj+R2+a9fcB9/4xiMHvr0xqCxcpS9/drmIcpqFjvurHd+TT2
UL5xcfVGIPtwAPFWCHYX86TBelvqvjNe8CdJHkMkxq9aYC9AX1xGiZ/n5ZsC6qP2
+UvLIzH1/pfisqI2Ir1Ljt0bJdDyhV+o8oVjxmAX81G3Ltfd2pQ8eepCFGbtZ+9V
CocnKvUeL5SI99Tl7MvstA/Nf5CAOlff5IRjdMid973KHGJ8JvxiszQrWql2LP6p
1MacHJ52vqYVqp2XXlmGdkWSAv0UWQ/Xc9zxgVPrJdWO4Qh+x7F6XuSNsDdIU4h3
QeFg7gpFnLLlF6f3qH/hjTd8PHWosxYNjFaz0EcEMtk2qnZiqrLFQJ3AqTSdNI72
AixNCF8c+yi68urWEY/VCscdk5dnzI10MYQH2Tn3edK0sllkwj5ONHEM0R19p28x
RbDVhNEE+ojiHAcU2ijNUd4N9jgKbSld6gjJz0c8ipyQn7wXtoBPvcwetf/odVFe
1yNbGwclPIVZp17E6qZEtAiRqg+5NiGMKOC6QaKhPYwF5e9vyb3XcpLRDx81K6lC
6e8tIe40zuw1OMh3u0A5PvyEPpQBPrAMaWHWeMr7KE030h9PdFGIcb9nZBdBtZca
It7vs5jY48KA3q77r8cD9kQwZRMMmtrweHbGsmvUzuU1WCK0B9uphgzK/XUCrpWz
xeR2YAEDdba4TBOVcsVCb7ihtBEba25xd/e+JbgHg/iCbDR6OtHdyf1XqAi+Hz3j
rx05qlHTtmmvCD9Y0x7RYSY2rlf/NybFfwNS72heS8pnmgb/YINvRrEShBgGxKs+
S4bFntxn88o7peIk/JvOwSjBfZvS4c0OySykRSln5YhGho2Ft/0UDUzXCUsK1M7U
23d5hQfgF1BhANucEMZU3omNemEUspCvQMCCooGclnUwAcYcLnMLNnQg9Lye24TP
eIiKxTc1OQbCU0OTJqET40kLFExvmkitk0a2tqLzsPZwey3XPXmov4M/4hpFb/Bd
gTYBdYLBFJEc8zNZbZPp/onCTZMQVdbyoUqmcrl/xnaTbbKDo9OhuloCvvAfi7bh
XIJUZGwulVPAfOR0HVm0aT3m25dr+Xwg5v3rS0TvEZU5e4Q8UW4R8P4BjDoFI/Jz
EKfvJYDgncsnkXWn+SgzpCY5jPfRkIyVb1iFRGwiRe2N3idtYU+Sw7rqNakcxfTd
XIeacj+28DAxjSm05a0RlNSembaC+z1lPR4SL+ZiptTjaAA2HqmfZsnyDke5VOmi
ReFDvGGwE1EUWZ3uv4slbPYBusMBKv+gDc9R1464nF1jvEdtaFlUFVgoIn/jK1pQ
7IGXaEObhzZVKfePm80zgpjWGwO6ARFPmEhAoWqkv5iVhq44ZukL2HYr6fgQWN6k
rBoCO5Msgogr+h+9jKvSRRQxn6dYGi29gZoCMLj47+DFb6gRLm0orGggvTBKNGyv
Tp2/8FNJvlSSmdYTJaY3bndqrxdToO4e9VhxX82F9PPEISo5+Xx7FuqQFl6fLnG8
RbuJ22Fe8W4tVoUJYD3o8SDMcWGD//jzf/E29vwttoe4foqoYfkHKyIoLMBRk5f+
6D1QMIXRUKDry/pfP3CjUWjsvlthfeSsBVNcH/Rt0lymTow85nC1+cjL3ztT44wD
VSFSO6+swz6M8r8ZC/6/sxK6z2v622t6Ruj/w0n8fJ6VBh4vOO8ixY55aF2IydnS
K0370yDm6/+ev1kBVUfaYqIMI9h3eU7qh6iudhWeSIJ2LslJ9MsnrQVD1eeqxBJP
GCsJ8dIcIybjUbITeBYtWbBP/A2OSaCyG/W1II2D1aakhJiIU0cH2yGqSUGVWt1f
kcOATMsUABRngVt0Uptk67VkQ45eQzu/rHRGIWQHDIYn+ElBLu2bHFJ7C2ZwtvId
3JUpJ/Bb/Phw/Ys9thKOmG76ZwjVsMaGEIyFRgP+8MeANp4ILvQBqwSXp+nH5bRS
fNWfAfNNeAgiNfzuQTuHPB+6hZXMHJAtwAuewOooylfk9awxTPFRGNitFVmKMsH1
QKPBwAoGlDhu94vKE+sM9hXCAGLQ4NR4KxYaD9Xk5F+uyQtymHB2dE2EVGVf1M13
gikA2fKFqAkcPpbnej+A7/0eLA5elT16VC2nBrN+voyYpY1khzdYg/SOR9SUTvBj
Y3GweUenp/AIpw9ahOgLntqWlfmad8BDNOcJta/0zKOdt8sNzw4937BO0dX8ae9Z
DnteNUPycz6IasRD8/hICJ5RYC/9goxfrB9SfKsVlUwGRyXNRO+p7Se8JSkS995z
dz/wPFEdEBxPkthGK4LXw/52c2YhtMENpsefoOZ35rJFnbQOVur54VRy/CLAkGBC
qJAO6xNrkDb4QyvejaP52LkGzjq4PYou/3/6IVSFxWgG5wVEDW00ZyssayRS9Egn
ccqF78n4MJHdNflJv88phpZZKZMZsGvGeOHhFWv0ImL1pDVdvjwAsEA9wMHRJsdR
SdBooO0WXTBooid83e9SucWY+0Tqkjn8J3e0a2ukrtVU8iA6qWZZCsxF5RF38I99
utheWhZJR0OYaXGE9syt52QEiJd5YHxEpGOeJUNQzTsz4I4xgIfclHgkeN9m2ynY
/7+Fi38FCoYbhh7XnJ03ZO6h7Wbi2PWuI3iYJPk5Ndoj7y9cEmyKpMddjWRhYf4l
hB0QbQ+1rm4P91giHZo23Krg8KPCjqLH69paku9Q3COFkzww4oFWxzWSucmeqhj3
/24e25BH6w88wL8U4PQFjsSgI/cz7opzwgWLyVS9/xv3mESL2zQzyXQgOZ+bD0/0
b9v9Mn1WpEpoz2ciGMp6pIrjqoVHZ9elrw6RUUozKptnqJkDrERb/c9hXvxf5oUr
PgWsiDdovRqz8261H7sC2PqRivZuQljOc0WDxGzaT8bY9AsP4M/bIbZdQBnDZUOM
sHLKVAkaSbIYvZjGHy/89O3d4En1/VK2Qaw4+vaqSL7R8Wxzy+uX2Anl+cJQg+Wa
ZZhP5Mb7PTu6q2cb3H4DLQ==
`pragma protect end_protected
