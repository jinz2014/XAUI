// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QuXCj0iE60O/8cTgV1D23nw13IhBgd9+AnPT8Qr9K9OtKWfSKwiEtLud4ZsQKgXz
D0c5dP28pla32uAosn8x0/kqcg1JGSsI2kB+HzCPeO8cxWq5hjz2wJN9acy5QFN+
DQst1lD/1Jt4tPAZ3Pj6VZW4oYPHN0OnIPjyOPMWkvI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15600)
RavlIXofV2DJDTKOf4tciWnlusufrdJ2WlYzPFWlnqSOL1KpAl/0GJrrTRSO5TJW
xjKR0l2S5/xsOryG389uWS1Zb1R9K0h5uaAs9CaTSFBPmqzydqOAAUWShsfT407b
d/Nq7yKg+7ZdHMRJj04DrET64+6llNNNARDLg6YzLo1EwAXGSKlM+1E2Qv3kAVJb
bAiFkhwvPsjfsbeGC0tt7kzdjPn3GSh9vkewEnDdWMGWIGRx23zLs4NI+7E+EJLF
tqpTRjY5b2Z35FPru3MEnp55Z99wYVAIZRP6g63dRxNAIt2/MTKIo9DrN8nuVDn7
jxXcU9f9ezTJ2o1etkncT46QylhTpIFxf/ZG2eKg/cKUqF1AM81VMytctNYv0Fv9
zWvGHA5570h8NEIJCAYcvNm0U6PclUYnYPvXgdQI92C8BKAwUz+pY+ECK9b/uitk
mfmApyMzoLfVbDLLyiklSk9ah+UjyTn5d/+WJ4GA+sis+IEFoZX8ErLoRIvMjlG6
J0W9+si/DO5Gdv/7XT4VjiclYgGgcTvIChyKvc32C/q/qzeUOGL9m3fmftAqZPHI
qfKkg1jJhxG/nzyxz0lDdXYMTaVbp5oKh2ZSSHY15BaUtHiD9WotTCrLULTnNQAX
l0BY0NgpMZpcNFTbdNHejwaPDYA6Y5kPEVJW+CTnJBksJ5fS8+mxgM+3lraw69iQ
OYhYommwrjzxPgRpyBJU60g1v5hoN49BXr6o/cZDpK4iKCsGsys1NO6mRgtO9pGY
9GapjCv5nzz2VuKDnujP0G+/dawfFM+0MkXcWgsBWESHhDakX/vi1gbZOiyr2fgC
bwUzMz5jwWYz4Lp74eeyL/ezKa1bSAnGuIYypx1v49+NHOdxhcHquLfcjE6EkZU/
exxgMJB6pn4cF4LbwfojP9oTXskQ9vwvAzwpM6cylV/WGmY5UWCoa/c+Z7Vt/m7S
5T22NY2VG5WG3lerXCQUBUZ6ZwNyNigzvrTNXYDDVQJ2HnWhQh/AFY1deLgi9tZH
CebtDUHvinkOXF6xmpdh7GyfQn7zWLpWN8eSWuu1R12rHm4fXqA2X29uhQqkxXhT
a2FryiYJmKrU9N23+MPhONF5sDHE6Hxt5Xgi9FMBMhAodqb7j0/YNdWYOkxX7tG5
tvNW0LnfKZyJJCHVRYbHyeO+MbEcI52U5pJj1OKWR08Q2VcxQKJ6fQja0kKKAQ2Z
JqHR7fsePCBYJ/SvZfvDFGxVWnY5lzsIbiwQoW5TR0Y2V4ONSNmNKbv9ha+zi3z2
vQzOM7g2hj09XxGPgtg9UDuCKkVMX05pT0ErbWH/k6OSo+q096jV7Vzgglw4h77D
p0xqag9GyVH8V2JrWD/g3HVEiwZMjUT+Cg8DA8WgIPPF8mLlViBbqG1Xr72KQOLW
tvfEuG8NechbfXIwEqT63k8PNtDEgcQf0oQNd1YcTei1QguujQ/ZCzHr4HoVHBJi
ZayaCFd/IdOXzEN37ACJlV82XMz6h4dyhnBs3Nxw3LTwEHM0tSJS5gToOYjY56vm
T2limLjiHV/IIyYWMJAhtIXhhu0FHoPoBjYYKjZknoxel+PwTGfVT7eylhAV5Gms
2CcsfYXR37THw5opt2fEHdMs8AeSiQAxtIZQ1SKh5Bpp26qmwhpL10FbbRWbVb0j
viOXkaDC5VsOmAAtLe9Uq2Czq+pko12Gpxp8Qi66ggHkBtLnmWuQLCrLiaz6QsVK
8tgvULaKOlToIFmna3hA3ZB+YkR6TDNr8zIGuInaBMcdOpSI0e4VfNi3L2dS/95k
kq5eSCKo2xoBILHrgchCpAD+ixotwSRaAdsFuWoR5isV4bMWIBF3+Ns50hOR3tMK
ramgzQdQwSm6efZDktQSD6x+1S0ZGr1yErNQm9bIKIm2JGV522BoK3thK8KMICNm
DViMKJZz08pmL0m96h1NEMQlUnqebTwE9yb25Nf8f81t6JLfhyezxmZUt50NQ/+J
EXbQakm+FtlQpudH6A/Xa/N+HhIYn+9KxVilmKicXW+o4NAcDpXgUwYm8VqElNB3
xFUffiKe2shWrxiHcVxdH83p/kOWADiNjrvsxKO4znae2ThE14poNKgGYdBgwnEn
MJDcZdoFIGrvbSuo7bMoVDtd4VFIT19vL6XGslDiVCnI6e+D5sLxYOCoVYYR+60w
IERwzVDG1ZSrb+xmrtsRbHP1ZG8I+DIQ0T0IvYtWQNnCZ1vJxa0Mx1mUSfJOab4x
gbXB91DomxhLCnBMP3kdSUkeb1pwEhrzUlPexp24w9hsl2wBWoW7+sAObkGTBVjL
myrg0J45KQSYYZaRC7vOsQd9dejqJgt6Tr9sGvKsWq7/qymDiPesUwF2lCPuYYcK
lLj2qK3oXktxeTQZa7yhReC2T18NSXjv/0Rvd/VJN/lSvtCxhvviKiwilr+DXZk8
59Gs6jUeKa/lIp5LDb2dhfmYb2ODNw+ltgsPVg4Qs4KixxeuCciVYWmXcclV8D9L
B/PFo82NvHrjNWEgf7e/5ypowqfC/2B3zzkEP6zZ/LOoOOROoNvfKvHdgARURB8b
nkIZoN/gSTFe8ZM6J6tSlW2Yy4qfJ60vo5Ce2/6Fdx2m5gnI5XGQB/U/EvjV96ig
8jersD0pzqko6XB14RxgoBgffR/Ip0VnW3OO958CaRDYk0bvG+MgBg9N60QnFMiM
qv448aRJA+5znEVJACyQMqvNaPHrrocNec4Zr4mKoP7pagBu86NxjZ6seNujWLfR
5ufJTTMm0Zr9Ys/CrYy30+L4qD+2MRfH4+P17jmjoBaJnNkPBaTGWuDThTMbBeXl
T0PoBS2JvKyiyRvVRlncN/SXoyoO4WkFzfmrZL/FhI/2iEHb3a6Js6RKJOoe3pX8
cxEzvXYw1/mJisyRmwG1gSy0wCizsiGGJeHihAqzuHgrpLL0cZWk3/aAJX2xygXJ
OOSDowmksOF+zlxsKzpcsLkUVUBEZgTAHtah1DUZC2F1CqDX5Sj35Cs+cteaKX5x
rm2pLTp7UfKaAqdmFD/bv7CeBMLdc+99yEqhlcyy35Ui9BUF2e9Q8o3MYrLPp2md
9ya+EhZf710Xm7ddyOLql1gkdWwSlCDEoevB8jN92+1z4xWT393AAvYO/unQIqKH
mnkc3v2LOqkDz/oaeU89ka6y7Xr1I0P4k+mAwutx9pFz352aAFEwKF4NMy3oAtwq
uATLPE45fNHWutVWkHSPraZVmyz1QTdK9MQgT3GESw7nmrVuOtKWm7eAz90iBXYt
u+86K9IfMbvWGAek0jjN8c6Sg0s8adKUD9zXEgWKySOWGAsi6ZHWVa4Ujyruf387
V9GHS1yjsJcWQGM2EAEs/rh/aY2HPCOhV9AhErK+yvLIZAroQa0EpPrmjpDG4aP8
OWoDzR4qalOy6cnXLhclnFIZaAD45HAsDA91EnWfEIi+SzbkRDDq/xQb7PEKG4p/
alehyFMa9icfuYSMWSEjxziJTsn41KGtYYvZ2/kzUnmlUg02PIKNDXcIM2rOZARM
A3TpX39AECruBR4PvffJtj1jIrwKqFHC+xg9AlhMikCGsDQflxDURPzEooZcgU1S
pB3wwHat6yXjzX3WsnnQ19BJPpT6dIhhNVcZ8XilE7GC8f+r06AVQXiphitLZiyN
69o3L1yDAjYSx8o+jlI9mC9hwKvxhkkSkku9v+3oc607GaPMlZYARjZ0IyyoNuzl
/Y7/BHZm4KKp0yZKFxODTq2M7vIDVo9bZD8dZQNwAOjBjdNypzA+UwYGt/+BXWKd
BccFfJSzoYaiJgxNM5+4jJh2+GmpzQbOr6dF9INF+ZCcCSbRlp98Dz7O+ip1nXHH
48NcohfIKJkYcLsrLZt5vcDmxef3XUullIqjNN2qCgzycidnQcK6oGNAwIu5JouE
UDssKW4J0Vcv95dt2T72S8Ry1k/xW/IidoB/cdSl5Q29s1a6E09GfoyOJLGd7EYG
MuEuOtUYE1DuWlgNs3e3wDMTUbAFFmO3za4XPaJLtKbUQdm60FGwlXVHZUalLrah
TQ7srVwyzNDCoW5UqxIIXRMmHwZxh9/AklP6xiwCdDx/vKnS3WhvEife8ODX497O
TuuoziR1S51ztl9cQJN9MK7YDaJd+cAYypPQM71RBPz+qR6MOe7ZIIMWF3tRB/K1
58UnwP/5b319n/9ssp3ytBtylQRnmlSwfYVp8jatYsNGHfQZyvnqGuhIyc+SMwfX
tSl5K8OSFclFrh+5jAasemvyrV+Lsh4ndGoVzHpHHIgNC/reP1XpaWN3Ns1+u+yo
EW7cIAMzXqQ+Dsuel7i+Pyc2m2dLuR25fMFcQZH90GUXFkifkYYE6X7pD2M7sH0R
CByUJwnzR7rd1bPo3fRHNKIeka1cRzvPvaj3pqXF62zTL/0NAhKuDDHop19zv/Qm
QBivynxGNE90v5PbWKuv77GC0j2NOwNa12m9DKfUyckGkUG+XI89nLJKmA9EhoOG
OluPOBIAhJ/QKAOg5vP4tPR/4pAX2lTtDnnIJpwBJ6DAqcB2Eb69KRiiL1caI6mR
Jjz7lEOogeU7tzqDqZJ+UgRlIqkUvOqUOwhn9ONc6BhHUzpGdL47SqYiKDA14iWz
UsvvjQmVCZ48kV3pTiSJ3smxyNLKjTjWHysGZYBIgyhwV+6/MB+4SH7KOQdoLWJH
QATQnxCIjlDLkxm5md5Az47MQGAoGYlG/DrhfkMQcOVUXFGCSxRGkWJVegk0dljy
oua4hJ/Gsj+eBOzLP8J6P+W9wkhz8FiQBTahZTEqvMll290rfQa+MgbyQES4n4MB
HIBj8cmyl6Ow3+sfQJKAVqeptVK8mJZ0HapPlOWMHqx4fLvf2tcCMtkEhz/yJnxY
7EMpuVQVvyewonnAUoLzuqecEUpXT5dtlOO6tOb9Ojf3aNYRGY49UJo6pIqAE/S/
dNhgxkiL+KKTmdsyJEjpbQNbbN2OUczeT98iHQc+AZRavmb70Zo2ZcfRrhM5+onB
zW6NhjqswQwY42g1NvBjKku3nsvn+h9jT/z8mWyTqwwJAdt0ByN7Vb+kp2Ir3pNV
7KIVUSShkCZkI/T4r30jXiVs9N29SrH6zzQe9FCf1u2eUXI7OFSYZfNNj9/KAD3B
XF1Ofr6J6O5J9GZlMTa/934roiRrCF+Tg6qSlOVgkTVEH0PfsTHODYv4Ul3t5Y3u
RiQrZtWu4rMf1MlfIajeXXbrBHF7xkeXlSUoqFF1QigqUfEXvJWBaPYA6zy9UI76
sQPdjjJ6+6ULv5BxAKx0Q1J6D2OZEjojVs8kY/bXT101uFbyzMWX8bmgzmzc3DR0
306o6nvFAil9h/qqBoenje+55q5bNQCMP58fkAfkS3RYB4vdrgsixY9pIHHVokfh
3Jx1ajZNPtBAcTE2Mnu3tX7kJzAld9xHAyMbe9T1GumyZPA9JRKK3V2zNzNL+Y4i
H11sW1gzyAVu0TCgaqGEKDamQIxIPSayM6CPOlWaijbdvqdSHV4IQoMOTs1gr7Zy
VL9OWUsBFTECria13uZ1V/xE3cZvWbVlv4unzKWYP0RPqxs6Z3Q8Tt4NIcXitwiN
KxZJQFyMmwgebTWGavW8aZCvQaH3AXgm+NvcM7PXrDo4nF26no1buoakglMZ1Xzj
ZHbP3dse/87ptgss2zXEZcKFefn61lhKmUJoYwnvSNDhDzYlZKK9QJuF697jv3NT
xJpIVW6opziN6I66jqHLaA5BxUTLbEeZwx1pwNLJjbjxROeyT3vn3yi61ojP7SLX
hPquR3yTTf58dksoaGOQHfzRr59RkFKhKcNat3kIIRVywZVgFYJ1azeZH64bq7Rg
Ul/edvPpKv1f2bbFotzV6AfLaB2Wk+Pthq8KJSC8pxtYKxGNoeMTwUcsh/zrRkSB
8e6lenVb/Bxdatfl799r8GJx1OdiroXBrM+ANEDVsWjG948zoObDgY85qyUKM6dZ
wJIVSXTiNeRU7+TB/5E7+YfGIlsAo688E7sqWk8FQdOewICf7Yt+8QAyusZBMTjf
cHuJmGk+lWRAitvEYJjSmyrUbEiPTIQy1KeZvd+zA5h5RNvGfiawvwaKPPVogYF0
YgnTXDQy59htDv2t7f4cvsf4wyDSgTXg55W+3LT8Flyei/jJrUQMNjZhn/rzK5CQ
T8BGeJQKtIvuES06YlGnAHoAHuStnrk5UQNmUKRh+ER03SZlffJsQPMNmXyK6pTX
MyzuFrHtBL9kEKlsBBhMIhfY+lK71MUeJv2GMiXEWNMIlKUwvGCba7dXv3upKYOR
iXTYINfqIHtHCgb6SY6XX0Cd/mex20mokGF6qZAt06iFkKSsuiUBE2rtb/zl6OpS
KF/8Ya0dp6tTAI7f1hcThd/xQWMTLInaFru5QO3UAW7UK3QV9yk4BW1VL8P3NjsJ
zTTHsnY9n1x4qxi2hVxUMkEe7KJz2CRMV4OHnV354kreJ3QyVYcS0sFsUTXJz9OO
TSSXFv9K/PxKL59L2ufF23oQSbZwIxHTVCysF5OPqXvZraa9+ReOiw2KN7WTHqBy
975EQz/lcBogCd+PD5swsqBxL5rgSvTaerlU5pBOgzIPu7CQvD1cW66qp4L8AqSI
NfXs2p1iDa9a2hZDH1wNqLYj18o9NoGAze94eFew+chvvoOt5mSIff1s6Yo1QNut
MIEgk8TC7jXHF/F/jLVKNqGnun7OmkC0cNJf/g3QgYwtebXnTDBc8hJuWHhEaHkY
SxbuwzjfcjEuUcmrdx+eqGJQCDCk4qN+2bS/6ZeVAhc9TzO2Z5mRugoxX4RRNdE/
GlTyPa44krop/WRikdilUKBcAeuOapJmt9ftFqSAaxTYmYtwatpeIRM9TnV4ywbz
xy/TXNZPKEmQ8DDOK1YjhxHJhUvEu9PX+iXjduNAmC0Rm5V+WQXqLlAKUsFY6tKh
uzsFN/vqL/lhTchZpnH7vdpcQSH/KUquPzqZYHeL3V7c3oXJ0xwKM5nGoTEEedHs
T20a2E3LuXJtR7VBFNYUlRMUlkI7TZ4khmxbVRztNALdiL/GyrKLS43XXbgBkNA1
jV+xtNMFp4oOqxGDWUcoBvneFUafGSbtja6IIKcMYJAc7gJg1ZgbvocntfHGdCRN
N0TPAI754pwp5xEDECGXXe7WxHFaL6Gk49fvRfbIZojHrWECdDi4rgcBso0EXpCa
AUzrI+oW+ALELSciS1kfw3H1xIfqnf7QRy6th4yBaCxNdmxMowY5OAnzqjemQA6d
pwIlocB19+E6cWRCL24P/OlaBmaKsR4uW5+koEm1mnY1YAI6uZScibLDFEFfn31Z
hQkeNG62mjtu+QKa4l74JBeGqTmQ4rNE+1Zetmzeu3TPGa98bG2Qhn0Qy1H41wbQ
VajY5TrI+AjMnt5hVxgLviZVWFksilGXM+tNjzp494Fo+z7vyK2eyrvtjLIYAJAE
UEyO3tmiiINaj1E9Quo9HNk8iy8na2Ef+W+lyg32z+qJDMcUEPF7+eXH+mhe3RY+
g+o87G5RV2psbxOcd/Hcz535yrrLeeef530hEhvXwt2ve1hTyFCPapiaGtwihIwH
mu0u+otK3mfHqdPM716b2JrDoSdponbwK+m6Gmlozxn0G5rLg8vW0jmzMIySqLVO
2HwjwDcNuhMwkwpTMsgfrQnB5nfNE/qgVbnim6FAysABPbFRmRCqpR8BJQ1CHUlY
cbxM3qjDBB//NY/aauJqKObPjsAE069YqwEExeOVGNlK9jPgjuJvX22KynuAm0aB
05eD2qzybA19eWdG4GnPY6Am0lbtzgqtssbL/VVcufL+4h0pWv9yTcULjInidVnn
Ilrq5B+zoJCkrIYbGV4+k4/uIm8OdOKaHV1WGEbG4yXGAx20jJkZO1Zj3/vV1OCK
kMdfePz2qgTwKbQcWoA22cNqyX9BGG20PhEwAJFBPpc/TqoLrbBIH4ECcFGgC43b
Nh4A5lVj62Vkn8NZh98MW31CPIjpxEAZ48w95Mn8xNXOj6UN7ydpsNMVqHXwlIDi
JCANpZfpGOauXAPOYVFRwvdorMSakl+WfNWcoJ/yJdRifFvZjjnsKkK7VHFiBrQv
40MHppDXC2VxTWq6pxfe5CLh2Ih+D5Mz/1Fy3j8cWMWyADZQuZIurMbuSHxuTjEd
kckxebVd1rlZ/c7x03C1h87gWSi3XLLwoYuNEX3GLjI98y55hBxCZF0Tsihh5utP
iAjQIqh4fKzL0vA5pVyE6bf38zMzcbsfIHI4+ZwzkaVil0OlKa7y2nh74Lxf5ou1
BRxeLJ1P+zogdiO4AnPkF7CKQ3I1RDVhnt7aqw5r1TcjHLVkggAZbJE8A4zZea2k
nEEUMAzHL13FCtaALyCXlqaDEKwBUGBdeAj00D5I/pF+X/wEJOlUV+khLMlV19za
F6F9FFtdUJ1PCuKp8Hb/zFQioQLv+UEW0TXdaT0s1LL/HqiYP4yD2abUmHVyj6KG
blhEoLnE7XlvOfjZYlYDlN+lDqy3Xrl3P9Y6I8qQKxe4bim3vaXECyHnRflH0PiL
oSr7yme6PhdOCAwbkz66255xDizd5eDwENXZk+VH0PgAdwbHtfghTKFaMo1eL44p
VTongzqSqG2g5WD488Mf8PrmMVds+zE3kKDi1bY1P/RwB9hKE1RB3UnNg4bsvbs3
cQTGOtWlS7FGkYYphTNDKFUlBLKeho1flbPq5ne3f4CoCtUFNRQvXOSRH7nvJymN
HWbCKToJv9hBIzICBAB1YruqbmxbOTJqiwiWHEIpJTkc8CgNhAzy7GPHMk9/tG/y
vy0XZFPjb6fY6nNPsBWNjeiOQ0WnNnp65e3wJoDh3ViqRwvVYPqwHIUMOd5wxf8Y
6vHm7DFFlZj0To/jsy95a1HWOVocDD2nz+Eym0hGaIOSmGamM90Z7Ob/fQQ9X9KX
kRw3AwvHsZLO3RQlhIOydiXeaG68DaCY2F19RMhlV6xCU5UCtafTfuubX3euv+jC
cVKPk1cyuBy+sMaQljDI3ApUjGQzJIJqZf7ph/AAAJVuBQOyP0katzqA+kkZ1m+X
i8Bp9TPwo+JOV4P0ze+WgUm/2REXJ6nXcx/2Rqdm904fc6/SWnw+En+1F00yloT2
zwmgcEpqC8SyOL/ySkq9HD0nR/qeMaoSAoitcA9X+gQP3TmPHSQtz2Dyr3MWSPf3
8XwV0Jn/qe7Z7wfO6lZti2VmhfukG9yeB9tlktPDA50I/DFaVjzckuZZb+zmN4kE
4qBe5h6UJ+G0Sfr/KNyOK0CpCgxJ+0VAwaPIkCj9KTNEi0+NCdHBVVUs4UOOJCss
QYTjZLrbs9POEykTjs8QO2cOt1AyA4+s659tbGgTDduNu5OUvFnqhUzp+jONHBqK
BYiF0ppjFIy48ohIPpRN/eEuv7oaDsqz/cD4eW+/f2E4wwDAaCpz8PledZmCu6Kx
Q663HdCNplMFpb8EeKPSN07CiQf8Raed7EJyQii932SqcMd2EIw/isczTVMhCmKs
ge+fd3gtHmKGuL1+LZxk7FMOANj6fSpop1NukFXS5w0E5/lGHmenx+sUkJxUtoI2
wG8F95JlC1DK2w9rWDueYFH+3a4QvSeoOsO653bWRw5gm4YMu3ciGpcw58A6Hmf3
aFflaWQk0+eG9X3nirm5W9bWFT8cJoHn+6hhpm/JZ8mySQQbZZSgkk1Dvd+99soi
871CkpbPqu4LyJxspz2JFcqDMmOAwLxsaGmD5EJCxt9mD3IhiYk5KTOt5luQgls9
dbCa1hM01SSrUh32QtZf0vnXzenG7jaWQMLmhOfNrJC2KJRE2wOPHl5LdJJzsWXV
gtSEp0TH5KinRySPHY6Yz+WEkgvGQm34SlE0u6hG562TCj6od0sI54GqlfczOCsY
Hwr3mxnKX+Qdg96yCzvzPu9B5dx0zKzx8p4tjp7j9eUQLtcBGcjj5w+rIoeYd2+T
6D5+P19BQZcx3NuZV52m0mJ4QAGsCWHRu3XacYYyA1elektVzwrsP8evrcowRs6n
k/Bpd99dGmuCXTpnZFirKXXCc4N2AZIuxEI8RNMBIRj9S+t3FVmcSA53c2149JoY
nGbOowuUgUepveQKsmVtU9cbouHf0LOxxXROwFF4Fbk7NrSxOT8ku9D3NqNbXJV4
UGy/42hOawcVJQ9yYoWZmG51r4li7sFb5lXs5Ey5SgyfsoC/IstknVtpYGED1tvm
19MDQd4yLF/wmy2GvbT7zv12s979OOPHoC8hG8bTYkrjXw9rB86iWXJQ7JguGiw6
OhdNFhd8E0tEW8L0UPCuFZ1UoyzQzjSQkZnvp4XdOpAz6gNUZ89mx1AvdxD19lmY
TjIoFwEUUV9MSBJpesL4aiJRjf7yfD2o1WGqgtNkK/EvPQ6x5RtIznM3cQooK1SR
hyHzbBV/5WY7oN2oNjCTv13cH2oAvyBHGUASbqUVWtZu9vWOMTFze0VCOL1bbVZ5
/3RPiA5vg0ISO06OV+6Wn3S709TCOXQRLp4heO5EBcHe37cwsIFcPDwRnUNme5qf
iFvHTQUKz6w4Xpf85Czz+QsEa2UlF9srk64akN2G6BnDzf9RZpMrAWzHjzr3jH9T
uNCWit/B+Ds4IR7E1JHy2Zmvitmfc4LUJ9Ep/rsbxSSplO4v1/iZi7ACfvPylQWZ
mU+lOXjfn9iUjBFvY1m1l3msvMHCKtYVwF72zzdQS0/RvY2rt2ao/3W1Q1w40QoB
Qvp+9t/RMR0CkIczVt2faoi+/KSyhlpBxeXp4hpeVNFWfBzYO2jk5/8SZglj/BPm
9OxM+TCzjsFVJL7m8KyAsfswB6Vd+qaSseXQiJCKlGKZSCNZH3cWSkJaECY8Qsf5
jdj7xA7P35QVM/aywC1+cbLTpVUGueUNHPXtUXEaMvG621ohv2Duo6xYFkoJtX5D
6JKm6sS1jeSkkvNpmvx0JIrBhDm5Ceyc5NfPVYcL0KcX3mTimnl7M0guYyG76V1v
S1Hp6/9cB76c0hI5L0fuw0Ti/kc3nqUwrtjNcjrWWCjqJ4GzMWmipKvOmZth1DCm
FiOCtgzthtikAwkOneLBc55xRmpVgMCefFIe52RaYrJHCwOmS1npKmoBfnAQGbQW
JUUwIHDWgRK0lqlW7hpKntG8ZVxtApzH8M2/RmAmMziZSuKuUXSHjYVSc/WLASW9
MDPrmwClzl9g89V5DUf9abGobbSXDNlUUQNZlXuJn5T8I2T4uO/2lKVeuqGtTkd/
/eM5mtrRcC8/2CblwDdrfp9/1Dg7a1qr/AC0GrfrsTf8NSAlJo2n+DkUzgKpfwfl
pKYF6fun+tiotg6GiV4HHWwJtPRLtJpYnwcjHz89y4+gEPVwGoTYNUozSgMgafyl
iOmOJmHBiDZEozj4wT1bmPlGh8szqfxgY3Xm2xsbzUmfQZSLBShXRvd53ZtJ+8+g
uxxEy/arbza0BMwNVJ8PD3Ci1p0FqR9SRR2rJYQuH3o9/K5AIJd3e5thxBfJUoS/
GpcOsgHi4mweYhS4FKfyUeC6GF/zZn+AJxI0QsSwNcf7zD6tb+zkK15o6ct3jpVO
RSSTZ4+pCzEWzdg9QFfGofRsw9YSpFWEatllr8g9bYlhz4wGiBrA05+8U2lMrDi4
ECbHnR+ykJkW44EzGR/VTPSjRrp34hQF6eelmDO9pLxZhKnUaFpNQkkNCL/sS7ha
4r+BcYFrYorWJ0yTBUi6U3DiEyxg5iVg182ILwSXTSxU1Y76hyNtzuaODkDJ6Jft
PTLsCaSEmVO72vtwx9BnqpMTPAOHL8LmFG4pq49Wf8QFIS2+Vs7OVc6pXZ4+eCSC
FZtbkQssDArcYgsdgfNBeygSzaqo7PE1Z/H7eF11mthhV27PN4shX4UqzzMxSRRQ
N0n8HtQA4IlxOUP2Zh4caFCeLuXX4RyRq94k7nIuowWdJvC3J7XwIrT7/zIjMYXT
wGC6DsV/bTJ5oUKx4o7XoEsN1j2on+YPdZkL1UfN2uqievtXH1/fbalX87ZgCWhy
zNUTlbISy3abMe5CBuu9EUCJ73bIYnx711+aNlTyz7xnAImOEZObMFezHGiZZjQc
+aDS3gtdX3b6EVr9P1ya4Ui2Qlhm1ereeA+UTzNZ6oXBdIMUmo5xDGpBkK3936jz
lJF7chAU4R0DD2hZQGcWtinfzfqH0kJ3iHt0m9ZMu8uMEQVeyr2NM3MHFGWBRhnH
qW49MJ3F5+gQ4teLHxgLZEPYtr5hAk/xJR6pRI0AJAr0t0wwwfjunA8wwzXplMUi
Q+aI7xwQleeRfl1w0kBwxT+ubGoKJrAKDb6QWAj24FB8JvsDBU9/p5ANIGRGESIn
Jccxv0/T3rs7W9+YKp/wPkqcump2k/TZbP1Oq6H02MP2fcolE4ptaZyike15f/mG
kkkfmSDNSJaH5mMpZtKmFh9eZGQGE46mPzwbK4Xpow3c9RicEqBPd7VP6q+QN7Ra
q1vbZ2rzscm8LxixjERofKbBQdDQ5aSJvnHtCz4cTMGPBGqQaWdWQrld19ShWrUL
IMGPewO/4nW0awXhIMksjTBq5DAll3j5dbGulcF9COjouD9gTqCRHVKgq6pDSjT8
Z5wEJEQzbMoPDDNlVGlhhG7bCTUMXRsEb6kOZzLrfQhAl1rhiKdJZVU9zBobSYHe
dt5j9Z/4pViPhRiYX2eDZHxIOHRfJRxGmCjlhiv+n36R5aQQ2LL2AHYW+hCd+xly
2Qi0krXK7dKi5x13XB44IzEBYzM6egZUQyWsMCDKg40i8LPjbAWjvb0PvH5xMJ2Q
JpKJn2k8VapvRlpIHQ6IHzhKIBdBclRZtWIwMA10ipYKHDvivyBgeCQtF8UON6A+
n/nKgXBsBqllKM7HwtN2BKU5/HrEdcUKG2xwaCNbVDm8Qo2jqzrNZV5k7+iasius
GTF0vVS6Z9CnzRie+g14nmz8sxq0ZWHkeicrBNt0rbpVtDfBBjfdYPp42sMEadGI
m5tGCwIS3bVmlJMSnl2NW7W6xBbTL5zx0UYjA0HKJG7z5OMcBP8yV7GzWFrJPAyH
4sL6e6r63ptU1BTsE6jDOG6GDVKcDRxQq6IRlfMSnghx0Q7P6nlZi9+yOSljiHoc
y/jXMQNmZmT6y8dYjb4vhffr57C20NpfnzYBqZrKl2dYrwe0sxiDXhXZW51HWkut
DTfNKup9YsFy8zgwCdsQumGOfz0dj7eNYt+YNKIj4c+mDPyNot6E4/hPqjtIjSvN
kVh8VUjvexNfZbjNbdo8/VVsFpSx5YYm1BYX2ppQHe87wEUude+/llHdtU8/LhLq
lU42C/hDRXO31N2pK2VjjM91Ua3BYNm6IAOZa+3yJSymf3GSDk8enkLGNqhMm/ZN
upF41jUXhtN0OVs3wfD6e46Wi0tCh6vWmmqZHLsdCk+Vpvh2W2oREVx5JKAaVimj
7SFd3uLrq6ploe4mOeSQIcXrBx78cxooBYymqjYrYfyZEvCe904IYtr78dWRB26t
bsvOZXEUJ9BMy5m5Xz1gIMXNopAp+M7m0NhPMXQGaulDv4dsL1XpaMPoicm1Yues
fK9pVtVITK96K1CFGILwYSP0Udt8LoMXH7xBKiFTa7P7SttmSiER9VQdnUG4/pGF
lBJbPHDKQFfpZ6SRXqDpYx3euLGECZZYJhr40+h3ySoCHvIDuAGyIKZGVHqET4Bh
O8gTDsWVMJ/0rvMo5SDxRupu2A8LHaMI4oFXFVNsvULre37K4UtAiT73jLUoisLC
yj9/QZ8UJ5sYZXpyPN0UQaSc0w612MYP+fYrqCR+UKwUl01/w1IZjHxwrbAVEyGV
yqjo/T1dsTYdaN2ABmkfhxj8Bb9iemt/OP2R50TsW7WEzRDw28f2tKn0hEG20k64
3iYjEMY0Vov8y5v7szbN3zEZ69NaYQ9aNjHB1IWUxwF5Qq4XKU9ZC7Zc9tWfJx2V
ldhQIZar1FA4qOzCUqITpAsMk09LEXkGDItWKn08EFhmL7uRa+ZEynZNHebb+8ji
VTRQuGoCYctb6uLsJPz+Z/csnYVVIrTS1Zh0g0wQLLDhw0bFvW1YEkl5xOL80RtH
CjWZ3Pt/EYSKA0JMZRh9DW4h9GdDX14Q9kKwJOv6uQAqeByMEQmTIvgix8TnkqSR
tzZa9EeyvSUordoieeOmR/JvYtZBzDdRbIDE4szfUz8zN9JivOIY5BWdVg68Rl0g
C1Pk51ekmndnyZKkVkH8lIsB0FaSXPDXdNlTjKC9Q9zzIz3HHgjvBzafJbG59cSU
stx5zusS3l0aMy95LW6IObOrmL9MRpXDexSy0dcCZ3A/9tjVLNwwemkqOEGcJlkY
5nZZ1lfYoBkUDz8SN0hFW060BUcsDAaPw1btv3FaephB/TcMCHs+ZU92A681fE0V
l2GvRQx2aF6ON08Gi6zQABU9Zcn0N+RyeFaUX2YE5NkrVjuf6Eswx7epg4gGXNaf
6/AUpgG4NO16fTwws0/vgRfKExlxHA40U9Hj24+uq9ZMIIPpAuW7DT/Uv4YlUQw6
DZ7FbXErDnsCA9HTY4v6a/BQ/QJYodZYEXLZkc4hr7IaFGiye0KtqqLMXFcqe9SW
YuLjLBRRKUyCIC0cUVsEcGid5KG1G3wrcW8bwf+6UsdAmSB/Zhc3jjmJcM51AnEC
cDREpZbMrZpZVB3BLn+s2SUBxyV+RR4hQaHaHD+N4keWFtRijQHig0iu+vRZBNAf
6fQwyljKUga4gbA2/ZneV6Xstg4WnbeH41MRJBBQVSgEKDvcBf3Az8AHwKCL//OL
AsQ/uPfR+yn1r3JLxWcT0thntxD4VzwLC3MZ2rwbrx5ZzXDcCufhY27/yv4Hzr/0
T/wZFmxQXl3kUmM01/Q3yu/ZKImYv0b7mZjZo4TFLXPvLvrvmNG0LrRi2XN3VFsM
SQrwugVhya/GqPK6UbSmVcn6dT1s8UtHMmBVsD39uvDlHysbQ+f5cFTazutJ7lko
SzTcKoLT35fZAfy82POXWgzTC1rpz8NRmfjQFCxN2qQ7jLEhLyx0PgT4YwYcKJof
vThu5mrgqy5dPg05hB7UQ2bCMxuXUa3egYPjIvxMX5KLvM/FMpJkk8TX7QmGiIFM
vrR8MZ2+Kr5IFBSkhJy02FuHr5U+yevGFel5IIPlxDC1vPhMKKxPD6o7TnSlAGw5
NWa30yVrlCEI2GsM9tBj68RGYAJpZbx3+QMx88t8SFWAnkjNioTM9ZRfu3mLa0aV
EYXbj1JA1gDh6xluQ1cWlKGdJj99Sff31m6lrS25kuArFus7GCudBIYVlL9NtRxw
UbYZqcjJx5/xyjJg31+6TWUNY9w97umVEpsv+DLEnazGdwF9LFhy3mGUWPs2YE3N
GnxekP73/SYpKcEtATRQf1X/imSqnu4EakK4SgWZ/EnWXmvUGc7WPMIOpk/eh4/n
8IttoijYVdtTDKNdmTp+Imkhh1FssAux3b1L9zn0JlQzBxPpv7/QCxmTjbZ+AsYL
S13N+ldfgZh4R8ITgzguDqDFdFAoIfbSAELqjVHJz0a5XZGDLDwZuWDd0WelBPcn
kvg+3Zn55D0oaP5ayNpXqjKgQLEEL+1gKlctdAgk6OI9G2qGOTaWzYMpF62NWx/k
kIzXxXBbe6y04E5J1vV8x603dv8iFFZPYtTuzIjnBbVUs3xOQ/nzqbx2H902nLa0
I+iPaGONGlBgaES2LbohmlQba25QTCO4Asvo/m3rKqpJZSwSDqxVJHzb/Bd3/jg1
vLO9NY7YR3lpvuI+IiXOeru+XkOTgDn4Kt7Ls8uO9AtvxSHTZ/6w1VEh5YMANPPO
BbTRvHhREi5m1z9ZNESk68xTSuRXtpWw3fBafLUE7qt1BXMwhEyiSK+NgN5V6Pgy
TFkBmdxZz939u52sWeFY8bAQwmobMqoHvy5/13HPLgTbqW/uDYKjKHMfjL/v0L+E
OBkGF3WJWnGXdHqpO89PHq0L4RDh5zF03GaEeQciX0qW/czXLqzd5o33jy78R5YJ
4hqxsFo0TnTM3CpgocfOT9Js/WW38Ji6dRbAgckyoZVI4xmXqlA9RvWAxUkmZq4C
8/d/viixk2mmcxSxriMcmShCX/QlJ88xomBTCHtqwOaZTxeQNN4GLLiT5EqXWbh+
rfFVcEDI3/RtTKuUyViuIntzbg86bhLvDIZf6Tf1m0mPMix78YQgM3bPDAgnsttW
X0u854xx5u5wXWteeGx0YYtQdiEkE45KY6tXtuDjSW3Tu077b4giQ65D0xNVZ0YF
5P9jJMMM/SvefsyuiOK1ktxXLs1H3ZuTPj0SYqL+BquGgi2t9PGYEM4dIZhNk8NR
59dxF6GlP5mBT88MuppCgc5UE1S9o6Mh5PArRjaDenhL+naejT+yc7y0hRIAi8Ql
RqYWyNmJWy/+iWeFgfgv1Q5yMOE/wPRCjIqDGwLVPm7WQiENAn+3YPWdIrQmCN0F
ggbH7KnFBh73KxBHPpPMXRa5L1uE0I+IPxKlHuUcAzxp9cyyLGiVwMNkS/juPkce
ZfS26pwX0pISGMhEyE1OyLrOA0dHv46Gksfysog+YXd9GXSEXojkV2Y58AwJzmPo
bHAtrpI+B5DQ8elBLmjvHrJTL29Dj5+ru3xH9oE72WWPucKE8VvM0uWVomScpY6T
jJ2j1bQnzpLJqpT23kEB9u4zAB1+4gJvl2Cu1H4wyD4O7RAjeBDZJwoEl/up1Fpb
gmr31Wx3/pSf/6XEnbo/1vUv38I6XsUcxubtpCXzi1riqzpfqXVmRX09Z0XKUUnu
qehxt/HJactRxmrmVGfQIfvWb1nwQiYCe6805hyUv7iST67fRkeDQ19Dq4GNd4c8
fifLrIS2IBERtUQ2ZMGDf4StwrFePWiG5qfKkNxZ/+TUDzM99b6wMLW7I0FgcgJg
92A/OCmQ6+zxUxeTbmGGRMB29Qmh9fm1gxGw/AYZvl598W3S6efx0Y0dMZ4zZHe5
QhrrDFNvWhkuIZDuzWBmgNq7Vac/KQcyGArRJx/X1sr/gb4iXfoacOlomxYJ0/Yf
aSXWgZuob/twhgE3nIA5jNU6gihjBbnARrDMRUAnDzfnOZK1CxFqnj3w72dcgtBy
KDkAFbWSTyrKmamASOBX1guCEbw72EF/UeC3JfAflLEQUGfYujEPNJoEXDvcBObK
hZ5b1Cj3wUTTPfyRyZur+2gBieCPeV0WBH6xAsAtUfoOS3cAQB4ajxyqJK1xaQha
QjU+FGsvViTo7f6SOc8S2yPv1oiFNLEQsJ48Y2wThYtgrubMyyi3Dlx9P9Pt2HzO
q+XsVWcPy/LUOvmrA4VqlpH9oazFHFK1mJhPlj9VJDacxv8TIpYlCt1KPXAHAOsz
igkFNqSgF3KyAd8tym8hbA8OREW7maj8pTZA+9yDrCQrqrwruwlQGJ/LqTvFcTRw
9jb3GtsM92gaarRbGMkQGsswzDBR3UyvFc3ThpHzGEmk7FEZYo4bI9kKnsn1Dzq6
K3zN4LVp24bEepAIBkI7curIpM7feKYxxoVTQjtK4ZegPHv5b8M6BZHcHdO2kyMK
JWNC4bDkBBiPkPqxbrdwSdP8CbOOPXvhDCDbtJd5GcN5inAeSQ61PZBhsCmscOMJ
mEAPGq5Xsezp8ib2iG9wiB1e3XdHKI4O8mr6+3NclCwHz+N+gdZqiwcYpvoULjgk
0hY3Luy35R4Dao7CRiDn1iJDvwqsNoeXt8MNjDW07dyMC5dcfdQlDP3ZAboprtn8
++gQZphIXKU9OHhVNGxygd0d3xWvo/nC6KoETuIe7OZEavOED51qk0tlFMtBlWt3
sS9QFMmXy/6HxVHioMW+EXmCmGf+GblI5dUbjCNSg6n4ucUfR4aOfthUhJ1EvZiH
2STyYo1xIjPENGSAIovP+BeTFDsKByYRlZViJ6R3PWHr7h/NSafTCM2yK5lPPF1G
iafZlrcxphYjen7LFjt/v9qtWcPszShwWkxHhF2X5XJoTREuE2BJ/pNZaWT+C0gg
Phl/RmVOwiUIXW71hMzDTXwKt7YEb2ssRRpjcBBEpJ6+S3ECziRq6DOBH+Gb9h0V
vuUUdakyDgw403oMuYZsapjSFgMrkDYPpmRQM3BCO1DGSbK4oHA0Kvdpd7hCeqzX
Lwjipl7OHyyQwy9uDHFI5gOn05HlgjblTZeTbePyRJFnhfAsCR/sbVodaCFBzFVn
SNGax2T490WJzmooZHszfSpSKtqGPXe3qLYWMVHI/ZhRWe6YAdUJphvEMZ+G3fl1
cgV5dtAdeLWs5zZfnMeV1Xn675EDMoQdU3K0nzAPeajgDFeU5M/XfcI8Y8g9WELR
w5SvQFSHeRQ4pyk6ewv2XvSCh+gvbiymcJtNCXkVOJvCFp4/MyLCTJOwx3lPYnP+
W84W676JfF3h+HvkCsiw63XNdOf/MkpQBbiUKcOfLv4OgfjpcQKk9XTRTTTH+L1Y
uv27fvZy7cTIvDIdGoL/Jlr4+3i/cbEU2Z2FdNBNiejGCQtsfAUt8j0S2CzdEAAY
z+j8GfscMkXL6tJi16fn9UDoD/BBtfyLiDg1wOyqulL9ljSs2zWCCBPlSbhLnbAB
hLcUijMVGVPTQmZKIELz9vkARdpHjlTDq6h1zs7JAXc9NravvbaGjWE9/qnDvF0p
NIhiNBBD49C6HWTtqyMtXi+0Mtbm+VDpa1QloJ07wikn5+Z67WHoml+cUnQRObA0
ozqCFNF9Wqm6+3KBQDaiLEjVB+gEFgdULIR1ISoQXhVe1yxvHoqLHDHUYZgAz+NG
qJb4Nq/MPDrMa0ITLTzySvcY7tisT8TMBXQgpNG57lCuZhF3Aqv0lsu27J8QUPX1
77ksaJDF8NUa6bFyhFlDzR0iR8NcLugV4z8u5dW0YCD/PR+1+cSOeHEtQtDcYigi
wiIHOoAD5VV65rpxMisrAodE7ZeNc7DDmJtQ7d4z9RlG4fgnXtIYYN43QjwUMMdy
QZ+Kf2NPaDM1E/7fqrm9sXzPcx46p1DIBK6OF4t9Rt8Q4/pI7+151O6nTCwx9DXl
I2fi0mxmvKWffe8EwarjIzt2tGtIQrTXWydPXyrDoYWjklPR/54YWzCIWrfnMYRy
0QEJ/utGLNJpJLz6YMoTPav8NZI0SYicGdfEcfZCwkCix/YAqnHl7accjSLZOXar
EiW2pDmThqPmCRzQ6/y33T6OQKiEqRRy7ISSooiiEDKlxj+aFrw/h6Wgnrm6zL20
i9amLzOVLzsjZ5TT3821TqlG2hmD+9/to2VjzUiyytD+lGW5TTQlG5s2yG5S8c3Q
IL+8o4pblX6C+CA3ryjpFmdjs5cqX7tQyE/4KCUE4MDWDxscfqMOfEyElRq454CN
B2iJROgZhMsqNEEKqD11j9BL/sUPW9ee47beh3n+UM3DDxT782km3eK0qTtLcXJR
w9UkfGcUx48UBKZKYuI7I8rtbEoEwSN1cbdJvlgECJyteJ+dwerERV22VDEhbeId
GrcdkupWJbTx3zVVCBusM1caKMfSfZuEuBOmhZUIMoZdGkCiWZ58Hj0MGfv1862a
O5QilbLFK6oo5rHKM6nqmPyEhOAcRbkqWXJ7fcxMoz3FS2fjPO7IMnRY1qL2Th+z
0f4CpeAEr+GIDqTEAPguTyj2Z3NtW39hjoz/H3AQbIqwZRD4Sa6KaJ8WOKIGhwRy
/yQHQcg0oPl0+J3MWicV43nrytCgZnLINakGPtjw4rz+3wmFUj6l1yTB7oTi5Jel
qFwGqlWoY4jIB05RZhC5iZf8JOaR3KtFXMSwrIsKrEfp9Pinh2W5Zru+apyFC5PF
/khyHkR+XEyvRJ1N/iuRnBC+xOsWAsGlQt4TvmjDhMEqD2lWprJVVWI20JbHKUbQ
xsaJeLTNOOnuc95xC9OBQbxmpJJnSI+bfBnmIDSfaTO45F9H3TTk6AGpK1Q7Rl0w
mH5H6mZjKEcK9dYFrgfqu54FpPoRJ7H9qhff/O4nA2FzkaZuHRt+ay6sWNLb6GRs
mmbgUXS9KUgZ8J55qYK6y49nXis94037pxht1WdmUVo4MlT9kl+3rp4JWHNea46n
nJNdKgUvPXYWVokDrLAdRwxdC+UB8Hv2OyF0lhzuIck190uvkCKK2hGw3F2fn65v
9uEEsYVQqDpJC6duYd72Gq2mWsPZM+O+gjxPQKnm36ggE7ko+lOEWJIg2HyUvyrF
TmTCcenUmfOnxPEb5zqtFI6J36Can3YRkE0MZyK0jPU9ufJer0aT+BEt3e2dUO2K
x4PzDFIBMLO9qEGzgdjr7eOKBL4GXTCbBjoWKbm38Y6hKfBbBEXjucYKwsMwAYGe
UyZ/PFrzQ3pE4CpQWe40TEX4/3YvtsAdPFgtV0p5R2G7Kzf+SFwMmQ1I7CRhMlRK
650O26uFPuY+aVMfudMJ2ZtzuDs3NENnOO3rfVO78xK6LKSLfqNnm7YL+A4OSHN+
EjQHSXSxSw/1LtfkWsrWiFRL0g5YT/GyTBPn4Ykkw9e9R4BXj2kSJOBf3sbz2KFK
rsQcVQ3G8C4eE31cvJ4kqSTaP7rdFrB5J9cs2qSPZwNQPWRw+DHasvnys0WoDXs9
UiGd4pRFtUU3o9FyAaxvIa6ebSr1zHsNgntubVpYnRjgSZeLIhABvnC1b58dlR1S
Y8dN0p23Rc528nMqt/znn3DKs2WLxuXACLB5NeRi2REEosMELw1WUJhErURA+sC5
8GjXQzxLtRL8QQAeTc/T64KDzWvgVnxC6jRrUFKMZIWJQRChOmSlN4pUVPVuxhhw
Eubv3oVwYYQmCzeyXpxe5/e1fSWpyTu9VZJyEBy4mgrvTrjYQvvAdT5SdUFWVMDQ
S6uzbbwKmDnktKL7gUPuIBurrXjXfwLl9JOopLypV2Yo70x/3hjRGh8OGnonn4Jo
`pragma protect end_protected
