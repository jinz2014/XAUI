// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GdMwlDfWi7V+k7uTH29XD5QYlO4xpg0o68G5IgxbqUAk+FNEp4ApT+FwLdP1RGse
qQhbFVBG6fY9LRo+daHzrR/69xms6Qq3PAGZlNYLjsJPh2LfmMIVnldL9SJfFRO1
6uFAuIZPbG5lM4z6o89w4appk+St234MHA7a0M/e5lo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11744)
SbG9CXs7BPIEC0E8YNvFfqId2PBA4SSFE4DH5XUQ+wpvldME1ooPx6OQ3OBCazsu
MKtDmjaCWmqmPGuIZF1sXJ/2qepeAbjM2J6t0P5cqPT0XD8kBySc/HbnRT3fY/xm
FOC8uliocbUT/0MVJKZsEw0CZEP+FQSi54sZgsqYdngU6anwx/Czl+EIYVN3LLqy
wHStU6a/4p7Sh7b29jNTb9m9+vovOG21uu86Zxem+rwWUYyd1rWTPmNX9j04cvmy
PUXzM/ytVGemgBR2YEOyPhv+7t9O0+TitUGw9GsxPC/x9rZ+D5v/Q4CDsik6OaTt
ID1YVpzlAgaanWNkRwbyTBPL9vEIQKG9zHbcnvScrKUGMlFoqrYrvseqO6pwP78n
1DEVya0zbBOwQSNebH1RTL4ih/cT3RQmWYYMKPcQK4IlFWSbQ2JjFA20FTVY2VVr
uvdaKDBRrSGZeLk9CdO2x74bB6mrnkBig5NqIsFefMvs118HPTRke73Akyq1P8ZJ
FPqPW5wizTjSHPwY9and4q2l5OcamLE9KnD5iKJQFr7KoTTLXmztVvKYxnvyZSqd
1PXSBwbDF/PwW2DxcfbpYdDHpQ1YRF21LAPFeRbol8K/zc2pbGZopWhfrSo0HIRo
O/VGyjhgDSRn0f32ArziVBTtMlQeVOJnjXpmJBYOUxhKecE+UTxOQwFiqea/haLP
I9kA2BiP/Lf8HfJk6pPmND5wjzA/OHu7wUtRBU+nVWTbBiWsE4xDqBVmnxSE9xub
nM48wzRcJgaKWdbViRxZ+ls3vA6YmTGHhsif7pBJYCE52HisRCWcS1PSOC94F7jG
hB0Qc+JUFS4x8sLC1H8HUp59XGgEcB2XF+po/XgDDWPfHAqMWG5cX/5A1CWl56Rf
g0MRt07pgWfxtoZCnSHKTv5A0G5RqeqYClscsBK9N3U3QW8DaNfnKitOBNzCfIyS
EB8jPahQQvYA7QTPLtTgTe4c4FsywAUtlx2mqdXIuHTiKAaGpaADLXn14mjIx+uq
39cKfoqfZSWGu4z5frPWIh1AViTL83S0z9S8BST0RbPiD/G9OeAez1xgsbVdsCt0
4O4xhBcDcvbHBAn9nd+zt3rgPKE1e0J7cVLVP0+H2zqsZocA1XpTdUkoYfXnRo3p
pi82CjDvxLNFrJt6UE6Q32DoQQX4ynropJ6t6nWsX8dXmXexoT7BfAvpmu4dYy+0
OazTerD8FecvzHIHMcUapRx+QPQlJ1N4XXlQHJ3CwMlw/JJyGad2OH8/yBFQjN6O
xtusKTC68G2nmPbKbYR+cqjvlYBmL+WLXlt2QdFHnxq3CC/hwF4OuC5GChoY5Iia
Q67tvtHYp4tp96HsNApEdtswtOmH3d5Ny/QTK5D+xo+Gvc5+/Pb75BpamBBohzHR
H8X+OqT9YhLnZD/PYoo/D/wUkRzIn6V4oYpQN5gtZMz6A63GeuEst1qqyqMVbbV3
if25vNmmdYgco+iKqkVqsblkhzbG9Sln0H4A9W8QnlsYHBe53t5BgYvx21+7Crdj
xxUmwoO+2D2STfeIufgDbiV6deLAm/2Q/R+WGvTP46RkJRGbByFSPZnGCGvOibmT
5+4OPsCK1E+9q+raUMIOS8zE6W4EHOQpwnhUCTMwKZw+r9ZKwzSPl+cu6UMJ/kCF
or7P3HEHy/dH8egAByCzJsQn2LLrEvjry7gL4WcZrv9t+Z9e2s29kvGsJlMZLCv1
XPdVhwePE4mCekEufs8z6XABlqMHuZveM5MjTBu6smj1qgofjo8hNvn2iG9g0yrp
ginZRx5P1+PLNqyKdmTau6AEnxNmEBh2fDAKs9MxtesHK+6OoPF/SuQnsAmvVmi/
BhUo8H87iI9UaUgWjx9p8ZPtSsg7rbBKNpgaH+WpN8jRbgmliNCKTyB2NE/3QFr5
kT+YANtDtGXpiEiFn9j9NBrjNzg34tCXVu5h0Gil7vj/FMCaIYQQGoreAfhwXEz8
f5xR3QRvddnSFmzvEFHrBA6J7lVB9YIBN9sIMgoFuhKUYeLQS99q0p2tORuzTLWN
p4wHMKCQebzf5iZOtbUaTLaTyUeH+B+IGUg1S6nXjXlpvyR6fzhg4PqRPE2OYmVS
H82qFCjViP7ZPJ8ijYeii1A+CgU0m9ZjyS8fRT3ySHX1y/FhmhCL7mrDGhp76ozi
9gBKn+019AdgLHpd/IvYESUFcGqUY39LX71w30aVrnNmJwU7LRq4rndjyxPU8mtF
SXTRsQwmmUPfInLpmDceshU89qUqBSwVRtObCZcW4FTovR/Bo4Q7ZgzikTTImGfR
JjJlsnxZUMnsC5MSCnNjben7zT0cCN9oRyvKYov6575t1qkhS8P+WNExXthtpV+r
zkIEJ74xmKUuEX/VDh05u3D07JC9y+kWc2Rp5jHjU/Ylcc7X7N8VQA0O32xJwauk
9ki+tx4b1wrrhJfIKWmgvVBC1GRCP+BAUhDr9+P3o09PQLFkQdxj6iaNatuLW0yE
DNeD1+YAZH96jnEQ/Q8LK6pGubcZkoZJhHdKgL2xhfDGtuySEBWZMJhFy+mAQWfO
+7m5J9bp5nvcgxRzFF28BZ0y3RUvrJwZI/3UW3vldN+HkKih2YF4wSlA7n+edt3k
N5Cj9a2NgITCU2FylqX0WnVRLMNQUf/UouBlu4/OpiESzyRuPkvor0iCCLWKHdrR
9CY1r33PNcgIa/xZ+NLiwyBBsqjCNbH6H/8zbPcevf5mlfiGoUtsjV/5VLBBgtyN
CGwPcCdTXfdqyCxILbki9C5fd9oC+f3RehM81XHCh2HWz3kiBhXqRia6mfKJPODE
lK3g48g4+SDenNcLCcc8cbWbTBZ9QdvAB2vvUzHhvmnjxpco5UkETZVrXJz0hBPh
Qj6cE48QHcjm0kEmC52MhQqsm9jKcNX2DMU8tzrzTVHQOcGQSwap6HBQRzdgTEMY
RcKc5rcWXGNUfbNNtjlZBPUvLEyqnApnkV+7P04WXMqxRZyQ+E1xxJoVdOvP5GXY
FvsMqFMW8m3ZxCCypWayQMNEsWoXf27omI0/CgtkckySyN4VQVzivMifUv3FzzNG
na8MVM2PP+S6L/wgUOuqgfoe4+L2sxknLCZtzyq0p1tCCXi1lZwaxMjZTp8/zn0a
lgBf2dcHiBXf/LaeMn15jKfY4pf3qxFbeP0eySrcyV2yFRJabg6PqQHV3sSHq5KM
ikfwqSpDanUHxmlFl1VDnXmt24x6PhTZzM043heOM4oHPyi/wsJzCA02Qcn577Q+
RMpac6qZzdCs9hHdZ1hpP0XzTghGfZyCD8BjyWSu1ZqfykGvcYPdLA1yEmFouWhR
i0vMTRkMNjkK4xLk4YC/LyKaPyn3BlgaH1VaFiXvp7RQTRoeYVk750kxU71nYlJU
yCCLtDkVNgwqxJ/h8Z6JY0MrJ3jWmPiiM0kb47oTfaKlQzdxIzYifCdyFrLR3uB7
1n9+1kdCksMu5KHUFftKdISpwulKDHP3bh+wSnQrRTAeAW/e7RBPY3EunFJ8PcJR
oxghWyDdAcFEEzHtfzJQ3UQjgceHouQXx8mBuQwi1ZzTlB36j0nb2KWttJfQUTtT
rPobYxy4GzWlWhsrkPuw1bXLuru8Cbrb4ACTEvCXTZ+YbihdUEKJOBbFp8YfIBxM
2epZIEG0fNvyznWS5d0PkXeuFZnTmN4OE3g0HqLJSPMzzlcf/wGLfCYXRlkqsRRq
LrlVg6xRNbe7v/b2bRnxn0OhmTLRu8AxkeYH09RpwlrIZIofJRnnEe2JA5IZq1me
+vNiBCT9n06FUuOCFwVm2HYChSV049/hvdiwHSYtDIWJejhLTaA1dttfe0Hq1WGj
BUTDyOWQFD7IdpjwqloQLo9xxm65y32nrwGNqCjTMx4OUVQBOLbHBmkFt/vqh2hn
GzkF8XGN6sjxTjR8GFXQiH3rsmTeNt6Zisfxe6aHXosqY3xWKF9Jv9ELqGurZJ+7
Hud7xxyRSibR5WwcvMLwrJov0IfRSWhzE4wiiTAzY4UOEktLcEZvlMqrZ6yN/yBY
/CxfsYtvNVkr0BjsRQkDjC9+qWzA7MkRP7WC35mE0NQSoRM+r40o0+FFPgmc4Zuo
oAcXdzO/xoHlQIU5rdV5UABUG3YJvhy0maUoIXsdVsNIOMI42qwjFAWh0K93e+Tt
8AM5c7JqfIFQrVNK1dj2Tanx7iF6a5lzExqNzQm0JSDGoZKiuXrnjl3MCJWuLs1O
ljtjkOH/GTjWAVUZ5aSWk+2lFpYbF21ef77U9E9eMmCyeZgMdgqYbYPILmr8kDmF
c6djBW9VdDyeBxBOzDtqD4F710spTBDG2AzLjk5Tbatg/KtracgservJosAP5cJe
VhYGWWam0rFkg4q03w+mZkZn4Cdh6hx+1hy4DpN57DJSEspmeEppHyh1NKmlHsaI
iXQmvMpzTpc3gXsaXJPg2tlyCpjSlNJP0yVTPLfyioXFPBcNdK7nXHz2+4mj9TD8
3Tv4GAngfgnpKEsB+zm1XSMgUN/EPZEYh51hA9ADzuxLFIMv2yV4EwOXkGwrNG3B
62Qf1V5MRQ24R6bjnO+myBpB7+LwhI04DB12ffcAya34CDOInyDMapcjfYjoRQ65
20KgC8nAfrhsawB09tDqEdYrz3xXfJCJsKwsfrnByvAisI9laCDmlLAW9K+RuSjk
D7gRDGpgyRacnSNhG9RJACLVD0/6E2cOIDs9T0HAyv/9JbYFkQQz/ujT7fx0+YfM
ABeYa1dZUAVB8JU5eJEFsvkzF/VDc+50XDnrxEMDQekPQ1qfFy7SGUJFX8BqZkXT
Ics8FIFavh4sOhaPYyzIeR0Odh2OhNDaW6agAaVKRWNMva3MsizYbTTIZgHOhVR2
oVQezn7xFeAQ7SQ8u6tbSW3KlOh7t+XekI3bL+Wy48w49eusFiEb1XEMZxMNuxaB
B9i+gOkOiNTxmBPAy9qpx+sOJ0Rf8I2IiuHIMiOrdKs9VvXs6SMFYZog/XbZayos
7JPmmgnzpdkKwQPhagksfpcnqBHMxBfhGo8mVgu8tJbzoeUJYP1XFKqRqsI83QTL
JLfhWVDjkRl4xlkUeWfXjoin/NwPkLBmMJUrMnB++GjcislAmlRJme8L+/im8ZSG
r3kyB8Tu4lXkSKgBMJrlzcUvd/fMMWLPXa4rz+CMVqAKu6O5y5nwpvm95oxo5ErM
14v5di0HTqgZbPsuF0S2oBrSHU3iBrujSxBmsiDsuAuP4i+BDaHjbatAC0TJcDTI
CLETnuKc/30kiw99wlrJf4fP+N7+AJfxj0TL43zO9/TJPV+uBE631O5UqFAgn//c
yysmYuSuJjjaPgSxyqSik0oMsgVKL2g2XIuHRgHW10QKo32LS/brN6UBFWvp4l7E
heespwk51g0SNwouqg0wgCaLHw4zE4/19POFQNWliAUkLwAADcQm6COkYJ0KtCJz
eVYk57ocYkEyPliMdTXAxv07Vk8Tw7qaQheGzOxkJ1I2ER1NocFzPzjSrRiPzQQm
NYYlb2S3bYgXyhnVBsJNplOFZuimKua2KEZa6aOT18SdnVDCOnBeFOzpEmlpTU4I
eAPfAzF4ypPqVhIEs2pe1Se061hsGEmp69gbjEhZeFnu1RIEAkghlQrKvGE91dGD
bf7YKiiuD6xadZxlpEhQaOoKSN8bFZHaDlTmp40A3s82fw6TAubM0SYaV30YZ/76
shvxUMI6IlO8ynGTn4N8uthrnUn6qWb1R324flA3E3z/omoIVjP7/dSPkaz28N4x
cNjB7otEtJx4w+CzN111qdCyT7px7uV4hO/+wLxheYxLGPCdsG+8OsLrjfWq2CsH
MdcKOzcvyTfEI7S6ZIJpgGuGI4NAxVb2AS3fDF0nynnnfdUC8uLoZqIE8nWvVilk
iD6K5mC/wt+u04m1qp2R1wCfTfP62dEOphsQrhlBkEFHJ8I3BG5wkeHFiOx6GADZ
Ai7Q8VG+l3Bq3J2N1mTMZaqhGZ36/Cft+St44OJkaAg4DJLk7RfPSppn5q2RpoHu
Ec7M6kcz8zil575aX7Zrf+m7ZtrlNE5FLuIHKXOD2aNf9Q1IQytjdkM8zf0Q+dIf
HxSDbla4vRF+Rz+iD22eXr9/sfUT/tmpJe6Vo5XprL7v3aTIe2Vf4nNkNR8Jnbyr
K0H9pls/0U9axCB1q8GtAmS4yIVrS5W3tp2Y0jAn04c0bBzSuDmRAPYQ6JTWlrOs
xZAlLzILZSDMmuM0mpsJ3kcQCFnonQGdPbrCUG4BjUfpHf0nZn+QGNmW8cYY0Ilu
Xxx6D2/XDCZlu2XYyQ55mEDFW7NYkvp97lq5JwYYDl5VVnZLdvRx/FGIQNACBEaF
nrww6ZzfwPkLfyH5bgvGPS2H0axPDGVgheVjaemsYduuG+3hjKcKPL9gmeSr1qG+
EGt2m5WdOZ3M+VM7dXyGnd7Rjdd35FFXSgE9Q4ABiOAnKUbUArCMlV3YPiCAho0+
y8Jd1wD8D4EvUDomt8/eKf5FIA2SPglVi0Zpr26u9t+InIr9Id4lVAJYWJk/C6Qk
YricN6vrPB9FwA4U0FdKhMmiipQmF2BVKprSv6X3XJhsxT1SC7ID5iizvsMPb07w
jxnwEykquZH3nH3h0Gh2FGGYi9pteLweUSnvPRCcNANfw3vrds/ZQ5DE0nWhKN0S
lYnylDrLDlAd0rxGAEJLSU617yHXM5S1yQVZ0Z41qBYtZVAQW0vXKRKCJsJG1K9q
43LKBIxVf/9YI4Xk7aA/O1U7uMKEK/6hehVTxjrmQLgMpRV8KOzLauNtTi+DiVjy
TJp0sBfUuEsu3qL7B/1sSTGmxGD8WvkAoNUMi8umd/mz+74AIoQcEDjPaiSpHKeA
tjkcGRJhNYUIWglLWJR2Cr/7mX2pWt8m5jQG12e6Hini/2xwey7XZ5Vg9ilMcHQk
zOP9WIqnXmYyWc0ytlIb5zf9EGHA5Shkjoo+RkBiSyfhnG8f7GgyPC/+nZjVCckr
fYHvi6Gq0fmqq8K6tHVuuyc2YKoJx/WvnoMarebhIdQgNRwx8H+Kru2VFghxk2gU
IY9dNVC6+uSlaVkvFdt97C7/eBmNZXuPL1T20M0hmXyMpN4kUfSlMWMuh5HaoLYg
vtzMaS1zJ25c/0l6GMfjNwLMcjpTW7a0AMs/Cqjxb6BQmlh7bqIr+nIVdNAPwwpw
C/Ood/+k6odV67uzBX5j9zuDE6727bcwBbdyYJgw5GGmF9rzkKahxa254GBx6QzD
c9Eic1BqhZi2aZapm/mpwOZncW0CyI/aIKwwl60x8E8XZ+ZhRi/80dKcpfpzlxdZ
l64aj0iRWkjgGVyB9pk+ICHUn+8AuUZC2M+WsUQ9nNpZwu98cSLwDOVuOX9bGi3o
BBQW/LzWKxexVWEKL7uEU32MU5CTyd4dK+5ZczIrC8nH/gSEh/9lKd5TPe2fqdLm
YgKuXmCKaFGefJ/CA5XpGBs+OpQQH/pbJ7dBKZUalcE+a0hcV2OX7/QrU3qXlrHL
NsBFqT0JrX313R3ky0FgPHxtuSLDw6hhVEPpONC5sdbbYDmGMo19uN5hme0hCmn4
7i88Dhp3r3NMwWOpGIFGP3X9vbtpZEGN3KwIbgpWaOkAsQgMvv7KtWtxCNrCx5lK
gROIo8vFstyWaDYAZZeCEnqfrIlks8djPOhzgQ1yrmyBU+HZs1E90GwMPdJSlVPR
w2Y4GCavhNmuCPUTdwWA+IHN3pVk1XaJSrvFP9qu0L6d+dz4jdbiEL0+s/8pfrjL
cpMn7X3dhg5ZsfsDST4kVGXIkayupm+SbNPAT6GX8yU9uMEAxTN6YZq0oFwFgGhe
jfgR2g/Y/NLUTjKx6BveBLEZwQhNWrNz4osrzsCLAFKKrxEs7dm/3pGtAdvd/ERn
3rO7Ti93NUOhmGNmBD5J4JipS98hMIsmDVMdOPASzFnHJd0ynj5/JyFjuLGXQwTU
6Itr+8iP2QeHhxoUnt1uJUmNSrQvhxIRIA45Rt1alGCWrA96MW86NAoX11YaMqbn
+DnUuCKNdeniVN0RhM0w7PQ5AhvRpqBqqh+xj3cHqwEReU4HEH4VVKUkuKaRkJwk
vDea9xZmWZdQU/iuXtl8pSXsmltxqrzoqihB1iOZuqe+IDNrzzdKBucFouJR76NC
cWkBnVzq24AMVyiKhYoucMkJIJLb0NMCil2c8y6EE4DAa4rkZM/Ubb+2NDWIyMTL
h28xrAsDUvTkm3cZenL525U4d1gSSpaiEfzet5h2/LB8lcBmjiek1fnBgxxtowE8
KTR/mXmlDU7W8r0HDbA5IxzulTFRWjVmKJoetILXFgCLiYBorN8cABMkUbeh4//I
srPD8PGbXYn3jDptNWj5KygAiW94Ccl0Wk0fEN1gftF2wG1tp3cui5Z8GbbQa0g8
gWVEkz7QKahuwlJS4OenRyYk543NkXtNiPGKGKSvMD/3zFZiLDDeGcoKCDZv0sqL
1YfmfCeKy1rEAqRfPgG/RSFcc0ue2j6gFbedRrlYVBo6Kkouf3Qx5wkBx6YMy75U
6LyPSrh2RFKQN+hkwMGnjYC/pooYxmnrwI7H+RXJkUCRg50bH8vGEg5g9R0Ya13x
OCt7hALPv6aJhHyXTxQKzzIitr+TmOYQas5nuZKfsFWqu9QUYCdG5OVIHlQ5moB8
yveGEVnqSIlfZvYHMErKxp7NbAKN56fMh+9w0dInnFC5MpkweMSriSIdP4RDv8j/
ZBVClT2Ic2iA6SI555U+lQDtH67RDF/LKhxhjX5tOsdN5Ktl2EvSfdU8WEKeyFte
EuhrciYcyRC/dHjZxcySlQBAERbzmmRE0yVsuu5901YM2qzQoWpxs8Ruacp9KU01
7Nvv+iwzIo3vkX5GGyBJ4CZaH5d2uDswrvuDvmywCGyWQt9CnlGqyVeTnsHc0Snf
cZS2OLLi4eS8L4AMIm+dl8YfrBC0EUnyWTF/HAnz6pNsIGN3HrlFV0KHmYM8coyH
BxPpFbqpjrp/LbzMPQKWPiJJ/NQHNPCaCPDENvZz/TsrCezLMYOambFbkw0xGBi7
mtuXJBJlUdJf1C5Piidtlp7kr99UcSvUD+Gjc7I0G++XrU+B6p4L8rcyax2AcGjf
SrFh9Vdf2pRfCE4jQykx2tgjkZJxkchACZ+nNXOdOLtuNlPHuC5eT8hIxEtogelO
6eipE/khnkdummhNOmrXNA76jw2C7iTYiB5LwjNjBG176/SsQIc8KgjyDngVCPZj
H7rUJXzJTSgKIpw0EC5KMhF8YusvOfiyMRxJdTzOr00P78V5J7lzyh7/u8Pcdb0b
vZOHk8ZAWixd8JyZp2wPSaVhLI4j0MtM4KhOXQxlNXgy8861RTxUzrkCFS+C/0nf
bx6aantZxqB58VT39f2zK3kmFjmZfpco4ZyZ1s+mNU2wbPP8zIMkZ3wixLrFobP1
K3d6MBdN+fMod1Kv6e+tACBaL5D7DAsQTe1RPfg63a8fDL7rWnWo35fyvRefp+1J
HB1qq/efSuQ2Nn8lZHAROc60N9VsUK2vH2/kwgEmfYpNKoPpOApwRQhL62Ig/UCz
AXX8H38frL9NFFad0f0nVpeS0fWrHbWDDCd1UYSXKIExF2XTuYroqR5fVPQ8WfFJ
h/Fe1o+awzWp9jvsoXWx2DouqjsEnCIeMlcLaSs3UyB3/PJllaXqBOcZuR7FMnEo
wAPif9VERF2IeL+vwhAY73YAFcX/LKIc1dd2xJLHZTzzA/U8O423Fog3aDXg3iNf
2Llq6YYyoyRb68w9J20CueK0uOzjoqdlzuIsFEgU/YVt1FtCM1/rNEd1VS1rdH9Q
61Mq+JGCHHKr4QwOuHduV1BinC/+43ewAfNGCw0ABJ9whC627hKWjO5BHAcxYGt6
bEf0JvmbhdQ2pQUsmTpEkF+csspD9HKynfsnKvAXLDrCNinuDrNMTf4KAz6YV5pc
qV38LMnmxkmwgMjY9qCh9cyvlvWFtaO7QQgInwg+HL1fk8hqO/3OM3necm6t+g7u
ESUzTL8T7moyU+l2r2NQQ5onElgVw9IcEQiBMLmv5/7HUs3lx6To8mYk08VZKDFl
vDbqrPMnI3ukp6mSg9Jr2/0uMKmBgTXP08t3dkQLiRrf5Uo1X5A0IPnmo1w0d+Ri
WQZZ0qulnizg08jY+ydiKaAUSKGtHU6nBBlttievD7PmkS8ogWO1WtCp2zguf2xt
/wzK7nLdf/nsQ4OKDStGma1vMRWdrPJ5DMpb2P43I7R7lWWmJ62P+4QNAGLZh6C6
mJkGuTDrZ9ryTGpHCg9NL6kCJYyuRCBzoRTgzpp1HM1XTWIITGAJB1dV3PkLQP/a
RteIfun+YSFOfulok6ftHanb6OnKEiXjZX+fmylPPOFytXihUzZv5uPaWHqLkPpl
8s+YNpDID8XYMj96809du+3io7ah9JaGUiu9x1TgDs8nAZatNhO9Sf6usX5K8yEs
PfqkJuPB6GnVqCw3H9ZC7KJhjjz/diMusF/3w2ZKHuz83ijhCHOuNTaPQRkG3WWe
vtwCn5r7E1bdlpzEDxNSCckGZTj8zKWTsnHuNNL4tvEGKoFZYEt+eeHC3rsWQlWa
wdtRlQS+hFY+bf8Hd/7t8cqDO1g7JcCNaXCM6ViuzZ3ur+gWD4/ZljUFThil6IMy
/1H4n0jQ/J91YXpHXzGmw1jZv7n0CtxqLoXTvdtmpyU55B8CoedLu4rA1Tq9jfvb
T7cgzfYL1yQEp9DNOrzwDL3YcwrSqmLpZaBdhaTgKukh1IVUSk8l9CtvBvEYYVKc
Shy2BsAYI6fLKO0Bd4smwfjR5/pugp9HT+Is5opnd+ZfXXJ+p6MvVfcpiLPwRqHo
YeM0u+IvpUq1mVXxBYR2VXTLXiNHn2Tf4RKOmKpYmltuMsbYxZut3ROy9+zp4Dbf
WA09M3uGzNCN8TcQldr0w7/1v8Qpfc8MBl9o+GBnbxpOcTdgnPjttC4PffhaaMJU
mNKtJ6nvOVcSPiUQibgLKyjKPvXqhELPrpj1QpSkzNX3UUvcXy8zwylGFYIygMpE
zPFLiroCazUgpXHVZWrVWGDR3qLWpKCF5EXRHpn5Z5pzx5p8Lg4qQBBluEzoZEt9
e6fvcyVK6Cbmw+20D6cFr0mSl63twZMDmLrG0lDeauE11Yw0gFtf7saUi74K6rJO
t2RUGgJ3t7AhW+lm6b7CHw2AP4jdAtez1nCK1cl8vva9oFLq0na4tuEGxeX501JO
RkFjrWBc/xN8BWVTO4T6qnK5suk5loCwTqtVMYJrEtuXkLPjta8csYKSHw3PJaJj
/tF/d6XQlvepUS8uoeIkI5sDqdI7qKtU+IMYeeVOe/a6WEfNRsufbg8LGAwudGpK
y9TzyF3gvG48nmZySBCgxNtCwz6S7w3KHO14RYMEXe8SEuz0Km1tuwvt7+fkKDDb
MZC6ni5ZlwX4hXyQ0JkrdH8j1976cQwLsu6OtkYRFP1Q8IcWVttPR3BLZ7drPbH+
29nLsySQG/5XNKbSRn2nAG99qI9KB0grI3AWuwt8CLxO5R5e30jf0RVVJlpoGD31
g1w4AEx6GDzwjc7EGRcwWBAWhNFwGzU85YxRZgMwuto9PtCymCdHu4I76gaX1ydd
ty1yQHWKc2yajt0gzpp8cRyXM+HlqKz8cGiP0RHPONu18uXzWrN7qECE17TQomuw
++4HQjiwL1Gh+znM8nqSRRtWCj+/+DcMdOusFPsvUOTA6WPU5dkE6zyTf2DllAbC
bNMtpk86CiboP07Ab05qbR39JIAFUCMxH3V3NPKZDHzB6aayK4gKT57TFzBxW+NW
NdSnaIUXwpOLzng6HuVt4kuVSLo0qJtiork7cecc+BjYcdi4FPnHY8KqdZxpHvwE
7k+HscyuW56fK/ByEb0uaoHqUdlfceHdgZ3gCGRIsS+uD4h6QizyxdG0bGo/PSf3
6VRM5GEoicS2nIepcdAjMsLcs1lAJh0zKkZlWzCDpdgTtdOv8NutEHXDtnmggtDP
baUkt1lfWGiNrw2OL6d7uvrbcNmJeWEudEVwoxF1tVykzMyJuBarFw8hiGbGkk3r
cb0liwmxaf3Ah57e8XqWbRTugnb/QPg4yBVBvmzflcM3MX+/cjFhNaS7P5fYc44L
RXGs5pUpD1KuOCcSU6LeJTdfFZO/AJAT9A34NopjYDd80s4gv/7yp+w4l+Q77B14
ukE2EsQRV14uIrW/6lewPcgvzzFQW0RY5qbezgCD6JW59ahZhMIpFlQiiHHR/zPA
1XtNDJv1Rdr1wZT5WbUHD6dQVuVpv49raDzkA0Zcpz50iPNFTiGuav/74r1exgWG
piIkS1AGSsMirCpHKx2eEaYWhpaNG3RI69oWe8SYNySUODrhKIcw7LY+6jbl/ZxN
oyAv9KNQscynw/Uz7aw3ZOVF+mn8a3QBVRt2aUMEJ1teWur+Dg15YcXQ5U/ymAy5
01zfeusZvUhPOZL6eP/drkPfEn6Q5ANWZsCLUZdZ0pJxuErp9EoUXpQOL+7safV7
hzr1ZyCXISdJF6z27qeYllrWPJ4gwWq7UeX0vOLDQrcPTaPkby5zMGFGSDOBtoSf
kYZPqCBUANAoYUyf60azllfj6Bnw7LWxkE4deCTj8wYweslXgMaKp0wNFPaKilaO
XJ+6bvB57NFiS+ZfNLQfHtuCdkEMuEPm32Z5zVC+syUPj1Ow9aMbARnrYVQWFbTv
3872I1jlXja3VvvEWiyJ1i13CQk2UwumU9tUhTc3c9Osi87RSaGWq8DggH5cn8Qp
sHnrfo1zKAUknOmpa9TMudBIlmDDHvB7Jw70/O8Er45nyBU555WyKQOZhhdCC5Eb
pEObRgszq06jDhVqjyOsJJ10XT6GTbkexqvW87jC5R2m7EQZW95iXKFDrg9aW9Uy
x+IB5KYfP1MiY/pnldYBJ9mGqRA7YK5NnH2m6m0IcDm59Bw9nbBsoSPISBgkjmY4
rkCTfh3VBCv/q8YSB2L9xHoG7H+32iMg6u+/ZYKWQydHhqZRFaPWHrJY9zbAJ1m4
jdua+54UBsAVb6cQuh54JiStwV0GwhUPxkabI+xH/HIekaDzLFrKrYKfUwgIiZlY
H1bbMtMpaZRZB3Xcbx1Ctlru8/hIVlAJnq+wgZhrQxg4DsaDEolAuXCt1KiLIBmQ
Hq090WOkjnkhCus0AKCjaEEDskWeKYFrZYau41rVsv05lDRJkUtj4yri7MHHULny
RqVJ0lkTf46n4u5eaUrLMf1EO4SthE6l65yLphR9Sv8/mR+VLjOn5Dwpphty1yXh
fD1k6nyq+aa0MkkK09IxN3A93AHPthjoCH5sRoc5x1bivXMIZIgAhzLBC6zso6e5
otxzw+sN6tcnO73SbStETlANtftbHSzUmqoWJn4ik8RWke33/yipPjldKzsqNTKg
61q5fcraDxu4iu/bNPUborsncAV6INaSIzpEjNjnhm/MCDysMb0ZphRcnxoZTy9a
/5YpQHdH231SX2qW6fUEmiuzi/se0cJAbcCMzmZq3FxAmKx0mhLYAfPSaW4u5cqH
URyjUpes6ncTbP8qFQRYCqxNgVE9qUmQjQiykXQem+mXLVQi2ZIVNdShO3z8jyTe
Ri6vgClEHwDx/afNpgCUcttQaT8V04z3ih27dLtYxC419iNz86kuqs7UqCC/sVNe
GOnTCBG+mwWexqwfW4zWaiOsAiYx6a5YwkU9XtrVZxvOTCxs6ZwnzNxveUVfxAsz
6hSRVxRxIAM1GS2qMPguKFf9S0oXcQ1/uNHTcVog8geQsJkJEUyCsiEbwbs3a4X4
dVgov9wh6qkkPil5nsALg02Ov6iaB/AgU+zX78SvhpUV2ZR0kmVnIIGh3+SVI33S
EW8HEW2SXYXBnReXMfLk9joBlnzhg8CofbBp3sGMpj45fIOv276iySTfDsbfa/cK
nrgRj44z+gdLTjjoSi2ykEB6dETGZMVuG6UYQnF/AkY6IsAf83IviGszf3+vX21Q
/pTT4rWZA2pyq0A5DNF9xSvq/YAvuan+dYXtgphvRV4ksIEeW7iPwdBojpWeSXkp
MW8RTadf+TKUOm+pOBFdIimg0B6aEXWv8J1bZzex34fy+ZcnoiNzYEfZmARiKa1x
zZA0nsi7GZXJl60MHiZ8mdjU45FwAcuQdKEjTfNQOgxpKl0FD9vvJz+BPoRsklWX
0InGuy59IMnp0wgt3PEq3hqGGQ3+1C4V3sob3xGIJNk1Yju+0076kxHnw5dSw8Hi
zAkcsJ70+hNzBCkHjaK5j/z4sVnC16BUfedRJGau/vcQY0cPE3i4G5eoKwSMBL1j
o8olq40zlqU8uLG3eyFSTciGKZDKUSUq/ywVmh+g4UCBz+7hHUiam3iJyVq48XGY
Wa9tplDNVngLtlP6vd+6e5baUwN1FHP8zbNVx9ug+MeJSbn4eKij7TcHdg7W8ppz
n0zn4eoOw9dp2wFhw3oyU2ABYbXK4//7cqZYfgILYUajnlvnmSKdjGIXSH/D3Pkm
dt5xg8OOARUBpHWvVBGFRlbtGWuWkhUS5ojd73StX6ibyDMjTOGTsvKH+anpGkQh
us3wV0MkygqFE8lP2X/VFkjtKj0QL71LMMjVKUKPtiTUH4wkYo2c2y5q4v06DdsJ
Eusa+CElo+vlnYKKrGCFR86nmJHqeLVSWZdJx3nlM1hNAGDgcwuWloVpDmJ8U1gw
Vu0MqIr9ZSbG65ADIE8HqzcC4EWz934Aby/Qim3ii/RUlmdgOWrHjCOoRgE11o69
+pjAISFBy/dTYCEERbeGVQMDivRx+sZ9AutjlZ9XRCk+5D3y+tTJAtP+n0jWb3RT
OvjikRJx3wplqmx1ryJpbKJ2GYwbddrwgKsCG6yvienSwBHUDyUvF21WVH7N5DTo
7naQBvvvQoGTodZc9g9w77AuC+KuEc6zlKjDZdH3oOkn7q/6Cl6ZdMolT/cd0TwG
e3ZZyvyclNMirxOhU5C9MeWcd8JeFoozhEgDdx5h5tVv/aZYx4tWpuIpHbBEdrwr
i3N9sCdguGzpDMbbsE9vUsVFwyytBu379AezaZRXp9xYQ06XJ4oQ7iQJOTiImvRQ
F4/payCahrLJjN/9Jz6W3Aza8HAMx9oDaQF57+IPX9+zgv43CiGCfLEF2hCPmBhH
CCTfgJlUMqLi/SYvyXNXS3PA15q/X6SKYRSNWtt/HoXT5EPb1POSnptpDdeYwYLO
58LndjjhLEAyvEKXc9wrkV8kPbrZ4xpRQBQSRzQR0xhanmXL+Qej52ixvopl1NAc
Y0rgVMZeCDXGg5o3HhRsH0+tK5YdwA0vNJVm37lekn0OtIwRRBPwjWEoMzWNmm9I
PduC7gQcB+Ja9b2WyZDD7v44q5HzIjpOeZ7XjAH1nBcGaOHqjWs53QKODz188ri5
uyV1k4WrvnSFDugxhWvpNy1xzoPqPKb8XqO4CwlHaacrYzr9KYJydr6DE907M6qY
RfRF33bIZKXsG6QiiKFxzWVAXWZEJqMqgDrfsRcNscplZ/Pliipl0xEiKhUpRJI7
OEOUv0WnJljWoHSOD14i17eRB+4PTYeTgCkXPhktWdC+K6FA5R++SeGfcSz5wwND
OtGqJGQEIdoM2HaLGjz+9BMsfzXO7qUqHXeEzLbAFiU34WCky5e6UqxxL5QeztWy
x8N7EqSkHnv6Xz2uOn23IxYr+vdJQZpf7hMRGgzN4O8=
`pragma protect end_protected
