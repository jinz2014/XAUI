// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EZ5MdnWYEq/xH+E3D5ZQEeD2i2ki381SGxZDazAoDjc3Dy+vnJJDFzXK70iFMrGK
DBsQon69htd1OS5DuCkES+fBSey841rVmnwVLz0nRcUPM9FmrBK699KBrqpChjB1
CjrA+I+GJc1sFy3xn3438T+xIrabOpp4Lko3kLmYF/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 126848)
4LppdFI9Wnu7mRsZLAPlMzmLvjBdNgjDUmu1s0j3h7SapJLKQX8ahpCYA5MsdN4L
pai6zNoo4mWWX3KRJBcukTzEnKKetFAa3JmYD3G2efCcPyQaL+8H3f0ZexfcpHkr
27KwCBmBof0dBBP0hh/bqtSlpHqaq2FevrJsyMydt5zqEknksoCVwsP1rklajxt7
eMoZyhesN34yGo+j2F/Vd8JThgC1GhL4YVstQC767IkdCDc5mp3w0aiHO+lKZhv0
nRrgVWLe5GJwN6zQ+bKM8yL2cDoCyuqk0lEY1KrUhFX6M++GIZsyJqA9eox4tZWj
C7jhAm41qbI5GBHahIT5fAydgP+8Df2sY6YddCIgwAgum6ghWNt420P6FwVwwTPU
OOu9yUCOe9qLvQvFxQGcXQ2Vld9mzyp9XgGyt8pips74FSIoarXUqvURhjWjo0+f
Wno7pjb8hn3xsCS9rwUuOkJzZndn4Zg0poEHFbxB2IeTSv5qOzNb25lcl/lKWjnu
IVwFJ03dxCCjg8f/Ip6U7e3bfsHgw8URxWVfbkYtEYlhwYIYRlvEeZf6+W8x2/KL
oalqXZwMRDZrsJMTKSC5hk7CuP5UWk7/tiakfvRzsVzZK84LhS/hySlOfaRMraBh
NgQt0GnIsKUo31IVZekFSg8qRIA8HmoSnDd6l6uX1wZ0H33lqO6nVjZKek4H+VCX
ZbXlaKaHxiJDi5psTj3E3BPVbdsWFTgLtvFsDD5+petEti+kygmPFsmd4ZA4K08s
FGRwDuAuVOkM2xRwaSetkG/pTgZRMD6JAFcZSEckVgLitFZjBBsmEdQ61ejlRpRF
VgyDxfB+soMRGEm/sxXtmi/pKVudhd3B/yrIqNxHdJM/wQCSW6JJlUk5pfFF3533
oKw7GBmS1Y/uIivHotJQmpLcYYLVi8fRIatiQIj95zfsvqNaFKXEG1mX092Jiq8X
NhMXOSum4P5JolpXvTJhOEx/W3anC8Ii9xobQNuhswlh+tk0zGQoryPXv+cY+qSk
cP+UeZbcFUMvFI/jH8AwnLA/ZVh1IXfCvDs1Sd/HrbMBXZjJsaadUGaZfVnzI0Ru
bNQLpaPvk7SCp6B7ATjcha8V1abKXLO+3ZAbEAvOdzLXchWDuu1wpeABpI1X1+3Y
nhtC+fYOWu88d9C1qaCn3EkjAvlWnBs1VI1y8exgHODdIDcxZDWgnbCibaoTNqTI
oSuyFcNpD2wJzSMlpzDeSSHOWig6dTQJvvnLnERIq7vCGhyTs1seL5WcUcUH3JYB
SxrFvRX3AvgdsdRsJ5x6tD3llviOreU+iyaHwBzdAVGJ1ey1IBVQcoOwJI2BW+Dp
8pEu0NfFv+lAc6l8j7gkgkicge9i/pmHNLoLOW3OUtrpciIU7SRLAsC0MFEbqTYK
zonGUo/Jmf5/6ZYVf7883Tp43fRYAzrxBSJiTMqWLxWYe+mx0ITP35rMu1scxjse
95ZnQRKLXlYFOKnYLVreggKS/HQ/eGqIWZ8DQnPtWmKj42RQqCldRG7uJkjLqPIh
lbJLYbezP+fbm5KMBXQM2XeCALfiJ0VLeo+T9fDkTh5NVBeVIpWkPQK6qv1hYwm2
PRvZgg5kx/6s+zVTWYK8YCmQPqFb7YqTpSydFVzqjoVFcsDzxSkJXQ4NjEi7lqQE
Wp/FTD32OqbALoowzqBkXdRBjhs1MLa9SKWTqCWrglYmmnk1hUQI09cwNKVdTVL3
gWXhe3yGEsYbSgZDlefPIn8yGpI/S78ijEbOMFCYIhrkP/CGjAqqrsa71QB0Mdbv
hcir3vRKQgNx2lP8FeHuISxycnauVJKAOkC+9q1FYj7l8V4yCoDqFpiRXoCxGxPU
+lPST30/jRZyRejAzUPYQcPcDDCp5jVJsD+b0eubp6PoSC77XbE7D+Rd1rNJwBhI
Nw3KnWP4svmZjDEphBBOkXHev03ks5w2xo6rKLA9XHhF49gg73tpRlUHa60ZJChC
5sT87EC7xlMB3Qtormq+OeC2zbXm//7PMS1eNQWc3UyzGSu0wjerq5FTlttzNvc/
54MPX3b8Z9YZ12BD688YbvggUi3tOyLXHUGZvf3Jtytsh6aVUBifyoL9+tlSVamh
zdur0kOxZkghup3Vd5fQAiiO6KFwrEdddGpA1r6GOa4WOCz/jpcaq8PMFFULyH4S
F2jVG3Y+HxZ0I8n71/Mqk1yoLKma0kJWfGr+PMl5/tpM4SJUnZqVY/nbxa3I3LVL
iyIifCFFSrNNcJHrH8YI2Dc8hrkt51tX6fDAKf7vUHD3O45mR0tVb9AY/hcLmO7F
DnztlW+1NAjwqHlHCjOhJdI7mRmV0dOILisyotgTOwnxSv05N+VuuYHzyvnsCt+C
M1mmPkZg9q2X/rkpKTZ5D2W+4H95ICrGdpnDVSZkaTUFA+Uf3iJNLpezsFdNqZN2
PenT7+3bX3D2V76m+llgcEx+ROI70xeiVmRY4davbADuNa5kOxWwSPkFtKtpUazQ
Lq6afyFHiAfYNwMepNJS0gsxGUENmPWicUuVQz+nbNHStp1GiMO3wXtnvTh7K5dq
qpPKCQeDyBBv7dQVD+gKU5RbtDV/bxtSna1vkd4atnhF0x3nFwWgE07VzNznW8RC
5FY2bUDMaWlNXBV3nskYP35fKwQ+xTFCvNT3//uVnQJD78bqC7etCLo8ynWN3RFp
CRnB3eAw/CuzCNTiih97P/AOKeVIgfbPUIwdP6L6JegXuCEPKaVG52VihU4Fcx9P
e2fDBWc/brcgVOJKK8X+LxQNa5KBrC92JsaeLDdAD5voahWcHp9Jjrc89XqmRY2Z
yUHI3NN1Xpm3nUhJHN20aSMyTII8rWFrFUl6v52tHS5TzojAz4XH1uYDUxE2KAHB
Yo+RMfuCSYq9Yge8BuEH/GGPXkvzPcxT2EMef7lmw2yZaNEEYlU8iYzr63d47Qlb
FDHnqKJN1kzWp36oeOdObNdikLt2puX5ttwmyS76zj5mtL/yjnLbkffPth4ZhI9B
JWLaMb+5l3jYNrKsQ64WnXwatv3ZmeJoUxgm7RNBvkPAYPERBN0JzPEishHtANCM
3kmqly9cVJr1Ci+5fveccMmWi9eK3Nx6V181TSfCgbNFRV+uUjPipzotsMB2iSWB
NKXQr+L7TKPyuRDIPw0Ud0F2m3PvIUUFamtBqBNKjMUQvJKY4ZbnUP5WZSJ8rQVY
g3RjjjxmaPMos0M0E1MWxSQJDayXfm/hAP8DQfyP4GK1wszBxLMSAzUe5Em9oamw
LvklWUoUzprQd2RFqErVi38QaI+5rFvK2iHLY60dH7QLUVGFit/NeXawcvLZyGDH
urd6lHj3lMu2ojoPnaCrflzaaoVy+GaOBvckq5l7etzupa0V2B8l6Sp/VzAMPXro
QGV9TYCrOw1VRPXk7YhD1YwPubVHZvS8O3lYeF8fSiy9Dnexg1/tUoOnFxQtO1zf
Mnadh+6BSb2m7G10LWrto2Luh7uBVK+bKWoQXwweLIj5Xsp1kmAeiksaE5h+4p16
u4sCIovFE03sm01AA2sgM1Dzr9mY8MDow9ltDDxqa+ql5rYwnymaAEUh+0j0s29g
eJOsjo0MImuTfyEOJA45XRiMxOtPXBbYsowictGKazjInCDzlHm77k5QWs3ZD1aA
Z+h9tT4nuTXAYNeeZ11cDDzl2SZ/n5JRVGGcIMwZKibMl0fky6NWGkJ83D+V5LBt
vohnH6jDV41DuqUAoOlFULDhHL/W2rvwbtcumPh37Abd3FIlP664JTMjMkfCENKz
uki+MlKNER4R9oBGgDl8EFr/vGs0r9DY7q4J9OTR5TJ9722Ucur1cUUl9bxO20Af
WQ/6prQkEVud/BEKL7SJ5Av8G6zFs2M5+w79Q3+IaVtRz355EgvV+1Qa36CxMFH9
Ng/q/uFSWXlxosN+55s0GnTqKZggDrnSEpm5PT7ghbO12+2ApZKXvA8aoyk4HGsi
3YljEdO+VDG34xZTm5RwdHZ6X0k6/dorfviJZM9174Gs4qthTBAmWL4nP9ZvLVQP
1I4E0ECUZDT26+dSrFNZ2U79W6DKgBCESYhXeWIBwqwVxqdN5V7blQkFlk+4FVyN
tzBTBVYJNJnQJ+RmvwJTau2gcvlAeOnhYKCZIDWCZUXgKWXC4AzRIScJL7QM9E/j
vnvlIaVvwGRtKPOhYgs02kcLfAZanK58u/HWiWJOF938P8250T0gSUt0xrJNqax/
xT09GoxHO6HQeh3Yc5K2vrOmSzZDJ3MvaKYAY+qTYX02dat2o/4dy8ZBq7j1mp+G
18jWyBw9pW2wAwmMqzqC9Aqp7oT87E4pFsKzV5jfUQHC8/Pz6k3PjNG6GeXymas6
cq/PPESs2UlK8wdDCOs71pyEDAkC4klaIAmD5SK2l+83MPLASfyCoqXq8LUCoWK3
IpXnEJHb6ZNwHEfynBIqRESh80JJc94tag7Wle1o0eFvzU3Y6j1ZA7GiJ9No5Udb
Z9IpG2tlbJDEPqgiI5x1SG4M4EtYpiNqLPez7F018eXy+rzU2wiO8vD4BXVlUL+2
o1qjsqGP250vVJ9UEFmxhKl5EkprU9rbVu1fgZ0Nz6FpHCbaZ+H3+7OvIo/8J6fx
I+L08YHS7PpJRa6bZ+0Oot33mhlaEmDQpm6RAfPV4gXfXMpZby8Ad1uyz2jJ1GrI
jEX/izy8sSWo+l9Mx8NuJ4842/YXgjyApJitf412+RxUJL8e2SiSf6nRY9Knr5Ez
aYNhTz5SYt/zhGHGU1UTrymm5bzbXi1LaKqdPK8GB0syQgk0nY9GK6DXqtj6lZxl
a4MexcYk9XDUfsBnDlToRHnuCK/6jr3ZOQQR1dvpcfyHQ1CkYRHo3E44gt+ltLFo
Q2Y3rlZOHOIl28GpnMgAqVsVrzUFB9tRsQtjMvZkK2M/+3rTq04MbuG3njX7eq35
lVvHpaZLmZnDAVXEgYO38KZunEBYskA+uaPPxdE5byQHmMUgVmVofQvdPtQUd5F+
xY73OP9K+iqFfrZFX4z6PFm6D5BvpGIH9sKSC/getcYwluZ0MdTeDU7TjBHxcv9D
ERtfr13D863chrl8M+AzdDiSEoAg8vyRrZsErkoXX0vmcHhG2WtQPY8eu6Bv++Ez
/a0CeHJbjgmex/GR5EOC7Kjmg6RpLhHxP0Nw1DViWtCqbOhVJoJezsVrg9+h3JB/
X8QE3krkmDSyxg/xYgnP9M05R5lPzS3V99bxfEhZS2TkPBiRxc0Cvu+x/H0Fj9zu
2fNSU6YdCFSTeYKZKFJcOtGaY/9t4vjb97+igQxhjEx8SxIEHfjNp4gXsu9ZueD0
+AoGz1kTWKcYBxwBpZV/9nubVcvBWnRtJsweZMAfUgRwP0ZdG6fhYo7iq+ULSoJb
GpLXIKFLCG5ZF/iNstReBzmyuJDVMi8DVYCK6ICjoQAgSjjUNaWRfDNDZEx+9amX
AUeevC9fjJ6GbYq76AhPUKQMQd8GRXc5cs94PVKVseJ2kBGcKUIvIt6aa+xOcgDT
1NpeYb6Y+JbiZpgqLVbGa44MaUzAUABjTKcF4oAKgrdQrPwZskUEghanyUrc8q3K
9/6IBPLEHX/r8+Mhxd5v5r9BiHz8JRVQ8pY3G6t1mdYSWLaqD1UJnAPHhYVS2zqA
X/945ZaTMUqZvRBORpFONO+yDdO6eNANyf+zCyBVzrqn2tPj5Gf8L115smHh7ybX
ADUjcMZflKb935EYvcc3wDKIRXUmqxPvzYsX+sNUnH9Lv74qlpSeDmwDipBBRsAT
QV2bVNLnXFP/p3LyA0p+NFAkwfxBq6MqiKR+dPUd2XEt77XzX+O0Id5MQHYl48Cf
BTke747E53VLCBHu5uHOuA9/4JUO4Y/t8etVYzOwUFWY1OQ8tGmeC73gh1SsbPjI
Ft9pLboo6eoue49laF5SvjRj+5GUOU+UHJL5zvMHTHnxgXi57Jqgb3tQAlY/hREI
szoWUyDy60GmL1VJZ5yBaEfVkTBu2VKeLc+EXCMCrFiqbpjt7GFLmlnyWG3C/z6j
v4Hy20HVb5U40xS3F1abaW/136GH4yYn2aYatpb82F60OT0ccsLADuCReKdNpWMP
K/MuKPEUtcSBxtLSH57k+a8d7odqhRgvXHN8wmsn5sIfBw5ph64e9A2WHSlWaYDc
XvDIuIHwofk+NwKfg4N1CTs748LYtdvt0CfwbEplWM7M6VQ8v1t8rJYRC4c++W5U
NlrkbLfyg/ZDKJFsC6aOZPZCUl32HffFlmJa3AgTqQX0laFZa7l4QKWZJMPAwuQ4
l0dDubZn8tAQt3fvftdRzVev0sSjhFpvY6GVDUU6V9mJglr84lRc4IaiH+cJQxnQ
sqDfm12lFF6xBZZeHG/fM6le7IMLJTJvAEgYRODMMKDZTWrng2kKCWG1jM9/YE2K
Pki64aeJtFqgSSe3L7W/mevl5qNoB1WnDTBV7VRwiM3G/ZNeTEqEZtdfefzxYl4B
Vo5/5z0EUEI3dhWtc/bcHIxvVoTridMWDsAgGetMDqxn3CwQjjse0wAhoorSDhR5
ttxIowFmYYTWiXIq4h8WidW37v3vTvt/GIOBWys9my2dU0QekzbE6eISk0hFKdl0
3YoOz3SgtGwtqsFa1cgr6EDfLn9iJ8OYFsVKIWtl+/yo80y5blgb5c/pqug4MRV7
zvm27BBjYNR+Y0yHOpkUQ9+SNX/mdVMs/zkTXFiDOgICNmIJbxH3TvMcEyO8RpVw
nVKimbXYiP+FAtaGWnT0EOvKeMSGHo14J29/WE+3962+ebYTqYkdIe3HrEFZcOQC
bJhr/m2L7Y3kykF+JTAk+6cafBV34tyC2Vi9KrYS8NfBkHOxxoOkEBll+toNnWEp
tkXzm8HAMqk1hHcrpG+FzXpLCeYD+shekaQSHkolX8ZOAAaaxZF6tUTWN3CuJ396
WoqGgT8USgkxO3IntWXjusVYzvBuGe/HqEfGKKefk1mMUfy5iO2CoOXP5Wb/D6e3
3/6Ezr7tw+NkuTUf/YJkkMzalFgv+CBvhXn8WO+/mwBJeCE0GoUIYhBiT/u94oKg
N0dMGL9MrToL4cpNfzz5UWVrXSKYtaXAS54VDHBdkvVnbTPNKaRhUKPFBRjZc3uj
U6eR0sdWx5ujZsNvsIhJzT0JlE0Br6M5R99b9WXzn/a1Wmp3MEVwpN7dylFXp+8t
B3+BCSkmP0QObbXuaAsvdTUPKx6edK/UqGTkmMZfwT4YG8XNXii0NTevvnW7mHZ1
dTFZBsYZuhWuNkUKK0Zr2IeGaphj0HoZQDGIMepoKGqP7P/38ouBClR6ehpn/mww
D9tnAK+88nkMgeXyY++y8u940XBObfJc/HabXG2WJZuPjSyN+MJk4n7L5OnMegp8
7cWnR4vDrzgEHwpo6eANPwIiiAA0pleiNp3KXtX7yczDZqmqgtuu4kuOXtKox2v/
OywP8JyEtFoqiw8wk0dzHAZvH5+oluORlLzl3YvtyxXVwGSNFCejfqklp4lTNKov
YROg7tcYh8Cba9NWj9+rPtYbXsDcC1JtvbYJhRUQ1mgTf88cuiBPLMVO1R+ktMnA
Xg7V6qRsKTTgY2cEfE4AdOC5aJPi8bGhnVAyiCJpIkXSSoU0D5QEwOZ71Jv4C5lU
uPXY8D4nTfYntFti4zTj/u27csjXiwI/+8z96wBSzw0gfyrKt0P3qKtKVK5pZMeT
9uGNKfX7VvymmwtkUNZGz+PMFXEp1wvyo1MRmwg6HGUYUlaO96lkOTF4IFQG8hRo
ipSSgmDAxzgKS3gEO9+1b3Q1xa8IUbKKuQ32jTzdba0/OHZ29XPJcMqwQTDJames
L7PE4dPeSJJYiygfZt+7/0odqBTommXJb5lc5gzGPtTNK96LoOUbbLayo8rHaCft
+mn7PTn1Gp7Juk6FYPyMcJU/l33Okz10oqp3J4qrK4lLiLdK+kdM507p598Pl10/
ZF8GED8nR+wNi9eEhHVnBhIy2R+SkNw1geEC+sNlpArLjOaguDyDYWb060/NlgVP
pIi+K/eQ2BB2NB8ZCIyGZ2zTAY3LG88ATj3dQ/9aW7y9e2jVYb2dXDo/aClpXq9+
DOh/f+YZgurq+z9MF7m5+wIOvqE/gBPdqUR3u7K1j86vbwvbs0MfM7p3VhFdh1CL
WrbDqFI8b1yskLTto+eCviAArxY73059WgVAeeZuHLlo5Uz+D5mSWkohujPIumUT
3B8JQP/AoyPor/yi0XwlgG2m29lRBfHQzGkIZWhajlKGIhSoRHepDhq00m9TPBpt
rk6RuDPrp0GvKb8+C9EO5SLJFOUWDmY/LcagmI9RmLAzYxgK29gJELSow8ZROzBS
Y3wZDNz8JI2PEijv6yT4wYazVR9EfVkGYokhsD5qzGu0Gp3YWe+KyObgneLmhiUQ
puCFD0zUpasEgMz2b/lqRCHxX8FTfqOJys16eI5HOWMNYNwqXZbQuUUHR3ODuoK8
I1Qs1NybyAORINXhqc9IakFU2Fqb2ZvH3CkmC1dDo/KXmyd4IGbIWdVQICXNIrNZ
pQqGHmh2ficCW7rqRfP0KBN9uefphybaL38XOzvGgjdE9eRnpAsQulAZsPhlYub0
z48yc8JzySgSul16qtLRcl0Pv0OIP4ZB6tIYgiRjqXo7RHuPFZ0p0mcEoHUVmDCL
DjniTJcOWqZPhCj9rrBwAmn3aEbFsJXs8XA2MmCIx+WRkmNjunvxOG3CLKJKzg0o
RdjZa9CQu6fZ8r29hF5WhG3s3Vvs0MgWURgvcWRXLvDNRz1qnqkyqhBybprovohk
/lLkf4slreSwA7CmGoEIf9dkEhUvQak3+fUG8TDjvPe0HlJHbhzAlAdp7Xd2HPqu
UdYFFunB3PpT6XcfSA6biOHnTCM2mgDFaiJNKPfeIxOdKyBPzTY5y5IbYGQTO8/T
3SNUMMST+hw/hCurY7WuDtAgguI1P5ikP8YKbngGg5yXlyShW5Ds5RGXvxWLLkdE
q5qBRr1+oFEYxAfY8apkayV/StlqpSoB4MB8/ibOCW3kesyPMKLlvaomUGdQOodY
wYzr70l2YKNgmVek6na1/NjE/U/G8ynX3VVsgCfmQVeL6JiJU6NbD81Wo47l2Tp4
B6aEn4f4qTACR144JH/T4TkSr2WOaDH8bsV9SOklla8odXcltzoyFWQSbciW4nrr
W6txz8MVnQjd3p/ucLrHZ/MeOQT1wsjRHNyd/ToVvEasnjw55hnHty5e4mWW3uju
IOgYWWK5NObKmF/1dOT+FNc612uil8lDu11siJXok/wTkOfQZTQh1r1jIqChIQ1M
3M8QZ5HWnj2+NFpuQx7XtMxY7l/4alvb4buDFgd72ossnDTvK3vG9zrZIMv14fyX
kaBKvIxpKQzjfFJs0kl4+M7tETrrcFJsoaC439+L7Mf2qsZuVEIvakDKlcZC0IPX
kHPoA48xwau4WMcu8s5dbx2nZbOv844pnWlzOeQC177FyjqpG70rxGn2DTnPHHd7
P9dwxv0k4ozn/vkG1nxmZaH4Kva7y8Y2Om+BpEv9JtM9IuvNgj+/ikJIw/yrNStk
KiEYKEXqi0mvXcPcMqVgReB14lsRmJCLOq/iUn46XtMfSZWrPchuBHy96oIHZxeD
OiQdB3lMnLYgT7XaOMY5ogJ+u8xs6dbayIkkvyQtoKuNu4ostGQ+2i7sV6WGtBrw
eX+ccPoi6xHUKPsl0LyARowdJsld/tiSs8l6LawxbQzaI7plcoa9PO3Uc0Y35AZd
kCYWsOmLriR9oDWVwhl+zhoB/6fRApHeBvd8I73aHWF/Xx+4JTRa8+RWJJ28soFn
/eDdmsUmGw+d5oKso9EHwyz+yCA5bFF0upm/NnFIOOtUf+k+pPCzvrGOC7O5Wig2
eeZK+SK3h95w5RHnBfuRQ+2wvJ8PP3fxd6m0BJBqVI4webDFwWemG8PiUXvXQtES
xLm2IWCOC1xtt4whrL6yphIGxK665vQUaCmwr+0mjr62RzkHml3CJirs9h9lj7y7
91tn6zjyrJ9G/UsWLmtHyXhcDhju8nH3QlIllJy8KZrIKE1rHXn0mC2ivvZoslu1
BQsyJzNixmhLSshCpgPKpO/HWaUuP4mmYPc4yD+x5ITLupcEouQWZx8lZ4+Wg/7Z
260l/e9M9P2Mdpjl3z9FgIBFxBiA1RganRC/CXH/J97fk6EH51rR9SFgmRYf63Co
Iw5mkOaExwoNz2cNanNLf8Pnr84l21qPWHEJ0UWZ0OcdBOSslH9mT/cJAgJrZ7FF
B5uBSQEodeq0s9CWO1drFdepDFWXmOZZEJqfddsivDJT3SJmT3DkwwCGW9X6Ikg8
sReGJ0wTmsKKm8vZIaNuJIfYteNCM44j2uHkzKrccafEqCaa9l80G+9HRxCV8gwW
Bu23gsg594si7qx0+j6uBJfHuU+dDxHTj1tasv4mhz2AaieQMupxs7B8uIKqTrVW
Sg+pRWIe/xaEnsGj6b9LHnYaWXPzoFUq1EFBKOYD7RchvVL0KJyd8EM/XddkrT9o
FOM/1kUA2nvUrdrl/HU2OqY2L1yt3RJUs3H5BA/Y9XfyDCY2+33zanT2/sveUsqQ
xqDQUFnjgVU9LYs0pNg9ZTKpI1uBzVxgH8oqcWh1XvSvGNnNuKPPRwmA4/uFaRYN
b9GE4rqe84Kp8ZK8EafYEglCKpLu+pl6ZtW09zm3AEMXshcEhh0+dm8S8lwRubex
2d8Li30LzRte96i/GoEcpeKda0xmkaJKsAwbNYsYWDSMxaa3kdB8DeskuHK8zaYN
ljjnwBS5CDbtHYXE4vrwhkIMYMGTzWgyPRvXAGSPufxhkcb7gcEEjJd9TNaUu/B8
+usSI6tOmhMxeVO+vxaTjN8qsXgPOqelVDCK3JtChlQ17uAUak18v282Yz1j7twA
fj5IxhvjJ+JXLtnURDgeolshR1iUfUOuq1ez0wC+Are4Op4EENRe+TrfqlGOkkvI
fDfCkQ9CyLsW/byXbgeY6STNYhX/X7NjaFxKHp9CSzUBIQXcWciOkElw37qEeKWA
66oa9ClNN4FhglIyo4D5/wBt/TKP5xgJIY+BZuttzueGkvFsmNA1IhN6DB3OX39b
QK9XDl1IQk7UWS/z0qmCHXBBmo+x+Xi1X3qniJ+j2s9e8DxBzY/r6lJfpexeNGZh
+AM+StLUe+HG6HKCddMF7Rc8B25/IzSYJy0BH0u2PN/34W79UF5Q0L/HSTiOjdnq
bEuuo/se+4fSu7SkRmCuqebcpjQdkzplN8IptP3aSJ8WKejxcEW9k7tjaReZqgNb
wj0w/GHFdItatpxiSO1bzDsSMC5NGMeIgN9g34ifHcPV+GVzi5X3tcqfV7HrRYOo
K/Lchr83Wu3NIsZgt6u0eOFU/sVSPPQz7IxM8KZc3LiCxysHMfzMc8lVTo+ELeKr
0rNJmdL+59RI+wXiePgekw3Z7UinI6pC4quSWg1hd8mwSkQpqHRJj6mg+h9blYvz
79rQqgVM95NnhIULe6W7cTrbitfQyjbTGalmJsdV+VhYqfPmY0vZqbyaihOgA+Ou
T03BsOfAh15yMfTHJRZ6em1iEyDj9mB0k4FYbDXKvLZ6IG6coh9wyFSHTK1GbX2Q
J64pKTYylG0eWsy6n8UuROaP2BaKwOxfDZaUR/L6XRo/EO1XCVwU3Wdm5p9sv+Zw
d3UrGiDBNXC6P66YwVHHZ9z470btufQ+LNR4mNW36FLw+a3wAvfyg6G0FQJvaOGu
DyqRkv9cifWqcZMHfH3xwyAtNZfiBXpr8Y7KQhKyZHabcNjG+Vbpu976at5QPIcW
ewza0Of28sTRA1Ehdkqw1G8RsFdJkwEe9Ru6C5PAM2fvKKUnsmQMe+pzMweqkSrV
/ipprEwJG+SbSw5Ep4IJyN845BY3+yvphTUW1jqZiqSp1yNERgw0Idsd5OrgYfd3
IsQI+qjsQTVCtI2PNbLD0uHajx4jDe3WwlCXrkROj5EHsOaJleQ8BcLuSwBxvVd3
VXIxS0LRAm/JS7YxIKR9Va+6rTae/7gn18WvCS37gC3LToThl74Wi2/jaosInZ7H
fZWbunL/T6DU7xIe/gHBMCZ5RaptsXJ3bERzYKtDndKEGlJ+pCyR0jwNyWQObyQ7
RdM1DLFF0BdzCxJeg8VuMVZ/zH8le3JxexI24lcVkt9vUN4nH8Uug6RDb6vGvc91
vkIOIGjNHkILU9fP8VqdYhX7Jhsp86QoElV0/HZ4MmOuFwRL+NfYcDwXpoOUsx9v
wHmMHWsYRhNn3I2SxfH8lED+SqILpin3K5asQG9ZPjhdgn+RQ5r9o3jpBO55bIZz
hUjMZUyn0HKjuZbEL2Y39aan90ZN4sWtDOOmL5+rmmTYe7/p+sgzvcMq97rrL4Sz
71iMgm5Mjm2+QspIRoWYVlK329HLfy53eFQ7Xtop1I15o/2tjhGWsOeRZ5JgwOE+
ugciWrwiRNhcZ5NbzayqI02AtP2n+Lse/MbjViqEcIO6yiRszbplrjNYEQ8fcUlu
Kt7GRNjsoKbFHsJ0zYADjOhdo38O6OfYPKP35HcpzeM1VmcKUwdPWuxLUEFsrA3l
l+/jqFJTBto3kxFDMcRTHKSbwei0O0UeTFbHOzGQLjIz90GMi65IsPTPTAYMIgVj
WLRu+ZENfeylKjGBweNLavuW0YNj/o31tXs1IrMhH2oEzBGCsUePH2E75DndgWqG
8IbdQ6volZx9xDBrGrMoBHXnueoSapeDDK7OqwYylPQ9gXtEO5MO2Th3FnK2IXqV
V1WmP0b2Xj0qkTZ+HesqeC/zmnsy8T4C6fMlGaleHGDGbKDhSplXRgUuz55BI+DC
KgpNHOgHXa/FsPKvzwj9d9fnb0RMfkAzbSJhy8TbVq0cOo2a6ns/gHGRabXeNakm
I5UoW0/1jkvU9znoMyTyuysil7a5utBLIeZKQHrwX2f9gqzGLSvYuxb8H7Q/1HuX
fsFGag8I4MfWNSW3gcF95ftSbBv5UzHgQgUs7yqYYbX24SWBO+6JflZenqjQzQf7
5D9W//zFuUxopdraYe+tzCsmVzN1JjbKOjG6QUzOcQmY0FimX0U1yyNJJfD4oI0e
F2dQEMcnkaf3oPZduEjDQLUo2PW4a82wO/upNXAwbhxurH33UIsJA+QSzAYazqHv
uTiPtk+ZoD5me9nlbx/V4+f07G6h2AxJ6LYDTPVsNMb+2Jpypc/lN3H0nbtgOkOo
Q99zJ5ZHgiy1aZ0K77CUjbDWYV8U5ZDL5eT+tw5mPSCEDRFqfvONpFNQq3g7EZqQ
Wxag6Wwq3EB+J5DtL2J99CJiIvU86zYjXNaWXKuz5XZr2yM4Gw/FH1KA4Yhnzf6E
lrDKA5aJzTj77CeZvwdAJz0df/eDrSG8iwdqwJxtVwx1xprSKz3CmHeQxPQidTc3
x63ANWsRhf5GRsS1QQKgG2IlcjaKbn44XuA2Qt7Pd0mTh7uGsIFCygtu0+PvO2VZ
BJVsZjsrx5WC2q3totMCE2Zir+xtaYFaECFtbrSwKpSWfodlRhwK2lgtJxmIGess
FvnVUMeueAiR0YUvJR493QfgGkVG04h0pWxS9DvcnDBCP7mVcer6ga9x8VpKLMpl
VjG03PDZEcXeaupP4hyKd+ap3xWDAs+ta1zzkddRcPDgRJsW4TxHlm3qr0DtBEqL
GuGibAqgtfK+3DijVfzq0qVegvqcQXdE3zRPylDYhiuiTmnInjCBdSC0rGoNiN1l
tjsVKfVzSsYIY7D1PRlYzaNMG9Ia0t7pNuYPD3GnmptoIxprV/QcZQnyds9OGXk2
35VXcFJmWCGOnBCWDve+8EpWuljSR3OKYx7s1B0XTM5N5BHZfcofJWARUGgqyg9w
CADCwVmWcDbLkrgS4349uwFK2giW2X4nhoOo8l86GTC0Q12Ia9zqS7sIC/7/vi4J
DHDd1k+U6o28eoGz3iE8YDJp/UaftJ4twRJeGv3trs6eZeTD+d3PXKPZCP0aw6TG
tuhexIXsu0SFaEKRVvlHJ3wKm6x7XRW5cMZEQgUHilOyuj4N4YRC9yZ1VS6uYicC
fCMxEyryxnjsrOvOEJoBr7XeurBYxzCA2LGvzvgdjfNfWuSLHZKonEzEa8Qeh3Vw
lmW6jrt72bOAvHoWURTaumUGTm7U6youvugPjRvvAwhtPm0k5FdQBKfpfi/izbxR
qxdbdoRe5B/60r9i1oA5GSAYIccrdLrPuV+B4QRDHwlnm6DcGt0IIcDpHFmLTpwG
cKJapUXCCgKqBZ/sfkJjjoeRG8MHZCpjLKo7atQknQP/KRPMb4J90ZevRUyDUb0J
MYgPXl5b4llOSi68qeqajxPK1PEUiYCt8E14Uf9xdVoys9hnYHi732S4Knzsgxqx
wm40qV47Mg45sC61hB3qs2UT8NuLpp9aByYa8aadF3AlZVjmgpiHhyhbCKUITnu+
D3AH6FzVJJYDVz6//jy2jH1D1Go8rDuAnRsv1GVTGLtMBrvjO6dEmP4YnOWNjlRa
oSIHgDYEgAT1kbd3pTYOItca4t81IrPJ2Som9/m0G/t8viWyZRrdfTI+7HOjcjYT
B9Hjt5DmM9ERQEC6A2Jj7e8jeHVpQrHSnHbB3FKKepxo8vwmTjWXYJxP4o/Enu8t
/mOIlAgEJliKjANYXVcISNhqPmaw4hpZlFFXcSQcZakT5fDlfCj+dr98/BafE4my
Ofty4PcCwdW6S0Z1F29kPjbBpSmWYjr0iwPOt09VEjaIho9+Cik4IUl8Lft55YkM
632OKY/gQ5+opYudNV7hevtPstQEhfgYGzemqdmPmS0amIOn7+UDZI3Ep+iOSGjk
VCvpHoZpZX6Cl56pvk6b3yRUx+5nNy2j3t6FVx19+qGZufWZR7309jo/c3iIXFWz
EOM0cRaQmsrnCnzWC4k3VE14IzE3UCbam4P6+4Xp40e5XhLrwmSIyLDtEZCZ8ah5
uDYnPdcjrnuS5DtKmfXhhpIFknT4kjDVKLVvrV/31nCXK6/7EIIrfPPS7A5k4N57
JdWl6+gjgDJW4XJgoz6iT8FNxE00Og4NVBD3AtIP1+Oixh2LB1kL6V4R4gFKAJ3g
CDGEZbfA+usk9zBDQpnyG+NsaTnRko3+NQCJLGxurme9cr03Dc5YdX1DklYeKlyS
3c7doZNn3ZfRJQr71ZovuYEo1RPyrEM7VMEoMdVvCwOuLAIbym6dlGtexxwyW+cQ
KLqC3vNPwyrMV/8wnE3Wpuav5D0HSgUuWqE/S2sTSbqfZwV2t05q/nBa9bhThpSf
EQU/hZA5RtyqK9n2WPJE8EmGv/fgMM/NoW4RKK/SoRK5Kg/8yuWfNOm6V+ZmXfQP
tLwRq9iNQI4qbwZwhGaIbYHGwRYHDchjWW89El3S1JktJini6MzWc/X4HzVCfTtY
bg4tzp7gEQ4VZulj5QmLra/rM5P607DYwz2JWja+G4l4Yza3Mcff1tfyFLGT54lc
/+eDVImwM3245i9KUmFn2SW7X4FjV0HAVvRgV/Y7byfPW/B6o+e4yKI7mnSzbMUz
NdF8LSb4qT+q6Ze8zWgrXLq6bfLikFxO/Nr8mDA3ekdxMTss9oH8wcwG//2jgClk
cO6R/1fE3T7TklAVie0IHJIbzMo4pljVANvIGgWYoWnYFzP2dL6oH8Egaa0FZKcB
I+DXBboAruuYa1hLXk0f9+CCi1/Db2wrgJv9lSBW/MHmB8naFQaPhDxQGktXZQpI
KPzMHU4MvlrYkTzVrBREKQY1vHHHIwVHIp1WuBFnSKAjx1hVIKdENJ8DksRWQtM7
TKhez3iLaJed6QlnT4I7420lbLX3MGlZFBt8LVVOB+LwqRHBHzXa+kcMYQyz0IRl
QG/7c5RZaoOYKp0O9DWA71hejaGRPaPoJ8nfVduxtN8aUjJCb4zuXcW5q9UJ4fBl
vt17qHFgh+g/ZCg/u+p/3CWPJVTMRalrzQh7N9F0TquZYE+yo0+IdrSZLCv9phXC
uxUos7xxYCGRHYM0srK4fRRemimYNYHzTW+bbQF1fKFaZ4CMOsnaTU0dineTPFfr
VddYIxxH6lUCaJRvuwlz9lVvEuEhzIeSH0HybF02LI49QseM9RdWy8/HXeIVIFvD
UmedsMDd7fUS6kLaGiWg3oMZjYPtXMTxj3aXub9+tNf2RRIo4Qec+4dWQGIj8qZv
bMRFDY5mL6pNWXg9NvFM/FesjANKemEkpQl1feiRp1QLHPHRt4qmCouOPmCK9/Ca
+l6WhlZw33VjOzXaNre2qjlSX1vg7W5rnniD8i7STROgidDRRudS/bGN9K7q+6Al
Oxm460DxqtP/sggChB5efFsJuTz/XNnMkZJ5wUVbPytOHgAqGU/X/Je0QRNMgSdP
PXbiJtAbfIesug/h/kWcA4XW/3DMojpypXOAwO1Ypjr0rsuhi/hf1iTVLtEDGfmv
TIkqPnyr5KAE6kiVe4/EPMccziJSFhvQkcsRkiTBkDAEs1zs9lVfVdHWny++Qf1J
vXEfYrk0Xmh9dSjh8b2Lh/yQw7Bf+jMc62ZJmLsOxSVES3jMEi4gF1GQSr9Xe2be
UK9O+HRxI/qS1mP9dhr3z+d1hdVAV9HkMZ/PQ6ap8i9n2uDHoVvHqhg18ISPTnTi
nEyJIE39u/PbjrvHRdrwaYBb5ImyuHM6jJlJCi+9Df8Vd1vHFJ5yhk6qe+ZaiZvU
RmMUlBF14cWLdwutGCu4CyQRCL+Xz3yLAkMbaPSsWs/thh2JR9AfeO3SfjpH053h
akNcpGgLqmcdWdUrAGPe1elFaXl4CwoOOtzpYgRg+4Tez663f0J/iiwsL70BlwpO
OqwxXEjkzjW4QR7QXW5lx/T+MBim953Mv0VSHqae2aWF0YMqnaSKBfb5VwQxwf11
fvl2JpXXTbrk7eZ5xSwsWM4HL2rJ06I4g1XsQOg8OA3ylUoCjWnPLAX21jp4VbvX
9mtQxWWQkuFFm3KJysO+HrHEObJhwFsMblya3QfKx/rbeVh6oba9OmDmd2hHeGSS
4JmdHEV70ZS2SRiEdzH9osW/YYtxZeR95B1oZDH/A4pylMK7aXk6kFF45ZB7+l/d
W+LnnUv1mQRsikgHxVZB0tY3DFGWEULLDIERmH2xy3rN4i+G/JgTc6s8fe9Yj0or
VdUe+KGF+WDvcs4pQ7zv78T7f5VVbNP6Wbmb4+kRcK7i3vSuiua8jXWQpGS4iEht
YT5PtxkkmB3Mva8SCkk02r7WHiacd4wJCxlWSUgCaYOkCVq/Pj1oYlMqAzgXj7S7
JTGj4BswgK/TIioPDSnWB2ihWYQ1RTpSvB2IBA8DvIUHBjeqwWeeBLZ6E8o5dbt7
jSz+T9HqAiBT9vSRxkJuQVrASUV7LtI/TBQ8XzpupUr7cGs+/MJ/10kP6LwflJeW
eKCH20AuTUzC2rabER8ctCaxxL8Rg0SjN+0A/NKbw+1zRnd6+slfUFnttVdIRM6a
wqKH2Zvm30G87B4s5o4DXSmCc09jQxFQgfmm5XgYNPXIjF3bVmyWjpucbMKNpwzi
cybdcvc3eeNhatDcYSgCLE8VCvfbTAJHzn2gMOABR6zgSSb8HHbXz7W/I860hTeg
T4uemxZWt3yBQ9mT/zyBja4/mLixXF6fgKbOAZadt9tNFufJT+jqiPoLPb2tcsoW
sVrakt7nZtCaqGAA/rW9WuDBFmvI+TyFzrJ61doAQMfLzj8ZYxas5ETvv3C4t+bp
xtoWqiy9qNPuN6v8XUz1KiMKu/aGtooGwgkvF7FkPfBccyyoPqyTlOPJghSvkzxz
7Z+HuH650OAnVGCwbLqhN5yOuI+nLOiAOXOYrS8lVJ9DtOPtA7/70XD0dIPsH9rS
MmijCr8uWr1vzq5FLA8eP2BD3VO142yrKO+Tph6CUnHuoGFlYMeV4CeRNqnatRR7
WzY+DBnyrZhEMUhetmjDEKxg8VcfgJLOH2d/KiAMa1dnjmlca2PtPSQGfpfrY+MV
Y6nuLv0umSccH5TrdGyEqLtL5hGTl7Z0gigQ/bvn31GqXn6L7v8qxbPR8RPdtZCY
kPej+M7bU2EzqFGGRb7P/JN41op7haH7bcs8FZBnQror9ILsU7FuXttb7bJPvBt1
5GfHiiQuEwQ4Gx5ctx/sKurAWwuENhEeLNwNoMjljPEDSnww5CL/pjjUSpe+3uCZ
3JNMqHWlQxpUxKrQUXWVvu0C5sjvxlog4xn6afjO/CC+cjR23h5xjd82P0rUGDqH
pFbvtWx4kG1DyPUj1QRoutIFG5bAlvIMRHjJ6U8x7KY+p/9sdOCDal5V0FHYH+Xe
1ZfqDcJLvSaaLdg2uxlkbOdER/dv/O63xFrAG+GFDBqWkVAs9EZlgezqyy+pDC23
nD/eUlA85xQxj4TMX1FWxHx2P6z7y02e4hmlG7iBzwXz24oxok/OD3PCWUP/9a6a
6TE2f5YwZQAo55iIAWXQQWlq/6jb1NsJbg4OvKxo94nFYxoXkIXcleQXHbfM+Dnj
kIOAeVe6vLI0INNs/1WLiq39VFfIG5gmI2C8glEEhyGfO91MQDUG6HImftf104BL
4SgG7sruslk11s/9ubdOTBTfVqo5qhlIb230pDxUYo/fsSEgOpxDnbBufqiArxl5
OUO6Js7embhE8s/E5Tj/LrJBbNygbM3be8V1Dv/sfa61ypmMWxAoRdjZLpuhe7+e
1Ml1PYaOSLcgNmK6Eh5mTr4aZAR8TJZQy9WKOm4jCLvsC/PdjVyLGqHdOk/60j0y
VpqYJUoMrmVrj/JZrBhYjh6v6U49S+uXpaQz1JZU6kXBQJDxwE5UkU7DVmXb8YlY
AG9I+pw6iTSzjoyWYgxp9FYdPyZGGhoth2ZFaVCLaZHkpno3NKh4uEtA2SWQOKCS
F+HmsEv9OPeH+WEe/jcYwLt/f7OP5wj2O6PnNZxDL9KHShmPUh5SvQf1ipdb498w
fWkF7NTjS1V1gRTIqgR9tlq0JMpUedrKecajFbzY+ovQU+i5UXzSLbkLCpsh+cTf
ClY/DduJ3oRp3S9vykWvrieMc8sYFesSQ7ZMg2I6LCnBeqE8h+gUKcQfTnyOz/m+
1VSILCejDubQyIGkQ/Ouo7/R0HM/CIzLs9/SRAGj5tHg6biCNTnSkSnlRW2VVVrG
BTGgq1V0Y5pBn/Y//o4o2+RKoWw45oppQ4km9tlGM/AuwgDoguENjFA+Fcx/6UwO
1Vfgdk5DfLI2nch5UGH6+x9C9qSOYrqsAgzr/TwZs/4DLOSD5k8Lf61kBQUZ1wYI
XQhxzQtenoVfqpqePCQ9kHmrs9vKCbahJVqamM37tkFdunkk05N6AgUhTzazIQhl
haONLy8kQSnW3ZVUDhFLFZOlRE3BfneaXhz9+oXg8Z9etLEXuEVqTQqwTG+xLB5K
XAFbMYEKWXhJL5UwYVbQPk1EP/9epe4IsNfAu+uGlSK8UIwyEab7xTReSE4g3p/C
SnxpkgtK4CsriJ+eCK7keg8NbhguLMA2evHlobgChFkgfbBU0JBIHZoJyTPdH+KP
vAi0ePLgOTdhRow7CaMjVTEN5yWmm3ZD6a/FQgiLsoI8nKNtWBUzlfUXw0oQ3XZJ
/+6wiH/Wql3rFfKDb6x3dm+QVD+SskKBMbrf/ZzC7bVyxdftyM0yCpWIMECPDCCh
6KO7DQTfBQ//1FzsbXFMuilxx5X6iQ1nAdeoIf3jxmk7Lr+feNKJ+adiQRoMTLD6
0uZxrkmVhSP9l24RzisBY+ojSawoAKSRiqVPJ/QlXqfyhqMb2nE1JCVZZs/og5O7
KA2phF1e37LWZmI2FZSBrl8qKad2Ouoo9vmTyDQSrRlignu8x4TxLNf066pdyZsB
4uOaEqpg+Lk2FaCHQlA6insp/aWX6FnICViMYpYZNEh75quoXCbwlGNemlKpqB8G
4XXdxKhH7KAcEg0vkBOAtmIX8lUUHeg4zaAIoJx6afCxlFEGhPL3x38toyh+/0s8
ABFBsiG/cgVvPqShnWR6iKG1gNAJTSANHVvgBNBB7dzuVPHakKy8LH9GtZBwUdHo
/c4bUGkq7qG5Oz9t9c/d4yKjifWKzcuaYMkTYQqi4I65fN/R0u/ayFdnUDk+A8pT
TiiUzXA9jzFMUKARRAlPPcquyOdMZzejwIhMIr2OessiUcAR4Q5UA5ZrBYSBg+rl
zRMTocR1vo4reKLFaszNoCVMye/oraJDvhuAUwJkFF3sPLHjFi5irDgWEjE6Q9oG
l20Q0RcvrYAL93aqZq2JJNgIsMMJ0ucKfSGZISK2b5FsBK1Av7Ub4iqHSuwVG6yS
CnsDkGObC+IIGgIPH5y74XEIgTunCv56Gl7PxY+iidqdSqIKP7linKx4PD5mPokO
FGHy/QQhu/PTNNHJ45K64BgwaQhiTwyHSSO4PCUX//L2sWX5o9fP8yHxpNyo36DB
eXpwRljaP5ZV+8F2OSdvVFC0CUFbbCfZqZ+acyGUMkurjptd3kexfMBoR2e9vTL+
ZMnEg6DQtKB2p3Ae9gQaKGzLFOlc9LGuCL2ymSPExJ9+CAiwBxKg4pJO3dptR9nq
AFFPN4BaAzLg9IeKtS3lPj4MW+wyeYrDYFIQ79O7hAmbava4a4+iW8T2ynGLO8hV
dYGQpI7SzeK63oRZmwksPC62xlKvbtyDSvDpihWrkuezfW70Qtb4YF67VZPcLZLf
E+JszdwrcdNjUTq4CeJ4Z2/juKBf+GdQMw8wnJZImiKM5S7ifo3WOZ9abnJiODq8
o4IFnisxLMWfC3ho/66o5V/aCDLgnmdglmq7xE38xust8dO8fbUV4delaN7gEg7J
qzxt37pIUzXBOR4itQ+vWQAFbQjSYfXWhCMe3M0ZErtViJtBprhTIdvpf5SDqis0
CgXUGmlE1BZHKHEISzNCeQ3oJuMdhx3VMPH7NVGAgEPR7Yz7HCh+S1mS5t0gOmj2
0Kejh7P970YkXbz8iFgnh+KLVcd+A/wPk+5aUhsZx4w1++1JckY/4b4m/VxzFaN7
vOvtb+IzG4gG0jMZM45STKW4MNVlYQkKZ+tDfXPPBaIMbvCIgroZI4fICgzsgmtP
k7rsvo9fhIRHfi4w9W8ylQdFvumll8hxhqUpKgo2FAWJgISXIF2oOPkRth+HJUfc
ljnctV7baP3lpARzFgUofExB8PjXFnBozPv8AoLcJ9OBquL2R7TKSraG/cmUfz76
qlzZP5f7rRCY6ltleeoDRxThA63nrEIDcufcS4p6UGlMEHb3mwQUrv9tOlXQq5vP
voQh0nsA/tLXT4AH/K3unxaJA3VfYY8OEwJ1pXrWOhQcy2kBuw6mqUbMMYqXEjVt
S8j29s1136RcIyoMfew0PWUppwWPucfm59ftuirmJDfvdTIkC07gREkMqV6Gjm8j
4PUaAj0CM8hWQk1q19a2PlE+7IV6VkXAgzoog3VBaZh91toKdGI+eEel4yQkibrN
hXMyolG2D6pbUryDQ5ayC1LNKpSbWUKSAJu5KggjHsQLKiJPpi/Xxw2lxpoBLhYz
fV4m27ACpFk60jI5nwNFWBqtXUyAVNZIg4mh9gHmh4vzoat3gR3p+ROrhWSlxwvt
XRTUdoan6HFKvf1EfwbFB6KeoVDrZTgG3ibD03qn2cQHJ8Ne9KAJgDkJKXc68RU4
kyaUPVkHnHKP5N9VhmaNB6wIOKD2CGMsRrNvImT3l//yzGot5xggqCL1koRe8/v5
trlDopWHorT0KrCX4MBFhoL1HDnTx+4GkVLpIaaQiX52+zktHD8drgGfl+mcEp5Q
r5OdZYMTse2gfR2cw5sOErGv9s7hgZhh6iXgTi12jKAoYSfUw/jjezQ4lMEsAjA3
PGpWNIs1vv3QPiDFBP7x1WEjPZ1BcFDlJUS9k37woL2eETKLhRI+wibQc7pNaMf0
HKry+pdGRB7lXKiffW8JdBCMd49LIS+uie3/xg5Q1JRg2WOD95+8qAVe5uHyWwiw
B5AVoqHnODPjZWWSVHNtTkZhL4NRKR495ybH20V38DTmj6VQLVkllqz4gt2qnqlT
dh11QG2qHl3clNnZ8ap9oCWCneNrOLMZVLSHAxh2Ayy2dBERCeaLA9tZX5EnOESY
YIxr2OwMRgm29Zoyf9aViBkw1EpCG8Ffm8tq/MiVBOBlI5uPqS+Ol8Yr9sE6+fMP
vK2M5LCdNmAbKhmhyZPG3hitmFmR8bXMgSCapR1I4IZWuX7F0q8QhVwCOHyfFhmn
te4hSmlEFLDHsBObzFWDtwfMmiYVif+2C3hC3u+1XPhGMX1YxJ1+cOAwyDBcRuNE
FP467PImoezv7HYzwe6ZegGCWWIx3L+IbY0r/XEWw8CG0ZEbvLv8QCySOoQpc77S
yGFn2rAgeKSrqFB59oYhM+NWmx59S5ql4O6756Jb3h9yMZ/w0V7yXuD0VqxEVqxE
qZ4JkqXQxQrR9l6qryjB3XTHIT6fTsMjgCaIeF17j/sVsF/AO8AxFNxHrzDf9xsn
R8/uHsUhf9WBqq/67xVABJIxK1ayKRnQWobqp8l4OYtj6Ya1w+xHMugJ6RmZ0IyB
/hQ2+JoGvsbOjavhVjIj8186n7swa5DcbuyeMnblW4ibgAlHh8EOhO97qp5Vd8PI
VGgbeZa9v3uiFEdoGs8Zjm3dcl7gkT4l9cTxdhqXSd4pM/8Jr4u593f/A2iS6d55
mC/babQb7xaYtlX6VfFTn8NvCMUUJ2O5UFBYS7hcLunDAMJyw3/BbYfVnNIA9CH4
YJBmj5gV7/qRx6dtTfmMIDxKawgKTjU1JhDvabyYd1h60zU3U+7qdbN+Lm8IfUuJ
wqmLdWEDcjrwTJlqZaF/iuiGRP5iZG8+Fux17LUdL69fe+v2sXZB2sL/iQdJu400
vHedHumLSUCzjj+8Um8iwaMROOVy308d8Ln9BtJ5VOHdBdCvL9u6cwPmn7wyUafO
peM8vaSxp/App3vTODaoL25OHhp251nifiAWmob/7NF82Y9NLOuKRJ4b2EQ06fjY
NCOHAD9yyCJTrD19zgkinlIW0oCScUkY2WSEBNzKsonoQP3237lVtU6dFL0NPUDK
DaVLruaxpqXvBIoo3Kg/7bgYCNfWxk1ms7kOLJmsgY0CwldUZtXHplVu0Clss9MU
55V3dTVbjiQ1BfK4HS/6wqhajhuttZgxSAsRU6L2EnT2AnxRieYPbse9ckY1ZA3R
l3u2MHdmI7SD88ibfNL2A52XN8QTxyq/C96r0mw/5LDY/TU+1Jn8dzhoN1LaYpID
B2JJ68ljY97JCeLelLY98komnjL1COiWg1gtIZSspbBbnXXejPzFgzEW3hLmmC6l
KRFok//zNbSyNPkQoEYOui/TAvHgzmcyEfJVANL5ZlOdHNfdSILjtOjGZaIjRl+k
c0yA4+9dIOwfSmMwuD2Ql7njqqcnVOizLJ67jCARVddOnXuERrPNPc8LmWkNgdR9
RySNpB0ERHrCAnyPrskH5eDrE+t2vSTk5TrDEcy6j5eDybk+t+Wx/6Uf/IKnGs/O
MHpWWdT+QzK2pox6keVpce7eJXw5NFUTG8eyLPd1tj8CCqJO8AbqSxwn1S+tx1w4
KfmjhOy06m0hDXY7ZssBNDLwGgT6dZP0mqO6gS1ni+eIegp4bg8tufmYv3ZZ1GKa
CRpMhtCiRaX6N8yzHDH9tZ21oRnY2mtQS2yovPnZSAsNie37qf32kjnQ2im6ZB/5
1XmvtMZ2TpR8QLQ8PDgD7XsHe9GzKxv1jp4MH3Re4qg1bJIC3vKubAvL5ROH4Nl1
/sGrnRfKcEbxj8uW+Act79a6TOsTBZBc/VjVMSGW/HZBx0boMMkpIBObRoRwX+it
OVI9Shqg6HeFBoxVmUlGwAvyAsvZb8NyEGLdhF/RabpiaToiHf1f0LDjE/55oEjP
YAFGo/yxiWTt5RJUFCM7Xl1QrhZQt6EBfReU9QuohHUYre/Z1DeV6tukJcWWQOb0
jAld6BCsxvyNblfhsikCq9DGW0CTn2EDkrrpal3Mlv2vGn5moQspN424W+rHxLaJ
synZPSgUEzUwoGlt8SMUGeuQ7yvKQFMwi9gJ2z7DRvcl/DfWKac6dzWf4Uuw5kWV
YWInAa/nI51xzUngaLKcFv3vELH+zZKzPjMQmWNc8oNOaK+StImEogGbR8wxb5Uq
vAgOAx55MyxDK8BxjxLx5mq9burrKw7GL/CN6thYUY6LBV7qaRmVxHKVCcNXrX6t
NqDldIkpks8dS6dt3ViiQdBkc+Ng8A9Cu3M1maBZtJk+XS6fnBv4VN+2xuM+1Ydv
hC50mvRUnOmGUgfNhYW3XSyRv2ndCY0/s+kXpaUQ1B0xsa2lUjXBRnZWkm2KkOPR
Aag0WItD8N0Xg1QO3gO+bBMqk0Rp2zgTQYvydqnw3jaqM9ikINikLWgWGELmnARx
TK6BfnK9TUpq/c5Uv+g4qG89xjkeSObrkkKgEyWfjxMMJrDbXDj/T+dW3UEuHxfU
9t8QEbQL/g70JHO6Gy7X7vsL9910BaGZ+YIemGVWwjySZEeaNL1reGVvywUetE8g
U9mqzmKnMMx41QZmN/J8Mwi7dys0xM5DKbRJK6E//swywfhHAgpdEMzUoXX2sYkm
Zi/0USg+sjkIq9heCzSQ+Y7sj51VsGVlZhAbA64XuglgwtTdK4jBjLOrnAJrAn4Y
13M6RbWQWqWnCQgy6OucSy4XGO1khV439/Ho7L+mWdB9bPNah7cZk5bhFLxV+kYO
gRMxfdflrcSlWIM4DbJKd4GPfS7gU5EARCVvDAGkNkB/iGcwTzvkvycxzZYW141v
uagWVM1bbjmdAYQlGM4f6jPi/g1MJXRy4ZWh/AQKVB2pH6ZFSIQVsMWKi+kKuxi+
ahuXw2oyHKAs3slsu4hEGnVipghDGuTRJIASjPVEa3LKmqCEQgHBYoNY6LcHxugo
fsqjaOlkuD/FxkCNQIjvR05e+SW8TKdFWGQgyVHw5uA92spoWEPok4S79TlJYUss
6lTL4W7nRhdMAkYKj1yBZarjDegl4ggNku9+9NitBLsRXY7sy7hl6VlrsEshnH+D
HNiq/lII7v2YIgGp+LKMUKCBi9SpeOFQjIFzZw4h0c0NwNy0KT1GT6gEahe6eCzt
nZUu21VIexvjmTI1aVT80nWS8eRbrkNGkAZrA3eJlXUaQv5xs4YLm2ZDvSyOEqUB
2BP6AOx/G4HVe8ss4BmKTUliydU3+37fnA8ltAOXOFMXmr7JH04wyBIpyKpvbGDG
k9FVoA52ieoqaXQBN6re0RL/Z+7sVKAtAThHSY9JxEut2liGPvgmZnkyCzQL+pj2
2i0WP9lg5V5SwnlMfI4zxvr23EPPmvfMmGpXvZRlZC/B8IBlpe+5++n6GpRA5Srz
/jh0ZkMxashVCbUjvo8nxDPPnbG4MuRGMViWGDBEtO/EvDMi9oN+axpHKWHJFUSH
1GW6OqmVwfgGXhwfN8kZM77ATENjeHERrmcfq/AwAtCHjdTADxHXARRwy6HWniFH
DBF78Bf7efc3zqHKQxUbDg9OzEEB0INUGqO+NPexOM3ChWHlt6H6YmHhCciXo4fc
0VFWRZxxZauQ+/UGdoBQJ8T7ZbojvTusD6iJsayp5iiDwuUFLwb5HqI25yJwttrj
nD5Cxf7TUkqCJ+aznAhF9cR4BY3jyKVMMcTg5+MrHcuZpJ6u3aYqgawuepSNNXb8
hL5TXYOXRP0tsrm8QbdlBODcdOOttGd2Ouq/n81EMsqVPF7O9d+pjmsVJ8874x1q
KRI2PVvCZXaP3qtQ2KLETLHU90w6AHS1jCfe4xaKa8I9T8YtvRpqODprAMKz57Xl
Tho/BJOA9YRnkXoLLqXD9GO9jBiFVaPW1DcT8I/KOG3kqe56fMS6OX1m6fjCt4bx
1N16wS1wPAwYRlTTvqKW6s7u4DPkaICWtxPAxKXVHtcd50L8r/ERrth5U+gTW9ov
ypB/LdgP+j6CjMOr76EjXYKtx2A/Ity+9KNWFEyt3yiC0Nf3ymXXKSfrHhLT8QVe
t/VqwHD+8lt3LyTyHLAqstXT/0hKlMMbsk59aPEpZk77ZTDJny7HiGwr24dGwULl
LmFpJyCfJOxI4TGiqEqHWt45FB+/r0do7AtdN51JyGQX7Ic8kHudI+mAll6fSChP
LrcGHUc4dkXuRJSq0PiOq6c1HUC+g6LGawseBX/ErJSe+mzg0ktHnyFmZconYA8b
MtuZQjqdZqmoGyIB0anvpoj6fbSA1mOroAF2ZDu15eyAKnqiR86FPi42hkr9UlJi
hargHOukf+XAuZ1knbYdelY6wb5mebvWx+5qd3SDCFqrZ16gN5hwzznPBiM82u7g
PmJsvVUlGyVpWltHFOYSYD5omTe6E5UT1CNPBg6x+tqnYNSddREjylP0LNRBHhak
6N8LlOqQMtBXQHdIDlJL7aljranMeYD0cX5u78Z5mVJDBkBfyvrilThHsMdhbRFw
gNqdyZ6wJizAlPRLopeLD7AYEn1/9S62vBHGm+DRZILJ671hm1DZmtrvWDXH0gHo
wI8YDQtT+mzXJ/hKWnDKKyfy9p871xJhOdIJ0GJhdXTE3RG/5k61LU+AIZbh1B32
NvcnaS0mC6PoWZ/MjmSZjRVR9zKT3vd83HKwi5bvFsz9LxedhCNbb5f7s7T7qKZz
4jjxHfBzrrxcUEe/3W3EJIZHfo/P8ytoBE2fpCfqKaOq8A7s6yNrIdjlAR5jSlD1
ygYI3non3Q3WKrUL/PGrsLaDdmMqUZT9ftVmD4Iu/igtJM10G7GqTDSqa5VSkGfo
nH/ydUcyeNAaF7A1F71lo9VIl2QTHc8c8a+f6Y7Mf4rdkecVXNQnlYOr2BYwP6C8
vqF2xar79DKMF6RQ68A5yFcktD5HXWItNMyFIyqNnJ18+B8pKFr7Zhf+9D/cnVwn
LQ0uadrDIrvLj1OYEL6RZKAw74u5X99/h/zNUlZFcLGdhrUrWi+wIkF0Nx9epGxL
WTuEglgmjKfEC1h9FZpLQtU3D3GI5SvZbHupoNlMDWTKGUCwk0XPMaGTQVFCuHEh
+q28P0f25SRn6FpCL7vZDYscxIKIMTTNS5ry5zKjZcsNBO7YziVtFEiPxV3d9p90
wYFLDM++mVYcidgawIuTTIPjCAj0V1Sykf5um5d18+jjdE9+YM6GF8gHqNnLYWjo
sxPolPyWJI/XYhBX2vmn/RSlmBnWAYNFt2jFZgBIf0UPWDfuzSIxp15mqJnwy7yY
8qoQTU5XMqid+mdK/QGqN8bEB1gwuuPmorO2G06D9eVlBSL+FO14W6H2u5dqwZXG
qF6SKfO8SXSFKpgHdNts1Ody9VPDDtJ1J4S1FCT4PDb+RuXswI50XzLN9frmrZ/z
7wJcu1rjpZA/cvEGrY/Z7YiFi+3rh385wpIeko2gQLEvWo6lYNZrlTEIAQlHeo2O
VxjLfqwtraj6pN3sPsmgPhTI0KPK4g9YRN8yR9Kjb+0nS4EzxRqV/0hDHX/6BkFS
h4GoF+G/0aPNCvgQ5f7hNvLrfI+uXhiMmDykOQ/gj0+8MElgPKzASqI4GX2xUgcL
9Xx8NqI+48yNqNNo90gy6sjISnkUZi8hxb6/SNQo1gEaociB6jXMTI1Y6XNX7nIf
najcpRkEhOVTakKmLDcyNxAk87j9Vu6UEx83GImXUj4LQ1cPoK/8mbuDCjG8FKy2
c2H5Mi1z+/XgnRqUiFtuTRO3c17+K2qAggBEw/VbSKShAOdJVAvcxGOCJAgYio3G
dO8XwtgBBD2NCORrUP6eRIAQ1U6PpKw8VKWVeqf4Qq9kOFHcuPneAn4G6e5kM9cM
qIOCwNgMF7Tt8CyU2VW+ms2uk4o8NSoAt4fFieZVcEO4Vpz/34tYpvj2P76no8aB
+FpSeLYz4BudePCQjeYRb5qfQ4y1/DuAUkv//dz9d9ARswGvJQul5J2+QqA9nveM
qnUyMzMYgWVFNkO4eqOGZuCEjiEZSOxtJwIE3F+lm3QsDsu+6d53zimVMlK2G15m
R/BQhOG2Q5+WIzsZNOPfUiLh3isHv0hlmB+znl8aUSvGq2nCAlmZWSx3jcRemEgF
xO2u/2qFJ6DimG2Cg8ymsGKJQ5Oty+MiIW2zh9Z2hNt90YzTmmRE0SqyowpT9RNh
cTd8MVfEkDbM84ueCNZxl/P4CBBMHgE6oLZFfpnlFVBnGxVr5WrljlftpSRRpWp7
BQovdCkagjRIJzmOTCrrhh0pEgG/MCMMZLgpOSVES7KleyC0fwYSjfQF5u7uEwYs
YkABvI6u5S6gBRnE2k1hGmhr8/Zeiqfwa/id1ps2bW3mhGA3pBgiGkMMzBjkrz1b
kya5QordYWnuR9+Xvfak74NDs08Pp5Tv691NhlN2i++m5xOuUJRY3MnERpVPQj7Z
liyCHba6yahwEhMou1gddyv3alnhpJ78EFcwBihzWUCixQ1SEgvgKG3+JIc8ocnF
yj8SA9JNHGYCDNaiNgCLygaTrq9Q0gXVPAhJe8hoVDDaAvs4RgqbOQfLptiGGwIS
XqpiZ5C5g7dUDkDHtcFnSpflACPLPLqrHfeDo+PLlT0a31lLapq5X0PROShkeUMB
5mDSOF7kZQv5/+n7sYof8hpciJ/+ScSpZqyZbY8H5dUAp55fIXLh0n79YzVe1Jz9
qe4eV6OoxYT5f12SGbPR1rk8V4cBooqXRBP808wVhZqZNzmgiwR0jI3YyuXpQ4iJ
UbUujm20Bz2qsQffyCZ0pXGLFkcP7ubxkZhA6NHUhdyDRo74kqXxDimAwOA8Jl4a
PyFEgsEPQe8EBxatEgdYo03h5/EwVzy4mFlO0OWIeSDFvKdVtcKkyWErJkLq8ULd
qrPEK0DSECnGq1cZiO6Uxf5Wqj99n16waqxVmaHIs7kRFOM537VTWLAtUnM96P1n
+Nyw4m3izF9ZR3duww8JzJkxZSAttZiBDSwd3zEozDQtbWnPPXqfiVEGGgueMxpI
vBgOHxZp0QebK5KXOKZ53p40cFypBjRqUWiutGltyXd4H9I4jYMTPyKTM5wO35Sk
7Moq3iwxsdOSF+NlQt64Dt0DakynnfHkk38ZMMwm7TfrCHCHY63ZfXw0zDLbXS1x
9FpqtRcM+MRfR7ZP6Q51uB7TEhmhtX07p6QjxKRBuMaSjaUzi+TniYHHQNtoLNm9
exKIvAkEnQkxolZJqf0LtRTgo7joyEVhxjQP+0RqUzI5QMRStWtmNwLTkmmIPFFu
OcDjaOAreMKD8PInPSLTP312k3OvUMp3My2G07TRgMQNtC+IDCWpe4AkiYXbp1JA
kT9hzih3wMAovkNnYzjIR8gvsMyXmub5afRBz2dUxbiCURLVr6FeWMcolb0DXAtA
SkEKiOHcXfB5s9xYGGpWLmxabWJLRIamSLcdZguViSWsQwxd8bAsoa0ZNuNmcGFR
h3WoH+H93QgYscNXhwbB5HFiXSiMt9cb7YziqVD2BCY9Rw9MFwYyRuASoGzZQdbf
nYOGUKNZHFVQ9WUKWTgE2xsSqroGACA2mezkUQ2l/a0VPHJLMvxj4Fe3gAsl2JDD
QZYV9fX7hVAdivFrY6hP1UFvddLB7sLBQS9f1BYeT4i0aZCRAVdkwOlYAFK6jChF
qmb7YNP8FlfmzGpwzD6M8pp+B9txcxv0TbQ5vIah0uv8hG6xQz//mHmgCc4zN3P6
3JNLq4Yxyx7abE1G+dTIJPKZ9OqFIOAaW4pGgH6UyY1EgFxqfxBSek/GHf3cOUsw
eu012P4XuMUpBBjt4y4P21DEonKEjJPxyMBUVMICv0icQqyrD7kFQYW7tfMeCbGH
9fjfNOKNRbf2RJLU8EcDOPWTasouwhRAS8GjBLIPeMBeyUGmHRNYAeYNC4HpiZHy
85N6TP2ldvW38K3n2UrUWRBrUXrSzUcuKidb+LhoH+ZS1DpamSrABR2Z764rHhYd
a3caDCXJOBqMgTi7ErQFFF6T/RqcjxhUFf9OfVcaAcdVG5hEF9jkvONEtFG2t9Yb
b+dDDm1l78x6ZYNngeXAE11g2ALwbJS1Qe6mNTLV+Qhi37fm2KT9aE7eXsIsTXzn
7WGy9byH2LbGUd3AjkJDwhgU6si+neGSZDt7hSVAy9Ts7rTaM9tCYIx6vQq6Veiq
uXtBn07hH7QM5d/oImLNrJGtiUNSL4GzvJln+njVPpeX/aa8n4S6071bfkkDD7G+
cABw+mjYXHdai2Ua0Gf+FJZjfO3h+SzMWBNYBkWMV4QNDOE7k92k6rDokybjjguK
Kx2RUk/UVvYvREY/LMGqPqPENaStDMG/JukfTbhQglLDZaIIe+NDEljQ1qhBCh+9
pbjecfIM/+K4Jo0vgePnyWTvxPmJXFNtA6Bc0D+T1JE4W0ESQR/2GZS+HpFXpVbp
qpdYv7BT7tsu0uoEwG4igSLY1RJREKU4ZYLjSzna75pPGS6w9bVkV9vGgggS1NpB
8hiBxvQTfnS5X+1xf+yjcjiTjt00yZBaFQkcbsEmV9SC03ddpk0Nt6x/HP1kkWGl
UhV0BbtW6HS4kHzbbpRP/tssgCRVDXF4nEwLh2kZE6100oQ5txSKjaB3vCX3YWdb
nzgZi2EYxL4w8M1ea373GZgoueM+MQxuNKJYKTrog11zzq0fOPNGRAslthLQM1u8
GUj8BbiRejfx3weYbkWRYphktFPYEnD4vlSszY3SDEPA+5xA2MUaWbU39a6BZTXi
GnrSzcWPm/OzM2Hbea6/Nvg4luscxR3MnXTkU6xQ93fF8HAfr+zyhNVxSn7u9P4n
OKT0U9kBW/eeg4tQcfcN8U+pdikDdqdV4WRFCisfgbLCJyReAfxg9Lv6Ekc431vq
vArInndUzLl1VeTT+k+y1tSeaPWXVhzJhYz1OQ/LzIS3jdCh4roPwNCDJV5YbtuS
PC+p8f+y83b4LvrgM6jbILjFit/OTbiG6DUqwkqpSpw1dGwLmxROP2TXIywieV+e
CcM9ejh+IGX7yGZXyN9KPM+0lf81aYQNGG8j1/Tdz9bSDE3tGHrwJycapkS0gsZF
V2JApWxLhF0Nt7x2JmQNwPw+h6oDIf5pRdkUr/sh4aMSbPGuR84DOV0N6OnBDB7U
gwBbq3WyZTROSByPk9qiQ67Zg7I6b55LtAF8rJ4hHn1kqTbuyWEgws61ajSyj6Ug
xIU0kEA35LaLpJOPnAZLfITKYsunQFHbPx6mOq3py8amPGBHzata8/qUmPOxrb04
BU3AiSYc5UmcTGTerCgm9Lf3AB8CMWfXMi7Kek9DdXhp0ag22FQASfbnAPvrpF6K
MndFI3OKKHLdyrNtC82ZiFSfPrWz0lHjhiD6CNKP/J7+y/OHzj4JT1W5ejJwkJxQ
fEYWM0nnlkGfp3jJsavabPICYm5onVi+DcsDlhzBhde+6AuUiN7ItzsMzUItUrng
pXi+S7mFUNnMHPQ13EY3Lid8+M1xN17wD1h9+l6focJXTtD+iBi8XqgEUMuexRkr
sGXCKmvz25hNgYmt+BZFnYd4m0bXEZ2844Nz6m9ktXbwkXvQ+9ukvf2gCz58X6EC
n3OE+JeKQrrCNBg4p399t7Eay7jpoMW1Ol0UiGg5FU2eZXkXNbXB3QOmtGoFPPfA
/rehR8jUcG91LicrTtRLXaFIJ36glDtsHNRzdWbbPQakUKmouqWglPus9LeA3mtt
FicHLBr/Qwxiqw8fObSjuUeThKpTKbCbOQicyPZQkfqMoR4HfVOHBVu6Qo/6yufF
FBlOqdId3hHIPJKarptYrpmRY/kZGAY5d0E3DjpoX2GAa+KAwQ6/z0kQIalSQgQd
haGWelQS5QsD8PLYhENqgqETF3nqBwVsggd1ujH9UszI17NW1Jd1Qhn3LrP+uvo4
iTaXsPxLZBEV0o4DqfnATq0qkBGGVb12P/4gX9nJrHT8VHcJ6gCv83T2TT53PmvC
MJ4x5uTRjBRi97Han42osMknFLgr7DgRJDLZoc2P+Uf24skyp4oWOmG1n5eYtGcF
j4S/3F3+tu5XzO82LpLKDpN8aJJzaBQW1mT1OpISEck9Onabe2kKaMBDPdZgnQL6
hEq6XGKRMdb29/XxgOIP8urdsjRe1CQUTTbtbrJx265ZlZRqrsArOtO5I6DI2r9o
hEdyI1bLMZabGffJq4eJ5mSkx4C+omEZkDUOvl4V8uflSA1NSvJWkEWGOdXIJchS
IEIxEwwn1RuVX0vaFU18vsOjB6TGx2HFNKG/uLkMIyXirEyqnCHiOIgo9c5XnTK6
tcWfz9J9MgBRAOY0riK7CmhDAoiF9yxnkMi+ILuxMylbmsKimtW0YJcEFq5a7KW+
M/reTuzpFQj7rk3s7AsT/3AlNQI3ZAPEOBP5AhjOeb5qGEUUadN5AvFWQ2qWsBcq
WuVRIe7c14265fn4Z67R5//nUWI8co7cQREEuIlD9mb+BzxbEO/uiDATMsCmoJtD
A60A7eZvM0xqdQ1Uyju9WxqtXzbsOzgD3ZGq0mrbBBQ9WXy9yV5VgcnW6f5lHOaL
D3zP/DUBJsa73jVR6pizfo/k01xejJ819p+DM2Q6Ng4qvqj9ufm8eNONE0OYLHCr
qbsp4LFMMGunmqZXacHsudzp25oyhJnc+eMd0lzoFVgg9VoRVRiOxekr1rs21fJi
Qs5rRde9lgMfITA+lCPFonIMrgMurPgWYuZr4KFuguRwptyParCat7nC9ZxVqyUP
fbPFb+ObKDNQMPVRYvcJwXR4jbJDEEm/xM6pkj3a5muW+yjcGm1YjYnsjl6ubg/H
pxwcJvVkFdQrEUGyaJL+YhHyDrEhH2kj/r8ot1MgUm6pnmYnWbUPz+Let/i5StSn
EN0lCjpF2PgUwEWginwoyWWfEvjma+DTCbZBL3rCl5UA14mjR/0zxCV+1cQCoMtt
TkgE/71yqdsGdL3oQgTylCh3oS6keUMkWfngevk3z3MmNgNywtEEf1hLdejy2PPr
akc41X9BoD5YtShqw2bxNjAGHcXxqbhz4AcvWbY89z8fDFxgr1Fn+vy+z5onxcKR
crhPFHhIAhMD4ketp2gFwpp1rQeuT78Dmvp5elBc80PlolLpcR8UqavFnxA1oWa6
sG/dIGHxgDtLtpnu5EksKr4OLMb+8Novo1j39e++K6h47KjvdqBuWBlUZGFQ/TTm
AXXLahZzSa66l4blgUjIqmzMv3DOCsPMOfyEVDHSkmPXHEhqxR2AHXhEXtMlOEnz
6CH821yOUklABxLPwetTO1GJmrjHui/3ox7eqHi9OUtrKty+xkgYIjSaTN3p+L9r
q+jqjI/JAhxeFmzAAG1udBJ5bxxLv5GzsAMD6OBLNQj1krfcu4nLiWJvnmUqQ68j
S8QtnKc+r3cc8V2pNeYt40poF/fVlsfBt2UjgZ4rY1yjlVgoRn0ZpqDfE5fuoak0
T/JBfiYUO2ZLG9qTI6Hi9ABtztNTlZgNOyZWI6gCXN5CgLGuxhh04wyuuXgEx/8P
ECP9bdB8yzjpSNoJHtkfN5jhQoAd/YhAY/1T1MSkOeAg2Ry6SDr+WQuhb/UtQBex
2NOnRRigx9Gp8H6aog79a3ilMI1iANXloFYHMJHadznROzmVHomCEulIQHwuknWL
dZI2SUn9G+yoQ274bSaDZl/XKQz30h5C0boZqkzrzrIVwuwh1OwEHX0wkgyiwYd5
ELen9j9v0Cv2cSaUrZgpvDRo86og34Cn573AU5dkAvy6TznBGYQE8jVrxRjQY7FK
TJdX6ekFCXs0Z1xA67tNhWFLqgHIkfFWPICF9UxSNW4q+/Di+m8uPdHSfVRqnO5B
X/jlpcvY1TYA1KLXTQmNsO1QnSSlRe0ujCpNIG/WefBighm5HTwSGVODkbq9adwr
GyS5YNM4dq2UspJkLtQ4G5WRlGk3Dgyj7Cq8nmmoEOWkjHOGM1Lmtt5e2tm2v2uO
Pz4uE58OshBYf4Xcsfwui7JMe2tNhco5K7TNo2RuQVeNcFQ6MBRImW62HFnQ5WaA
aqellSUbk+e4VPGSYdyVq5e8a7j4Ch1DBvNsviv8h8egsy4vcdbyiAU7dIRFEcOg
IzEXNt+aQHrl8RQcURLwY43OH/wqRFYwkoMhKD327AbNYKVIQG2AOq+7oL73lFFJ
SghISgbARj8EgSrtAJNSYb/Tlp5vHCeOo+qdNW4F8dsutJ3yzWKJVobqzRZGPrpp
ps4kExsLIMuZPzWnH4PXHaaED/famywwMdHZkSLWtz6eaeLRhTfCzxNZR5Z6rS3l
ddLWU+toDpaC5Cqdb0nXatkHFjiOJO2dYSzxLFEG4P3a7WfGIYEP+2/fTn3nIOeC
iCLYDPsfTMcVIWcG7Ppp5vHF0D0mZP2uNXBlCG7IiEJO/Hbpe0lwRtYqQt7m5RrH
E3fDWlodnFrPDZIBDo3XRE/TzgouYVRMticAU7LRZAdxFvOz/rJQm6mAq5gz2I19
90z3o7mJVtnebzluvcyztvFnJ0eWI/qvlNim43Y5PlCqx2JaWgcQluGwnWaSSUZY
8TA0plJaY9DIN4RUaJ2Osa0FnQSBVKrU17Ca6XcntLkdycIQH3pLYJGECV1tHgXv
v+9VWG+Ld7+J80C/rwiUhnOfeTEgTPwHzCgV4mrfl+1vgb9OYQVdJqyTK8jpqrK7
5EiSQrXiAWwrYBZHPxXuRBYmB7DskejgfhV4DptfPsIHp9FN5f10redYHl0pPBzY
ID28z13cb/bmvm8RuECR7xsHD8F8SV/42Rg8Nx7eQEPzONpSjxR50imSmY3U2DCD
fhDetuWr22AGSfInGagnHuaWCaxnXZixwb5T7xzbLFwalt4sNGdzl9DzzqyxNPKE
Wzjwbpce6LL1gX4A+sXFy0dxGI8mSP5kfqNufi9OrFRffPumgot1VyzhEYenrUZF
zrv2rO8zzY5/wEY/IoZnFsNUI0VKCWFo1y4D+I28bRYXHhVnqUMM0xohNXaoltXr
qiVyKKz7r5dNvPtOsNJxL0bjOtdJ3TDuf8mkOL6BLiQ80fjoQHrLonbYllOB3pXb
gEqpnUpPquLE+NghifEBFhqY/lW5mXbSdq5IymuJ8sLI9FtMSVTxC2dZ+3dMeEn6
Qvi7KrCOd59phjzXBAg3kEupGHROJd8MsgDGcJ/xgs97y7ImgdSbzUbVLCgU2+q8
qe5suAsf/01yqZV48dAfCy3CxMocKgPsZ9Y4c9NcTShHAuKIgZrXCrNsGF8y89Oj
aaV1j6vONJjb6yXrN+VnBV6vIPXmk4pxfSfDcHM9yGzHt8osx+CxjcMu09pBElu0
OW+79eUQ6U/+Dof6I/Su/pH3hKYsmwlELDvGO6XIjrDI91NcQxeGqGNCazfB1BZ3
9kgW26G+7hVTcS7g1bUJSSW+Ks6JsJHt/CkvGkfbAg7XlT1OEYcdgKeNKd5j3j6h
t8dvLk9C8M2/CaQo+e1Wrtdb00N0xIwhXjNTetnG36SnfWaeyWq/A7nonHOK5NHl
RgzfP2dB3Wez2JL2PxlX+gvRqJpYm8xLNP8NxFQlqEQUIMPAmE3O4lIEjtrZEAnP
84F226bPl4qkJWZd06R4idu35K5KPoXhfkHLbgfheaB2dHsb0J3raBzmrOERARHA
T+x245eR9+f+SgShSy2fT2giAPZFxDX3aqnOYqUPuQs9YvQ/h2+98DyNI18a9Yo/
c+G6UeHHetHZToSBBJ0KRp65qeqSy56qxT6840Zk6IQqzG2c5OG/DEL1a/fE3KON
YqJbuqTMd+sfMapXyBe+RvR2SbY8V7gWm656Mq56/yCYalr9I5gC71meli4Y1wk9
lE9sNdKYVHrHgeQ+wlm9we9hCmCc/0cf93Ob1hCB0sbDml2Lg+unIkHOrZta9HE9
6MyrA4icihxmTCpdWQVrvTHF4wLCZ6+Lug8PdxB0425dqG9ZKuAXz5q66pTCBk7K
uoCL/6MC7lO9IVtOCFw/KFXO+krZ6nTFBtCzNLWWkYmxY4FZ4FX/jcl0hfNEnKJm
IKHXQUpaD01kolKDv7C7UenaMXxQ1cqQ7Rm03BR96flQvd8R675NFU0ux/c0FaVS
EvrREVS+vbGEycw7KSCUKl9DUHYO8ixdyM6XQfqWT8QxQxYGObRL6D8jOtsgjU5s
Ub8/XhP2HK95qqIGAmYi4qCxDVHFpFDTRVWcVqn87VCP55v/XFGrElP1oS1DOZEm
15S5QHZgZ0kBOyFTnnrJhawzTDHvYaZ0CQIO9sywStfxEiiY88jTyP3KaI3zTvZg
iyOc5YMiXzTaVtjlVORBVZCZ/+IY0nbQSgb0SZdRB2gQIsuYZ5KTwPwdOkXkh5tK
1WFlFqm+4DLk6cqQ/JoQ02OfeRx6czqn1BqpzY714d/SCh0Vsl4Bu7IQ4mZhuj9w
KEpj8HDhxGVDlJ2IOofwKY8HybZeorsk3SQdbsQcZik0YTyBdAEOql9HwFHgLA/i
Q/fvWGyIB8doNeG4qrERImFtqa0QEsj7mRlTHEmb01gx+wGynjePag0ZY1mhAOoN
IznBkH3tZMJ7Dpx31y3vBI6cZ/Cr1Lp2nTtSxWV7X6fDT7qeW9zBqJKBnOJ0qzRa
18o9ZW+fS+FhmgG2KBMLlnW8e/cdGElSAY8dEQlg9k46gep0HU93H9htp3gjKeUM
ItkE/eUNbKgBNZr1t36Xu06FT5r/QQ2Hb03ah8hjahCNEG0dr0nBYEBXnjwrIkPN
YJx1IvaJQDEMvg8dUx9URywL5DEFcuXBxHfkPNQRmntaUfMLlnwseb1tS8meYvcw
/zvmTtJLuKdqA4YBgCPoY99XplY22XA4560J+DbNu5BTbKvhQuqRibs5cpNFnwcU
MG0Spjs1y+nohtbro4c4g/WwnNl2OMrkAUXVA/ia0xkw12YRY5q1pgqJWBbMkG03
9ToEtbfjunBVnpdIq647zF4+dwZpgWEzEnKrxlBXZuO5aFCnqB7K+L5eWtDD7KPU
p3i4osFcM0kIwgxGLvzhMCv4EdPKq3x8S6+2x6sB57MEt2/FveWMsPQuX0eIpJm3
W+2DMwfOwub0RrafNCc5Z+miEgUNepSdrs1SOVau+QvpkDK3ad+rC/vSVWu99V9z
XX3wFuLSdPgVT7wsx4Fa6xBWctAOqug+vjDp7l5l/F604x2XsYPFtLYyG4cJNb4M
upRGVx5GF2oKrwdwu8mAh8pmeSIxUocrsF3Ec1LhwiuuKyNKsEfO6Lc2kkE3IrG0
TN/c6xhSgigsA7H/vynDcv7edghOJL67w3dzP5W236P76CzEgxf3sTiSE6QvqPbD
hLuhuyo2MNHB6I6CYF+8nOx3lO4NQXzV2BQopDwshzhLqgURRdniN7xj/YRDm/3T
gwWgA1Lv/3wEFc9+uyWbkis9rGnZtQQFDidhLDKqhN2UT/JN9eMC6OC5A10j2b2n
2njyWnsAkLqUc+cnAAVVidUMsaN4wH1QF1yYMtzqNBevBOQ9kNwSYFnYz9fbr81G
C5iWO1clE0gYrne7rhM97ya6wY3jUD3DXuidwc9oCyIgJ21nP89qUoRo7XEFq+fH
Z/0499Z1dmPbWTCpMY2hfwk2+GeRp6s4Z9hZqfKro5/WQs58rQyopS/lq+KW458R
YZ4g0Qh51XYg8VYTaTk4oLxTGCa/GQWrJ1fEJCGuTlRzgMDHwxK21WpYpBOl9T5N
awaZamji8UoZ/cuykFShW96Yhftw5QsHldMqCeIuPYa5aywbJxK4Hx2t9l1o4xNY
286intfrY2ZH2eTisX4jFtsZp2tcUJClt7T1RVEQS1mhrVN8D/5JwLK7yA+jxs9g
PwXPnESmxd5YMWgU2lI6um4sQUSTX0ZxFY00gP9X2oI2w70K7XtKGnzbbEpnNzur
Gf4l/ooWFvwkjgOH/eN4n+ORmI+rX6lCTwPOkgOOI00P6UWq5Wa5JD7e2YTazpxl
Bj0q9YYflnj0cArowEngkZivMGAKfbL1WI2/cvl6KzivRGAg7IZpLS8okfuDye6W
aETNZ0jkcbfwB2SDco3FHjDOLL9kw1zGFJBnsg2bU0YGFw90NKWKeXms6JX/gp0+
OhqX9qiybLUerlGk66Q7QKJtgHAW57hTUCy4ckHkJO1F9pNxf56fQOn14ANaHMf/
xNt3ygg7gnVxKLbBa8DozUS3Fw6xtjnq+/xkbD7XVBivC3F+jhxrL+h2CmbtG9MO
of+7F8lkAiTfIXjJx7wyF1Yqt9dC4gCoYkLp9o2hVp+TmAiTxo5bkPNpMnu6Aetv
AT87Krv1/Xzo0Rb2dnX5dDcEtmPaL7gfkeaYxskwhEDo5WBGPSFJpkZU4B6w3q6u
JIZbsKD1Y8ilLIgC+1wNr+t/eK21p80FS0E/4d1Qsa3GIrfh9rLbG9U2fZWuovWR
kAXZlsGOQPVTbDeKuZ1UMldR/sYaD7d2c3aiGjzzm55IBfP3AJpEbjkN1zecwt7H
r0E3CuA5VS/FjFiVYsRqPN/CSSHeUZjQSSt5Q4/b2z0Zbb6SxAvKGiZZmX9vzyOm
913JHeRrX0sQUoeoYGeDvaNbjbwVA83hlrUP59I4JI+BYSURHf3Sd/gqHrsoPidm
TLMdKXB8n5rL8U0fSRh46TYI1XONWdF8nu+FMkO4ZE7u55dh5U5r5/04SsWQD4AH
g5K/BmOOfuA5QWdtZQWHi5R7ON6vBpA/EhO8hG+h+aSAKdLu/ffVPwMei4FsKHRE
vT5njx1wgW3527hyIsbDsuXIM/FQBPxmyf0LLwfrBiod80Qj78KLTla6IOPdAplx
cH9n+h3NnkNn9oawaOvZwfIkjmv3aHlk9ZJOawyFw/v9xvJK2SQS1wdHLg6JZIMw
XkSUD9RqmCBqLdislysrGVh5NGFG76xb2Z7rSPXtXaE8UaBH1SjMDXe52XKPi9Jc
55K2KZnVUstCgkN7CcL4a4gGmAOKDWcTfDehLtkNNJ/zlIvsiAlcuCEMfzArXh4S
e9k74oVi0q4KDP/FBHTI7kmVfGqAPbtkAiyj5+XAT4FAZi8Kgvy1bAECEtvwjrc/
BdWbgM/oX3mFItEKNQU6UkA+KXn7WrUpeERi1j5oU6USE9c2t3K1Hb2vhHfkQLk9
kPMv8Ou5M+kDQ5Dxhaid0QAaD8WdepZ9gM9y1wQP72aTgpq17c+mhWTizZsECw7U
M94IGvy5LMaA1yW8E5jPnnZc5dWhn7k/YI79BC3kzs4KdVrzSkJ9EvY91qzJus7h
56sShkMDHwFaHzDIavjecWkct2MeHpCud7GQ1ND1CE1o0QFCozkD90ZbjTeZ89RH
V9w58o7aWwMm34zjRTwvrAhlOr7PuvNvjvWr0IN5IYZoi9PpjLMNFO9wLHCV6hmC
Ji2rj3eWN9vO9liwuoOU7vGS0sJ7YIYs/G2MuP3Zi0AgFBjOa0yJGftJ7NFuK7I1
nYgIGzGlBO2KCWcVzq19GQevb+YUavbWKGgCu0YTUY/yAsbObwWF9i3eT6BZI/Jj
k4EHm+lU8rj8Mg9Vtxn+z1Gbql2TRcxH3zQAAkV7Fe6MpIk/sispbSU4c3a6/CL/
TqhjMgCDlCIkI3Td3eQHQaSPGYBzuYjI7LyEdMkMH6VhOAFyZLGFA7n/sYrz1xaU
ij7r8ilDieSHZY0of8XTtNh+1IiUpXZaRR5WwHt+kWdYXcGR9y5TIySA185BWIEu
etj45Yx2pK/QjNGIDB9qUYkFh0wpsSMWQ5fVhQXb8XRLfQm+N3VTEl4wSN6kQKQa
gdlzEGdP23cFq+DC3ykhaRsYrx+F8erzrxR5qrClC9RAvR5aR2OD/AhIKK9DVGbh
+YkhEefg8h2D8c96TbCvnFYXiq+JPlRcB7UAo7kTrgFigdRVE3wBmSpGK+xzsJHq
yDf5O4NA4bzsZKze0PjMdwobqZJmiHa6dh1nT6GV7bO1Tss2/vjDBpxAJ9p3VnIO
hs6BgqPM26ivmwMhK7SHXdMe0IbPcV58zciiP0PJdBlfXC6Bc2cK+U4DMIcBGDgr
2cQ5DLMQqGH8YTlCGqhxC0km90DeZT8CN6vuHAfs35RHeOhop4XIFFkqj2j+AXe5
Rl9iknGb9CHpZRv54Qve2iFKyyT2dYcqAvTmNr0dSz2TLfO3gaKd9Xy2Jx9+NWYS
aGuTIx/FBKrIMWubrN2O3XNSJaD+RUIlD7lkOz2zN81EmnPjg6Enzwhux1Gy1sRr
jHXruM1clb2ROPs6IR13rcZgUOZAKWRkqy0UDkgS3kNbJC4xMx/tK2Kx2CmAnodW
R05NTtEuGT7xfuuHIuUYT2ARA032aOgEnrknmdsY7EorUPH2OgqJjKbzPOzjknJK
OuUrcQtluP3umTWfmYUHL3o83OF1HVpRtUYCYFkqB9a2m3FOZnhdvTyPb+CMo+va
hiRZxSQeqT5Ypco7z4/P94DZRnj4FpCRZfU//ovMQiTTi8thr4+2e2ioBB6HPRUm
lX4iRSolPWHq3Rjshh/nZjB6Uqmkz3KOogcdgSMt5+uEVcv1nQd0ctzM1k43HR+P
8qcwO7dRHwWznEfXqa1AWkh0t1Jjv2M4Y7EUuPRBF+qpo5B3mzta4anJGJ2iPYLD
KYkKIJM/G/iuKfWwed/D3pI/xtr9tAX6+lCnrdzDoYXkgzb7KWBEqHXYmjYBErhL
8T1iMCnkSrts/DYBaQph1BcS+8nJLePEmdnSIITRgESWzVxksLKe/6Q+GoFbFz2O
GH2O/3ubwpn9+qkju1fO4dku5pLictiGtYio8xFjvhnrjpP736DobH0FAwx6krUh
Ejz73CanSSt9rRPpHlJU2p9OunZHYcwWXNWScwrZ6CMx8LifzsPRT0XOBZHqCeak
jwvMAtqgzKhD6BV1saVgq/xa+CC0/go0QdNIw1amrqLDUsOGTaQ33xr2dbqcqZXs
L8ejUKLpzW9bZBgrt4RWy1R8dAakGFq5UV3ekorHWMuDENLtgcY2g7CjSjicW9ru
+vm7qjyApPGL1R9v3I8s8AbtmxbRKIfSFKualFIlt9n1/eAa+DkZ70gcE6aNJpM1
zAajE1iRA/gmHk5MTP+uyJZx1vGzpEYnQ2kRPwRSoal2/OcP6og9ch8tSX+1hpuu
KsxChAKjQvpusDnqHeO2liPHDLzXRQyJ7ivuFAWCJpx5DuSgX7aGAvKVia/1p6y3
ltYs6ePBJN5avDSQqt7vnCsUL7TzC2gWfxkhIhHqdkiey6/LO4Cx4Rsl4LSbJvYz
vEmLHYSqOK6v2MPnJiz/b1XLbSivYql0nEjrpchhhbhGT/Rx8E1kI+HGkp0Dftoy
YpiI5YiSx9Ki+sZI67vFzFRPXWZbH8l/5gE2q7RMqSoTtwqSIJN+0gXeaAy03kPY
cbawKNxoTeqvwHL/1lVbdV6egwSHsOr8SbW2i9FRurMGkkedC6DV6OsLctqNiPAu
or5qBMq1nx1eFyfen4ERVrHNkZ52ZiM6sNW10JCuNhCR19eIQkHhWHIVmwJ04K/z
sYeixb+PSlAMTguSa1h7g5u5LRPfGfYdOGGI4cNIkxl/ygmq/RLfvnIg/n4lnK69
px6JeO6IFmNZcWFqN2VRyvxF7mjXt/zXDcZT/dD9SX1B+fujAZg7aj55rNBe4+qx
KHNW6tii4v8P+H6LqAoOEHdy1Q8uO22c92NJyIDjR3M0zXLbVOPqLOBAvgPKp1fe
7NgsRKOGCkRydeGy7Y0A8wqLga3GUEcfBiKgYH2PxFXr/3ZLALzQqIZe0JjpT7JS
01gq0wv4AByDlKJ9wksvu//luDsr64zYWqTdSr4zAAeA6ODIhyxPsR5P+oYreQtu
wxSV+9qbFSVy1qCwkpYvdGg/XivFNUDzTaY6nSq7RlFCxZ/6oiEajKljiFFvCRH6
Cu/ATgQwzYr6742+57JA2xeo9nB/w521nZj7ejMR6bGK+0ocjoifh2Tb8ER/4yKB
rMgXHgsOXRdkPBo/Cy+Dp0MRI5tLiKrMBh7+JxQIq4L4fs+47AAs2ZXbAaQa0de3
HO4D0vMVgArE+gu4iMqrO53U8/RnD+IBZS0hIDo86f+ftnFAOT/n0dYh7p1eCye6
7qrLPZ7bOVu9io8/U7ZjGvN1KnYk80n2qgq8nnt96vaVysr3d/MxdRoeCGGg9/cx
UwuMEcTfLWwJa0JVpP0tbjPFpUagGBDquJcxZAHCZBBhPUbElWa8l6f9718DwG+o
tO4yK5OzTe4pxrqrglHANr/15LiGMO63dCnLpidA+zhR/AAoEskK6csGuX03+Kdz
HliMxdbWbrzty6KAhFE1Ag48lDAYr3/dlPh+3yXWGWD9a/nsl8B78ZtdO0zjrmb6
yFUlQhU7m4EPwdhGwDt9aCF9sg4dbTtJSZQWu2br/DKY9tu1R6up9sVf4qyoCtkA
/BP5qu9XxgMOYJsqmS8DHUtD2iRNPKSKWKk0UXtGAulopsZ1AnGzhw66ww8FE+8M
YKSZA2BE3wf2iTxOuIJnEUEZh6oUV799rqnGstH1wbXeCz9pDNw5qQfDLhXx3CKg
eslwbxjj3wOfIY6qJHRy7RSdJHohbdjCI1Qkcfmww4jY7u7+lR6lA2kIjxYvfsUr
3DDxqMEHNNv48E8DsoGvVql3QdK2Z5nnSUYFTvQ6i3GQzIwHd2eUeN3rKsbJJCeB
ncB9bT4CLX+9uEFZQM+PnKj4MRv2pPxZ0dBbY1uAxuKrddXahaYQJZ8s/fxX0qnU
U/Zu4M58vDiIoAfNGKTqKJR+Dt2dJb/bsuGrpNmFn+Fjw4nTgqq/LZFbpJheSQfv
IoC+efcjJp08/a1GQbXMkPgn9d2p4Vs99YhVWl+cM7PpM5eg9x3glwOJNSLjIrn3
7h9gM8ar5hTx/EY9QvcUFT5qGGJiESpw/IVHT98GXvKCVmonLZ9gnY0klVRFkUg6
I0wPb0DzZrbOS79Md3P4fMyzvyLv2VlAemq/bRk3ir2ExflPIECunnP6wB9FLg81
Flf1L3/KGkEBgCyNGyLWOQKNxhWZLVJeJ0TpgR1cDc1KThoAKbdR0q1DdLmbFEQq
tLycefExyYTve7w2sHyY8T4h96dcH1TXNbAWHFgr7iP/i7NFRKfr1LT03aUkS2RY
GvjjVMlJjiqw3KczkB9iiRPJC7R7j3SdIYkpt9QGEPjzUGQdrZYCrqmcEOr8r1jK
kEXkcSJjXGYlVkgmbg/WHXECUaEIzMIpVY/TMjRevCmYiEUgOCk+4JffTWG916kk
DiARxuSuqLq6yopaZ6y5U5jniRnPTV8FV56m9ZAzOeiv+c0NaSLXRHSR9OrVbEwc
djIoHbyQrgnpVv/GEyVdLm1NiMh78zOtbEyjjozvcV0H1sbCwwXgHdD1sdtkWCrD
9THy1WoSmDct8XhDbhZH3KLja4hozG7D1lUyEzG8N2Mb8EL49N40xgi4LZH8w4hK
5VWjBOdqJhcDvg8UZvwJJmKr89uQlsy8O1BN0eEXR+HT2grcyOusYaoOLvsJdRXt
MkGYLok6caVBrJmZ3W2/W+w80sPRcYGCoGUsyIeuzQFYcngFNxOg4bwde4GRwA7/
z6puXfXuQpAYcSOlhB3fghWjBPW4OQ2UoZ8esDEXz0Lau89F9Ds/7sBs6ZoUfKxO
sViIKZ0XagYyBygKLGgvmOvT2kCPf2kmpXxmJM8ainqdxZf3lUpWBFmiJ/5gcWbl
hb/1GlS2wn3JHHBdbR+1GwHEXE1R8Ueq6imatz0HQRC9Mw4DN2s3+wk/QS28G2f2
EvxXAbAuYESTWrgpZtSEsCFHA1jZmprHdCg7n57C5LskC9b8WajGZp5ZNqETHDJv
WgaCD4B1hlcFk/g9qFWXAYUrMQ0430qf+danFfiv2PYnENKMQt5hS0EQgja+/ixm
eTs33u95kCEsBBWJ4Kncyc/Sf0Sp7qgl7ARLJtv6PwXQ80f9ppKh/fYhbQ/bW01Q
qyj+AyQ3geUrXio21GcxRMNu0HSIPxcROwiOUVb+kudty5Yk540vI8OSubfRF1mt
OYPBZDgkmdEm548obGrwntYCbXMf9zWx6qYfoOu/6LxwKIm0ZxScKMLUaHvi1Swo
tTBksYjtGzfyXu+/IIqHjwQBbBqm3DiDciQsxSQOhcZuItwROFTmhDtZErCyI4wl
eYfkAJ9Xg8PNtktcgHgE3at2xMZPJqLA1qBiXlRkd60GWaTs6kFPTNiOJ/rmws6R
Tj4hQJdG3vd9HNCg4Gxxvcl919zAXTE60CecpQ9uqLmVM80x+nOy4MPfrEr/yZ+Z
lSQSfJQtSVlIM5BzAVxJbbYtK0zu6zk2uJCfnMXVn9BKT2cCSdn5UpWPmaZXVKgv
4S1+8ETTcc26gGYMWbz24CqULAtEKqnP25xOM0KgR/MQ/xkfzx1zHeIy/bLxmw/9
v4n3UWhLUb5BlbtevKTm4igw66n/rLkB+pTuKr2Zdqo8EjBWlw9RiP03sjrvA9kN
J29R0oPM+QXXyTwkOvSCiZSpQ58ZjgwEYe7bBfkN9st2l4PPUyCrwI3gsWfYuinH
rh3YxvjXcuNS3iWG+H4DQ29Q3jISsNEEKigxar9xx+y7J/ytaeQ4zAayLtJXN1Ja
6o8Lh03PzAr/AUPufxH0mwA8BZu5hx+KuMgfIKo+sbU2mhoFb3HdDFTkCVk0yEvO
aUqnxwOh0r1/ZT9e9cffE9RtaHwaC9mzw9ZX7uMP/UrPfsNF7xpSsjBMfFHyBbel
nRpuJMalFz18SGyphAXaBJrA5KY07QLulo+OMo1sNI4QGj0L7s5eqDv1E2Z6U1Pz
kpRGirMHKXKFi+CbnAXyAa5dltQLrjyBNEsEu9YfwhFYLqs7l6rVS/a6FPzd/4jM
9g737jRaNgXaUI13glyZjp1C7JW10PU0qQboNofv21V0XjYpIIghueYRvFJzaQDl
Zgoj/8LhTGeszsznIuisRU9WEP5GDQvxYDuGCE91KOSkFRh6u8Jwa0Cr9FGxpli9
YFMycBe54DoBRgNeeb5eXBvDE1rvsNdm1a5nhJb2/aGVXPBxT2F/8z6D09a1bM2y
TUgq5ebWO3/R9SkyaidSHh6+QpnoiPpXBb5nYGCn/+AKQgI8U883uxbFBXKGnqh1
ngpP1j9oq6OQZDIYYg80ieYD5TcDtWMxxdls2bxeiNXq4eNCHvbtuewHrU/I0S/1
ZTbUPGcndr3v4b1dT7/nyO8TKVgVgXBO/zrrKL5iov5ffl2Of4K5ShO3uUc/Tkxk
tX8HshHjy8csT497lC2siIESV2HNeSyMlUz+tLn3wvTRIoV2SYEQM0YojnSBQrgu
59ZnsxkI5JbFr2fvQKvAHGHWjJ2y4nyXHKirAma2qCyQt7XDrD4RE2SoUFN50itg
FnX/ZMGTB3IhJK9+njyqmQ24F3Lg/xhQF0v3PTPDNagzETDlMGJ7PEURzQbNwrjs
p0Qz8Z8yWacep55ScafVrFFKvav/OItlOCPfCG9BGl5IAhzbjoLywOhZk/1cvUE6
wjkkrOXXikHqbzRwM016D3p3HO8ZkxRgHwsFLxY79oB/Bd2llOOFRNIa/bQ5kSWU
GiG+MM8HmYVGx3HjrFg5h/h/RB6sTNBr3HBkpl+fYSrzeC/0wlGsb8M4jRv0qOIY
iN0VYaRnuJ6oVPn8Iuzbtvi5hE0AeNJs+GklLv5kJSFwIOlylbSmk25nfSZpjdOw
duIGevDMYcEK7GnhmZD+y6K3c2+n11d7w0/dBLyfe7aA2pBV4H49cSjbFJWXzW5t
17z2TXVOd/EGZkBowbGIRqzhDOa7chC7yJDCpDGME5t3Qgyarv3SR4o/AkRs9xCK
iCl08tcWKnuB6UuaVXbaGaD+uQniCS6DBBQe0fvZbKeWMVsyndXnxgQuTTgLbG70
W9FwHLsEi8C/nCmoxYLAlkAFWNqXL5bRJ+tk2zPVpD4oVTuDj84kVxTFWVJhpsGI
dgeC5W28SQ76P3gAlQGcZI/OCxxIPowj7gqVo9eo3jYQqfFcAtVJOnuG4SZeS5mM
0TsETx9azlCtWA0/YVXKXgm53l4rjkask31hlolTKkKSYzIYsnc0LVGA37HCmreT
NjzPlrRDpB5sIH8tC3GQ1QRkBp/5fhepNx64LiomRxzHONT/LXnDT+4aHt5kWL69
uyK09+OIXQlh+8Y6pQBXUs8qn/Lsx3PlVEmsY0vpsFwXTDXlMt4PSLyXza0ndzQy
baQTHwQpFp2DI0mdRkyAsmBKh9JoZzch9eBVlWd5DMXeTC5Sxjom5NzQJa5m8woH
7J7KScXmiPLH+3EKUOJchuZL5deElE2my6Wm6xkc5EL4XMpNsTq8oMOp+n7cO+10
pvY9/SpL/KOfsrzSDvcJ0PKFF3BgzL/H/RoThIuef0ssbwlAMWIrs/fsBjWwTff5
obaIiEcCCXpXafyQXY2j+3nxL7knMerR2aTOzc4oP3m2FgvoQd/OOUT5HB1ilrxa
DiF6CPBgMC0/3AzkPvrCOxz8VHrm4ZLjGStyx4P4WQelvGbM889T0v6jlO+b2Ha4
8PUmpa2ztSYxfa34I1Aq2xNrAVsYqZsOcEjr+U5v433Pq9X0cgldN0aqW1zakYVM
X4HWEm90nVUVtg2PVHdY+WKMw+Eevdw/AyQs6uMayc1gFYiP7QNqaUSCaXPsLd3D
0wpad45AfQuCaVRFc4LmmZssiNW5kVAhi44RQEvUFT5+RFmHHJ0YZPd6rmVVSK8V
2Yj+SrOhxYOxNGeKEID59vbZ6jWS5OdQ3VNaaO6ofSWF7i6VW89DVoVgDMTR3p6W
g31w9zxDcKxXLLohy+GUAsBzluIXnMgd/G3SSUiZo3SiC6RBRGHZ8mNhvzbMgJbe
gd3NxQcg0gYhaQ1ECiWQODm85RkFAH1Yc2p0FunyQ4O9j1KJxPGu/kvWepgzE0z8
uw0cCHA7n42yZ4Z1Esc+/WbdywzP0YOLRrn37qp+9nXeZKGLc97A7BP3ThQa8spy
hICjhqWj7guerkkKB03luxb5l75eHjW4Z77112cNwFopW5Uyrj67WBPi5cA4UDqh
UPynSJ8h8tb4aXRZpTbaamevBv4F8eTTL+o96G1Y1hN4MAtsiPZUcDl+TL3jeGEC
NNa5ixmr1IKOrdE/M1nNKX1/s3IltW/ciOp6hmR6i7uQxXOq3Ul7WxaeDCx9mZnC
N9bwBTZw5o1e8AHg2ioar8dUedUcYr/HOvmlEBPyJ42gRcIbHaqS8UibPaMvYruB
95Z6DPtUFGpcQalAW6uWMiYlQ4jJHDRqtPVMrGX46N+SrX69S3xgzHBEwh76iPx9
FI5UJe0k6qsnXCbGgnbbxe/EXMoxsLB0XktNmeu8jVAGzGxSf/YnOlODSm1FC2Pe
t8glN37j0LBUzghZHk0SDjnu+NZXyVjEuSFZrHByLKKl0CmC3oY/sS+q73iT2V2W
SVOtrQkkqSp4rNOezrmae+Um12qcH/3d7cceYCd8QKpueQIM6QQNHc6ju/u1zPM7
Y0wbWyls14uHoKa47xJeHMuVN2CeW96nvKSS12fthB33brIedk0DMfuEC0GP4guh
1hRzk3RDwFPTewTvEWlVtXs7Pbc5+Z+LO8lJdsjNwJynRRxykdyXzsmadzqUZil/
4YSL8uXEzzCwNR6/gaGsSCybAq7HgHAAhf6CKZlq3m5dsnmIJ38AmKdGO4ySNjKh
mrooooZbhSgjE9ZU22XvK4uhitW0cqrx9GdT3abaaU55Dr7ZiGTYWKJR/oNLnf4p
FU/zcXMABJP/EeEnnt8oQP2A2Q8SWp30bXj2Y9Mg83e/gNNX9Er0Bo0Mz+i2hTnD
L/MQFjGP/CbALCQ05wIGhaGQCWHJWxkiNxNTdF0uHDM52WBcoGSlq2EssoMxhIAI
yJtcaoAbNpDww+lgzi9qCr77hC57c9OQJknhye7tpJ81Kp8SmU7s1ADVp8f/IMn3
ezBAkaHj28QytA80ClkSM/cJX1VvLO8ltq1rBtdk+H/pnZqxujz7uKtaT3Em33PX
YRVZh5z+NrtPzWLGYY4nvq/UsN+0Y1zhZYdVax4e13N4NJSQ8+bRTFceoD85gFx3
SPp6UqQFox3Vo4+H+xesj8a9W5bRWq4AAfgFy+dQW59vjXYkm0+lnbbTA7ugzVDb
2O6AY4crhjTH03T31+lB1gw6IoAsadbu9Fg/SMdEd2bJKuxtomPGQaxz8asID9y/
fJI1Ukw7r7krfDzctPfeUJtg3HbtEmfgdVjf5rtxWnUE2aOkWmGjWPEqKYfIOsGI
H3hZh2tCe4FQCtaVRkRaw6MefMOQzt/+lb++Nu1zqVx5wyWgX7zZYMz1NdiP+1Ln
fU1B1sDSYnme+lcbS7LWjl1Bw8qaz36IB/iRFVM7ls9eLGbsdV04921RrnTN4fXh
1Xm3NbAUjA0DE/PN2Y2yoW2aZEIFD963ell4X5D9Ekf/g2MZ8tYiRgct5/qhxhSf
ZofNGlOnIGqvg4ZD4kk20fsDW6VliPPNs5/VwNfSI+DL/fIKeRzgNuz0QY3E5MgN
gFr8INVvUKNgolKvfc3Zp8EAQKH5FtmxyYiUW1cuoSTt+x/uFiEZ1OaHCL9W1RNt
MVJ0tAPhGgSn3tFs5lL0PIaMGSwlGtBASgmZdcHsBS0mleAluKRmlo+uiD1QaO6e
l52keGhwT8Oc4AMsr2WFz0gVqBruon9aDps+aHESwhBzfBVtxo/6aa42Fc8LGzBd
bCtibBtEvYLkSc6vAhFfMZG05CJiCdp4z8Gt35NtPnGb2zCLN9wVyNvjS/nLjtO0
BGmkT0ABwK7R3VWrUKrsaQYC2svd9TIJzqux2nCxkRbYGff0I7+3ENRr8/gdNxaT
EmOPQF0e52g0/8RyZ6dFGCfNNoeLPYwCGQJDjjQlueZJij4/djo5wMorzqjHJOo6
qEGWaVdRbOC/B3YoHNscsewuiCiJ4G9fo8xenB9U33lkiM6nyVI9011S4nilpasP
xjheDrCqbzjtFwKuBNBVYlO1drQW/AdNbbgX+3kVCZtl5rP8fTu/iWL/d90YzrVF
PmdepkiuFGAa2xp/glW2v01HkDsip+4dc1KNk53gU3PrP5odrlGX4W3WgoAJiYH4
ruV1EMC63wmW2JF/aOWtykVDR8QnrpxyYXHqKyvguh5+W5YNhjbbN8dH+rVxLozo
PIY9iQTXYaCUL50KE03HOrh36O9THbpGceLt7T6SHdekCV8hnCqjP/fy9E3eqYZd
scoFUUVGtA2WDE0GpX792kTxZXlagrbYwiOsMYT+fHURLYLGKfsg2PKO1X7jIw6w
3CsHhkbzhMKbbo3sECN5eF5jbetPc20X9FVbSPMNlPkek+3k17ANirKVrbW5nefV
LtH+GkwSjMMr12L7+ykeNlOAHVijYSa5w159lokm62Y1cm/3DHm69MVwsm0i7mJl
COu0a9Iy4Bi5H0G7nI3Eq5cvkLqQzdpd99SErM1smDMjEmsj7ji8ajIfjzPouHYb
vKs7gdmTQMcOy8M8ixVN/62yABy84GEwBXu8Exfven4LrN9fR3JBO6wvXZkl8EoE
BHbLUtWTcTtLZ0oX1lhdOvxzl1yjH5SEVFLrdwCGsAi6ZhPaizAuFk4icrUS0Rzi
vpLuWXY/xDXtQFKKu77GjJ3nZlZbiLeaoVe5eV0CTSiSJqWgSmKdOLuMjhtnjR6d
GrFG8ybmOe9k7lRsIIYucvnHTQJfaZ/box6L5q7wRmFUNadnQj+DYocsYPF/CWkM
NBo9lrG09+0mJC+9TX1fmeQ9rYTxWTlXMRbG4TsGFcuZJa3YfWvmN/fjTgXqZVcW
oD6tyKCcxGzMBg8w6ggn2x0jkuNGFXuh894anjvGd/sYBtXG77z4vxIAHLkanC7o
q3s97SFS5yg6hKwd/1uEykzfiNXgqqlSlkGi7fdLu0bg25/gK1kFIGf4H0JEMdDO
vQKVXEB7pkwcvohm5JDxoPFUAoiSpI1AwV/YwC/XH0XSGePlSpOG7yQiYQ46tEt8
duBsLz3/cT0Hy6fzIGjnp42nKU59pbJo0rJgy+PcZuFR9i9zVjklF41NG7k2aiE+
CpvXwY0YwQRDWO10pJMzNACUl7nkRcT2dPBBQhAEDPqNQMOuBvpUYh4sTViSTetl
tfKU/2sZhwdGzYq6MEdk1hTWqxsssPCN/KzROFjR7HH2qdQ//fKcylrXufAbbdf5
RplobtT+DhnVJR2rZWBMId7ECvhFU4qy/U29vznWjkxaYj6f72BPhA87OP/xz6Yd
lHoAV1yAHN6dZH3jmgcyMDSpblPfltxA7WscisPDXEmAAfhHpk+GrDJbbLqaQYUT
zZdHs5E1c5C6d/RlAHVfwGnOWw+0XGRmankfDe5/A6WYpfL0/Hl9Sk6iJEMCe/k3
pLnfqF/xLrMMDxpfKZPtajir2VZf9XoIrW34k2NNto54EE7KZXvwr3f1MT8NL6JN
GCYCDDeJQHq8TPVZMgplpU2EfzuTD5C2jSvHCmRT+A2zHPdyPBHIhB+pztCcBSuH
/MEJes8EDuDqHpVm9kyHZJ1xMXxGnR3yjVpJ446cqKiR+uN9bzzIk2sMCT3kBt1D
TsBMv4BUlj9dDeriscN+pGw2eskiZ/Y8gmGBWbtK62x6+bCQW1jPplq7DGLhk5/4
dURMO75p+cAv5e2/lOyc2ZPhVIbnrTu+lNGckDvKum/s0EyxabUSmXLWi3gFGwrA
PVnzVXb79/z45sgku8JwpWjvJSLp8YHb7J5wRXq5Vt3G2JQipeEqW/kjWmxtUMHM
c5W+IlSBE191/LT2EBTshJOui8sndnMvA+bQVhDxaTwFaFLula9pZGVroHda+8ao
aZ8TEvjcqE6MMX6s1aVxQgCJ8km0e1ztTeJKiwEXn0O/5zLlu+xol34ZPdWK12Nd
RvPjIUncEdIgf/IgqcHu3sHV83/o1fF74KwYs3ABl4GZdoyBb9sCFyHCJgzIjw3D
MgvWVw0EeuEgNRwoVzYr141fDdL02O4RGXT4d/Fe4UR/JAwbr3wD4yX+Sc0UWvUz
bHFyO3qj1+XLQZix62m6SXaoQlAo/ytBAxsqoM4ELDyQq4V5/Il3c07JABmSdcrR
ZFuDlogsZKfERpTsRYSDLUth+8jlDisM7a06dqu6dDR4cn65cMhTQTI8WPPhCqZm
6MPhrRDAlNIx54xJ65gxaOHndTgsGUkdb+/7mtgYpu3Yh4Q3JxGXiPyAXcuVLVzs
8F0v/b4yOD4lcWcwhpXOFAsP9TvLyjULVAk/jRgp9XwgzyEf/IOqMvvHIiLV4eBb
hw97+Fl1Jgnk9dCRwwOi3LbuuMJiUtDTCsKNITHKHYATylyn6p1/8S1ZqgWTKz3w
F3kjH/bR1uIaJZUlaj+MWHoGlVlTskFIjy7pU6fNs/rkQEu4NDUR+pT6ya4VyCo2
7pnHNdjkMPEDvyvKMBte5e5IxQUgCQYdHa7PaGMIpS7CH7Esqija3USrXt9DzemD
y1G3Zk1uGa4tks6MNU7LaRNDAgU3hawoSpHNHxvQAKzJdGlQYXpcwy/A+mv819QO
Cjxf4fPg2BdhtHAVz9i7RS2Y24vVXLRq4Dex9D4BMkf5DZHr8z6ZPZUi+ewxoni7
ZmRelEUv2pV9UISVk4WbCQjSlhnV4CSyYf4nJsIT1JxiFvbidlg7gi5gpR8cCNV5
tBlAQ77m3/Vpkhr8wCCGGuxIoJ+6mvRl1ectiRTLJ3LfoG5rZ1k8g6PEk0J2fOTC
C73pmG46zvdHtwmte43leETwIshArNXJ1Ib4dUaN3bhszSOrGVBLS9YA3jEclwmM
Eo+gdD1wfIo/CCAOHSuHqUWWSj+0J6CkEp3SW7HfBD6EVVP6090bq1854pIdTgah
wVh8uTGXTaPE5afQmmpr9pTVckMbMnLxG8wOFkDPvhQlQjsAYaGYbdyqbTo+OV1S
MsRJ1FCKLJfjrxuXo/RcCQj3YMxTd7vj01+GOILVUaU783eUpxxjcj6hBzJC7yot
DX95kgdkc9AyCFFpfKfHJdQGPrwtVuP270wMvW7JqgT/wEByE+H5JHso7hoPX6Zt
mykoe21V7XfgYZGh/nz9Hx+fy96qiGsOgG5WemjTz9451LODz8ugl3hPmhWLoLTd
0VfwdYjKOdK7shgIgDu9wQkQ4TB7n5T1gegbqyM09r3+dlibCwWWHDNPkLLvV3A3
Cb1DtQr8xgZHTPe4fHpTbYEU4Qse39ew5BiK8JzVqrA8ewcgGRbt7cEHaAfr1YYL
yMnbeaRAKTn+DrpqyMaSvFXP6288ST33QtAFvfbRBLEfTpjUUkd4B7Kg91a+RpVh
dHdLFq/mcOOWkkfd/CCYBc+z47N84Z/oDa/fSnJDeVKaeGqaMNAQx3sdV2qJHBDj
kdpTZEAfIblsdJ4tOFFTa/RYinRSuIY/E15rm1GKNU56FpsIvRgWLTm+JBIMBqNm
2by+LuU4qF3O71T6e7hkDherpOJNnxgU86tirGo79XcJDqqzinj3X2AJmbdNy6s+
jIpjKed4SJ9FmPDntpaAioSktrQSKcCU4Cz8ITHQbewgznORbAhTEZXtlHoMgg6E
hTP48NBEnfbGIBbfjAUvney400A4kKs9NeeMf4IsqPw/a80Xxil27m9lJxkm+NGZ
M5jQDZUwdRG3R3MKrEAlkyTzAh74vT6d1DGZMbk+sJuaAf5udhNLPger0dgVg+o7
3BJocs9JXucIHtXJsFzJ6kjyLOpY5Kp8BWpm0CnUqisxTtD11nIllQwyca2ZpE00
KP5XYHvtkKYkNLXYE/DncIwibD+Jf9j79wdV0Xeuxu7Khh40EgG3qcgav3Bv+wA3
BaSzY75sWkch6HMgM+HvnYcKg7N/Vww4gSvzmmb0r4t9rgVkCDs652LcwViT0svI
hxm8Ba8WcyvDUyHLyN01lDZVjcdUuBIZJ/htW5VmSyoakT5RSf65C00JypCb8eqo
ro+jZE3U8YhFP57q9jJ8aZpfuy4NGZyx3DR/cgv2N16E27T8UdXRH4fxNK2knAgA
I08OkUulvC7wsxPcK4SzhSagghDT9sxFBafB0ioabXINCAgrMr1Y+hta/moE45Em
s79hWUclj11fK+vSLIQ5i8uTB94fFLuDOO0Ow2ENep0uZJzBdASrYgLtyMLPZP8d
+Lx6k7iYGdA9TE5uWjZv+FayePDeMLIxScaWW3U7ixz4trlbeUqIAWTMzwjEmEZR
v/awYrKQWuYyqNef/jh2tYHSHkkkvZ6p82FoGi1Psi9m1rZNjVrZcWgJ3ODUX8cZ
FwT9NFTh76lj4Sq435GiTPp+q5kspq3lpJvrj4MDqia0fewM0/EqcARybgcrqeo6
RShFQKiLTERflQPY3vNWKxiOFdzGphO9CQGujK4gVT94JrAata2f8h8uL6lN5Gfl
qN14iZmKi9180lLEPm8pnWrXcg/Wz49aotE5LP8ZKwsDNRuVjaOtuS5n9OG6LS3f
p1qUrEJHtyQx+Oh7u2jXd0CyaZaTIN4WnCLzIucrzWlhoImK6wpQGOh0Yhdj8nmP
Mw9tiL9Qje0te1Mx5R0W0y8N8+KXk9eibLt+ky4YuEmls28cLFBxmCYDFthuxw/G
FIgyqRx3T7w6hQJ1aQpw5R/xAFtD0TMAYQhIVVRyTpEPG+xD66LXAsybxG/qMOcg
1DeBkSKrcmyV2OR6K/1yc/3Q0rNwE0yf1XuUDA1pWfnbw2E6Lu5g/S4Izdh3jIFM
aAxADVKXNh06x+PSQCnZkrjxInMg/S/Y+3ydbn5RC4T3Yf/CuSeUpKwnSSKHQhT2
KTiJ9wK2o6sFipa1mvBlsgsx3kAbVzs+gMG1s06d4BWge4xf+Qc94t49bu/2PAQJ
gerWVKXqL0g2XRpXLQ1TUbiRyV7bfZm++Khe8r3DfzC40s2GHnPEsixVTddtE2CU
BMYA17C+iAl8xRw3T2C3G+9I6xSUSXxx3UnZbEKn3qDBgTQGAvmGh0JeLtydztj5
WlgbKOOHLMWwKeCzf493hQbSg0xkfoxd9MMQS87I9U5R8Ge3+maH42BKtHdTekDF
Brb3J0FrXcalQlYz71fTCnFIkA3OeiFi4Zp/tT86/r70l3BEU31NNWWko9xbutZF
nPNbu838xpGw2OaPlg1/MbnAmdjscWkvTO/x0SKK4sBOdGMME7DEWOHC8DR9j684
K5KvRqpF5PcHgK1aUdWHjH+/KKnQDDId2nvZey1TGQ17jgCq7gPuUiNHQ2qoXHZx
u5qioVLx1fr9JG0RLMy7UBNwYa5aMeGpXqdyZdTrbZA6N/keHTI5R0vV4u9jftnb
l6ll5rFX438b5hMVt6Zyc/eVqnjKZBZIAjXxev2AjzEAX6Y+NDB0Fb8dCUwYXd6A
vZYtEfQOjGpoS/427yzjbrDJ/7L/72C0IabultEhfMfdsxhQsz59WpeW4+ymXyU1
bFH83pqBrT+3wROtWOurbb5b1dr49Pa6ux59nOItFEAKA2B82Ruqoh//Tb4VIbXW
n593gfJxJmVCwhUUC6nh14j+trGd8heWiX1lMMeV3RoiO4SC6JzPr+lDwLO7dLQW
f3IU5qpY+XASsiUoFDhSxpXabC1bNudYDrAJQEGHTzw0pE+hSzEL7H6fQBOPqLe9
5ozq6bx4HFxeaYSfD03E7Maf+U2am+adUiLTZCC64rZRN25pMcfiWu8lGi9iUWZ1
G7iOTsDWsUYTanZxab4Q0pfT2RSIMPbwyzLmfZtVqgAJv9ufWbkOPp5DkcjRXaOV
XiKbaBjOmOFz/6Qlj38UMR15+oqdyl+Vw3pZx6tcE48Rn9xwOXxY+yHBam5OmcuM
zq1ngR09jI1oohvCLocL1JZ9QsClriUOsYz/Mj217bhyH7cmXN2MIfP+2Rq3jmZD
aPbMo10SKYr1z023bTbrDhN9sxG72AXM6jAvaPYLCOYeIylrdtBB4E8DhTENfMn3
Dft++Uz/IczA42GNxS6xWGRf3QVM7FHhC12sCS1fgn68r+SCD+fVR30iVY2go/3N
CFlIRKnjRPuxTzu6J40qmDGjDHQPRcFlUtKMbQUfmVUyJ3VW4UQi7Ebgocz8ScXm
iRLtKUau+bUU2e+qE2lr8W58HQspDzKQw08N/8kIBF/ULM5UgCofrWUfIBo1I7ez
UMrj957/LhZugrTDCcFZDZKIUORvGP0gEREWamu1OzXQAZ+CJ3UEP2cWoSpJL2Do
IgtuU2GIuvjXzsRh2QWH+EkqSKFrjXWtZbSSID6P1YMJrdnAPu1/JIdAXPtq3Okz
cGW6XZXHqHLW1Fv7nkDwFLG23OvOvBL6KviS2EdVAR1TgKfDLs5wkpV9RK8Kzjy3
AmEtQlMJPRUJ5WgfKN81ANpgpQAppIF5EalKlwH8UNaTtP7/3r4T3DwuNdxT7diX
b6wzjKXAPwJNSmBaOup7vauSsTb63HLsnWaC0NpUrrST8J6ennaG0wOvWsYrhArh
dGbSF6aUx5u1+TiQ+sMCa38mVWXa7SPI+f2FlJ8kyvVGO9dxQwFL1iWM7m44WsMt
OOqcfNa9nB9WSxoV3Wn4EYblXP3VAiRWsnKrHlE8mal6nFCjweEKxwcPg2UIAdvC
NAPjkVV8RW7j8mnD6MAn8S4U5EQ5g2kes+UF2arBjOaPZ0LOHU8CTN4ZimWF5K/6
IbA1N3VfEfDOQ0Ki3vqqccgXYFOivrJTHSD6d4dsS3Jdf6a6q0GOo9TdNot8mG7K
zhrgcM2NFltzak/1eOGFo9D3h7/Wur9o0aUnzBM1egKPyHDh8nD2GN2xYUKsy+g1
EDRjPpKkkTnXtAmMbT25eAQwsa7uWgX1xa1HIOhM12HlvlG6XcqebxVwko1DX0eT
wnJRQDodtb2mGxmy3paVkiL1hUQRLWIFBnNRjMFYgLXj6JaPP1i+6+tuAj58VNjI
k3ldYM/ElZ4WaYKRz8ByGhYp+kX99GjTLbsIslxOCjEa2iYES8i0+zBfd4RqZXu9
4mVmC3VU+tVm5x6eUSqIutPN3lSormjdn8kVIisiVVjz/ryfsGlfackQp3JMg6xR
sGHJrgU+03T+HUSvAER5RPby0hjoMRRjDXijhNETbrM+MbuXXNB5UizRVLn4Ot7O
7mnsOS72p2Us7IsK6UsOJA7yUGjTvtzDWabF9ubBzupMCFP9z6hu5zqVKc0ZW1jB
NZEWWzo9K48dCGK7S6ivFZn7E5P/f5nxmiae9RbCvVf6054d0Fm5ArvpimRMwy2Z
pu3ASV8UYm+cn79d/2yBZ/GvfkY49N1bsOkWjAVkm+/5Cu1qmwXK5uUdd/YKG53M
3/y+tiAuBcFhKE5HOO2JvJLPAA+/jhLEHi1ppKU0YcCc3vv+xVNdJlV6vf31vkYu
FtgILdIcxp0stuER8emmbli7yDdJxtgyZSqxGeSerHatF+I8wHZDmA7gfMDuGsL4
hGCLPw7Y45l5NLCzqKC1I3GCTkANpjufejWKBgDHuyaRGGReYPfoZgrCpdHdXwDD
Q+M34zcN3Oi1QJeYX7a5AOGKVJ4i4+ug6+OnJXGiOwHtW9NuOSzm1s6Go1CP+D1U
ZFTtYd+GUGiqzKCftPJ1RdTUm+OX1ECwAEvQTtmZVnRww5lD+59Yui0nxANs7jPa
xW4bqcyag1FdRH498qnkY/TzHxISfpuM84CQFjWTTUPpqIiz25mdQbeNYa4+dpiv
VMnfxSFym3i3hTN5YuHVE6o3xS8n73pVDaxV0K4wCLYl5vhHIzZblUU9OA+kPPOq
KiTTg2yU9rJ54nmwWBhhBGSRW5Cn6DkvOs/wsuroYZGQMyp9qX7FlDlk3RXo5cpa
YtiknjfQsZAcGAQPezbL6saLB/RPun80j8YQ61ZTETjibyhomeOYS+6yDMuJa9m5
ud5YYCKdNt5hHAeJRVHOr59LeErhIXbF80/YVN91iOQW7lm2d8K2qGHrJwiXb+LA
WrCp1eSiH1uEQZelbqAD+789o+jauF5YxPjnX+/3bXWUrCSk/0vDN/GGqjYVG35h
iE/OvH31Db1B8DfTSHdMsCd3aao3lD/0hjliAzDQnbcIRGGlDl1oWhGOWH1B/VEi
lpZv+98yE9y4hhNdg9adoLd//pkkz9KtBwi4PByx3FqdrkgIvcXs+9/r4oTs2n/U
jHJErMlDQJ3d7yZR/iD6aJPhQSdAa8WFlV/cjM6n92YahJzMTluZ8RPa9tdypwTF
tRelOvR6M4NEAs07VTtDzK1mlzNG610YHOtuoP+HhAHY0n+Zh7YGDRHGSgjhQL2D
WRt8+mj2tip3Ld1N03xQ26aEd+1jdI7aklRLVIfwpOnzWBLVR6yNnL8+hVM20vDL
B+uZEIWq5wMZuumdGVjRNt+fv9yQz/jnQWUl100XLziPbzpxxkdDHh6b6/u+XG7q
EgveJCtHdtqzPIXOjcyQNhguwMcDv5xA05U4XS7Gls1uVDOefSq7a5woRHNHR9kv
RIFoDzxNdALC7gElsJxpNxbU8yOuEBJCbNSD5FScAvWEZftU2sOk97+CCpZe1wcX
H2iu87Oo0kxctG0JyzLNhU98d54OoI1s6PIQP1RZJqloHu+PUPe1/QrQ9+vvm15s
4lnMQJ6le8INX/OAn8nuV0khyPij8AwjbratKrXa8K04p8EGyU/be/bAzwH5HnOu
BHUlEmkJZ1KkqLD+1TBDBovcOIJTtKgliOHCevx+C8QALgjMSYxO6ovn667TpRT+
wWeTYMGAPHs+KjUkfrYy70RH1+E4/dQrWfRpGQQLDrB909rTy00RowDLVdiB3qD9
H2HP3WGyysjQrZp39FRGe07z8lEPL4LnY0KVxBRdbvWrVmq/B9GPsPtn/KRWajps
QXS6WNtmzUE0m0Xl+BE3zZ8lu3lWS5M57ENW62dKg5tuktKZkLxQM6fi+VCm7QBl
SkFoRqogel8rMeJ26zNpW4Krlv+1NrOnm7wx4I/qitRm+CY2Or6K8Wsx4JN2oAmA
2w1qkAbkp5E+9CeOjfbotmJxEY/RvmRx0LLKNpbq5keasAWyv93xy1JhR1iqjE6o
sVKH85d9yybtjQMlmNas9rPWeuBlDRLWuElE1k8V0ECUI5H7pPJTAaKcgekpSa+J
53SkMWynGyorQb4ql2KjLJKvfe2JueTNFyUQV6zlgeNIE7x9/e0vbNIjYbYWeJXz
IefFOqKG2Ge5bQ4PRvrRakvSDB+1XzegbvfdwLNx87mADW3bBPbqtk6oT8ARWirw
NMsCEZdFsFGeuaAbNvVG/KemlM7agwRaWg069OXMYAaHAdseSeMZbJF6ktZ8zKV0
9yUKVq/aRr3PJ7ZIx9WEAmFUT23f7Z5h/mHoL9mRfi529WtLTW7hskpKa6p53b0/
H2BG+tV+oGDD7IZ6h+MMYSz7xlpc9cTEosSJCrjqd9Et6KNps/ZMS2350AJGfGUd
D0UeqB8cKhlGZ7bt3rpUIiCMAMPe3pNIMFLzXm8PAn2eah589wy6KYJcWAghsO29
EWJZcxW+OSwWkVr2mn3/+B32EySBezzL04dAGjAWEKlwmgPQSw+w65wo0scPbqSp
gV/lOvWG4j4knVctYf0EGEUvgj0pCbJQsl5vsdQBqM3bqQwnEo12XZe/SZVCM1hZ
FTz2kRSN4eXpcyBxUEXK5YV8Ef/m3JiGdRrUF+Ns4wl9NWA5FKO91IAZMcYZDoBO
KFKHieSYU2P42EW48Om2LL9WFr9iW8OQhVaLPZ3CHwADypVgdnLyfcjOIqg70VBm
r8ThGUGDvj5VfH0VMJDUrMlIfhONxTZhboO42cQmGL9FeP1xeR4PVvSOoKPRbUd/
jzGKIgDzbDBPLPshM0J0q31mhFnz2uCca0Q2rxmmr75Ge3eAAeEX9kanviM1y7E4
rhc3Z967rzyiTObF49y6C8Mj1yYdfMsVMCSCYj/H20qvo778eanf0eRrfyQ4KRXo
XvjgRZL8gju30465UVFuc0RULjNJ9tCLl2TyKohXhrG0jNaiCdfYIR5J9G4/AxcA
UxdklCGAqzuWHafNgfvc39K0DKDY2hcGHIPu1XdbrA4ZsvKNmUjw6X+gbMmB4ZCa
o53uXxa5z9kVYOK6Vl1QuMS2PxhkK2ZzDD6rNbivcUvO7j2bdcRofWNwadDaEE7P
nmICsB3Y0LiwpCNF3CqpNoCtVcl+yP8AgYgZAhtmcC1pw6YjO14MEm3xypYIidqK
0EuCmaVeOtpH7PI1dzEjUygY/3s/QI7g3Pflb/hcZvZTabGaZXajo0BCPSIJPS2H
kHEZFP5V0kDz2OEh2k6trbngKRZlL4vKWe0s3cyjFwTYcI1q5P8K45MoJplS0UGk
X106RkFiUe9sC28ia5wK6gDToYSsWyU8dBIC9lzrH6cPCtoD2H8Mn6VtnI/7nFZb
Gm8VEY4Is1t8yXCjm6XEYprPj4Y9oV+pgO1KsNaZxQV4CLxCqKVnUfqzUKblD1bL
xUpGk4/nLdVQLaro3jIUCfe97YH4Inw6m+pYhWohwJ5Di1Jx3KnXk+5Umsyj2lI0
0VLjfDIeXsczEgO2Lu4V4uJbLv7cfaTbKohEerSW189jyM9oxGrWHj02vfV4zupP
hZLqYSRoGlhaYNpYNVY6WAc4QWiUsg1MPMFMteG9Mhi44m8XCBuH17HrWnFI6ZNy
R8HQwAOlRJTHNgE6Lfdad284eX5QwHLyJrUdjyTs/cXvZsjMjnyrtSltkWaibUD4
qlbbqF9OXbwxZsj9tvDNM3VtV1oL3V3XvJeQSOrvPesTic3KOefgQXAWVJkw6DFd
kFLFrlA253S4/OSrktAYMsVRNGTiVKRaLSmX07E2uJHI4s2O3UQLgYlKzo2aPhIG
FgPDfm0/mAkc7nICxe1xT4Krc6BzOwep4s/jTPfZQg6aQdqXj5atRiioJ6JjctvI
BqvuXr4C3+Iy2dc3qpe/a/Bv/Nxjmsid3YEWFjg/cCwiCwsSBpU1unCrfRu8nEyW
+zglmtAUId5O4LnpsRoBwjb9Pnyjru+PWzo/X4Cpgyh56JunyMl0VHOfRV+dS8jd
UP3zThfpZ79N0CmoYLpvRqbF2v4bHeyf0y7o8ymTvkieqNRQhslm6oNXBlvVmfA1
2AevS//m8dyHTdS5BwemSJfO6If3+LwUHq/WyFvWpbvTNKo/Vu8+5eTfD7sh1lZ2
vq1FgwkNG80TMjpiu6LD08ot4P/7gD85Q8jAXa/u3WTm38VAbt9se354j5+o5cAq
mLBWTexTOzsjw5yfvmls3Xkyhns7OesYmITfK+fO2yPVScXkOSpfdI5QV4mrbzw+
UEItB06sr/H2j1O4x32xQDHpJV+jqcfg7VL2Ut0h7F3DZN2RqYREhU8gZ2QidGNU
7ASKK33v+V+VArPyRBZDwQ8vuzs5uRTS/eOvKEv/JoAUrsnozGpW9paUuxROUVnz
klt0kSiiHgHU8ZAJQt0g0A+0PWTeH+Ly72HeJcWMmMD3RbyUDseb8HU9TyGUGaLb
IOSicc7xeEgxMBlbEx3SPuWOR1AsdwnkNvn21L2HKqmFCd3pJM+OtuQJ2Fzo/sjM
n94kG9sEId9CIjQpK+VTZZjIp8vLBduivAANE9Kdeal9UOLMJYRetYYc/NRw+pCS
l6q3kiMneCjADiMFjwaTs6UYcepTOeM2Mjy3tWi+txy4QFbJ9RF8nkrcFwhQCZLt
CkZtQxTR7TSWY1M4NCXkoUzOov58jAud1geSQWZsWBNDrnyHQu6a9+fflNzGr2Ax
Z+8fsU41kfExkO59DWVk9v7lapDEN42JEDKOPBqAiBDnQv3sa1Y6bqqz8uz3Ya4T
pLTVJmebdic39DRGwINn+fkA+RYoaGPIgaMGX1QLFX8KFWa9FsXVsRxLFhCvDti6
06dHf7YghvaQ5hJwk8NBv8KIiHDfA1z1oJNIpwj0YqBxl8YawT2Jy2w5SjgwrZQB
W0pZ7Bo8Nhh+rgLot+XacmgssKuGS/CDFQCDXiuLpT4e98yy5Vl+HpVIaddwR90a
2ZGXAugywL7fLFiFD7Pre+M6gxF/HQtzLqzdYr7PjJ3Oh8ctTqmCfpz7uDVdKb3l
Hmy5pLnG8HV25c3KYxyre6Zrs0KEB+8pdNuKtUwbZ4GZ9FsakKfHywWosCqg3psJ
Os3mHeT0DPDoPaV1egHIIncHAY18z3uhovyYl9hULarEw19Z5DhpqnZurpub2e0m
AY+oP3dFMpGcjD6bJaAtJq+Y6vQJ/vuCHvs6Ooauj3UhPwBtpTk7dZHzrDLYgLFv
3Yu13OCBsTi1PhVkDoUo7ce3FEZh0iQmgHBp2zgyUOEVYzkzWx1s95rGDOdAJi0p
Py3dT+Rm+vWBIMjCQBn/u1c+oyFPu03e/CdqAmY8hWf6JntbdqrYNR1LiZwW9TiY
qjByraYzgPMS/e9XW9oV/jtEB4ZFZX8/BdYCnmFIFPuYzDgNO8Bwuc9NYQmtclSy
J0OLZiukrf/ST+ypT6J8A3NpvNqb8oh144AeoByajVxGtN7fetmIt4zCULVnR+zk
LfEAVYF4bWovj0/H59ShZV3mqFx7WT6TkEJywsiXxliS4elKOsEzY47EVWCg0kwI
lkmvQteRfFr3Vsr3nVHCHXcTs1/c3ogxMQoA19wuBv3xXETTfISCduqjnhRRIwO2
kKaguZ903vyKzOSTEetp34hbzluLCpvs5lNOh7+zOipkCwewWqpqF/DNL2AjoG10
RFsoHedRvDkBmT//FlCiY81Dm8MB0BlLGewI/CWkA525+Ts3MNsfehFxkj4Dp4k4
xaWQxSzIzxq351xBl6HE8Ph5ojM0JO3RWOQFb541s0ZkH8THnDTqWPlSsh3C9BjK
p9uTqOphu7iocvC1ARG3YAVgvoT0Nyo/NpiWbvv8/KppdWnCquxA0P0FbL0nngGD
4a442qqhemUWxNIt8vnsJFrJa9qDknh92s9lq+J9azW1hOMnqtz8IjGddo3yuOyj
j61VAXiAlk4eAkWtU3DM0Qq4xLH4evIm//rnnXmh4Nt8H0W83HlborSYbYxHtBru
olhamqm3Xe5cszt7x2PTvcqZGOcvAV7Jeg0V6+G/jAAY2n2UJxa0CA3QQdUkt4aU
KQ2K0/1F0NMPrY16n1WI5YmsyPczQgs4CI8W35v3MamUjhAp0tm5j90yXrzmkdSq
+b1LmcJRvWykIrmKapl84hwbNrkP1xInc4D6ZtA8icU+VAFjDRtoXtdoMSRqd5i/
bT2Hga5NrI8zl96LFI3aLkqgbpXDNvYoTERVSWtoE8BYwKqHr+qJyr+FSX2o/Q6d
zy4PQNd8h1b3QZSjy9JY73Jv0mqYVbTzxCz1+SU3TNbTWhDQqajoSMajKhM17IoM
xPsXAbVQT0vg1V6NdjZnSgio4hOzZHHe8X3rRVvtxmu3SNmy/bcD/xa4CsSog8lW
qH1G9Z0gnv6xWj8XYKX1aW5WXgEjAxRZjzj4f2gDeOkctcIbRBK6125F3zySSC0X
v3BxIZJ817XA/rTrhrND8tWll0t/RLv6CTeysi5cEKMg5B6HbomzzvoFowLOSyzp
mhXgpYovutDBYbQv5P1C/DDUCCLNKW1zWhQ1j1UgOy64hNJAZncftswNNNuBr+nT
tg5y/MbXRyRb/irJuxMecXDOkyGuCOiN1Yuwglho1sJ7uceR+Xack+6GN8nCFOzo
JeTn8XnYY3Cjvfl4K9aFFw58VlFKY6+tAQf3MzU9jWqzSM+M7jCxpQKifMjqssbZ
pQXoUJHvs1Z9ujxVGNxNamC6GufWOWKMa53iNM4veEHc7IagCFvoldb7igVIK/Mc
Irhpm5Cty8sx/YG5tYdG3KD9pTjLqWe1/6sufUb0TNo6oKOPwsoaH8Q50RVNIDyu
GT/Bn0MJPZ0dJAAvHUFIGQ43o6Jzdom5zUpVfl5mwZLCg5KM1hTMeOLD2I8Cu3fq
mqVuKlP/jBmGdrPKiGwlRjvTz8ioVjvKZ+SZYoC8Erc2ZhugwNYr8H1GqZxGnnFH
FBYYb23DDQdvcXvKkacxLajnf5y0UL42lY1LYP+RWbMXNFXfHq2pzsQFGxqVU9MJ
K5AgOpo9gnHexvLx/ezoFYSWzp9P5lW+kq6HrecxS6t+V1M3QXxWC7JHvAO/Gj8N
T1qmGcwXNXmu1T8n6JJJZyOao5jgz6f8sNzMtpWDVbFEZIXJyh/VYEz6f618PVJe
6iy5bEbd83cT8WgdFCHnnAj1AyLYJL/EOwHyBGEiEXe0GExzjjQKF8gpo7Mol4Kc
3dw7HT1/Fun3fZQgOggnWzV9vrtNd36BtL0P9oX5mGfGfPZJVAKaaOiYM+k4rclc
EtUwaT3I5k/c1RiEpV7CZ7SA7vAHL00qFox2Jqx76BlGLj1hNbwUpbwmsvCqB7XE
MW+b9jFSBsYub3g99KFtsesbMXGtVxrVfb4WHihZfcrTy/VOezSkTKjWB512cNYh
moCuJto2pLRHgaSmDIQv460wRlOVe9VZF2IbQ5/9Msdz+2TJ7D64n/oeNtopneBP
9qtXefhCS2jm1wTncX7cbstNYq1wenz8DXGYhjD+1cYIc5hwBceJgNTbmarGOvcq
fn4vbsbsH+OpATtWUsoXCLPsyE/JYCTm12p1px3dREpcu1mD+y2ovPVzra9Myj5l
U5BF5jJFh7SNEoURjVU0J+srmldqweMkJ7490Uje3aokbjT4lVaTd0orRXDPBLPG
ynaWJby3awvfWcguQQFapz9llWQDhOlzuCzUAOVug5XzQfGJBP0ICYqqenuWdYX5
J83lEiew149BTJdkrTMwvwMFF5UL3y53zGAPfWnpc7k08fslkd2iR8NnoYcK9vll
RC0T3GtVo5QrePic6rZzgszn+Qb033PZ7ZrXeKcRYFFRXTRjQPEIvYxTyYSbhSDd
7AQN4p2iWd2faCgMQCdGR53yV70X/2kcPmfbs8HLk0o8iDDeqCt/CKNADJEhXjSz
KaI79pN4DhLThTyoXXhkMB3wILSWjKx6cIv8GWGxUbE1sqxTRMhDEWQ9vgrkGA+q
XuDN7isECGGqxH4Igs/kWBw6GX9Q3kX04mSSQdQkiUKhTGtUK3zmcyMAbBV/1YWX
oa4xlY4OVGIQ+7T21XP4ebkGc/QwOFONvcepqM3uDSSBC6MekE/vyq/DCjsInFna
MMFV9Z8CCxZ5L04iAZ+SxfSr+yB6hobImtwbHkH9ug07NSp5vSUVPmPvac/fmxky
MetE2PUQMFubMgfQo4tNeF3Ey/7PARa4YhNNyD473HCfVBzwgjOz2uM3Bs109Nuf
0cydj27ITrEGgpY9Poa4OY+qhKPUc9oU0Fh9T8F5JK1PbY/3vIBNwprhJTwyeUbe
+9rnrx6ds5MrLJXr5nVGAm5vQOED61irtCPuoMVrOrcSlm9C17kwPsLGkPlV430V
JQZnzKH+4DQHgow8upxgbCmCGTcxGzsXGd+ILqHNA6guynxQ8tYUAva//mmAlScf
EsAabY+tqqYh7FumVUd5eWCVU8iMmReBQhRtNKdemrVLCd8xImGDO/87I8vVWT2H
xY/XjdvEMcUPhj7BCJKIzI/SV0twFOgWFNZvJ9TjKadBdMeGS6T3+3ryBKPBp6qQ
l3taHkiSo1Qj4H/kLk6hs7SR7Oxbign46t7gC14LPqoZL5vj/GCDKnurbPaCQTCf
9TJnKbE91UwJwjKpJd7oJWHmR8RbtgdXUoG8MI6OcjYMxQVp/s97AFEEDDTI8WCu
X6XDQ0yUdCA47SEjGRTLATkidTTvhOFuYPwMbBJIX/qReFmJpS0ngPv9siZhfaNT
H53yQYRNh8KrlsgvWqImkJhLCestNwESQJ9+xIPZ8dwjJji/wBycjOdCeJ1BiUNY
Tc8XdFUKYgVwUnYU/c5tqWcwPCD6Q81BAJxWWbh+bc1dEPV4TlGNLQit9ryGRizz
ot+pRiV4O+28frkI0p8xslfrWvJxS8PAeBMv5TJiGTjYo+14XWDf+qY/HGUIAjOW
Pl676eqTS4SzqsQwLRIBlu4HAjnkB6KS+VOVfg6Rj6E5wGF0CXqjc0GqLADU+F7Z
yRYfSr6qxB1GmsdqUzNGvPeFStfMFOfFIFyn+w03bxlKul6HPEzsBeD9S9WMpkQh
CR0ELHfPV8tGHHfSRlyzjd2trGxWBd71t5OopjDAKOZW2LIVw+gEUl0TOc5g46BH
wta3Q7QhGMqwHMqbWQ3oqVvDvb1u0sL8ZIgfv0QFkCoRzB7tx7nwjK2tfZlyKArY
wOUfmCRAk69ZB9MNuISdf6rxHAIoQakfn/90ofVwKF869dfelKpZ7ZY7x17bMQVi
twPmjG3M9R0QzH1gUI5A2gQvPnVzE9SEtoS/3+TjJ0JU56M2ZXa6LS2DKmQcsQZr
kvOw9kcgfwFR30SGn9hYO097GHiy9z5jFCSv5fnBigqEEs9b7AmLUHH5X4d8T52K
EJchiCYaVhwjq+8ZGYZk6BrPRbaniTAgbhAIZp26OZ/xLC/kh+cIPtA9W+SgGxOy
+v0vfefAr3R3FWbukaOPlvuZT7WqvOSiSfDDpB11ey3pJRIV9r8S35saj0UEakCl
Q3v7f7nXDV2H10k1pDDbVRn6jUS4YR8WX0FAnLu+i1eLT6TR5v+/vJ8mh7vMWCxl
XGiFoMNWIY4rIKMEV8yrWPhwwiUAPS/1OOy2GL6qSqenaAE5dOs/jaXsNnS6yJ7S
b/7AWaTdKVS8Z09vJTO3EOZfsQ4iXKkO9ZC12JzZ15YQY2jr8qqLHcYWyB4zyyKb
a/kgoG0nfD1Qt1peFFkJgMtvqOuJFw7cOfcggUTzuDOtdZdipr8DauTwslv5Mpqh
O1tkpD2R1HBYvGdy/BpAfC9nZXLdmyRtaB3LP/h2rc0K4DU8CWfhszKQpKKeOHmL
leL2jHOaydpzUBi8Gz65V/BO/ZaH+VYjIdWBEQdnUdHWnH7p4plPrtGycnRH1zoZ
nV095lxWxAoncyxE3Ka3MmO/q8kfg1Qnlj0rm+lCpukZcS0tOzhX+US0ZCFr2RBi
SxSbwDny3EdYimsPSGwowjup6ZMRU5Go827q957dGzadSf497v0UgXhkpH0hTYJA
a3/EgXT6cWHk9+yxLINem5uZd/itNKbZP9oRyACcHNSTDm8K+eZVv5NUjqGGyaeT
vmhlVDATZFRv8LIZi0Cc0tKEGzoaKRKfRBfngE7O0co6XBdkFcfGeuhnvoWfVcwn
rf9YZ/Mf9RZVlI+AZmoTBo+6eFNDUwjSrhXNbIAaISSQU+ALXE8BoxXn82m1QSsP
wlKHoNU5jVVSmvRdA80TLNaRtihbbaqx3jxUbdmCxQMz9n8VnUJEXZwQVy9jUkZN
S+C+ktHYWJrNSbpOnVVC7hq15NC/iUI9ECEAvpgEKWUJ6wRK8q3YGxuvPARTxXDc
tfmwQ5dPMS1YommTfIx6C7wpZXxRj/pji2Kim/bxkEuueBh7OoiGy0DpP3MVSTDo
URZ9RL2TNAVtb6LeZUgRjIY03ZT63CeAMX+IkgHIkO8AJf6xjTI7EJF86/MuVTgR
jT4WrOj3+NjRLgAme3ejC1U6sGwYju9yE+3wZavYBMd7ef34gbC4zPIeUlVmgPwL
Rk7KId8hETb1nIZuKpjByMHePxJURQU/OG8a0TmlwYQk+TozhpuSY+Ybuh84ZYH4
pbYp5OhuIW3p/PNuLjr/ekYU55GIFp89QokfeRmc+FOn6w93QoobvOWAB73U73iG
MmZI/fFYPEJUPrvTMeklpsgavo4/wNhQpLgfmLONeG23uGvJwX3Yv+W0Tvv/OSrE
QDrT0AXWMiwcSOsKWh0M/hAu4XVgo8ZXv1Ow97BGKJV/Ku99YcYODfdeGCmqDPuy
N+pA78ioGm7qqgZQoS5IP51FKGUbQ4L2ZLEVcmxE0a8LFibXq8zf8vuEJpDbSw73
08m0BMU0JsdnMyiQ6SF9JqNWkyDSAXOnBR2XidOA8uLQwY0noO5eEuznmX5HCnL2
wXid+y4kV0tHiNIHaEkVVX9zr9kMRnFK0e8LIjGurW9WwXh3cdMDBkprPuVfhzLx
KwrZ4jxpkZ8PCe9Zw4CIzWZyZBIjU/97IsrOlhK8ey5Ne8QZj5LvKNaQ2Ll4uhjT
/nuqVzg5rxLjttFovVz+yhPMmGRo6gzPL/DzvNrdSPNs04nno16oH4fWU2r9IJe/
1aHfdntiisPDdqNYoWdzaB8Z8u4XhyBQR8U+692RYNoaLogFm0ybTeRyBkKe0P6d
EmHvFJRoWN0k1yAggiKZ821zmjkW5D3TKV+LzGpgpH0xDeRkRfE8xaWbPehebn74
jEktYlufQP5tO079mE6ksBAmZx6LgTvOk47SGa0RugW0267ooUtxYZ9OPLsTJers
Hawu2KlXJu4SXWSGla3umpSV0lvn4LWa+OCHwa9YWRCPdMOIH6jG+Drr9aKwjG8F
5Z9xcjv7aIsXfot/r/NCwBSy5xm0PYShSi4aLtVMOeyb25tcNOY3qU2kGv6dde81
GjM4tApjHxfnxR3bZgXgP88ldrv9fy1mLN0DSUfYkThdEjFn/pnmdYrSqKN1DG9f
AsHzsl19ZyQVYOQE3N4a8HUCdnTloj8JbdQC/uhaC3vHGBqMX7Po/Qy7enmyRTyd
uPPGL7GSwBC+i9+O7KY6HFB5EJorQTOlrceJxzSQbeRUZGalnNRUYd/XGHgT2bTo
qxwJpJCmK2bVve2aABDJCMAwbDuiDpfJOWbcqnblktnF+zQh5J9QSODZLngth04G
tg3PIRAbV/Me7BTYGYz/2eHxoNGq3ewTmWBoDyzWl/7PlNl5M29U+2D5wkrjRaMm
Mo5/cMC6ktEZBXBwU0mV9Ev6MjcZOFYyGZY3dWBRyM8AUn/76aJ5o+L1pqnMw075
dVa8zaQSNx9Jwa0vEZ2GojJ4bzQqwjwarcFLCNiC97H062DmcqdyqC6/QdyRlzE4
CkR2NqD/e7gX6WnxD2Fhesen5rX6o4SW0isy1i0ek5NQBLorgphSlnhHLWuSXkkn
NFln88Xwg/CHHN/oAixE2AAfL5Jon6Fvdzp8hvQW2+RI5tFxHBnANhWvfnEJmeLF
fsAZsmvLs1ATzibpLk4FhrNWXvPtOOZaForMOenp/uZpkf7Iy0YCsq7NyMPGXT+j
nG2hT/taSINQ+u2+W7B2GUlsxNGp4Gf0/LjUi+kseSW5uIU+y1i/lRI6SrHE4mIT
pPMLTWGexEkDZRbLZZrRCKzc++v5IsbJ5dTpPzKHFQLVe913LK8RquqL5tc2+Lub
2oqWnWB3tafC69tiRCstYX8TRkUrB1COmkx6nbnfGToTXMG28Bg/iYeFVK5YASO0
xR03n2FrdbAm/YGwAqRYIlrN/HPKAW1sal6iCjm3BRb5M8JyT5bK/maNpGqfkMJ5
c0aUqk/hn/jrGsJ730Xe7JzQPCnzci6pXPh8+dopQHtZN79LOz/5LCZouEWt4CnB
Sd+hEJ3GJY10gj9tPmI6hbRWZQIRp+oliPNoG7GBqMCRwDaYVk5Wk/ylopIi+/rV
C68JbQJLRlIY7uFti4P6y3++wf69wQeRYqF7N+bEU/bPBoYC95Py7DDRIa/Q4Ecv
QlBnnsxBnGFUbWt0d3SNcL8OHWpZx01pWqBFCa+xXJdZLEyoj1pIh7cdR+tHhj6H
J+Fk8htn59pUJyAf2PyYWijkwvkZcnpn4wJR6dfu2U8BR/bx8LWAfsviUgK2hA31
GUCX6NkGgb8Xg1fii6O5NoTQxUEmdqrV6tIawhK2Y4OS8tJ3BHM/FNS19zIWvEH1
8fK2a7jMdSVgi2Xm7/YH4/qmSpDeOixPiHZ2wtyjYLBGCQpeUHsai84Z14K4CTWl
unvOlRUlJi7VDZl7pqAK5PnR2if6rKeRYFoSXOldK/iEM3/yvcH6TDJH2yHXMWjs
LB4YDnJICxhGCj6ryCLDsIAkzN/4iG1P5o9vIhhQvhLyaCay9EW1bHo+xTOq0VvH
blQkgfI7o4h1TKFKsygQl+JY46eG+YN0oSvbk2Icvb74UIqyWq7pq6Er2WfkMXR7
vcaAhRkAHdoWzfNf27M+80M5oBSKvKWacuqCpPW+N+hb76KwHpSxwUcqF9eH91de
F0A9jR1ISfaoHN5/AhvfXXGM7tPyFh9JMf3MXcRvpmcdMH9YfbEbNILEovdXFEOO
MiC63btgumSIiybmcK6+KICD+j5gvaRz+PD6KsGKLL6Cdqb2y/ws8Z5QkNogkEnd
rJWzH5jaepTJ6RUt4jIwpgCnWPnRwrl4G/EjPjAFQGU8BjI6XeYAmDW7wO/yOaCk
5WthSxoz+AXJ9KoDnXF7Q8DFbf64jP2ko/dvKkVgokI6+yEHaDjrSei7LgG9+G2+
hrsv3VQ6+sidK1NuwKkUanGIjBVgDJ+53QcYCJR8+/IDMeQ26+HZwAL9CHOoKODh
lZ0jeP9CJ4vTQixn/TLo6/UYqkWxe3I+NIutiMtlXx/0nEdHG5l961lwwoAULNPS
3QEcegZyCegJ8WasvdVl3AU6FSxb+fd2qOuDQ0tKqEuy6nFURT6GTKeK0H5WfM1m
+k2Nj+JOPZ6NA4uYG8mNnBqvVqL18p1GslBPkL+TnGf3U458VlnwK6PJg+kYdUhL
ORU7dKYDs/HSSImFY29zG8yh5wWYns1Q4HLoveBOrcZNqHk7dA0zr/hg3l4UWtdx
cxHOZhYSX3eI/PbSNdjJV1KFHio9Z1lzrEXmIXlZ7mjzVmX5NEkQxOLO+nVXG3Nx
vbaLK5V/DEdW7BUjT+pHnG517pUPffpUfy82F+u3d2v3ypmwwddeMLp8P62Ki9EW
rbLl6YSRR4NFC5ldOx67c0GDGPqE6OMmJtDPU8oZq4QTfugcBU77R4d4Gu7k6E0f
mbBWO+9Cg6ujGgnpd38tUaKtqR2MffGLXP/cOK0Tn7jvS3alP5ziIHGQMLv9AMFh
mDRXkSGrWD2n0MC4dMlsJEPqPbaybiVGfhmTXShU8zr1wXW+1hWALQWT8CQ7fmh5
FmH/CuHD16xCWm8BoMlMR1I71jyI5O/AikLAGq3ZmvPJIwPhn5CflEg7XCS6EvLP
Ae/HbL2hAfmKbauqKlFFTO22jUqmFVaZDmIqrorC77g2GRZNDa1uzB7rabNJo7oI
OB8myt8cL83VIK2N1wPrzjBTWc9JsNuwRib5qwiJ0Vn6N5kdzT7NSQOUKKmV0txr
m+33eW7jySe9q5+Kl5cCrfvsF5h2Dch/lW+RrycCI8u03mgZE6bZD2HYJcm4iR8V
FhiqCy2m07LjIm75t4ZbaOVqo9+vurOV7rrf1q2VHpqj3ZbfN9LyLU0hR4wj2hV4
Px36W69SPWT5wDwLsefrOMWMMqf+7wQDx15HGdRIGse5l359RoUWmEDOq8zAUxHg
O2NsBb7DZbFpxVMfqbtKgqk/D0tDUGjBI2YYkVOTbWm97vVUuEbj9xY1dgNML7lT
CRuDS0LS2L1yVUPoAlFAPk6KiypbzPC1WhSvhZlCSaYkVuZ//shlN6pgoQ4eU9pi
h8Rjkv37a2/RyItjpAe7XlLgWiGDw4D/VInutTTzaTZs5873r1wyEhSJBuYASbYX
5cMtWiZyTts8mlQwZpB2BF97dB0vOyN39zzuGWu2+3CGfZkoafkfOrvW2YPfgxxd
7zDZNvAZj4uuh8u3jwIkKO+r5Va7Zv6VPeubFpjMQZAg92yzxvqmm44s0046FKgD
Kl4zC6lhyhmd2SOLvbxOx6I9AM45nPXMIytIL4Xo+ksQrIXnhHYx+iMYS9xGHLDB
lU1DCZLwpxmOAKUzkb0sW1lgZU8cwvEgUcsi4LvMynN4Y50mn/Haj5VyyAIsR+5U
MF87vLdY0jPb/c9TzGdmcZ6eDWzW5y33UVB5CiCimcJDlA9+XfNP6xW0UsC0CDUn
13RalVp+1GNjcR7JXwEx1c6eJMFoqFDyT20Ge7oeSrGCkbcVMxmREUOdkxnKRkcM
4pslUMLB2cI0lM8jRhdXuGoCRNG9vT80+n3faiNaZAMtcBb8UgtHE2PJjQOc3Ufc
T+HIFQO0QXXZkNuXpyNSCyfCaa7ITFtY2S0I8lbBJgwooLWKix41Eh/gj65kwJg9
7oj0zqvznD121+6kttdZRbXlHkrxZC4QvreOmtBZtyfasLIcNu86x8y6Wc0e7ceb
6FWSy914/XyC1WI0XN3qUGCI2lrMDWAEqbFeMZZJsfIJ+Az/20JL8nC1T1oJe0Cs
kBhmgkjm8IwqdKxcPFx8Wte59Na9+T90aGLBTibcTn0073mysU/Y5FEF1bWVf8+M
wgfpKyw6QA7YyxT6i8BIwfaoNW3IRJzkj97X0gYi/D44xxJAg2mIgTg6NAH+oG/v
hsvD2iX2VOdccZvBwKIzMYGIin3LeuyaW504wNZS7ysgGeyVox1MMEfOy5UJHaKK
LcIjCYfMLauvjSFuMiwjetTNnkF/IS5FaIfI/HaQNsiALlMS1VLeRp9LfPzSVLZf
l97x61mYra24jqq6EPAwNPlR2Im1PjDwHCxK30//aEqt1kKi1c78unY4+nmJhiET
poH6GiXwLKJ/zbLoCZmGkuZfXROlT0h8+C8AbOta/ZEkGzwNhyKKgOsOMjtBg54M
/kGZPZ76fOw2rR/XDOEiqTA6lLI0rc1f7B/9Ix8ytTlUJvqdojYEbCO9/NM/HdEw
LSmwfxEjUrk3+UC9ThHzrK98gyuqiS++0AQCbzAhOMXqtowLZ1IJnJZXSOsbU99D
K5uGK8dTwhOY3JEHJGwVGOF7puNe3sz2fbo4eTuZzjLSjQndL6pmU8F6dm1X65eZ
B9yvoL7mEGUEOQWL95jy8ZhfoxsWIv36rKG7LlfpRM1uRGGFSWVB+0gzFdLQHf5J
0bMm4XFugCIL1ZGYzZErkfZZd5HynqrVxGpm0sgHuuE4HXxye0KEeuLn19JCNMF4
2BLtpfg/eUg5Un8Ytd9Gd773rJbKCz3iQMnQbjySHcykYAsntnNnziX8bBN930L1
2dNWC8VVoPXnsAXa/2Zj2zjZAVVVkNEsKtK87vYtlxmUZFQsayauspZcfEBIs28j
UtZemyw4oBAuiarUJeqSrLSDIULPBWd9bqIDT10W8obOFn8peQ4GrclQ/pN2egdK
AN7Z2wcIszY+wH0gUjOq3USZPcrRnWg9TR0A8C7+SCovj8Q1ZS8nx5AgXZCtwLpQ
bvwG5LdHF7Ujyai6VyvT4cS3/Ao4ZNrsP0ebgQMKL3uCLAfmgfT8tQ6D3Bfzg2iX
kNtsg7sE0BbmSrbMVW1yQcl9RIpl4iwXDD1ZEdrN5dvcVo0XC3RNJH66A7fqCSFm
Z7F3KswC6O17rdFnhu3giyffvWH0yrQWTY1vWP0Wy0jNnzbU6GIxHLX4jnwDWYOE
heZAese1ApPj+o3N3dlXfi1aBErYmXyUQXESXPqz9fXPrGAecwE/UNnCw30wqhuQ
9H/cmbVuKVLpCgQTy5Rap6oUdbwe1uLdH8OefFDP/j1VmuSP0BbfcJin8tbb2X+J
rNErsrkco9/JhqZBsgxag9WM+l8c4MOz135jJmKvIRIrg5Vqx149MCXQZ02Na73q
kbujH8r+/TQvcOYnZKcMMfRJiEPZQruPDXawQXi9e0Fx1Hp/A+j4Yf8PUHMEazAM
LYeuFzudlBxmCYKr1Du+B+NNR+kx0Rjf4qnQ8y5tW1xonxKRfns/eLuoSO4zwhyy
6nTgDWmGWes3zQpnAKPuief45l34VRZR0VqxwJdnZD5Ay9zJRzUPgE4zQW6L4o18
Ue5bGuze+zEQBAWCNDZtsCj48hSp3cRLh0TJV583oPySwFt44siaWiHVVifHo098
fOdD5avsoGOGjZOpMAgCCpOsH+8IFE4V0EvMWqewO1sgtoEwjvNv/6ce7qLrunLF
3+sZnGe8rO38li8TD8raXNT4XtolO5jQ07yS+NhYhqc2YRHmVdYy5HexasPqUOoV
KqqoQnM1L5Xd+A75kur+lNw1Dj8pfgydK98x3MTNvK1PQLD5xHPl9c25pKBNjVXc
NsErCzzw6j/WFoiS+Pg2QdsQF2UvNZ3gVfOa0r+zCR3wdIrYc/taKvGZdqg2ETnQ
LQAiDowYJjxjdbOYhvcLJjfeVxnvBtpj+TMNml2S0kIRtpr4V0Dux1my+hKeK5Qp
rldeO1FixhSTqWExLq4tRwMIOePgciz9I7mnYOqnz/nS/6cMEzL050Rp5yfeWkAK
tuDJ6+KefRjDeO/3Fw77BPMuLhsed7h0Eho1VlPJOmqm8ebQ8Az0EAezJr0vY/4X
dZfaN4Dq4Tt6G2hHwoIOBZpuy2tql4RfNQLqddT7GPi7qcDUNDWV1n2JiPGpSKc6
600Bj++7G/dT8hhyAMRhjs1wpcU+uhVI0U/e27QylwlyuqBsP5UzpD4zkBXrvVge
+ia8+FBE14vb4ZHpZY+8wMCXwuj+YI7yWotyWVtIC++VfWR41PoC8x6VYFLw9h1b
mTyACgJyqiIU8i7g0H5IpYA2rmr91giRZ1Pfx2MZTN8WYXFgxZbjY0lJJP6Wxi/x
dVhb/0Jql0VcaEMDMXpvPqce1ZgaVwkjNxWvJ/TnPufFNgqdxuZbgKYqZg5I0eic
97QKdfdvuO3FKXJZdgTVEL7Ke2dFkrizpV4IKKluz0oHem/gpNHyifhfyEcRQ1bF
WsLIn1QyTdrvhFPhTsZjirPXV81tCpwX5Wnhw/T2zp2+1bx/vcYh61WTAh1LUSeM
sLcA7yj6UjQD2H+KHhxMbTOexjUJ7Mj0zE+qxIsNqRoTAtiEJkioRJcLMwZP9fhv
e6y34gNSAZTDydZVhXxrcN0Z485WJPQJN6UdyYitMnNXjibMGVCT7pdwbyx4IOig
0oDadbtrYiyZZnGBbTsBzC6RBx0KQ3nHwCisWcJn/AILLzHucPVTiJjQXYTx8T2J
qzgaV9XAtkYuv/+S18HoEze86JDVH0knQdAdcSP2ppl83E/Jn1UNZFlzrSodnJ9M
tMoGPKbw5hSBmJZETVsanBdeI1EeJl4skKu9wKgSY3hG6xVWJg4NU8va6sg377Cu
FO6VYdjZzZDon2UIN9xBkn6rroYAiDjnfj3J4oAP785IO6vKOxw2EWLjTIGqycVn
Atb6l02HF8rOh96QUEFYHzEyh0BIWlwvJq2MxcTEmcLTq+p2VPJzWcwFpF5t9wNa
2y0AbRFY51H3SYPscLMDxI2MKC2yS7PN+83Vd1gKDK5Ra/fxOezmP+OXh1QH2VXR
wsPHLkuSGN/1McfynYUghO6AJMp4zyIxcBUWGG4eEPMq97Osrv0DCDKUaWaM5gz5
r1aFK+Vtpv3WcKfPWHRiK+vBE/8ZClCVj/aPJDM0MWIOEIX3yqP+TRHRgS0raRuE
h/i22NETi+/WjDW0meCMSg8uGHcX8kEvDyFehtezyvmBsWuy4wKMACZ9pOqo2faF
9ouYn93vThVKGnThmuyWWFW5eCYtxOc1U/mGys90IkrpFRQXCuE8C9483mJwmtiP
z5Gh248Gra975tWFexNoJhiv+nnrDQ6QSWrVS1vCouf5UN037GkiLmK/LfrsqOoN
KBUp3kLY7AKnJMx+lv33ndEZggDoIJ7GPs5J/z1TTSr0ZEKvuVKd5S3LQrBGlgaL
F9HZ3mgF55csc6797ZXwimnaB+WizBbUy12TgQWXMJdtRWJcUSUAzpzk3nXJXKdc
/0KaDfX2cQs0EoxIgaRYfFiygEu3fdcWvV3L01EXBmWQvpPLEBA1G/ICVu1W39po
ROo4Lc3B/DAt8qG2uZ4GG58yBeImsSCudpVvLaAGWMxmBOPQwH8KorK34FEVVl7/
V1H9gFLavkJEJuP+0l0+j1Z+Vy676W9dCE+h4LokC5t8rsAGnMDrr8wdJzbD7lvK
YuI3DJE7dCgblSUcyw9PpTuW1Gj98VmbZ8noxppuFnQRQjtB5deuAasGiPYoD+qp
gewCXKbLMc+tXCKaY8eJilqR9vJhH6GsJSPxZ6EFPcNYrdQXjnFJUlKT2a5pwv+D
9w6jL0OafSbRcCjnJZJ4BpUTU7DdbisOJFPvcNK6WlMJbdIgJRTt6TFaOmWSMNSR
+vV/CE6FSZek96SrCa9Py119yH0fPWi564ySMReTx/XMFZyaFgx9rv+F/Yr26GL8
PfFSm5ZUMd3GL6PrRG76rpj/P2vaNesAOqob1u/+Eg+kMgZeXC5br05AtfI/PhsR
XnNkalsRbvQrd0RNYm1dRzWmyjD49xCwFg/el5aAfYe56f7zHMuw/iIwlM3A//WF
zGvt41GOw9MRdDcVBqJgUJJYtzxWrlJpJEcZ9+zooGh198J56BisJb2H0GnePrC6
1/py/GSo34vVVg7QOCGECfZcU4Cozx3dIkl94H7nGsKIrPg1ZN92xxB79DuDk6gl
1Oh3GUQG1hKvfRQmmEIY1K+GIPPsJOoPZRrrwLUYtGoZnuQhxuWAFlTSJxR37AMC
85blACTagYCDjjx7zggIhL8ATM/d3EfLe4L/q2bXRFi8QHVyIA4hPHUsOQGnvge7
DGHuQwpCjQk7qJDOV1mNl3ioXis0YO5IXDhUQlJCaEIQRrfXYpFNUCB2TtLRJaaq
WbzcYthFN2H0WQOpszmBueY/rNFYcnmrUkWYPMr58c7oTrT9hn8FEbHB/zPe+A+q
/S6tfepee4CE2kX8gOZ5olfHjhufJQHFvUFIBNh+bsWlAIqfvuV56xhqB4QD+wYh
mxtSVvjI1KAGBAOTj0dD9U4wzJc+P1/xriLMi5zD1Hc8PsAosi4UVQeD5Ngp0pjB
WviipIZJ9OXd6d12Z0gjPIzufBL9mcISZRKGW5W9qEYMULKrSOk15MV1tUWlEntz
WwFBg2xZU6wdgWWR9FhIWvViSgKuLplirWeYxqVwBpYLUJcSeM7CO+AkwW58k3a8
nMgn01bf9MMjF7Ub8/8mXNI0f9V15wSBmNtF4wnBZJRY4LuYEOc82D8i8uKggG22
Uhx6jFLgzzRvMKEBEt95V7x6He700qdGjI8Gnwp1fS8s1TnYVqFFZGYBxVVYnBkM
rcq8z17kYbn1gZ63VLu7k2UxmocNb4KmpUbQmvp/yDOvExDSZpEfPR2Tz+mWJ66A
Fpd45Q+jTAMpefWMx24XvrIJs9RRJh9LPsllbdYXYCsYtnNXbjeUWSurW4khTRv6
NyzGw20+aUNUxyrj1PUBZRk4P2aNeGPRsmbSitVgcycPuMyPmLhC0owg3nXiF4Ph
NzfI+fvzw+nRP+TD22nFN+4sMYjcRdiJqnqM/MagNKjWJlzbJ3f3jwlbSZcQ7Wjj
l8KHN0q/z6J+zwD1XzwIvBvf2l2jnbSftRbVpXQpJUxbhpm2BqspyH7ZTyxUlpet
ILoMho51tY4ecldJZOcN8pw+DzH9TxpWhrxn5Wfu4Logpmrylqs3HVhjCKtmNE0O
AhjAzYrYON5N6LXWHdXHJ+7sAo23JTDQZHRUuR4X7t0nOsUA04HnuQcCwYJorSF+
PJ4ssBrGWDWAJ0ESC+iNryUYibjyh4VeyMWuo3/jEy1qeDyrbBU8y6LV8IW3zT0V
YbghEhK60+CGwnOiKEl6zqeDhD39iYkA5ezuIqXlddkfjj6Z0YTNcnxrLQS5/mat
svifWA/A0IDfyLg7m0wdgzP/G72Q0rymScbZidCVHPPVSaJLvWZOLZkXve2c2m6R
zy3U9lSI1KJTp5YV3N38Be3nktpy33+7jTVDXk7CjuEhgXMdozMGTZZg95Mrxxph
WvB2EiimhTaohcA4RABeKoxspUjhm1HVR1bUklYoZga0Ewa6RYgT2e5GX8c1AQvi
btbCaKWqpc8s8aLIZ8qioKJDKxDxNJ1C14DY9Zcomctuj3rzk6uXGUQw3Tjb0Kwx
Ackufe76sdIKISDtwDuItCIUfN2tcAPhCONEGRbwQtNSmukjpiP+I8PGJXSpmq/z
tD4DWYRjoVgpLk1bKxEMYLTefDjJ/k3Ig0uQ6F87c98neEjxngahA6e+GkzUzHeW
AZpI5vJ+/8S3HMRoo6yqk/L5uf+C9uELD3ZS4Z7UMzaHxuUPHTUi35HOAI6j8ghn
qvXSFxN9ZW4xGU991fgr0/xPGCuXreIJhGvSniZtfEim8wv4e2KHyKSm0WqQcKR0
2J4x6GAM5v0jtbW3X9X9SJRLeucwsQ1pEYIWBS9AsDEVG0fZ4y2YOiJ/byXw8GZo
ezToU7bVF0K99uPFMbt+ONGdqitCI2tk9ewGt38jMVw02ecpVwyM76nLz1R6IVKO
g6T3T8wAEKM5dF87T/o7jte2gzRHzvOy9QbWEs83OW+Dy2zR+jt3swU19y0sbPQ7
ox9J5gT8LVwJJ+xbqZfe6DFq+AFz2QsPRNLzseSlvpxKPne5bZM5yjIiitb6AWSh
iu/PRMcW8kxjcX7f7rIWU4bkVh0eCgGKcdE6RTsxv3MTApKkS9WGPl7lgNE0mbFL
RF2706ZV0hNBisEc2dJ4NCSQYNpzUUz6VI7mYupupu02Kjg/O7FAexsr4lYKQWRo
FABCZh700ByWcupgc11W54jg6tFW01FTB7fJ46IwiAS7UOVXjZfINlqXTFGa3Xxt
0nBzmr2zQbykbl4cTmJ8x0WQ4MdHaL0J+6ZTFfqMoipIiT68io66iraJqk0wOG33
bO3v2wrEwLOJ/0UpVnRzvWveiZQC4qR3BcJxmoHqHab9fOxkRqVZ318meiFU99t6
1cVdOU3xWfPX9xm624XskUokJ00vsFfDaDFqfroL+7NC0nTeInIj1QjbyOhfHtEV
t7zO1to1u+wiQOXiTFCdDOF8hsgTSkMSQqh4fH6rzCdJNN8gJNja3VNaKnIAYd5V
5GG9YNYPRN4C5bRcaWIsTxLIwgwhQ1qLg8xCAlftnOjLpaPPqDRE68Z8lcogx4XE
P60CgleonFuBXk0sJ2Fu7QEiKvnYpD5s5ZYbyzsYVNgDrQhemOFn2As7JaWFtkYR
w1AvrtWrzkkuJM5jKksTGwLxKhLB9htKPalniyP6v71TNF0oEIkO0MeBnI9hHBZa
KuJpRyiXFKFv7WyMAbV0GLBz5CM/yHNQKjiB883a1xKNNlfOUozLyEcvFzldV0F+
I5TDgLzV9tWAT/PCbdw14M4FPMBpEzX/bOFnH731OGz3KabL+zWRttkO/mxucZeN
1uqNfH0bfHZBa4QYyYkF93typSqCWeiVc8l+NMpENTLphNjWVIDhfJu6FQyeuO/3
YnMiLi+rZkOWwJIUmMdffjJntck5h4Hk+kiiR/W6GjpJZPEL0bSLIF/5OoDFBBR8
4lut13qs29jb+IR+10UUzkzKDEJTX4o/eAQnq0QbKP5YHwgCkTs6nkGWnOfyXF4j
ZUxFvXcYNyDnPlnKfavyewA/JGb+5YRU8wKJx5yG9pV+KcLk8eN/q+6FwGxL49BJ
wHC0IIkBQzovlD6IaBlH/MSlpFd0t4EwYc5Klaz7aXD3MPm7fX7F/40Zunt+VzGa
BlnMMLgWh6KR1V/i4Hqxxo50pplra1XRwwrpQ6T3zQNC9Fm8RMaYz/eBfYUW3FLU
ozwqLL2H/BxXsxEQKdZCOc8jlmSz7N5QfkLITryOOzhQArWXHXe4BWa6+01tHalh
+tK2WAFKqLXrdyRzzh27koL4l/eirrJ6nXNIe2D5dPEYI9dDe7ZJpI7wk7YUXLtN
+W/+cD/gC0QuV9LsEzY7EzEFLWXQNR/KjZYbYsPK4Cn/HQExvIYQFl0q36iSScdL
/Xot0ktzWHi/2F/a6UUCw7ND1+DHPi5uH5e1YYeVsyExGgZboFcZR2uSJA1CAAA2
D5bpjCpLT1oI/MQxjyyvbpnYBpBPYIsvSLBxbPPULurx0KY9trs6D61kX4+nUI1S
ggubuzyPebVO2Ld4Lt01V1UbN4mes0hyRYeldVD622cYZst9C2Y2qoVpqwm3GRHQ
lQgFy2U1+AmIN0TxGjFCccz3BDQyFhQmASiccf2e7yb3RvWI/W3mI6OB9EUB3aPV
D02s5FNvgK8Hc2k801dCaJjLgrdH8xi0vl1fnm62xaMiXJ0P17fjfS8ozrldLPMs
qUydFf5mQT7WL1R31Yr0Zok5jdkAaGvCA09QBb8imlouk0uEQ0ZqE1SBXA4ISwo+
H007qY1wiQJnoqmdxRJfJP4eVDwhzsENuEPeeuDHryrVSxf3to6HiBams1rahhTW
NUC0/uabSs3i2rmCdBIGd01bKS4GkfJU8atZZ9GKq+9Ef2ylbw/jTyVg/vtJwRLK
dvHULS68O8nVM7QVEy7zIFYE62YXSNonCNY7A7LzqeWFAwHl7MyiNwuYjhloKnaA
By/72AAf0dS0rPetRqMWqHDVmeiWydDfmdzwF1aTbr/7JY02/zqWqMQ6JGsbbtZW
8sAMxc+IK/JWuq4tx+iMrh+ftuuXHL1Gzaxk/BakbLe1I3HwMyRdBI/2Fa8P2Zpk
GlV+adiS9zAVzG/mLHFAhz+aBYeT6Uuzu3jeSbkPOJdBWjcmobnbG9nvurD9NQa+
ET2IF3lJUQNbeF64/rP+p093RXxoLJ2qplZ+vdMxsOe0NIBidSJrBfkXlFoXKNkI
oLPUqWRro3aQ3j9VhdKSO0liHRTF40+J5nK7yuoXFCkuznmTgd2L19DY//2Ovj/A
BY+AhlZyjGZaUf/VMXWNFj7GW27PKmV69UHliBOEh6lpg6g6YF4AzmWZ/jO/ajjX
sgSOwxdl4dpRltNEvS0uHy44EPomRbMdsoTXlGCpyL4ezWH0Su2Y0y+FsTG9CTI/
RaU8SEs1vWN67fei8mNvZW0DoPl8gaEks4pAjQAXJelgTBdy5VKXx0Kg1G12yT/s
lP/p/MCM7QuW5WrAawWCoTDFMARAyW3kgsNP1wEpfTXiVVT3RQw0C4o2dvSo3uIv
r7UQALdTR9cSmzgbNNbhm1DKz6d8bRmwZKPa63Y4NSzWZm/+0zPFTZy3vVs1+Ulo
j4N36eeWkn8iuyd2BuESr91jP49S5ipBnWHREPAsAPf4SETDuFjcq7HkSljNGJwV
kUhUg56QiLZFQSITflU8B51MvClZXAL8Ww4tF/RfB8M0ncYXS6vH78wiU+Owl4lt
Lh913VPLCFiQKP2m7IrpN3FbYiBtvMURvU1ptiDWBymtjZwK0UjrFWz+DUZI+cJz
kWwbeD1aNzyyp0sJ4aF+7H4KLCKQsOPs6zbrGzcrGyazTMqfbXlhzqk6UzGRGnZR
Lx52bhwcInvpoOSCnX/mF9d3oKEYP9TKfbf/hx/mX3JqmB1ZEucG9ghJVB4PZNAj
ekKA8B3WiYNZxCnBvR55fJOE27K/aoTnhutR0SqcIfQ+RprCGGwRofOsnvItdYLI
P9vZluqv7eGTnJVsPy2x7y+J+7TTTzHIkZ8J8O2UZ9LizPo6Ob+rzs1qey5bT95w
rZHNPo0fkTgCVZsEkUOsK6unvR2IN9IJ8KfvG97UBDJNOQ9LvJVi+7QSVEZTyHfO
0bVAznnWQdYUkmZVn1eoPxQ0X1p1blacGYPvESvgpVF6PNKZaO+dZFPYghMB5869
ZNLS8cWD+JUy8XI9z2JKyceTz+FS7Icppe+ALG1tVOR4rIhx3Ib3R+2uN0fYcRmm
keLRa4cAcbZrSsMqIoBXUqOh9kjHiqbSuLLRum1C/14frmeT+oAQbqNBaXLewvfi
w/SoHjJZ5n0d259Fk/fCPoR0DKrzQEGj8CdHGN8GMuVdI3JI6ZtAHN6WOTZCb9rR
9KTU3wrho+OSWHzZMP6mB+9didBts+KHjg1fViEDPu8NPEXDtOTuYJt+X++WedOV
y/ba4HC3KuzONgYnIWNiPF/OKuOKXeWvvr+MNUkToxj9RGt/SEXWi1aDRLWKr1KU
1BLP8cBJZmpxwQjvs6oqbt4UBYbTO8NY6y/hiI347jHKZqMztCGGTeLdo4gDW9ST
XxlknFrWdX9i06Lv7vP+VDLMB3GhbXhFyqNKXa6/Szs8c+HM5d3TGiQGVEfGkJHV
VpLK0FYmmngmKOfB6mYJFQKz3lyfpQCikkJDLfU+PEtTwKze8fyw9qaH30yYTw/u
9vJp/PSSRoUJ+V5ejE0RJLBFQqAdMO9mAhBvbu9YBCBvSiAlpw7foDmEaIesMlI7
syXKMLljrc/kTa1E0M4sMKEEML2z6XPxoxf3NsnbmNy02TlYbzfr0X+BMGw9UXHH
pUQOE5MXbG9MMygSRXGQOqKJxA3nuTDAQSUvgwqpdaok+iKMUVrxDM4580TZS7Ds
n+B9KKkNWPLx2kFWaWaLOYYQEGpyJCXjKUQ+6YEOobG49hYMydHkGsfOri/LIesB
5JDy5fuQa8bvHuTsHL/ztR56gjOBnymt4tFo8A4uQ8QK0ObQEU51U9OJpqrnE2av
huuJj2O0uykxG9AIinLfspTSq+5AMzSZP9rdLnEv5eCYodTcIA7C9qptxF/CoXCx
eBpjnEMolLe3ykCzGX15aydiRgRk5YS5C2CnTM7p3hXg9aRCkgoes+WKzHb+v5Tl
5O0y/tLOU9XrILBD4LbnL/6lc5GAgejhcAHtCpP1reEfwq796TeVTA76bEcJ2PlU
cJMLffbvIAyJIhy3+RTmkim7tEAHI5PSDjxD9x/tamD1DENmcqzWh0xtcK4Jkl7e
L5IxjPvZFTzJ1MO+zD+oPZEjZMstThuJ4f3tVGUybgR1LSmBoH7nAVHHOin6GyE1
Kysa/9q8UIBRoGQmOm4GYW0vfhOD3eG6tzNhqdLCeuZON9nx5g0fXv1iXhkbTYfk
Rr3Xx3aXkbkWpUfDwfuPS1YcDNgoNb2ZGdp+5elzo5aroMcdowLzX7wLDcD6Wj2o
6j+e97MIWWunEnbfJXrGV2KJi3bpytkjR/LIGmputLDLRjP31qYEvBQJhB0DrMqg
7la52f9XzcbIjpIwdwQGFLiAM1dN8Qc2axuq6CEutbqilv+Ack1dZ0tFTV/et7UW
y1uzVDa4cLt/gE9bm6uup9gKH55ORqT1Y50EpCkm1EBD2wauMfXO3iPuWPjW3Ggr
rA0Uppks9t+twTHAFdN3pi0PWffv+HpHNX2PMjRuE5hh2O8SjE+WWOWkOMn40BjT
XzdCWOiLbv8mpZD2lFPfjBdOhVVZr+RYYnWTGTpbm+Ke9YjIJHNXeRg+WVJk+HjY
f05pNgBxOjsFg7l3WQ1Cgz213h4terXfS+c2l0JMgH1cKJqBaey2X+as9ZLNI8lR
KuKlAd+yUvTrZQUkR/O5INQlzHPsULAWAJX21iKsFsJi+D5YnOVNBu5bc+ibx7dO
bBdlgZCxWz70MXXMXHYUJEqr4EV1jpNf6vp8DJhMNmBnKXOBEtvgl0I6QW61BTwk
uv2LGoq99kll+7oO8d/t2Edx8IESwGr7Uo6IPvvI2+VCBS3P+gMYim+HITBsEBCD
o3TVlKk8WkFZVCeFVqBFBX9IBAPD3JxweNmH8L2JL94HbHpn+abbBqgbAqGhRlt0
FjjeOM1tiP2nYAaW6QODEhq4pF+R02DSRnr0NtwFLL7iTd7nTaXwyoGBjB+ZoHtW
/kbaIg3hx/2OgRJ7plAShqBbbq7S8e6eFJn9VcLZwx3b7TBgB16kro9U6zilTUar
9/KdfogrO/nA+Vlu306XfPkASBbSM35dVSO/ZIE9np2BMxLSUfJ2UwJ2dXRvaNbf
rRXIKTYeFCjTmiJHn80ReUbijIWRU1PtAWE1nHJnCkf2EMUnSBEzTxi08GW2eaKZ
diSzG4u62U4acB2yj2EG8xFuMM2EJ+KzHlPPVlePhl2rURwPJmsHnlnYLHGEZilm
69AMg4vGqfEK24LVp+hd8kBeiZ92yx4kzXedtOPFAZXh3ce3+Np7cTtr9ZMCj4yt
isOSYGeurKwqVuhTvEyifbrnDRoaqcalcPWFezWhjshGedeX/jiAJuro4+bGY0mh
aqfjQSOvIelPdQTJ7FISVs4o4SBcQHctMtHNX6lZuhYtlIS9BOadPIU6xp9h9xQ+
LnDUY7iGgyFu1Cr0ThOJvy6TIX2kCpesIhmv/BpbMZ0I0XKWaTpEj4wCNkJlFNFQ
HmlFt5xoSB3UXzpw1WkOirBMLngvL1HzB0xGojIWXIQnoliD/0gwOcICQKEWeF/V
RQ5n52TyibtP85t4H2Qt2ulTgPVqW5b3k78FJn4ikhchPbq/GYbVKl9cpt09mryr
p+lLRxTkNhNYgdYq0QUFbR2FT7OxT9BNdpoWL5KOjZiJsBmqrxYEffCSlU2fA6bY
vqCw6FswrTgcgxfvzbHmcVSpw3uYIsQ+mznykMQuFs5igT22W8BXRv1J/suiA75h
1OcNb20kXWfhQMDI9fuNkMW9zdapzzXeWaemLRjfj+T1Hk7mOZzZ11gKll/v5Vb/
k5ZhFl9prdoiTcMvIPh+hF7ZnNDbBvP7c+D9VGw5aIkDOXj0ZM40hwjjS7y50h1+
6146zUbs8FCnSTCijuJCrzPP878fn0JB7S80dPzNf2bd0lkZG7qfsF+jzbMxikb6
RYi5CSFUUXAqgO7qwOvCga2n66sTlGUvl9U4TXNEsxCcwDpftoDhkEulhWmAkqpK
uwX69GueUGV+sU7+/WAfjUx8D5qkZuI8GccbgyBRe6tzT7vIDZiFYuHnYqsXFdJg
eW9MCXc1lP/opBE4U15FepQZLWOsms/8BZ9mZsHMSrcFE2G1cQg1DvZu/aCtTqu+
zI53q02MhkqwyJU/XPsD6JyoY4uKiXnlDcPZ0WtSv7c4GRQWziDVxPVZh7xNA6hr
oNal2SSHVvNWBQC6rSU4iEJMjUSa5bwytm3qDpSku5icK9Ipi25f+wMveJ9Bt/Vy
ETyUFLzlcEo+JlyyxAhP0bnp2QTInWTSul41ZaAi0hvSCi2Xwws6rsYYXX/crHdI
ACxcsIq2oI4/LoH/yAslKCqN2TE1QiIPrCSvKqzbdKgjoFlaDZaHeaeKHAt+uoLO
ueBB0fQpFXXlz6XvRRkZ7Vz0X2bv19/nvh3vX0hj4eUmC5cdODBbTQzsVjtM0meD
AymF+cJ9uy1KtKNF/mY8woxuCN9hIDWgs5agA1LY+GXNC+jQiQmo0ykaueM0Lov0
/V+c7dBze0o9MScNw1Tq7Wd/YWjzxj0t0w6XakLyezsoGTt7CXtzDqhsCIXW/07w
TJRLXkSeDfxKufhKiawkDUOOVKJSGU0VhBT0Uepz9bWbqLDC57CyYIOe3T3s1MQl
tXJDYmITHSUmuf2/TInh4xNyKkBYccOiUaKO4hXHnPdOtbCMXR4gJYdn0paUQRnP
sYuFm/axAfPaDEcRq4TTBS5JSN0wttW0rQnZAaQ4k66o8nB51FftBRdcZuXm1rib
41FiELBCYJDwgxRQva9hJZNlmBAw2OlQAsuCFB47G3hUknHjmINxWOi6JeB+v6ZW
5NPhz84wE6eHkAfWB4GnEY+85wKic7wv9QeedxFhe5gtVTac7uF6ibN6FW+PBhNJ
tmiyS2b2hlc/28aR/VBae9BiJc49MAN5jwddMip2CblIzh1cdP2CzfE3JA9i5STb
Uwnx8IikkvTW8i7vpdb+g5mmpbA3h23FCsvIE3RW5mJW8JXSe8caNqAgK3gQPD5s
L19ho9vEnSTI6ZPyaRTdVlrzD8zampnjdjOFsKdUFq5OrtdZRKukklJIxHi/CUPN
gn6g39YPmrakQmZqYsbWs5+194LygDgT1jaCNyXS1vD67t+IuGBJHmYzeUwvz6HT
i4RFsjY5O8RjZsQfto7/nCbuITN5qYrItv7KWhyTybyACM0/An3lS0SHPGE0X9Zz
4Jj4vdPJC392BYCiPXAckd+xJYB6H/40BsZFIrT3vaCjFDy4zOYBV+JQ4AeD+XAK
pFZg7yo6WSTXK3cmxxqgSiukW9HzlTYIvwRaa/arhSIaanYAr8AivsaRCuPnwST0
jZ6vzlTRyVq8efsQDm3FHGDr0bkf3+adeGBU2McIR73RjfpFtXR4TyNjlEImvFP5
AisF2BYqBx5x3fkOg2jJ7hOrEw9mROHeIjH+4ioqqhbhD2wp0xYQyOkUI08Zog3C
o6HRrSXPmfmPVM76QvMZ4MuLwPb5k4OXoExZnBTpnaPS/McTqpW6M2+daXi2PAA8
0wQA/+TLIKiclEOZkfKd6EmCegAPErJ47SMOLth4IDvZtjTOPiBv10HTxeZGACiI
DC+h2TuhpOzbhRWS9ImiLBEfjX4XTWO6Q2BCxoQBRVt7N4TmZqDTfPEtIOB6Zi3s
zo9kodFOimvc3Y+GznExJ3Buhezt2WJQ5I0/C8w2pPOBK7AXDC3Gn9UnnMiYn8M3
pnsMVXsYtsn+rSqV9ucjbBCSqzaWWb4gDYYOCD4LMvBwsiE/VQWwLLHya99SG4pW
3dGMtPYpv7C46HPOrtTt4XEPPEpJnrqlEC1U37DT99Sqo5ADaFvyKeXVkzjkHKcV
j8BarkG1cAk/+kn6J/6Xq8VwsPhYsWFcrhaPqNTeHnc+8DT0eDGLQ+73AyHXWeE1
qb4P6JGDWLO2s0fq1PxaBI5+G0rZ/h1Fmsul+JsXLgIteZMT/SboEtU+iEX8nLt/
CcB9e3Uyi8mxMI5L6uLleenxXntHH1AqGuLpBO0hYEN/Vu8B1jJctTouNPY1R5cJ
wpyB5aldr3BlC+OTrR5eUs9AYShAutzCZ41wUPr+oDxBaVzEw+65T8dv6pJkHVAv
rAPLyixFI4XV1lMUvdLwHUpqIE0R8yGsDyOLrXEXvrmy7Nq+qkHxThoq1Hx+1MFT
BFOmXsKbx0lY9ibxSosH7yL/bGV/H2nAF7h+1FFooRku1A1L0oouUi+jX5UizVJM
ldHty9Awk9QLw/KTccOlRMxr0SDuZumKG6tSuEQWSpriaAESa4urfkK66plFEEtr
3i3VUFvqBFe/e48LG5Aul10JGbUyNkEI/AyI2V1fGcq12z1VZL/r7+7rarfb71yM
m/1BWGgMnB8ZyP1KWBvvldjfx1l0vNBon6VKLKZmwkGP95cixdv9WsbpS+8jUA1B
FPvwl50e0mtK4ogpy9aAE2iwm5CGaHgWF6f9BEHb9/T+YYK/UjOJVukgwTcBxddY
dnKwbbCUiDoB2scQKxXE542m2ZwbB8p4T0sDOKoH+ZbsV75HqCYM/9HXV7a8RKsC
Yj4IohhhFkZMF88I+qlVqHbRMBcb0/zOZNtR8TxhcA9Oyl+zyA+59p2ev38urEDu
aIqO7Mt+pBLiCJpyhoEuzA5k4GcQyejgpvI+0UMC7JPIgQtTS/QpnogDyFgojLvn
VhLxFVLfR0pYX6ieNbn6TIGBUC6qzP0VyJMAKHsSK+9z85JLlBTrYRoXuKRLtnJk
LFWHlhezvk1kRK7eaZWBikHUoU1SSxoP/lswdxc6cOEQ5U9AEXtNMrSpMB56NZbs
OQPGsRWgxQTUbX7HZ7lGbPjZCURJj9NK/HTyaH+aErT1Dt9tH+djM4FB54Hiu3aS
0A1NAyuTeMnJNVtw09Uj8xJN4vYWyJ4VQ0jI4SyGD52MXMogMc85yDGsGmipbXT9
RQCKpy/SPVo89qiKQf1k10cDJ6Q79dtmjBkW8kjV76WhvdxwumnKn9omptCp2yC/
5edSM41m8ssIXGL0L9zcuFEkOJlGP5bxBlIG06JtSBE7Fow0Ht6+qO9E5mgE4LO8
TeCCW5fDgLbHZPuRQvWQN5Fl7OMp9O31QX9/kBrd/kKxiRS0RqdWg8ZjGjAvumXu
Iwzq6UIxC0viAU02pPsM95QKy3Esr67WiOkLJ9ZxmTRO9HCf+HxEmhL10Dz2gaQb
arpIXA2hcMJxGtHYO5MNQDVnAB000qJE1mj7M8xrl6PTLHqzsTeXrIdch5lAbhic
4tk+KpABtxFGDdilnwx4f5k99OAdQd0NRvHF5B3Y1GDKKRNSN1ogqCzTDPC1HyDA
K8CJ+RW0gfLtAVxMh3AR54Nsa0h2wG11b/gxALm9QX9Lfa9lN7glsSGWswt+xGTA
MbApQ5JcMMwJ8EMYsM04tq9nXZS//ItOuiLFAqurUtC1QVfraQhJint0NK4kp3em
Mwq4Dy5y2OZfnA5FiCGk0gDitL+TmPXG/Dv8dqMq+cSQsx+MR8KUtZRBUcKK+X8s
zLvjobDw7intzpPLt0NokoSfhKPhLBpeWR63hXkOH5PipTg2l7qfgJTcpsjGZLw9
r9JMnalubesHnRbKeZ4SKBkv07/O84KchzcxOS1UnCAtD1oM4jcsReCd+jyNMT0b
K69yVHFmoiJdh2b/D7T/ylv9kIqzQ6Fk5O6xm9HiUIliuweZxaamKI/pWZ/Oh9Xs
1oHvFOk+4I1ILmRWrYY/+LgrtkE3XI3VhkyqVRSCcPZ+8OpZwK6IWLmch97XjBQl
6eOeeO2jLK2nwUKcFxafqrLyRTv7++alxUUg8BtPXGw93k9lsEIlEFGBEerFfIUs
LXAEceZHWxu8ozvrYeTLhoCakSnJyRlq9ez3FRrk+muzznFr0h7A6e2lSqYLqHqE
mDol08MNzxRxv4+aamHgXtJ0IA7Vrm92yOijKSjzAb/Kf56q5pAIscZmH45h5tqr
tEdH6vBMK3ZWNhbV23TzSPhDreNCJ4c8jcfb4k6Z3zHGwKhZMRESSz2uJ7TeWCKK
8WXRv5oGS2t0fJJQlvFIjicX/LYHDz6BjNFpWQYgF9W1pZdqnavAUM8+tuQqeBcq
7CSciIbNZwd2wd8T+YxwVAdlgOCjwhA2KNzpMyj4M7CPHJMkb3PpIJFtzxIG8vZT
zOCrD38+TuYdChm2AaCqyBUmBWLahi1O5L71RwZOc+cxTKv31heqjzGrJUGrp7vA
rAel2Uy3Er/0337/0C/FgAkbwvfMXamMS3xAL0cCNXAG7dRRUFpVTnJNkqF3o9Gn
L8TZSj2gIGbyWEeHBT6PXUnJctBDkCKO5hQGe5REvpdlZKgbuF5Y/GdjlddvG5uA
wtzF31BMacPvjybxsEif5LcJH6IetDeuKBuBnur5ehW5BeoUOhyiIfHF97zbh8Ta
qAAJCcOy50aPFQlhE6ok0G156MVMO5A9YmX4NZW5qSsQjyaXAauZ8nB04bSczlse
AM2S7979ZEAqgKOXijW3FsQ5Bf/4Fev2jUwhFjt+4a/IIRjz8jrQVZNQVj5aapdL
HASAd17wr4MGI3NrYbhDOXb39Em3w3NQW0pAGvlKPxEPfagKRsW46vp8DQsE9L9P
LxblxMFIHlbA/zHJkwhHBcfAGj2+0ld/wc8bnkRW6uDImIH5QK8h+7XMdnzBUDgL
nBqaAJqgl5FKBKQoiA1xff4jciaSB7+rEqgsER6l3aVajn/5pevMN7RcP6SDOo91
3JA324vPluInRWa2lfG6UcfoXsLOl93T1xq6IL3us27UzCQ20p5sWJAPdtvDiruj
+vV+vEhIrDyMgFu12qZVDnxPjsuB+Nk+D6Nj+w7CmZ+eZ2cSv27WORV9ZzOPvKpl
JzzDVyoqPlggXU6pGyQZg17z4vwTLon2zP14MWS30HqKBhnVT+VQQvg8dyMypPjm
qlEVC2yNhCpRgL47Ub6XwVISHSxaekLVQTMKh3J0nuGKnNisbPQd+cHBl43LZvAE
sIaK0K3K2rT3HJC4f0H+P8mCLIuV4k+J1/WVdY9Xy7mqzS2nSDkw0TYI/MWAUXep
FYTvS184ycDUdbOmybEhr8HfgjfxllBp5OOWU63AdA/RTHA7Gn4BvNiILisG8xnf
MoBD6d31WaVQXjENkKSwAZILEr9Zs/XS1OASD1zWO20bVOSD29Ia0KWLjcg3guQ8
Xc3HDmPTDmbjGzjx8rrCVnaxuhKSqbnl2jy3D/KBQYnUiDa0729+SBAtrkS23sjj
n3FtqppkQiLn4wwmIAK02esDXw/xzUr4xzXRHVxnbZYJwGTu4BwhP39PEzb5AWIk
bHFvUCFP+53gE/fEyBAzLo0joW3pcGyELoIVtPjd95X6s9wFX/S012Fz3aRwdXJ4
x7wnE6o/g8xS8ovEv9hkD1HRN68XJs9PpjtfHN5N0KDLXg30y/Xi+Xspa0KI1cMx
w+85g+9oHLcZ50y28x67LQCc1lAbtyB3u4KoFVIL1T+HHS4bWjo17FWU22Sfv6/s
Abxygbz51B1nBkyTgc6C+ftBxDcqgr2mcXVXo3ePZM6U/r8VTtZxkz/etT/W8rKc
YmdlFgrsm4uLCARWxCFU+UXxgQ/qFs/3SbD+IXvPGsXhY7lez9qTpF5tPDuUHJz1
DAntU1fAgmwtJsygAR9YxeVLKSf8chttnhbLHnGd2tyeks+8t1+iOUmtkBIvff0Z
gWQmdTHcMxWwqivW0p/GTwrNuUd1HNzPV1jXZwTsfUMm+K7oj9EyHHihqLHw9piT
oSusDtObwofeChhgDLMpucLI1dvJy15ZhBZJOHKjdg8VxZ+loY6LpnWqRL5D0P0z
2ebgPOjavAHtRpc0vl3zSiGL5r1ttMgblOtOhoIU0lPCY9PVKcoM4ZD5t8vBDkYJ
Wr0VUr90Iisx3sLgt8vZmXAtNz9mePUa707YbBjgL8UEkCffdb8FRs98CQ/CKh5+
AGXPg4f7tFIu+K+9J+9gqPls907oeAE7VIs/aDkc7cBzWGg6YfXbOL7YbkAWxGlM
EiRFbd/FLIf8Bwck/fjDgeHRCOnOWn7LLZyg5fBPUmH5aQk+uxYHzqp4Y20KGvSR
adWO9gBNFWgXdSNRZvm37dWO9x+9Sh9Wr1bHaDQyOZRQZvupL9fg3zXp3a0+bh3z
PZsOA8tncLfEfyfgtuVJuFJrArymod7quKcMo0oW2F1bUBQ/NNh4BM9qXF3AxAOr
voue9nfDwLP1gHBHzmh1r3/UXukRc1WoUllG1Z+tn7bpScuj6cwVVwPqaGaKVEGu
4DRsVKOy690i+q26giJWfd+a5J3WwxOwLeMZQpdfgaMB1Z103vcEzwoIOXD2Y4mC
KWTINXs9cMGXr8WUZvpOJqn9HugxSpwDdvB1wErtVkHcLJftEH0zlvvf6RpUTCq6
eSkWMSuyRkceJlGS5QcTV7ztDatI7y39WclS6t592SvSLJdgxIzP3AZMUXmCMKLu
Z6nriihhfvxHDk+yt9B6uI3ufPDJDTp7kbggpa2ozpnWXxI1RWorDqwqWQzwaMmT
MUPfislNFZk2E4oUSH11KyEJjFlsonL4GMS4L0VKv8At8RsbC06ey4hQm1qsc6Py
i4BAm/LURzgPTkNL6n0jiV+GqjOfmVuiVXIHPqgqrw4DsH1Y3+GTHVdrYmDFl5VV
oockRSg40acr9Y820u5fY+aco05V0X8PP+W0FcfX3KP1YcsP8nYecP+uBpha4eZc
8C7sTrq8C3DFfEuDTU7KBToYLDhSd08jsHdq09M93PXdrxc8XKtRqoJJOuvBjdjr
Q8bEjhkRpVabEFtz5EBKnCZgBmy8NB5GSsf8Cz/N3TLMdY3WCSbAKAXI1ntDf+gh
N0iA7yFZl/vMuOH5BDBEpgjcEWwCm6fzZRzutrNHb/8QoO59pu5hplSsYdH/+tUr
WaGX3JbmFvv3qnPL9bfvgebnupwVexkzc+WdRY71L1WUcuNKwFDvORSIIeqfcmuK
LSe+YgokIzIKVaA2V9+vKgb135HywLaIzKBtPp0S0dfs7YVaVXGm27q7rFi3QPHG
A7C9AjVSVxod3FzIHMPfFjDqFp50fNpdql0/hGe0pkVjDxJpOZVeRk8wJvmVnn50
dmnpYmsiTEU3n4MaU80JFgZkVMkGvOZ3xPmAhNiDP3To6CMBZxfpRNH6LoHL2/CY
TpcGJ9bf2Cw1Kzn4+7EnSrmpaZdI2sneURPzWoIVrpIm9qnG+wdapIO8WX1V/erz
huE0q5KY1KMA3qXUR7Tj8y/2W3m0Asu1zJEuQZbwWkUeraWCha/jMZi8lTAsu3B/
/PkOOQ/Dl2UyUST7HULY8z9BAu6JWev49ooe1LJHSRxxB7hU3qs7n2rNDySOMi+j
yz4OEoVgdaxUQQHf2ZapMJ+B23Z5GCOCXKFFpHcpswRfQMm9kPNtkK6Z3peYjet1
rpk5jdHLpI9Hb+koNzktcCDvUKuh3XlUGuDajXWDJAP5hW1TSh4vpU2loSJimUze
idQORmwZpAcLyTL77nHoSgloTy3l/6TTcMZCC7WQjaV2HFAgMUcYSmEy7UUDEgBd
YVXqmmYZu4ZRaDIWPPapnLUryOT7hpsBBybvsuTz8oWIzHhaSDcPN0LXCd6JS57i
mfhW5rvrUETe4UCapkYfFJl78evDvbK5CSEhxvCq3PoOrM6WKoJc4XaVfJFaF0vt
xcx7Yq894nDvqyeOp7qZGOXsrEo+RAU6uqz/nhGnzgfvcajNR7z2L1aYjjgGdTZA
eeV49DUQ/yQwVBxMlXc66ijiFXYlYwjfDinyMQP3mG6uf/1mhkzs3oM6TJNdi2G5
EOmuTn024SoZGAFEeC7/9OsD786CGUmG7VzDkxoedBj+NjdRM382t2Lvtm8rKH+7
Sq/BQU95IKcgEhTOCDQTXr/rGNAJ3OGZa6M0wqm2h9y2Lqn3ooVAkyis2rjh1YHD
5Rhb9E1qMCj9TglcJcSAkQ4ojMAIK4QE3GYhVZt2t/juA8x2xIH3TWQaimAlPUbl
q7VCBvqFdT8d64bFJ1I1LcE31bZLZ/fHbzRECk5Xi97SRU9UZYzVjLRmDtJF2RDK
4h5gnGcSBW1XFPUMW/uJLdBV004t0CcvYZT1nK3ALox6gXNoMhkL1A7Jjk1lkqzt
gHyu5Xa8Hrg2DaqSiDffynp7sfpH1Fs1KxK2U2t0ZpHi844YJYuN2gCWKV+S3yaj
dqqhBsGgAcSpPkLYPNcS/RMZ8XXKtSv8v9JCrO0zq7FG+EnPZeFZF+Z+MfsDlaKp
pE8BFjcqY8341Q+G3dhDqOtE8qoCjSzqDMvugJ2/IjLG7kaSokD9V9T7QvdeKrf5
Xpy2mvgFvDKFzflWaLMORUIPPaPMFfeODVeQapfIDYyfeu/zB8aaF3eb/okKews3
aOhETuir+u9/cNdFJZUIe4yVATkxyBCrpXLdJ9GTdXpuzZvNSPE9e3k2rA5Vn+7H
zhf2yqThDRuCsgMIMo6xxi9+1nkuqfxgdgygv8JpHhe4FaSlilKDf5w6WhIOvjtb
A5P9Pvgkq0C443sfjM5vk3uAggIqK06JnzTdjrf1X+LZQrNfJUEqTfn/FfNcfOmJ
H+zkg6vIqBTeyExz6TO733BQM5L+3LXL62paRPG4ivTKh1QxQrRz1ZF1c3dfQFJU
MM9lDwwbnE0x9j8mrQWyYX62zS9/egcpQuo2ZDSnMMs0nOHBgJdfWGOYS87JT/3p
b0qYz/G8orpYAiOQCKtag+7EFVeZqmFYE3gvttrfkPMDHjm42UU52KJ9Rvf7Fds7
P7neXSciI3vbg5eI+jTirnudEqHRg9VH1BkRRKD+6yr4k+YflC65vGsHKc2aZlHK
Qsr7agdCqX4CilR4XgM8Ue509ZFsuRWSgvTVuFs3liD/MCG+KJYncR0tqMLGIcy9
wNMWERjpD85AnHVDF/Ob9/oeP9F2myKLTCa267I8NuulEy5IkpXMPkJ5InQnEbHw
RaVlwYHEwrLBgGEzJ2A3aVQWXjbiOhCUmphefPZe54h5ytINkv7e0QfpcyhZPswu
iguSAwWoIYlamwgygz1r7VntgBqzHsCtA5A4iH11GV24dAGzgwE6RmaeaO0oLHbc
oJ34m1yBYIR8HeeqanNEEbAY20hEL+Ozm7A8pJI7sNi0IFOXOqCVAxxa8roPOEJh
VVEUMgOIEhft+NQ8h5j+i1HwQBT5eOUzmwBrBn7Jo0JlvUxnoeNo9c8lcBS7uNC4
mGVurjy/QyItAu2w+6ADnoyfCOSLnjbmggMzysV1Z6B7jI6mCLWHCn2ODKkxxDW1
QxDEPEUZzXb2N4Ds/bgVmlJBGfDzzeiHojyk3W7F2valq6o65zdMpiaP+8FxhVKU
ZLQqrOaMFIZcqE1pO76na4YFpKnqGwqERg4EA90XhwXxbhRKHf2i9ow2zCKwJZ+H
u1uuAACfwq+u/aUQn/b00SXrX01EKF8nAi9sUsFLNzhBgrECTIWdcVdAm9VeS9rp
MetD0HfzrTMedDU5Zde7IJ7W6QgTeKeyMe7jNZK+ahv9lD+udxYBOYMbV5DsweW6
33H5XqvnTfBqiTOnAQLbEGpFF+rQfu9+VbehYhySivPghv4PrAARKgwqokFBLtI0
oJE77xZDLkuu+HvGidXCwzGV+F/zRpW69teKD5zo1h3jlwFu45ZRRABi+pM1FSUZ
D2nnZgyX5WhRoAX16P9aHMfXb3bYIeHAz60rW5la1sCPQZ1gz4MLEHopic38R4SO
slhI2SvfI3HXPc6KPI3wZz2JTPPy43mXhFc1XZQKSLhk5h6HVQVOLZvBCWL4fz5z
s7V5AYbp3dRX1zBoJIja9uvfZKtU+ULhKYa6hCg4BQBMh3WKWiRBEO29BTcYbBjZ
L9NUlqgobek6Ndj8JW/sA+jXW8XXhNyyJJQNe0PwgAuoC3X4Amb51BogvftXQF0H
D6metT4YIrd7Kp+HebMKVvHThDvpnO1xZvRKTDBXfO40kZAQNLfNlCPlIVc4ZD2h
OthWcl+P5Ha0kl9AGTIXKUx8jqsRT5Hi2hrzFqIVSEvsAFXswEIZ7QbCI532UOr/
shu4BkXIOqKmL+rxc62utjodlcSPa0RTD8T+G4cSVB0vjNlkLfRw2h712oVm6M0K
Nw6X7dzCqvqgpjWNqnJER+BmQ99s636+RGfGQp1H9aZ2mbAUgx+xr/vNZ7lLqAz4
IF3FA575I4n14mmw31U1N1jmDBKCNbKgfRp+3tVtBbViM1T8/E3V6brHCV4HsriC
sCZnuXmqglMkrrvwe/EqNun7Lw1Pe3iGxzjCNB6R5acW+jyozWauMT/itL7ifLl9
GAdhsR97wJfkXY/Z9TvMfEDavZYAUBlPisKYZqMac5vvXCTM/dx4m4ySgkGy3iRw
xLobZbxWY+1TUAmYpidOaHM5GHb45qTVMiChEmiFTVWjWyk+7EIX0TjmlxvmjeW2
stZBv/Y44QTy/0E7TUY31v02G1bHO5Ws7Tg2kQpiAsha4pqW8yzmTzPwZ8xAA7Bc
kjPtUj7npviliq02exYqdq6LeWHyRUZyl6JLMAIUEdbDuk+DP7SQTBZZLOnZisi/
atGm/5o04C7GJrT4666tsJotufuYUwZcp7iTm5XupdmibASfJzuGbA7XarZUZf5r
iTldcZxkVbUL8LzHsrG/fT04lz2LZX87zCgkygEobNOoxzbz3gqFtNpDZLmuoiv8
YgXF5S19vLdh29sPNSFW2qC/NqquaFDsl/7zadSg/0RiAM+KJ3Ret5TmKl39pyXH
5QEHKAuemHM9aPaNYs6dFIwyInSVMqHGKWW8mgJS1gcIkPHr4HkgLI5ruM64urMc
Dp/PI/dxjRPd034swNUDTM+dLU1T23KHbE5dXwfehWBlbJHxWBW/gWNbc7D+wg5n
N2TdVDWvfk3e6UUsIfn9YAtQqPkAlJdLuvVWvRZccAGQIoaE//RLY9LCKBMreKOO
dbaI+PDw1WqzBIFsqsHmsXKvveDG4whcMcoU/4pe+1i7R2oqdxZWKyeJbnRRDkRw
sdeppxJlfoSBfx+aLqKicbHJwQMWOqzxWh2677a1IuUcbXg0RCqyWg2nYwyjyvBf
cX7hwZOBse9a6+ypaU9aKv3b8XQ/RjXHhwpR/eu8EasNDbxieA62caoGwvvk9DtF
znhtaQh1609Ql5p4sTf/jdrFCwrIBqdnqwmDLgiq3xIHwHN7hbDA5ixOO1WnTWvF
9dCQs0PhD04oafl8m3/4GkAHYiDqcCyc9C39yW+2yI1XItCbAd1kRSUAv/jNstqr
KFjYwGgtWwycXjYiy2ChLfWud8Ee8CRv99n/SSwqi08tOcM8uaBIY2AsqzbzloEo
Gj07BA+CgAd09GZZssgr3xLd+cxLpTgE5VMwg8wrT0DqrKkbwX9j2j3qWjkiGfOC
6Cx12wdA1g5YCvd+vpMF/WB2JjI+gvlrvmZrsummN47go4Bn3lKx9zw15skQLf/C
DEjZGrNsxIh3sioC9xR/RyI40e69YIeMYVdMuuDTmiUuLZ88svGvFYund/O6m5LD
bqFi7Im8cnEKRZroAv3rNqqrUkMmBoNdITH6uOw8YGQBb+FR/KlHUyf2SqDtb/qg
3rnomGkBv2+G0mgtGqCMQp8sHNT2YUaS+D77WVEnIAyBcLnAMSuj/AQ4kqKZ4PEA
e2ScvwuwetTPUUyXzU1RUJg0Pd+JeTEsmvExrNDKmDuwNKgjZDK6jZVP2W/EmFz3
Ac9OCTE7wns7VEwOiJzoeGfp/ukIQjr51gc5nzFHnqLLBMCu+un5DdVCjMmVHzUZ
A04nftldvnZgLB/amDljc32vBDKCqHDnEoG6QH4vN8V7LgD0rhfatoDDZ8+xRovc
4RlYZPd4HvimijWn3vHFJGP13FP5cojJE5qh4gZC4CKGgoVqK+1+sZSr07il38bN
02AsoPHi/ngl2j0QeHMM084ZAwSIMiyuahbZYmI3T+akLGAPj68S9a6oNmgJ+ww5
0SOMEq3gvldM9MPl4QhvKv3Y9FC8iWzGPAclhYQ7Nmktrg2p89jnJkrKpE8Qbe9Q
hGWSNcBZzmG+FzsMjPIsqe5wwNWnxlcWLMt+bzhigVc+GmzINF9bvJ+2z3fpS/7M
7qsYfhniNpYbqTNO8WKyNwTsPQIK+2Lj6gyNf0yClwbl+L4Hz9twSMCdb3JF8SK1
MPOMUsKDDcKGIzGlSZzvKdydao6rug1ijGxFyMAAIggoLTouBdTiMto3AIonPskT
Xj4l6x0+2EF0NkxfY9+Vf5LsYlqFvBBWQqQpTXKdBd6h6DIMoR8Ba6NppHqKWHfF
f173KbW6Kcmwje9WBSxSo/FxrGsSDPDhGVFWeEkBY62hwSMCmfY8ZZz9ikWiGEgH
3lCZ/5CE8uplpOC36+M8mF8qVphcxvqNTuYwtC/FborKxhpVvrWfBoo4WgW3OSWv
gE/NV5LlYP8oizp6TY833vgQ2E80VkA0Kg3I1AuMsstt5SCn1Sfpzd6Dv4A9PSuz
ZX2qLnRy6uoaVMTNCJ6XoaM2C92DINL3pcq1AI8PEtZ2LIlhWBmAAkdLiIcS+/iZ
mhNLA6tBW/IFFTSybg0PIjKJN6+SxiXV7vJLPbEPvLVT4DmOgWCnTxL4JQi81US+
68IS+AsT3tFqN2bTvf6pMxfKEhfbpWbwbGYrNzgUYBq/y4jm5rb8OmNIfv53jb3O
VaAO/OAVUCSISRXVFhHN/FHFTQ8ooP+VODVE70iBFL8YhJtfgYwZeQrWL+Lw35R5
riQMDMKVg0f6ziDgaIh33R4zY75SuFKUCpJ6SeZ9a3+pqS1nbk2C4nlM6SYyPhXO
bGOYphYVQuT8HujxdrevCkNpNlKqcnlDuQw+TPfgsgwG+RQN5ZPIqXjbU+3MfsB/
t7Sgba8vmWs6xl/ULvgJ2NgNhXdHw1dSxF7NuoueVcWLmh6yMoMc9kqTgtts6J8a
RTGZ9wxHZkXqOeRHgamInD088kmrm7GWUx5aispj8IXxGKH8SPc/GI609R1Jl3GF
QNSK6eEVPtW2zMUaAp4BWGoAoef4uHz7oZDil+faNB0fSLN2LjJdUZSVaxCvdKFN
McxCFcLgl3EQ5vnz47AUDCKSVO/TrAoxrJo/by9VINagweEqSt61KS0Vbt5nv+AB
4cRPIB5t8EW3SOk601fVx+f4jBFN44R7rHZC9i7W8dTCQltqZjcY08fZHEHJJiYR
TTY6TqIOglJZuNFbonxiEQzmvKpPjz3ASkn8ZtflOxakyGvG+X/ZxcgkcROHcOht
6MdypKaMzlfQ4KbRIptkkednzIUfzWZVHaz31m/VXRAa/aKmC6rUMXLTtdLD5UmR
3ml+4zYwBlP/BavkwG/YO221OvgO5hj0sFtSjXwbLCr/L2lcIxbgJ10NRzQz5Ysu
QtvGRvukEa3AE5X5WyAcWCazRQ0zAF8hZAXWLoFWe/SsHkcvPjdPirs/ZVNLwlsg
/kOspG0UqBkedLUTRMLzWL4qF36aoQehp/r5CApp38hsVXc3v7V+GVD+7mcpwPWM
/vTLijEJe6p1vZYO8FaEB/68lDhlPQR+puxLzsQgrByzy75DmsK7/UgQ+GedP/Xo
t1ikXXnypGp7vl29dQsDFucG4z5SPkWbrhWNAnlkl5hN6fYfWRWjv1tAB4rYett+
pJGaiC+na8lw4x4vRN/O3pB4VFPDrEgcO5q2pyNpUemmdXw244Vi+M2m/7TTWYL8
x2bpPpmrx3hgpscOmhoHgHx9LX31fShlRhWLsZXwZGkrjvfTk1cGTQI4snLUifDo
SxZ5ph+wBeZGM656iWT983d0uTaHyCahHT/ZbUMUt/jABFD/HDA3JzBcA1KPVoyd
ENwfIvDzMlUt7xX8e7CHA9W+IqsEi6c2OA9NNXSPUKBoYQ8OKJGMumeOzAtgW/3W
HhCeXNklDw8P7IhYRdoR3OG9/FTKFHghIpELELyAAd6GqwgCRRjdMYWPLuSOcaYO
xzrfuVELakhniVP9wAIB250MIHUh8Fo4c0tMf7wrtiAs1ATJFKFste9LJ+l53xCr
846QMXzkgPV6vXcD+wKF6IuYq69+8nogE660lS/bxhumQ6Ugt2Rs6u+QEW+p59oi
FK1EMVs85RvGTjqOjhDCVyXNVNtdq0S47tORLMbiqdjLKW1I+cdy5/rZzLM4IEH+
xaICgGW0sgmM6y10m999PXwBKeJ2Qum79h7lgNpPDzahiY8vZsJ51WWoaDl+NFeV
CYjbXl/ENFB16AzItm5tGRwGNSil5IMdLym28WQgMKQLhHJpVKJEu01Jdb7JyyJv
oZy+e2e5kx5dCub9cRw1MeawlHbmSywT3F3YKI+hX+W+M7f3o9w8KTTzkRM5UNZw
Mm7tvmjEolFNRHwYY+GXBbqkSFfsbwypStqalrowlREH97Z7sOkfzWXOVVmE8BVa
/WKfxxVo9IFatHUZr3JwxDSyEi6fvGxuhUCe5I+ov/gUD8jS4+NgJCoDI0cwivb4
qHNJVi8be4qS20bWFWHSNP+MiATz9KVCAns2zkKVIt+crhXY2jORIBiY/TnP22Z5
3bRwEMOfum3g0PLHAIQQrKpBczIc4sB2nlho2ES5+Sj9Aw7LGwVb9QGZG6lNjFyp
6ajqlhMD0y2YTzb+NRlf1mPCNX61LQFv0pSNDEIU0bx6jP0Qhm6X7rfRwUkMWE0B
UILqtXpYxH85xHjrihNZvKGABbzpIsc0A70nhbuBQwFG+5p3lm/CFK1BewVgt7cN
+3Yc6z7bBvefLIbz9JfWQ6ppgHnlb3xP+APcaJWR39q/9xS5Pz6zzXaziF8ZAUml
uArZDC1CEC1wZh4oqUU+h5qMzWRc5HoBT2aN4cExGRWY2WIpHC3QvlyERt0fl2MJ
XehsldkFa2iliN2D6YNjhJ/Ek6IXm5CukzH0UlihxwXaroPfko+MRDsYEPbMwJaJ
AHb61XUPTgh6FFNZ0ADTXZg2+ALqxZeov7BaQ+rmb0bxg6fytcr1xdqtzdt1ps8y
VLc+1b15N28fQdktye/TrijL66mkP1alDvSW8paxLrbXQBXroU3ZU7NqHpXJ0jJK
LHqsD/NaUQg83kmgIN9y6bNSgx2QvBWXhnLjcX6IduJLM+ziF+dC1ma90ytKWqn8
0MHFR0e1xQolgZvWjuYhdLL6C/uWX+bscsEAcRBBS8cpE47tSjyXGQti72Lf6eLK
cJ2WRtpbZXMi2aBoEEzlZPWwCQy3iIh0osgV/mlK0BHhOkNZ0lEgpMYAFvVhXJHt
q2F4UCXVLIQRH7uBrVXVWFyvOGTAAww+uQ11CpBF/uwawf5VDucBM6NwQML+A36L
WG4/e0kShbSWZyOo/oVqjiG32BpvlDKRzWreSUA8BESKB/O4rgi+nVTOJeZbQAIf
QgxmYTPI86AdOZJ/mXhAgmj+341+F7Rmisw4oa3bIIC950ILFZRoPuaxXG1JeNDU
Bt1xlDABUKMlY7w+fDKXj9+zemrhWxJjMngaDKStbSXKdNPCbuwT72pKTCyY7Rpk
XRZw4cfsHfZ04U+i8kA2fmzm2k8rjcdR92gUocjso3KD3Ex0vxCIPIrYdve9svSk
TGEHYBdXsV2q7FqrzafPkiMLu5bGOh5ubvEs7qb7NSMGflzuc8EuzrM9jVrMYAJM
oBJ9GVcyNXwLxd0PBbLQQ7M58/DR1wGzVcBKs9RPwVQUmxVNJvHcxxiAdBnDdKdZ
rXVTi0d7JnFpvOSLwJw23CmCA662CUBT3WpZPYXE9KMm85khP9f9SfmV7IEfvWgZ
HCNKOhT/Ua6EuKTpSy3COroISnw94dr7AENbEXNe11VJ0rFcCBxaWrEmyHDppaWp
8Mx9x3HftUqCHOFcJY3hgdZC5ywLBQ6IzzprHJoPAVuAP5ad5MoAOvdwtI8OgAuX
tLwoFIgoUoSQG5LaQwIBpRgGpTpuc4RyNkw9HmVM9/SVtK4VEQHMGIXzX4wUZPvH
gQaoOJoz9gFSivFh4cBTpzPV93D+R5Ch1VhmYIXt9QLYU0VYYc3WjvJyXbAqRjny
i4XHWvJrtLR7s2WcoAh5zUFy1jagI5edQLYEkauHMZuuWS/bz5B0DPacKlityHLd
ungwzvlUAL06ZfgyHq0ixtAY4LYtLnDH5DaNM2l89xdVroTHnkqG8gu1UtP0MtyD
uTZghmw2kLAOPfBoLa/CKBVUORtGWuYD1hkz+mCs73CpCKX0s/hjgvNNNvDLSWrq
F6+csA90JBsVcIQuTQOvnxnL3MOmBTy7OvAj022WuFxv+ep7IQIAmyY83ff78LMw
K4jDDDy52vQQsRBW8+9pantPxfvpkYinK0Iv0MTQ09Vgq2bwDneRWbyyS+uIu76r
PuO0tust7edUDO8BK0uo1uNrwTIGBxR5MGQ8cz/m+XrWJCFe7fMklbJI33p2G8Ge
SRMinmhdolLvqOmHgQhlgXZaxgR6qzBCBFBxMlaql33UT8/8UmM20cxDyh5IgHXh
9IC90ThaGe670RZGj1alDal0TFr4F6qp4BLLMIJOqid4cakd1oOQLbZe+gduc8gV
oZTjrjquDxU7W50iX1u1yTbKn1dQu5+DmKgoZ3iN+LrJxd8BgU/PgUDsJnWCNWJ0
lkoyJ9bDe87D9MX0YTaDqmIYeD5kmtKoJWuuFozuAN7u8zxsgf849MGy6uCq5ftK
JUpItc7GvC6AfOsz+Wq3VyRWzqyJkex+cO/HTZ4VLH/l5M05g4pnS8zw6lHXQt8J
San/Z6LIWne9wWTdZm/viXzmexPgGjeGQtPFTUQN2IvVgRKcD/6Hh4bp4DMMSue3
EcXgPrJlQeiJ2YvNmNxoXTPhYOuTZ0Z4tpk9/FN/QRIMbYgyiUohmphToNWMKsBv
jm2nUlpyFbX6EWJh/cXd42rzH3ER2/UTzvBNKDRvUSHUXmNM+qgwHKvRB9caP/Nh
1wLQ+gY3u0D0YXnRTIvJvdWhpCju34x4uY5p8Hk4WlsB76BsoRoQrqY9q/hIk9Rf
W9OOTULMfJ+mKhG0sATlCXkzjPCCNs3XBhZbWhsSmx3xBEof7uvUN2eYu9surjy7
5/FNoj2VUoohk/Vkec2rvE8CBGYQdwqg2sRhKVFNNuJgMQ76WyAemSOCmJLs4lOu
aA4J4kcNeMDRgeu9g5HtZzGbrsafveEAm31rQ5k07IG5YvDfq3DhiKHJERwXbGeh
nFhS7J+eqKpkkTu2P0JAkVcJwH/gvf6jDjyt+os42oEmE2kv1GH8dLL6Dsz+zuSk
c6AMF9+DdV0KdCj5u6Q73NDmMalbIHxX0MsSqHXFKMN2gPhOIPkrQhyfP0jxz7GZ
OqC5NKPUWlAj31cEMJCkuY2FeEMhGVmR6l4dj6W6aLHg6LCvLxpwIzREEkMqvMMR
U/h0DgI5Ufx6Wwq6ykWAZ8xK7BsNuSAsPVfyj4GHTfIb+rL1PweSNNSz18JmhJjo
C/nbnER6eR7XHSh29BjPbJNi2uN2iAoDlC+TRuV6UDMtAQtYkjCtuYRvqIvD1a61
KmOLwMbR3GE/k33iPwDENkM0FC6AvW0p5sSsGVG4DE5I94JROYF03CiDdOSNdTc2
42iRVChbM1+S6oY6+LVW67wjUWhraxxdH/hLIidPY18vaERFLqI9nHte+Xtu681C
uet9tAV4MyeJ/6KgFFRdteUrNe6D+Ku2nYkqNXQv0Qwf6L3g1Ql2qls6AZRIfs1g
gqNb83Xv7ikxckz7rZbSl0UrvJOcU/75/EOEtmmTd238QdInyI3dW/cQc8UwGt4o
h3CStlceGSYfyL7jnm2aLnRa0OLDwR3KhdJlEO9IytystswQ6o3X//wbXmblY3L5
DDfv1DoD0LwUPGQoZRqw3IBT10XgvD4QaTvSqJLkNy7jeSj9DRJvIj7bzRvchxLn
E8rRrGjT9L65o0X1LbFw4Exjb4pmJcYYo++aSKh7W1Hfn3pdcly999QLkB6hjgEv
u/RW4bJgT99NETwQYpwQTj0h0p1ImvHEQiUF2dOSF1q9R6E+Dj6YjrlvJ94vbmJd
JjktDyRWxAuPijD2b6DHxjNXkCK5+MPcAhJDCodZyaJ5V4HQc2owlP9mHJ7Pirtx
ljaUW3tuxM/paiSodb1/ZgPNDNZv4cBTSUDFc88246kV1awHj6dwgVBaeMhqviU/
hxiGGVOhYRb9Ndx34yuiF0c8uEj5lWQhVidSjdZx9Tl+QGFqRs27r4JbsvXIgXJo
+YuDH08wI0IbRcHedoH17b2IPnNklNm+ew0TSGvVEAxcoHbsg1Jkzh+l2ERBNchl
sSedGDIsHwfNudOg5MxxdZg1WxtQldVpUHt4N7jAi2voGvEUuGcPQ62TeeAM8nkj
EXzYw8OHV1TlJk3/E5KjUFoch524hjH87dI0FJsypOW0jUCGVXeb5GNpQ5dKH4sV
oblfW3Z103wLbSsT35NIyfWkZZqwqDzqJ0jZdZmW8PEFhWDhX50y4yEzYuuVhV1o
fdi/dNZakt7XZ1SzHxTGpTFACPbKrmNjylUIlNh8ZPaHaquh4r6DptpAmFMDSzfV
oD1pDIhUmJoURfq1Bxws6rOodCo9NL5FUbL0Z6gE+EfN17G2pylp0hlp0wjOVl12
zuhdRwY0EdTxMs0eF7ACGJemGSKz9fJu2YN6YK2IhxR6Tz6RA0hHlWGnRai06HUJ
omtZo3yuwZ40OSP9zwsJifyhl/ZX8qxUcPOr3hxkZSHOqdEZbbAlDwhP+PJyQ4rL
CDNPBsICmI+hvwGqVq9tbxm6JSod3x15PigCQmZwXUm5IwmCWamUYEBXDjv00OJR
2I8eQ2E3tVS1BSRANsBE9GxoxyzqDcyyLO12em1wtz6ma3JX64QKp+XV+wwZcZ5o
82bDM9GN2dIVZFCaLSVuLnuRg+GK4G4MkFPUJaVL3Pp85H/tSitW5ztYwEjjm2e+
hHoOsAyKR6TFcGASt7KVIWGvm8Pv7Lc3LL0ioB80oT+zrlQWOOUxSYNRRR24+P2s
4xmR7iZs710yRLx3S4Cxu4D/SOzETz0hI6WD4LFqNclPnnSWO+QBhWtvANbwkrAq
dpnJbfBs3NNi7XVzCKoUIuURYviUEp056tGpCZKZGjf6989uBK1/svQEfzLVtAVh
zCBHiAtveEActbucL4IKX+0V5S6Lguu0DSok/OPmjlLijZNZ5fw1jTTuKTarTG3h
UxY4Wxoem7YaPYQhb1kXJpe+bek2a8eZ0jGZK2fHxQu43kern3aOAnn3J0CTjKQQ
sx1Mrbu/il7+idgXvyw9sRapnqEYyf2RZISoJAGn57aXp8bK3UkrcnMuPc0/nKJT
9vJshxSOknOMvhk5O3ue0cdFvGHZDLpnrX5Xl87yzTVyy07jUGRrzXJCkdhSxYyv
N+/pO1k4WgQMh6QwiCnXWAot0YDuigxwqFIqRAQCE1GYe1Nf1fS9azGZHiVdDCzH
dCZBC5zHIHVxFHOtRbHvrn0VQ3zA7np5cqre44KW8CrKsFrp7iHRecwD4o6tq9jq
cjxKI/+sqfXbGuNtZc1NuZA0Wl5hrab5teH1lIILjTyNOJ9Ckcv37YLiHNqWH7CY
cqhWlh1AYkJBGQD44NZwBHE01WdXDwKgnOaB/XIB7URT+7udVrzT8GwYT8iIsVY+
ouTupUXEGBXbDe3DPw1fjqYgBY1/j+kI1X/5A4qiRUifCtF5xBA5n31zG0PldPJR
Wr/Yi9FTcL44g51ghpHK5hD4lnL3g6pLLDjhsZhxDUduPQJC0oKTow75sp2n4nUo
PTaNEyoq1HHeOKl2YzQQmmBo1SCSzMeG7hVUoEIpuflzzIyi7AeHRF6kZQfEVHsB
wT2a8a6ymreLF1lw0v/gslFZHriCtSqu6N2MgRLWzkDlYp7xFAFd7b1WB+KNHzET
0bas14Uh72kZI/tqlcQkZsrOFXPD9btuZgM5ajVHztkmAfV6vzpe10smG6e3wHtp
bDMehXcAU8zgNpw298d7cX+kHhN7W3EU9Buw7NPy2TB/Cxks2HM+Uqb7Ocqg+fpi
ZN/T7uVQAjdis5wDoea86rwywwUbC6IZQhuG4Fg74sw2zBEAuGtC1rWEU/QqctMs
NJjyk0CjtD3MtXPB13oOEGw9T1HvztLDqpu809d5lNTk8cMku0yKYeduhtqSPExs
8Ezfb2+wu4YrxyypCmJyZVUWOR9oyGm2hBFTWEYKczs/l1JnR62iwfy8OfkjuJKt
Gjv3Is4+NKQ9H2HvHzHcgM32rtlUuUPuNafx+Wbq5TMDudIlg5oVbTpjyDmSVG22
NwoKMGKxuWAL2A7Mndxo6ZFGFijYDpfdrDz9S+7aWtyijDjOeiJIHe/L/RXFe140
kyFhh+gGQn33LY0UYHhT69CpPDekpeeo4CXsXQ9NA9xaZni3Vmtn0OOk1N8+Zybd
r+g8N4/UVJ5SdXfOIK1SSdkHE+ypjbPhn8MbnsAJnI43hclb78iHAgwVHYdDFJdd
03dRzsl2RtYaJ3I4Tr1BKvNyD7R2d4U6M2OFVohJdxV8EtEIP3K3ytg1QhfGJ0k1
/v3Qr93p0W0gToNxPok7lnIms3BJvjrsgHh71POT+8m/1uZPwhr1IYF0XDKEc8yv
VQ3U5zT+wUQqfSWrPMcvLpPhVj7wmNKwXhHRDN5mjSop0EKj2lnxTfkZMbdvAwcC
W8fc5mW7S+wn43qCKWfjKlDkx6eFxqizH2jueJFcC0tkRGqnF9iYiJP1a4TiyzLT
sJ+Z21RP7n7HQkofZjURGgPl1Kd8FTMR9OYR/ZL3kzjhYi7NeXd7ItG3roaAcOxo
MEW6Oli1xac4Yqkbd5Gz89rdve1q2hiZuo8HEq4flFb36FuyQGKAAiVnc/O+Eoi0
/TG2kJ2CexLe29r2lzk4ZU9Sgd8UXYFMFBK8IjcXFpNxrCillFHJWbrc9Dk9aFgJ
P9ekL+EmdrTrbEJsZpTpDCcZRLVJ3tDNjZwTNIP7ZhqNNSW4Bj4dLgXip0etBwO2
5TilINtA7zjQ7bVHcIX9vaojkaki9cKR6EErWb8rsIDAG45EAyOwUB/4Dz45M9Cf
P3FTak1prn+dqB9vHKkClYhjFjqXzntdJAIi7BrtfLbnGWTDgzCQ9r/sL3nvLrzS
7MPBKV8J4+TsLPF9YZY4j00M7dcW+fWkPqrIHYpNIdQg2Hs0HdNX0oy1R05J097y
j2IJIplKywF8lfl49tZuk08zwy0GIJ7MSMxQaS3fct+H7QFWmH9Gl6WAw6g1Q3Oi
PxJxImBGZHYEpfCNFwUdL7yu0cwkVz/l8DfFa5K3ANYPB+gSX8GsOI/Pj4XlkKzU
CJymWlckyMlfRuCzEubfjxOJiyRXYmtH50eVxha/ECc+zVjNyaNCpve9c+CyEpmK
oP21hjZCZsXmC/VTZ2Gwb2H/hwTY/cqOfNWnaCgdl4klTQ4ZB/wCpd71+quo/BAv
9CBVYukiKwqXbwankEiqsz9QQ85BuXRNscqbKv0gEL9pQunASzPuwZ3yxKEB0Yri
uVL6N04jXgD4ZopiUJCXKvQg6RzhF7bHGMmc1XHIdFdTytEjvxBzdxWhUTsqKXZE
eVENpZVhDyTCzypJyAXmTvQCEkkhzPkk3QibosFGxigVCwztZmgb/7P0Ppph3TLk
IYd3WtvZQq2nSMqHqsnq4MRBTaNt6cixBMZOGtcHeI67CcjMGD4ReAtL3Jp92Z0H
89mgItD1bhaEazowrgjSnihFrc3ICXvVi0mgkJmtLXicbfwlnVCRTJ56wIZscln8
O12DYplKHKmmuBsM3okFFghjWQ4NbCrgfIlLP7q9oDUsMJaV3E+1QrtJA9t9sbfw
qjI4ihrX+TDcUTwD7TO4F2+2cCG0nq6p269vrTALp7lHiaQvFm6tj+H5vSfUwj7X
J3zaVK3ThAcMtfthowl80FWigUsVsySxjXr1Cw7WeG2uAe+KgLk3DLqdqZn/k/5U
PZIq7w3k8cJ3BZ6emhdreFjM/YX5hvWRiR2pqh7/hnPXXQfN5uyQ+ktdTq/U7L2s
x79dTugq2OcrVKmbofUZqb6tPGMV6O+4fsFff/hilEhuN8lvOd8owkhLq36lAYxI
eCMx4rTbXGKYPSBQro9u2iOWqGIugTr+f4fr+/FVjWuuRwzdqCgC5eYlDnDKmbAy
Vf+6tH3hlyJ0DNZRWzycf9oulRRn0eJWJ0MD/LXmDUf7EwD4CzFOaCc2zSkwahPR
NEOwYGrRk2tOGa2rugh9RZoBlb0uZneAmMtgIdHKbMqqVdydgmtwmJ1c53XxdSfZ
spXirykGsGr07UHQ96TAoHezsMyvL2/tfYAYkQZKfjQ+g7e7TgUPSIsGZ+KXhNNf
cGYkx6XKJmLtLH85FnTzNH66QPbxgIW8/JRdSHbx/ssJlE33J33o9H7kCbG9ttY8
IGkcOhZgFo2Ty2Z/ST2+nMJ5voxZaSykTkPrWRe+2FV9TzjgK7NcjZT3ZQuFWD7T
9vfSFLmUI9TnbGpA+fRqpSL6ddgU4gVCxdbyxIaWauiGG4Z2xSElEhq0+lMdNfNX
A+Asw2HhfzmBi8bi3KLPCcWTk0JdsUTcWQ4c34ePvRs4JsBp+pDiOY3cHbaj0YKG
DWZXIX3socLyWIpQ0zFv5iv/ZUCFoNZnBWin1n5TRTIxFwJBuxdxDKVcLOk0PkMO
P/fFX4OSlRrr3CyDIuayZfTSaokojkXbCmjldulxf01Wr+X4YUPnUfgNCz965VDj
03rxsAVRSDyEHJWnu5w/sLYX/8gxTSkfnxCBdpu3YBr/4nAGfj4yocGBcEf//bTf
2rUH+nys2+EFwoUq/w1pfZ4nPNAZ/y7HZPZ3I7N8s1ix7SDzDMf11BjCfhpTCQav
PmLQQRYrZPNpsihWKuUCWIbw87zhLdcbNtPCqKxjMhVOnRgLu//ZI7rwrMfT3mrD
8aMJaUJetplVvFsHFDNf0iE/DS9YSs8xEsVy5QaKfdXgvfEIkmi8TLCqK8secisJ
r+LNQgcdk9HxWL1PSIeiUtgQrtxb7EmrFpDfAAWwyD02xXx6G+AWTkq9O0mL7Sti
nGXU0y0zi1uLPFnZnfKbtH79D8DB5405dPeE0VE9GfalKM/uo1j2ZC4A1NyihYVN
I1FtlNwhMcBvwgNdTZEuQJDukQeeBYgQ9foLHLnJ9SBM0/AOPFn/BJm24C//Zla6
pTtrDQi91eM9/uDncBoghsxCDUX1t43uRxExEHMl+uaNopOs4ujkbw8p/Kz7KJTF
LdzhhOxknUFJ0JDuB3wEAqEHoZQQqiS+QknRqDhB24XxPV+H+KPKGazrKMBkRxZV
lKl3nHR6hMYwsRZ0vSFXN0AOQxWIQd83urCU+QzFo/GY+9VOk5N/COTEPbyuCPqY
1ek0dBKgnhY4YmwhAEDKE9Nz7ymyrfR1QzEJv075U2vihAhr/sGyosQhHvIft1zN
i8WM8md2oCgk9je+A6LnEJEjhxOsjF0XaWdCNfx5WcF8KBW5FsVL8cWX1yMRCn28
OWxput/qw0gpiDQiXUyF0P+XRuV5AxFn0cxCrydGoiuMO9IDXJiq13/NDQv4O5R9
1MaSS8CgFNhDugXtPjKilUFUEW00vEsexSnROFc+2KLzjPf/E8DTQ1dAPqfORUhQ
xeAv3KZtiyFd0MohViVNObZ7c21X6BUCZRxeGV0kvtPRmHjoHkR9LBNsN6troQ36
Ohst5UWAm1NEojdHtS0jmd/8vyWNNiHfUZPrmDFtWBGiEuXAOF0lfSNCV/gTCyjh
Q6V3FuvhnTpbIjCH8UC6quCg9lNwMMFrkINTDNjrPI4Vm3aV7BeOfy4q8MvcvcYY
EhBtK+56h8dBgkfig+JGYTiQKhcNw6TofkFcAcPp3ORoSezEI0SUp21SYa2G2z2U
M2bLjl3SdrWbwBE+OihQNuBL4E1gM1CZYa29iWk97gJ8xMF+YAsHVGrIR/cCQTKD
IxN9rW6to/Ti+YrEBh+EiLCX84UjjHsHpbfB/w67GEd0fdIvzMpdQQpvN7g/O2Pv
PLp7OsZvW6ljx9B94Fr7XwXPWzCI+mBkTbfwrsvX1ydyjNAWfv+KNq+11v3wDpcy
dsUpl7GDxoNUdLfWIzvcbkiI0T6nIScLWAgfvHePN3e3ZLAN+d9bHbrTPPbbjZbE
5cHAgA5DakbbbQKOMZ4ixzM5UMeS7/q7bIDQfzuorGoqh57KBvooqYh9Nf87FpN+
zx27hLqKpdd0xOWjn3SWQp7Xz/Zen9SM+PED7pYBz6VAwIZAuIL1myuplWGGpjuy
FoOZtFy4z8coNAobUFR4JnUD2W1TzthuzDdsmaFhruCCniTn5zgbwt7oulOCTc0P
7Vyw6/a6uIdWNH0af7T3APeJ8yEYwDInpqlv/qBupQJp5yX6HBu71DjhTD7Zklph
abDN+TDyESJdjgkYH/x4oVcWBNZaMudfJiYrpi5UuFsPXsXhqk9zXPrZa1fcBeUR
X1RtiKGfHYpwrLiWb5UhSA/YbcI9+6+FugqFv9Nv9xwb3/rhfIqYWtsCh+hSEr9R
mQDIsPiS59drL44Oaf48pyZjpKw/f2x51xBY7b7FkFiN+FXfHpgACGcyyc0+XM37
zn3BHSG6y/UrgzO7h6FIfBEpVBs225DqI4jQ+GJ28bO06j6kHYp1hk58wcIgvceu
ZeBPkeDnFFnPHYkbi/NY83p7P9EUiNTI0L01krSjpfmWMBAS6pI3ObA04dsNbnBO
+XWOS1zqG0cv+GlAQ3oFQpm1moEMAsf3qKXn3PI860R/UIAh/ww/osKUhQhD8BYB
Kkz8WZelEqi6+TLlGUHcuqTmvBXbslKjKY4JSuD7RtBa0yWW4yWtfJH//VtppT+N
wNEV6OAyJFKmhn6jbnumO95B9SG1IzRHyHTk6HLMpQOs9/pEltqUcgWKYT8C+k4M
X8QTdq4R3VtjFBbZf37EFt/3WhNX0PlpvrasisrlfeQZRATd+nsvKbs6U2VK5RjH
IjjQZKpbg3pcBR5lzLxU2zjffh+Yng3wEBhtJyEljoJ4ydWY8OTLJJ6tQ8cH/RSr
tdudSkzGnOOeK2LK37Aw3GeOQ3vNyhL8Bn3Pv9200PoF4NmhcqKQT3PQgAm57NbP
O4Ia8F+oKUyEQy4LKNamaS4xoZLzgpRQtzeI6tCfpDvkUbRd1GCLHbal6zDMDviz
70sAU+GmH/EL5MkLCzbF47Ryn3hwi7l150bS03X3YeJ0lYalr+fiBLbxIW6gcxB/
YB12FUoUHnVwFHXna1SyI3dx05i7XLcupFZXGlNx+YyvTnh77iuY1A6l/P/ydBKL
JsN7r3cuZzsIh+7u15B+cbW7/v2d0Qe1zj1lh/ivCel2/o3e3hoSc3l62H7yrHv9
LqWrVZ5C1SroK8TdUhvz/XyUWr4ePc6uxnijEgVjvReHpSFOTXAkh3B8Y49z0lwL
ngFQ+waxAk8LHBOHonDknORwj2nIy1l5Jb0QbuNVqd199xmrW4AkFj1sFCkyEalo
TFoeGDn86IwNsYwIrfrjEROa6OquiBZOsXmimGmnLFqJhrOn5CI40SqGDNVHkZ16
Kt8e3UVfChuS3fV2r5gqdXojEz5lMG8vxJJ/m6rxdCtO6DdelyjzRW4EI9HgojmC
cPP219i11KUGIRi75FPT2+gEaFhiREOcgkD01vlC+zTQjt4oe0P4WE1uKBopZG0h
QnMsQijckhU9JvV5CS8WTyE9QetjCLlcVs2iIeFy46xgQtJBCzsSeKD0nw3T9YKI
0ZsLF3qbMFP/TG7HEqSsazwGDzeCpLIt+0ZVl5y933iWeDXnfaXHG6X7sZwpZ6zT
30wNVX19e1tHD82eZ1Iwl+PBqzFiMaBd8DcU12nxmn9Jbco0FdtXHbx4tT0Pfkwv
Q9ZoZKQmoCPEC3KtIWafaPHqpa1o2gzgE2ZvdWKf3EMKQgXMGdtxsCft/R1bSEnW
trTz4UJTYf/4c0w5gQ7lou7nX7SFyj9NIyBliDNAH3m3j5yC3rCK+KFp/m9o4qnT
NNAr1Q94MBnFk3CgFTLsAS5h5MDBUNiGLMJ04+hyFnu4GEc7UyUmdl+yMtECOKvo
ikhe64vR4HwDmiAZvkfbl7V9x7o7yDVAuBVILit1NKLfq3XZP69TnbJD82kb7A/3
8s3qUAz20zrl5LMi01HnaPDh/UTX4hXznzId3tuRno5kXpKU1vJTsy1MTrBlpCrw
Z+PQuZUbvIFUAWwYtlHypLefKP6+TgOvkmEvjR0aR4zdc+ktyeKHmw3fMRa4tI7y
IPsB4QkrUJHVacVsA9u1CCRY6LOFck6lvc0ijyJsyZ7ic9qGutCDIkgTqfCea1VF
8PL9inbjlWG8s7mmJM4a7nC2H3kmVwv6IPNKXEZ//QNpmfP2Y95q8iOXQOHt010j
Wl2jT8dpCtHdasU34CB0ASfmUHXUNQNhbfmOYrKxUlOQlCTW7jaXit/NZMRfAMvC
vKfQbkhap/2MsN7wCym1ylBs7flwHMlNGfnzzQXskiJITkOUrPvieA6tLiZ99txX
jLG8o6gA3OEg7QSUhm7x/qKjDlZDMW2JkicZ3+TSrbDViK85r4Z3JcciAPcjMc/S
Knu+GCNafeHZBqW/AhQ7uAGKrpF3ttRDYelgC2IhAMzVB0WTJWiH7GOeyglPkFVx
WhA+mQXHKEpbo4X1ZOntLGKjhXS5cxqGaSXfWXEOvgB7VrGt/ka5XyHVek8WAhyV
WexYtlP9jAVxIEU8h0R7sTPZ5jyAiHQr4tOVPE12Q0OKshw+DZqheT8iy09CoiWl
MNffQNwMcZd3zlsn5nu4oswSjXP7gLqKTQhgFkAxk8wzfkbesO3BNc2wQ5bfWCVg
8mB+mNcC0vParvqBavAV8j+4F9cyumCeyR1GgxMY6rFtin0ygAKjI7dg88lzLkHO
yNzRR227fgktp1EUEF1ieB9ysvNV9Q2xZzcF2zTJ7wdo37Xn95fIFCTWi8WeceHC
lYLfNOWgvwKwtadwug/l00d9dGcOoO6hLlMRZOVKlRdyyqklN7EgDVqS5ZBeLaWX
zentJ3BYdeLSBwJegIyZUmoCydY91YpPT97KDCNYLzBiBqd2htItqsF0ukq9/NWE
hCAKdUg4epBean5xf3Cnl5NfUrgknZjhu9kjwdSBdEU6QXBW0hak2UZahqnUa8xA
SCd7KTFlrPHJ3V19+nvlij7H4g+GRfJ08+y2z8VpceP9YWJiXJgVDwidRNAfmiec
BfBl0agquBw2u+0lkthCf+dBcTjEmRuldHiGWJn3a9rs+zJYJJfUfsS1E4tsOPNq
8kka1QtND8u0pPdAJlW5z0hMAqXiKyV/MziJLjL23XQutdaHNytBrTde+yBC7FO3
joTtoTURDQVSjIEg/dVvo7NtILSO6+yqpRazjLkMrbrKy8Px6mmQyLcBqmhLsytu
IXL/aK8EUXHpl581eFZ5EJuzTNU27KXtql14GByic6dhasyM/bX7qVzUGyOe9Rh0
OBVV2o36uVdhzJA45mHoxuK49kEufL42yDqoudJx28aTYNDtad4lF/fEvoJISTjr
/o69pwHEyd5MMT5t0PENtCSz8aOvbPu+Ul4P2jqUoLdgCLbo40FUBkr4kzXtn1uB
dX2oFD7KO13A49RVDNxqbRt56G79EvgQJFFbMqqkiCIGyIQdfaqdkuNEPbrnfzZ6
ai4Fpqq+MzzihvcOVhfWBKWruNEjmDkIhoxU2uxrajMeCqMn4Wet1/IdJ4ZLs6ql
/pNI3Az7FrMG1BndxbED3UtXE3rdM0P6JH+mCjQr/HnK1ra6KE+RNM/IbczjHmvE
3XG00/1O6ZLJWTNiJ3ddVjSYWlurEo3WnrKWepfEYmD0je4TVjIiYqY9fLxitkhX
n+m656b70N08LVtATfx6K3Kn/j5ezM/PZ2daGNO7SfoudV+kxN+n3PaIEnpZF0FJ
GIZH43bIbPv1q0QWwjQas0ReWaqDcLUp3Rdm/43+uyebR6rTcprPWagTaBnkmvGY
1V7ImiiQYPp29KZkh7uBBZS6XQy/D1gT0We3ResoNVd6HzBDlCWOpVyBrSr9bDgi
f/ZVBC/K/uvhTO2v45mc4LcTfqfvtZ20nMSEIDF/xfCw60+EApkVWXFuEqNEwVIj
hEdD+rtiTjsOrsbvOAVZtPpk7MdOr3ub4QfbP5mNMJHHTnNhoraQ4auFjsOUstE1
Lqzfxa+lCo4LPvbzBz/50/1m/VnCUHBdQpr/H0cqy7Vtq79PdSVQfPaleG2vmNjq
MrE3WozA+cCAtE5hvHMYaj4FIHhq7uLEltEjlT1HS1A+tAhNvOT9Fd6nzhbicarB
tA6/b+W6Ay5YeSuPchITE/aE6RlMP+bTYpbSyWOrNUKCUyMRxYIDcoYhLoHD5BKu
oUz6G4mRJtGCnabkVo5D20mFudMTd5bWDQ+xnkHRmhCKumsuZnxqgxZOPk9GxtSI
kqL+88GAMaoSXUvfb4epd2DVH9Cy4jO27DdyEopsM0KSw0GiF7GKziYFT8ZVFX0Z
J1klP4wgeFSLR7kxFQ/D4Gob514RNhIecOMBdMyRwFEjb3eT6Bww4flC/F2mqpdz
E+aCmKdutU+fan6K4HrN8sl1zDQ6DGvM9hN2sv86kLbZK4kdVm81aqsfeBN3l+o+
/y3xgCUaRMa/c7SRyGtAJbghJcfzMInmaM3BLRNfPushkMHsg9p3s4Nrl1EAZkO8
jM609yTWpCb5scOTe26iwocSG/BRIGbZGQ9GW54mBjp58kxaaHjZY9QE/ETPnNBQ
k0Xv7KGiofkQRQiZg2GmYd8Ps33l79EycP0UVSrBiuqdtcIcb9Pt5zyJtOHCkJpg
z37cOtixFBUKJWDs1IRDjONvX9R1bZqKDGS2vh3CRMw6TveDDSgW6qww4jp2FtXo
cEhFe6VVdEZ4Ys9a3YNwbhbnFijP7Jk48uTINQztDoUfF/xIRmJxvk6rBpOAqaXn
s3pJnga7axcyDV0ioY5lDja2FXkCtLJBX82t3iKcbq6Sv5sFGybpGp3p2+f5zoci
aUqJBMbB2Nh54zbl8ozeBLLkkTEaIAIHYLm0s8yBoWzwOoHaxNuQq1YWiTpUeyzB
TpeJGOf+qjP1M8ZbhZYwrRnd55takCq0SH2H0kdmE1VkBo4lySZdw58IvRyYcQal
DE7b+vdmnNmp1cKYmwQLfmXWt63IV6mKA6ZyZSo0BbuFFhyDwgn3XhYwTVB3VcBV
2/Yuf/gl0dUJOVvanDe+TFPfhcgpAWUClaoROQ8CK8zn4UYr6Oseu9a4jEVsU4tV
j/K4VSAsTimXZpiR7GJCZbxBnyHdI+bhz8mSbBPS3RsSSjlg+Xspjf+ICrKXZfEU
Q3eWE//rZU5JeXnKdCVQEC2VyhW0/qUFq1twIBM8E8cxryGcL3JVT1tEtgV2rE0k
vPZy0TmuQ+RrDRVQ+slfJgL6VVb4yna7Gu7VteHCFnqGYrK9q4c7YOuIA+CjBLQw
5N2JK0mMgBwv0we+/wbYiG41xTqG9Xc0TMjnW0T2WOlR9ukZg0LSp8rWzIRIADO/
8jaqiaj/Vyao8yMQDwKK4WUbs0XCkWECRpr1TsY2n8hFf0gAr0o+S/NabPKOiXKC
J8XOVARiLabr/lDOp9ujl347Vmp9ifh8cfXus/2ENhta6NM3UnIpywqZLb3fCRpq
4603S4RbEUnMJ65Bu4Z2+XPKCjiqYByZ+2ua49JMTnLsp9UcH1wFE+TacJNlVao7
Y3CiojoUldWAI2E/lbiO+iv36d2tXweRB0pbSKJgaFJPdJ07dSAc38gXbKbzaOhS
PJMW314igy8dFg/O7jETWsrH3ro9KTq07ofVe36QqHrbPjAqdFG++IjJ5GdcpeUu
S1Uy24HUBpzKpZcnnE2DkUOWbD3kCX0dHmSl1dpgUBo32PtXoQrBAYP2VFcn605l
sb0LcGQjOB3m4O2bAqy6XAm6Tinc7YJaiy2M9Rp9nielzfq862XF9bwp3zwRHt0m
IEju2s9sFX0MLPVL0dmXYFF86sXu/j27vDkK40fsH7Ovp9YD5ncIrqEDS0BS/Q1Q
yo32AAhm29gkbYSro6AfxfV1cecBr5xecv5UosKqC65S7YNwqUj3QRubdcNVz96I
Y4Vs5mozOGTTzsVY7ZBKdPxCajgz9KmfaCD+9itkLlOYdBTMQJu5FBoBXAGyyhpo
elDEvagiYgRvVBcTKrBPoo6g+FLtMog5pFeHGQqCYSeXyRcFeiiGyrgjQpSbtIp0
XM4tPapk+DiFcZlm0KnC44Nc8763YzqzD1jdEzBoV66l8HVyxhY4BzZYLApt5xHg
0aK6GooO+vqBoTQqDYT9cUZ1rjy59LXKxAJXi9vL+LCq6fcIa1abYWlzj9oS8FvH
3t+AjZMuky2rzc5XaUNrhSrfhEU1TTYweEiXz595pL67u+D13tVc+JISTiDSWKy6
Mj/qFqqfhFvzSJoSzr58/Xr8DguvKbQVOKTsNVg+H3w6UBJmJ5KYB5FkCBilkrZa
o+8tSDbekTPmSO9/tHvT2SwH1gWFEoHIQpQqVraoJ00OOmaovDSbJjMxzhjCHfq3
1PC5NyY8ppUNrDTS9egD8VhSjD1HJUucw4HPzfzjW18Ez/pzAKSQnVlRG43Oft3P
qJkt3P/NnKu3dRbBZFmDhbiaiBc6UkMOYa82OXrzjKzyfZQv82EOLF0Pws4fQb52
hrtUYqlOtbYwE1cS5hzZOj6AQ1Sw/f3m5fUBUOVZggUe0XLeSpQME9k23C5c6n2u
OfQGBL2gUb3+T/6Qw8zSiZpshZiDpm79wTvSD9Ms+Lh0xtzf5Sp8YuNxEIR5yjiA
LVv1pcg4rq9mLGbJi7Wb282G92pGMTu5yVjoViDpM/UMf+XbTL/ZFzd/YTOhch8j
VwohObXuaFUPnLY9/fI++abTFdDZVIU9dY00oGotde4+yjW14sILhem+coIID/0u
rTnhdcwJs4jNz7/+fx6glzzDh7rUO9vfydBNq0QDGjt/uXFzK88es+wg3s/SYO5Z
KObp47zD/S51s9d7i0AnhmuyMC3zfP1UPvfATvXkU1+v4XSQcB8rW78OG7a6pt3O
/NwPPxltFNNEJx7HIkYkB0/T0c+naA8fhq75f4ScPRikKSDcRWLSsPFWBQkh50I6
tugT38zNXuaVyp8fJnPMuNEkIJkqjESprqeRpXtsgT4k3FEvO5IaLUiflqwSP6yp
oeNE+n7iVeW15uzZXTChRZuTpqVc9SgIR5z0EIIkqPIWBA8dGEH4J0fKKPQkt+QZ
bNX42Itq7xdkim3OjA7zwRZj9dUE6zWyQeaCIQMNNi6IuGyXT2H7SUJTU2qNZdDE
/b8usxMFTKH2joRIsnYMSm1FmOuCNxIKi7gD+OxD9msfpuSnFVr2b+faEi+nWaQp
WSX8Ff172Xb84k6UTHLfvwyeqK1NqRXWEiaF7gFJBHnjn/m0cpN8Obm+N5QY/zu+
t1E+NM8MdBN2DjQ3acw4J+0tEvfIR8nExNl6cjb6/ZHh/nMlBqF0BjOun7EiKJpO
8PkNbngcyCFBn8bh9YJb3PEc+vs2sFfw18yfSrgwqQxTXHWLf9en7Si8r76jZQcD
r9TxtGiYipkeVVa5/gi2bIBPQWZhm8m87dVL7YYykh+WZe0RS/SqxqUQ6p+wINTe
vmn9hnkm41MYFogCuBIRjtNur7UqTtL27ogoi+RKsKqF9mVNbF1yTWiqsLs8G99N
rYRaQzk1+F3tK5+fBTlrVT6eEmoRVTmlOzNJ8SOSE0Q2yvmx0MYi64+ZzzrEGz/K
g1ZwXqlYH+5o04SirQdKrkNoEw4CB1Lcvfdb1dt1HdCpD5U5TyQa2VtEU9UGRhkX
qZ6u45BzyQy7r2qZFWny7cWFKshjrstkcRZz1ZBNE6RVPK1x1ycT/8Nma+BBFIeY
thPl88+jEsfo2veF7PfrzhobF/3peGsyjDvQZkzhzOvHKzpFWZ2usoFutpfon8Mk
MvjwQl1Tueoys8ggcCS4U0wHoqIQMY3c3Cy8dqYmN4QX78iHLnowrinDNNXJ2svq
Z0S9IPocwi6ia0b4RwG5/JZaFZtZiDpz5EZ31rKVJlCbwvo8QuFjEc0oj+6JAHNM
HEcqNL2b/ediNivZonb4XYCgXwJ8BgKU6zfQeNbetLAhzz42Tok634RD+mxCdwbM
bWj+qEJQe7Zbb78C7tlGw5RabnYA/jxHwgJ0113XHDhKzdLkQ34IKOJppIQ/Wz20
WPd8cP++ft1rU2HdBXsz5mKmOy36U/8MZrk+MBeys1VyOPym7f50tFF/t35G6K59
P5h6Rz6d+RLUKTSXvg/3J/1sxPnDLnNMu5TgJLMjeSUvWG3zCjyF9xuLbTkRMUDD
+4/RXCYkOsi25nMsA3Iyow1S0Rx5hnoV4ShK3ECg+4NebwY2YwWuAycMhf1pEgMW
2EzbNazwgpp6YsTqPQMuos6K1poYh5pbtxe/QiIPbZO+c5qPmXbPUnwan2aOvMr7
cG2nUxJ6JzAko8cuDVK4LZXz5OFbSZwuNnByN8oKoJSiPXWI0a2lon+xKI2Eh/zN
fDw8I8XQ9aPNxiFxp+MTOB1K5+OUQUItmqXSXC21ttG9wIPeg/bVuN2RSiT3zmWD
4B23ZZ1m3NtoeK7nUrgutFILKUMRsu5yNXYeGWTekIuqjgH++aD4jybXTV9i1TgH
fhnExFznqHmg9v4lyUjkIHN+o530N9rKizeyB6mMaX/aivnWdf6OkKkH+CAGqI3W
VIrQaq9aDC52zhEM227KpuozLiq73aJtxULp/TQXAMA6G51E162y9Xo6PMfUTNcu
jfg2V6pn3SgjQ55eadQNnyDzyjT6dYS1DDvzzajen/dTgG+ECRbVLaZyK3NGk9Yb
prEK4pGT0+QcrmMluuI9epgsswS8HH1XmIJX4wqQgNYyrC+F+VsRCDHBb2/6frNV
FFlTZ5vZk98S7hAhTNt59hzKmC7xhL+VZak4jc+v8j2qwGkMAK71rr3BR3UtrJoD
BCuRkPv1G4t2V/VlD+leU4x/PHysPrETH7cgR+doCeqVLU4GwdOn+I3eHenk09HQ
Qh+3Pgdk80hFD5wx9EDswLGfJfqN33jD4H1GG12gewumpBw3cQB9/VOuj2twptch
7GgJSeo3Rqi11slB77lfaeIR/QtDx+kPgsX6v46+F1FPHi+WG6V0oWxcw5aXAI5c
k2bXcBcEMxhU4Q3Hwmw2mSq5CK1w2p0K8nGcc0+UL22ZjzryynprwKzOtLhoUNeO
eyt+o1Z3oUOwin89OnsBfWWSSgAH5gM5ulKn3ESzjqQfQnJms8VTq4Pec0o5JVJ7
eoxJgbh66uFqc6IMU+twjcmxNqvKwS24JCaURmTTnS8vSnRWqHJPHYCMUi7feDve
a5/d1M29F/MiKb9v3n3uy8e83SkquAkNujnlFviKgczm16Tit1Tv9jxBbkuV2KF4
yVOCGl8w2J6QC6FL6YdHR+tkUGFTMtn8KLiS+Y/E2OQyyEa68zHjHaTF+u3J9m2d
YZcstpAi8fVRbDxbhjwHaD2KyUSArplGI0CektEUVgvRA9cfOcS7jxmLLue+CSzf
gK5K27JvbDryU3z899MmNn22+MlqOdVG3TnWhVI1bzZigz6758iy/Rgfg09wjhTh
adqrPUxDQ9vkDddGhavgXnWYJF2o1cIcfooTD1SS9g++aQiD7kNH6/lzdkaDF2BD
dfAVpLJ7CHAcGxYNOp0tZq0AsY2hQYeqzOYbRLIfgI20fys+xfKOv9jqip9Gkvml
qXD7WBeo0RzkvUc1D9nuEXVRrsUEgK0aVoq+8xtTT9ZLVwBmTZf0BCcuN+Rp+OLN
x8o0SofU6Grb3Hf2Ke6pJhpj/0rTKEZKF6nfWKfFx7bQMttKSLTRHjB13PF/VYx+
bJvC2kTCyCcFqAcPN9Hl+0WA+sKh7topHd0pTpPEJV6CSLycxbJVA+f+PnXmz05Z
OyjeOTXu3yGRLTKW0XXjeJyVAIBeLutFiL7Y+PJ7byP41XKydMb29l8DldqE59Tt
rcQK5vknHXWbGmhFOoZ91oNjQKkVHhSBo//oZJfrVvyyUSS8qviKWZlfouCm3dX/
IG35XlcpoHAxNJLNzzybzLahve1qzv3RJJeRxTWvWLpuXP381VvGODHu3dpi9ewR
i+v5XeDJMYupurfLazawX/Tg8lgyTfHxxI0taRZFiSfG6fTFdFucIUnES8ZMcJKR
KxhDno9k55K+4xMy6aPmBtgjnDyw3ow1Z7R8OblMl8+tXj+wvSo4lkwBKU7KK1b/
F+0PzhWROqlTdxpbStXXh37do507euAl6qUA3RYiYS4P0RKlaYOMce1Rcc7a5gd2
yUCzjiNiRwND9qttBrw0i5nqUA58K9uop2uMF4wS3lgdKNke5gKxJmsw8n+kEgJG
vMIY9kEPtWinNoj52EAY3bk9a95pvWFssT2e0y/bzRHkXWzb6xbSEe8FYWsNXJux
SEoyRQ7ja5WOZdVUlwa6wEL5N7w34km3QmRDIoZc4JdWs/s/s8HUbSBRRzIuERiY
FKIwMgMRUgqHih4Jiho4DQJicaJ8dN96Te8OlY5x6Lh/Z2S9P2lGGfWd8p8uPbkj
o5ySYUck3CHjnUuh5oZj1ne9S5W0/bejBhMgVCBSD7lUjbPwUBO6KvI9Qek+OYmW
v/G/IoFBFnK37SEQzrQLaQeuzS6uFlN3XseK8tHdYbctIe37JoPWh21qUq7RniOI
Mys2Lpt8UT6ROZRtZ3h8Yp3XtLbr6xJr0OLAtHLbBu4d7UejHzyLKwyEir6zwCcF
FQ5ZBfBVEyOtDY+bIyCDjVK4R40+WvxazEhchLiTrbQspbi4PzAFC+KtHxCa3nuu
/w7hKnypUai8Oa2rwpcRBUOyQhLU/8hoJ08cFyHsms6TefWGqTXYGX4/GcjJA94c
8YUAsW67NbhHuLOk+hzKjvtVKNZQQMeIKbtGpkJtw5yiPi8MlamR8xVZdjnlsA3b
fnoRK1sVk3HR1BsiKXCkyFFqIZZwAp9dPGJDlj8rXhdrpm2AI+OSGRN5xDxAcmAZ
RZKIQWddOcEB7uW7DBiKiKt/1WhxvwTYaTsPNg2JcRE4Ioa8UlEEWBzlWPuoZS1U
naC6u0Q0EGIgvpx6jl9vS3FyxFB9NWtL1Pkevu1U7inT5cEhQF8/Tu9SpSl4JcK+
qb4aQG1V9yg83w0dHJfR9syU9gztmmxa1cuDt6lcSobdWhLUpqIFkiXQvtenkH3l
dBP2DNo4K3bVhwToo1R5Al+IHBxrfoB1VBdu4GDT5+oghlm0iHIT/Jz5wsUva7mZ
tjoojH5MB2tOSNHzbTKXw+8FnOXVRsH/TK4YTSq1B1MkPBYYvh9QJWdfqVftJf0+
L0dpuVzYPRCVR6tSNkQnjfoiD6muWgB/rxO3bnTxTcMBVPkA87fRClzha0ITMqYC
k9WPPFjaoPg7DsEBAkXuBpMYUe7Yxfb2OZr4PnFABgZZsS7zn7aboYWH6QQNfIHd
gt8FoQM9pFOXXvkkMekV2m6vft9jlrPUXOti2k/sSFyrEzj37Xvd6TU9Z0cj6SJC
9KRxf3Ayp5g+C5pHSeZErf5pw+GwRTyLqltoFAawJSgpuiumT1r6lncPjDiNDqN5
iqAQ/JhN6cV+erOTmFe5V3Mlbuq62Xbs2HXoogibQauaRF/oagyrGnUbx7OLPSFr
YeSqjUgl26k4zSLmSosfpMxtuZVn5AnFqmjZ2slpqffn9d8prQMVmJMWM5Ksi95O
fh3gkTrcks7j+KDf8/Wno0Yn91HcoBhO/DJ4bIw7mdO81KhmpOMgVBW/ix6vjtZk
Vz6hfMsdS8iT5LH2Gtsu3UvrpLPoNEw+6F+uB1h5RHhJBi59q7TGOU5IA7cZZDNI
DIP0ZqiwIxMBHDbNrmb2vghhg5p/mP0ylQabCurq/GftC4k7R4txNwtSUkHQj36M
utRXWKIomcCV/gaBcRrKIol/FiEodPYstKdlocN+90xm/UNWGKSYTa1CW1KpDMGK
/VYC++JnLGaRVUhxpUHmxtL8zKiOZ4v5A2WZAS6K4DjBLlIasmArYj1FjztX8fSQ
/rZKwv2fYmL6ehf5y7YsVxfSAttbUI82cqOWFghlBcI/eaxj48/DZNZJl6ksivYH
UiyqRorc0mO6Vxck/hcSuT5FLEJzs/t8hOEUhaYob43mAEfThjqrVIpiYryKJEYY
ITBv6wbGMxNev/6/qyTHtscLALvah8ktY00lnUpuTqCp6zsjA0Pvz0vUf5t1VMk+
0pf30D42l5s4bKzE9e6JPgeudN5R8o92kiPapyyMKqD/YH4i063s+PH/clbXIrVr
4ud4MDMC6FWm4IoTqnIO9cx2ATdC6ShJRtQIxK8hERNBR/9RgE9qyQwER5OB9pzg
q+Q6NDdKQ0b5bG2RYxhIMAWYOc1cGWUDFl8UGCB+bBXqDnwRhaurVxsF0r8zzf4s
B6fzo1ZMUj57T9bBwCbNPjgmlS47Y/IBwiqUPrzpEg42BWn09Mc8zt4hYQIg9uxX
lfR3tI2TGtweZwJ/xJUVNiQiLMC8pXAGFwjns/wbeGzZKxgbbat7mEIeAd2PWNQk
0YUuoVR2YliyseNqqVyZy80TzkYaXwfvoRDDi1w3j8TSl2K8U6B3d1TWLbuxLulE
cWAdzj7GPrj2m08Yj1mKQG8JvVZIO2Hl6JQ7sS5kUqBa25N9xZbOioFoF4gIfsR6
9UO4xJBxO0IczUEes95ekdiMbgIJlQzDwKciZbYwXhlu3ez7qmUrUSUGmnfAVXo9
zvxzg9+OTsL4R0Pc9HvwMFtcSM1VJnJz0qnJVKnJWhNt9o1zjm3os7zFwjgeP4iu
6Y7WGgSBwzmdo81bAM2LDANJBBadMjkLnZSBuyGr5SNoj1nxnOMnMtDaf+HCjeag
T5qcnNXxBDYnqSNV8jDnC3KsvFuKVSp7/LI79+VRDmtGluJB/mPwuOOWcxyRLYpx
XchekCch2K98UzytlxDPraCUOX0jnup3Cm/M1aRRN0mA75ufldMiGBnDz0vwVSk3
6ZmY7Q1IBiNOmQW7OEM0ylZMjSijrtTTKi+GeGP9vcDetuob6f25DpuoNytruunp
CtRkSSdfaBraXIVOB2U88JeGnSFZvJVZB1m3O0A2ugk1YqdPaqIZDx0rW7Cpmx0J
KnSJi3ec6+mGiSzsw2iUCSElGciZ1uhXS/rhCzF6VRmFDkkJZM2UZtXIs148YbWC
mGah104gevTQ7U1uivbUVgLOus+OXKj2yU5vh1qqEvYwKEPN3prPPOcjvs+YkH53
LUGXJnrASXsAufjIO5AR3+hxr/rV7fj4fChSdtQS936znWxnLs+pRVsa7r7+dcKA
b/6xBaUqT607Hbj9gFwJe4NeDePjx2epqyGv/+HjHLaDKsGMGlW166I3BkaSAEAa
/T0wMtLY6Hi/YHYx0eKD3/ngBCZU0Z+JGxtXa35O/x+ETS/6ZebBN6QUumLcoIBJ
bzP9NWFuAgpXAN9v5czJ8pChzCFJroiZkdtaiKkzKUOM+dObGyKNpVc7DPYhpNCD
O12V4LIaxhoEsP2uGtAbdHIuCtufRmbpOMcYmts/GQakbCf2qHayz1Dc6aw6I5Os
X6GF4MyAJOQ1Jf6TXWVXCocXh6uCx9pZoan2mxRHC7lQTOyg+rpZ5RGacABdbPxy
ths+y5kUX46A2zCZXIiEcwaj4TQ+4Ug9rX5U+eli1DqOa0XMe0R8vx/pxLNcnDyC
hdDLFJRbsaiqu1zdFSGeD23/0LxSAgK+z67hiBiIps0VkBnPhsW/+tzxABzUi4BR
O00NiNfbi4OGGdNvkw3/BRUxJo5Fdai8rEHw1eSChaQ9G7kh5lkDEXmH/vXnN6xf
9xZPRf/6dOJclcYhG4xYTQENeNGdMctpu08GXhcebwX0qAKORj/+KYf4mlD8sudb
lr2eYsg0ZWhHd/0hCzuaVy4axt3ispd34gRV82fUj7oGdNLww5+v+XTWjynPVZZR
OU7MJculaAbaiOMOF3MGwgLry+tVyAsAxZTsy9tXqsOgpx2kHFREd3zrnwDj6ffq
xzCgXQ7UWhmTtThamIy8wgmBw0w+TWWwhhXjQaC5XxAj9oitoE+OcJrNJvBi46Kq
hY/xphQhmuRAZnJ3cYDV7/K6R0CwEv7JQXYSpfXxFZfThBE3GGKXz70FoJf+HqTD
We9SZN3TD/F9KQmPCrcMC+u7kDjWaQ/dCA0qZ9ovsvJGGr7l5SCJCqqO8o8cUO/k
eWOqNpIfugjP1eTV4B6dV5U1p5QeEELaz33QPk8KGSgXRD6rhtr1bQEifmQsgZzC
nsDQ57BfIXHRQ26M05toEkLRSgWvpc9FXLKC6pXcEyskyAvwDh9D2zMOlRFxMG9y
CA2J5yqbYaZjaxnhFyLOSTBDQGpPiWapH5lqPeUMjau069h8NDFqLw1wEEVRxjXp
fy/DApiGAiiqc9ICrJ92vDctYOM3iVpgcQsSLXdOx0WHWB+F9f6Tchd4g29WLHN4
+fkiNgZqPOmEfOp07+LjRzkxHF6niVmRg5Xx54tQ0EfdACr6rAsdDSTaHbhBDbhL
9Fm62bHFQXMNWj/psrmLuC5DIkmPmJsh6Ct0Bkm5rQ0bg+UPOrPKAnH4VAhMwi70
a6JVBGdg0X/Js4qKoEGcdk4wlJ02VByXamp4rcWHeJQclV719NTAhgvD8ivPjB3v
RYtgM4v3dyh54GZZrb4JFRx2vTBx3C94pxSzdcUNseiym0NrVjIpKQW0bbl7ry9a
Sg27VjFVxmhSwQOK/vejABQAh/+XT6y69zYpPUVrlPDrABy3RzgkrQpS6lfv+SPH
dRzdB7zqxEHgstOswd19emyFfPySgRLtNM3WY1ItRWilBQ/sJTHIUb03vUUe0dxY
iUggTHMJXDG5aOXu5T5BPn9MsIurGD/2ncS/+Y+8gwn2eH50MnmA0sQYpVuMZ/SK
csUHgrCUZ2gxMW9TpA6dUixfTWXzCWiV18TgEvCO+p8hvvS63CQf6RuvzoRRzSr0
Op1m3KpIsr7XT8XwKpCoxo/dl2eonxbubDacMRDc4khkQNdDd9QgB04h40N9mk9Q
F3h9uF6YSkqP5u+h1nsT7uFDuhjXMTbiUWm2wHgjm40MEl0On9Nc+V5INmBD7a+Y
s61ZAGeTZwNGq2aCLeCNXN1kUUTmWJV7xPOLTHWI5fwr4Ow30wbLm0PnyBeszfx3
cLAz9dqG7aeTyrmREWgUudcOOgx8mIQtZ1OM59cKsKnOVSsXoL2KV5iBIGsZhLkw
G8FVDPpWB6ZHpCCRQSM4eEfpfSTPO403Qn9y0M3HYV+oyyIlTWa4HdTHuM7GWSWH
MsfgIWsKB1MCjjOHy1ZKBnNnURV6Rb//kpu8/JhBcRpjYZW8N7vWkBv/6iM+EVLT
DTpuPy8U9AQ7Qbewux7AxMupEvdPRgPoISn5ThdQnRpODRlVbaWq4Sptbgm6k64J
yfi+jG7duUdtvKuKfgh41t17hVaGMGMHyEFf5x4bZxRSpqBUHDdb/cP/DsP2CIBe
33hnsg/ZuDrKn4Jf/+ewTdFHbi0svzMAqG2b8uMju8RoNeBfKgNFaFxiQFf1rMK5
VwA330kLMz162NW7WyQ1rX/2xYEyhvoHmmOD8bwCj2cR/R0RfdzlGOqXNBBZnrYZ
02yLoDsjP09OjHJLvmeGfhFFtcJn7rbh74IUz8LbIDu80VnIFmKY924BIsIdLNvP
80+2mPILOvn9E3KcN8skt01Mcxv+mFtcBbzq9Qct2PoIXjMCwaobXzEenWNNBYGX
3LetyswsFuh1wCgk/4uCbsiRC73v7QIN3TsG39zvaID9dvEN6wagTI84BvmzedmX
T7TQE7o+jnTnqJG8Bqo/cKhLFI9rLmse6QjHHRSWZEm0Blp8s/Nww3+EdWRjrqTA
PJPzvIAmv7Ko5CyechKAiY6EsyxUpUCsTdFRR8N1hpb1O8x1cIa4KiSG7D+nnBM6
lqkaqRMuoQ1G33OWHXXMiHA8YTEM85fA4PWRDkhg+7hEx1s6r9GQWrodPvyGq8ep
s3Ap186/m18MCmcfqTW2kH0nM3Uampw8CiKo7Ap22+73dSCislF6ViY5x6esXg5E
uk7x9gOSqMcx3sSJbUSu/1Ii4ZYM8cndX3Fps83xXdDRJ3bK+9vTm33wiv4B0UBn
fHd8t2KlcLDTLJDzIQLrDLIvTq+Gs5p4dpt/E0CIVagX+aqxsbi/nkuhDu/Hmt/G
jUYzDtPxJGIoD6MrhAwkfP4K+0rqr9PlmL3l3aA3lpWQf7TH8limrLHBDSf20jIx
OqiBPsV4vSTUtArOBzBm9jHLyPKupmlp5tbTO+badDqp5FnG2VhEqUZeWkIrX5TW
AEGXuU5X/w18M9oEvtN/95czczjmPcJaU/7xH0P3HYS6KwQA6Ts0yGAlHOInXDOC
f0r97A/pObUIqt2u3USNDyF9orZyMv+Pyzo5z7vDEjjPWUXkOa4X1SvDitFoRGXP
yx9W908qTPDYPBIBXFVLXaOG57gBkVnXxFQyiGnYcJ5upqvB2w+jzs/yM2i7ATYO
Th30/ukl2cjoq8uKJO6DK5hWtl9El35ec2pXddS0GTgLG5ARQuCqNbBhZmv9xGFA
+adBagWj02F2iT1r5OmvoSqvKlzCDGigczN8v9Y7RjS7Kg+uqV96qG6kVYIhdQZp
3GW4DOu4RvEtFawdU/q4FdFrq12MUjLyk77P7TnbFPq4+aGsVLqhAlqdmq5QPD1m
TCc9ZKoJjgIrIGXRe9GBl73x5Gjy4sUY3IhINAfxYokFbzX1WPgzsiRE/dY9s0y3
aBll1As1buB0sNS73F2+Zt5RuXZKl3VnyWoTdQy5Y9ri4zaEaIxl8LpG/yAf++hy
xLvM5wEbdKQfN6eQRIwgWMAfuEWuUFFo2xlOHuGAYk+oSNdkz8e93VOzrbxTBygY
3sYSYFU//DvpUMJYiiM+zMCgzoM5AuH7/ARllmQyxLhSKC77eAFliyEhXnt1HD16
CWHtZmz9XevU4dHd6cYxwa8X35JHriqruWbZbA9zF9njbB9nHsM7j+MLDd34wmWa
hZejMgzHUuAxg8ZTiouRqJVLERe6MP++IXGpjVHNUuh0EJjSJ93lJjZwPGGcs0f5
G0VYLTda5NWlqL24re67/yUoQGPepb+5ANw8SmoYLmtynbU07UDqQX8FTqYHtUHe
2h49stfLfHmiJQo0j+lVoO+Fb4y0IyaPLFRxVWQGijkaq/wT9rX6gmaA7MexoSOZ
TuNOTTkaB6orEzGzG3gpfXKK1Vi8LXO8YgFYUZuY5PEFmANx6uecVAKHuhGR9Qkv
QwlVAD2BeKRDKkCbJ+cQ9yZmIAq1CkRKoIHEt1LwzbfF+KvcavmX9j0an90TGGOZ
vlpeBJM2pIqlzDHVMEHL7QhXnEq4BMavfF4Gof2buyfqm/Dowh7wkkiggNlZEVCl
TYOxl7d3cVZE+EYncnYAs1V1e/5Y4rAOGlr3JRKDdkM03QyOgLSQlQ+n/mKt8GJs
WzFs//fFqo2KyBgPGyI1MOQZzuE7eb0JfjEwDuR5uDHjfMSOONEAzz0dDXXIGNrV
Bnsxu7uyiirZtD2ESM2xkXTJcwGPDxxkP629RECcJLrswrXeYvSD1Fcj4rtSzIqj
bDvTje2ElZcMNaFVr0Q5QsnZmiGLdJ0fmyw2DLGzIIzJa8VjLVkp6jZ/iNihUVnu
cVPoeHKmJ6o6LmYfkCD01nUHnqweK2DdxAm42RsJ/tur1DGgBJ8QZa/miiLokdMu
p7y4n74oEkI9Ro8AK425dR1V3a3MKsZF5sfXITkRDY9gfSaUNA++mKEBx1XAiuj6
zto4byelEVTrEyni1q01adaYyEdxssmkoqAQhOB5CJxfrZAlJ9bwt38dBTCehWav
HH4gCw6/gYLl+WLg5uFJi/8ysqLkl/EpeelyuUiorPcR63U2TOfoyDfuWx2LdoHD
zFuD1US01B4eAvkx9uSeQ4yxCZwZPWpKQMemLOOC/TgV7gJVyr9xDyjgiGpqPoeA
ubessq1p4/fsy6yWP0Ak4D8OfRPYc2jfHfhBmyG/GCah+yHCDzjI1FrXX8PfOU0d
zKWhGqTxMU3q1QTfd2opH8GE2N66h3BjrAQDznMbF1wT1CsstM8Xwq86eNBLWbVn
IpQrF/AYABtVO8R8ymjQt2jNsEaV+RXvi+dyH81OXmeUgSaM0qJGDWvaMV2pI+cW
IjUFOSLT9kg52keDy7xV5rmF3hfQ1l9sn78+nWZ2szCdlZhRLPxwnTRl3jN0+zp4
fRwobYsMDUpSx+GmNFCJekBy0JK12JYFgXmqFwIu+NeqGyPjrnfpNrkkJCNwT83T
0bWgCCU3ltkSk3cbExpE2mEnow0CwKagx44k385OnR0PSSs15t0i8QchTOzSRXae
VH0lt6sxhesOkN3NIRzQfiJedWqVtjSknYxQPqk5qu5avQAhbx3/LYG+/ms1ek2v
xEXXiG9QziGO1qm0WP6Praz3ahcTO10MTJy33x3Smnv3+LXymjzRiKUtQC+FgvYu
/Owaqjmm+ncVDeT6fFEIPvbT4Z+Zt2vDPzZCB4FXmTtzhkxYtFFFjXa5BcYWpbfN
kh2OGrJuhOgbBMPyIQX5OGB7ImmK5H0Oadz2TTRjJ7v0S422HlTI+UzOM9cHZFEv
vmWGYVKVFypF1+vXlV1uUWj/kY/62BmTpDforMkmi8ZyWBKFiuhPQ41iecTvgson
ApGa3S6I8HRX4xAWOQM7yF9rwPMl4u1p8l2CaiEPr8O5RyicTk6ON8GW7UQ/Sb9q
75+ds4hPckwIrDWMO3ssm70qq5c/BfWWjKvpeaUJdttzQqo/IVVsvXnSpgjrwjfq
BcxluC4P0Wl8Ue4A3iPWhHBFnveh939NYom8C0cIj8r1G1pCm7YQ74yefQ3mcxhC
zQcFQapfon+Ioan4KENYEor8g9yTcqnIOeIB2tMQP5Oirfz3390NZqELVY2qFAfN
O88C/7BH35LAxu76FCNj5sZg5oPXUElZ9gL/tLzFL6P90sxP0JRg+pdTALDEdNMG
9ogHF4mCsKkPppIbXdI8nBaIiS9WSnAQ3th+I/62zK+JEag6QvFtuiFAbStaUIVZ
ArTkaqndDUJT9kHIzYnVh/a3WL+qLFX5UEOUbnQdORN5srEueaXejEwNGN0wBkNr
Vi0Pqir03vO6FiCIEIRnRNjQpnknXx8y/vveM1nLpwvXIewBAFT4+o+w0Gi8mk3k
V3pCMEIVJzDuwRiEUn6qeGuw4LqtxxGnpP2x57dS0WjMIdetVYo7XqkTBvrAQV/1
65FesiAz8KeKpfkgBQ7hmqSVsI8C9RgbY3HbOUgGrhsqtKIiN4YzVM9R97p1RxX3
odhfIEomeykBsdWqlb77UU8ggMm0STwKe9QNhJ8v6z6u8APXkiem3LlQ0bRG8twE
L5HH0NiXNw23Qg1Nii8C5qAq3f3emYp+1GT8YnuLh3nQ/Gv9/mTIInchpKbUElqf
TlHIj63NwKUJ03sLC2ZfIWxc+Iy8d/dLhkTX7qIVtkzc1gszsDZ/1/5QqiVFKblI
Q6b8jmUMCkXwr62Vbd1UNcvqwvjV1nLY2//mLuLcd4n8w3/obrJZHdCX6Cm1Sjal
3xbGGiWqw7mxKsywDI1R/Su+3XJVxzK3W+QjyV2H9lyoag6qCWjk4CG5SmcRYYkl
l6U4BVv0s/WTxopxPCL5nq1ztFNMTGnYyYZ19FGpYxoyL8rGxRTlgjb7NsopPWjP
GlzMg2qZ8FcO8prYYdY3i6kCmSh8cbxE9yCDLTqaGgk3bdEqu5aqCdSzl77EGsLo
eA589HYf0nhRfiIma32665G+S0lGYYUOUielKLAnqjgT9fG6DW6z0rkLRhywBS4n
ud4uoKMtSFNgYqW885lyH0cZ9je/qU2/D+ReAh/UbbmBJhDqsr4y08QR+AymOGGn
h/c46oVL+KleSCRdbO62aB0pHT3Mk+aTDtRdhXSj2VenYDvOfkDYfNGzeHz3ZH1m
SUjbphb9BuGqDX5FB678Rudp3Fz5PuuL3MUgy3+tfL3WOwMEQoeV1ltOqbyFwCqR
q+3ILJYOpqCOOepMYf9ZHBiuCc1v+5VUholYhs8v9nupjGV7g94rG68SGm+uhAvX
q5f53TauwYGUvyslTdqEJJcs2CE+fPCFyw+FZ5USu7SeJ5lAxmPd5QkjdI65hzcV
7mfzoxC7RzE00Kr+sEVs1x/WbTjqittrZf8fbGc4GJqiHIu35WzfydyUjckAu3so
OlT2dYWkZg2xIuq3VAvhIv9NTeKMEkHaFQZP1ID7vdHgew60JlSM1bj3UV0aFdl1
Jp6EC1FTexNw3faFoStdLWikBuTQQoM1+eN3MYYzw3QXKd4TFiwD2yNmezsGmr/e
HrEl2e5IRWUWzpslGWrGRXNf7loPfEdJ8KYz54GqmcSnYdElrTDHP4zQPLmRsw8F
wbX43E9Rzu1GH1EKvJv7wuGnxVFf19nsOYjr2QCTci7gYDHkpxGZv2qBs7MwJStr
5U3bRO9H8DHAxU67MRC+X/zbQ5EZ0QVJxx4RW0EXKH8kwH+arahzWinrjsjlW8D7
juDFUJml7c8OWRyz008/cCJO2pHa/77Urjq2FwBlv4AG/m+99u3aWpevsFtEGLmo
JEjUbhAV/YP2nudRXb9DGdiZ0PhjrucbCW0/9/VSSC4q7xCF/9xugmGODnxmv2K/
2aJkjyrSW5feV6sxIvCHpA1FOJWBLG7mm5gpm15F6yEUik/2VoLjItwqh5eImVUW
bSe6Ly15+I2ot5Y22LZiBE0vA1f88K0OPfbQc1LpeRJTHpU/dYamDXbPsnne4u/3
BV5zeVY7w0QDDT9DGhbjabQ3S9EVGSiusuEUV52Ub5nmGshScK+4cNWuYvXoU3+m
przh4EIyw31N5rs0Apfnt8E96UptUnbCIZGAPVtDmjZCUZPp0S/EYoRmaZBRL34z
aajkWkzw53H8jMGUEanMAGOz1h0p/nd66rLahr4l/3c1u+9/n/zi9ESBMSQ4rZ1w
ypSOSkLzxIbphUXhsE+lsbTMmi4PweNbrrzUVws9wruFZ6vLtfI90qLilyZNNQwu
1DPj3gyt5T88CnOQQCwaqTSQqa3gc4uC+ba0ZJKC87MPZjd/p+ZKl+UDSRwuGy2d
KiHd/hjSPNii+yzcPbmvmoKotu/6XUMKzO0u3turvppKzOqIFEfcseLp0ZiezYhG
o6gdaeIN6Kdqt9sM+Ps9vGydU93dQZAV2kWqz1MulY2cmYnlNwj1Atv1kGS7xA35
3Hb0z8mxnRrytR6UW6GyTFLXYrE5X+7hyWj4c0//13l6Uk02mACPUwMoHieEanEh
HggUIrI/M89OqExnOyNCxlAt8rvHEqa9cWn3i6rb1eozZiZXitcrlgWe0EQwbaC7
PmSTJP8scsnc/8VsX8ymvnQONg9sOiaseARwlS46vAMnHjJK2CZYqUQ53bX9XU8Q
rBNmQA5xbE75mxELvkvB710tZN973k0nfrp9+jxSKcdRzV8s0zOwZGKlQPyE9ULX
HdkdiI0dG1l/wWvj34V9+xeapltFhiHDqaeKKiEmtGY7wzcPCjSgXwHvGXJymgJu
g+aac3zHtCrbO/FYq1CQO9WsVZJu1PUhOH/X6EvFH+y5zGG4kSwApyOaIzvbyLtl
sWS40zaX+M1iQWNrqblJf9YNea+LbqF2BXgOosbqAGsWI2A9G7cVvvUx7IJ9HR15
7S47bNJVj974mG4ie9EW/KOBb8xIR++UkWTbXtbhUnV9FYg5timKxMpdct6WfALc
45XpB6QFe7WxST0DuSAU9XFw1AHJI7HJYXMLj3ijhXuKx5BtFgUySn3cqF2+fTss
tarhzFD/hUZZ5ZI70ad9Ca11xqLhvf9VHZJLQ/bQKVIRQzD9I9jlHUi0PottZ2BK
fUzZSZJ4zBDNRzcyGkzRhVeSSV2e70F1pf27Vce7wWFl4b5kNXYzcM7dTo9DCr+q
GHUCkHk8HzQpz9wMghlSySo7tQViYtYQuFtdvnuofDbs5pTu6FMHgeh0bi9EgoAI
R/es/TXkpNMHppedTWGA5xff3LvzBZ2UP263ZB9R7ADkVYFcfaOAf2P0tZmGCHqz
bDXM7ufX9ISFeFJslecv8Ng1/6cPLOhRD7OAa/jdU4np1TAMnXOkilwRCQJIvk3M
s3RK0xdfbc98ohncz/4AGVFdDGZAknG3szk7AaD3zQym5BPEmvXBk0GdYPkRytdD
9qtzAfg3Xm0JoAgRMr2+NR51Oz/maklIv2HHHID9mB7StjKn391jXRFq9OyTL+34
i9161UwPiLM9MkLlRVVl1WvRryT30XrU9g99fJ1yYaTFLSVjWkKBWU1R4xpeGCe5
ZXXspNyzUAAOAxvdaDOUaQ+pQLVuRoQ+UE0ORC6VTdXqDAD8yv0YP/7qXpJ+0Nqc
xmcxhtiE/r9cZGNE4oc980Ne53zPdm7QnoHp4MbU61u7Xg80UdkUIPndqdviWJUI
S839rQP7Z8hOG5i193xMY/tRFin9sVl5sL54/fM43bxC70KdepDGtb3v5jx3y3vj
KedPRoBumr40ckGa+qHtWjNg3Sd5ngyDjJ+oF/dWTGs6Vtocf6SYsHz2B3pf7pgH
M3ZbCoK+axGEAuy4c+4VME3xJ5kCZ2KgJMi/ZOX/K8CXiAiebfzTZv5oG7ZY4o7b
E7nC4zoNmFyJ/ZGnCg/x/mQk+x9T64MN7aHRcACS5AFuE4D29Byf7rvNGTe62q6B
5X0cDYOlhZ6E5WE1de77PafdxB+dYBGU4UcuYXqFo8DiA/3TuseOwL2BQrbTwITT
PnAX5XlUF4zbmJvScvR+pQs5DyRyRrtaAKXCw+0rDuCPgVs9xxOblwhCT321OOhs
tC7/8nz8wokxXWE4rf014oA7TzBRnOO80J7jyIgws0P/hMLs70A6Nv32YVXuOWFY
w5V24czrwu9SsGfXffUUvek06zg76Vz6RxrpPP1GVlxP7YRpOOs7vqhsXc8xcuKC
PrtXDS/KxuCqARtLsdRDiAgkKtddONLz5mISnkpGETP9wg9ou5BEP93QkBNDKu4j
g2SFQZ0bO7abW62AN8uxctyQcmz8nuqXgNeRtkbQiSpCaTBrolN0oZj2kGwQH23R
KOMEFshFTdVZXzuJAbj9yF/79gmP3g8jN1uAr0A+Z2l4HJ56mbcoaflksEI6iua5
M+utvbEIEsqEmc1nJ/Yi4F2T2xV75c/uv7FhY2D+oh2eU628FihHsNcIsZIiPwoP
bc1rNk+eymsx0st7SYit6kX6uVaYwbyIlrxbI4mEjVz0ZMetY1wD2Z5+SFpj7G2v
Xcf1HOspVxdIp6/cyXeexsjkI3mQzYj9K0AU9h0EdH7ZUC7MGcuRhJpBPlO1tqm9
DX0WGFLw8Wes6MUGKA5eXua/D6QerXo/OTXf0OfA2EynzhzHFaiGP8+ovOODAzCU
BmRJOU4hZ71YSt1LvW8Ue8zUj33w5EtP+9MBgEgri6yPYEGhlRGyFe4CCWWEW/sy
6kSnEsSnKrOuWmJJ8H9dEPuk3It3GIuSoP4fA/idrvRBI9MkjUnk4u0FEnCmeDwE
vC0Z1Qf3U13yRhlRbe/LWUXFBWIUgZU69Y7OeylWp3i9OTCENrehJ99aWsivJD1F
NoiKEasQosr+8uvlO2lIIEh60tpwB8vFaqe+tinW3ZDuH6dyH65h5acmrsR8+oW9
9C8J48LToHvWDOkp3sw/qeVhKncrtf5TLoYaztauksBsnyOJtmXhry7ktRCajoo5
PW0qGBXDevR/aYJaU5MQs6IOFvna2g/rRoXW2NRkR6jretrqzX9+wFdRhbyh5Gdd
ZDcgqy1q0VBh5rSP8NiGhdTFPJ7F0Mcy9ElCjFK4ibsh1V8fWVp6cTFCXYnWNQVh
AUPF1dTn7JxmZP1iCiZtZ6ntwC+vR5DTq4YWMFJ6MvWiQBbrf7aID+UHfAq6QOU6
LMJmTzURmwsgqlmok/a0tuElsAOm1OOoFgHFLEVtT+dR+ODmghX7rQr+ZxXaTtG8
VTC5sS+LvV+idgA1S+mNz4qYM/XFzDPggppqLU4Pc0dkEXypikpfeMv0u1zVD7BB
5M+jTciXcWlUfRpj+qNE5pP3m8Mx189RBN/dk/FMaEsZS8aFJgkgFIk9J4ze16U0
VWom3FAhqKqI+GsVvyjgh8BPjZJMXfALIqj5zF3lPed80MrJKJCu46onepd6f/Vb
pvrCpIXMGrlyLqoz3aLWSS26O/naB5HT1w14U3Td6EIGVJm9kwS/+4a6VW8Pgxx9
OT0wTK8As4kXRFGOht39nUqRQrdJ37A0qqFK2X3zKeawttpdUqPfjn1IW7gjCLGC
sK8hcQRWa2wnMXLeWU07BHNmyKxk9KsTWo695T5oYfqjvCKUf7BVNp5OF+i2wJgN
CDJnvGE8+eorvz5x9so++Zh+POZGFMRnDeflgNcxJJ8HRry7xUC9FEMEHZdh9zRV
y3U49ARSzvtRbBCbg7DnEHdqOnNb2IIXbi1Y8g4+O6pZZDpFkRqUNleZkB+4+Uf7
Ua/rKN86u6dD9nZJxadS5LW2SDXniofMmTQOlgwY9pmEdghC9FiVz7Fe3duB5nxg
wxyS+qIwI/fWFyql4c1RB7wJJRJYZa51OGdAszbS8eXGKiD3UsYoNa5CTXPLVQTr
XVT+nZqpUYgTyIuLPc2Brzwre9xPUqXrI5Ncdr76gt0gJGG3Cr7WuREKmkVqcgIm
eEhc7zO2w1hFEo70XB/dUVhB9MsjsjTzmGI0+OBxeJKvuJmEX21Vif995sHqDkVh
MZnEnatoBSIz4X5hR1mA9iiPLCaz+qmJmEFiPsYkGlDjxROy+tgkpYnO3SLgse/n
Kr4/BuLjyEUld8W9t4ZMONGXP1U2uUP3WzuIOa3RIyo09bheyAwRLeFYtz3Et6nn
QtYU83RsEkW2bSuQh02VxvRs82MyLVCuGS685b/a/cW/6KetYHbA7SnbxUGNCCrd
bFQwy1eS004bHtS3RCN1NJA48YgslzbLotSF0hIgn9c6VI52uCeoMZBWoDLIS7Kd
/B9Oe45qvCf2iJ0nsrkOpfeVoiv7Aezb2uyYr2+3tw2ovvkCnthkNYNs8mSOjJZi
Qf2eFifM1kjEjyr57+LIYvOTxz5ItCieGXUk4ymTO/zbCT/j7k1IkdqWUHCReO5+
sF5kfxgZoJByLx+5HyXEPtGkrcJ+jLpdSb6uGVJyrPQpNc67Hs45tdtdltRB2mro
zJL8FkUO63ES973x04lu1IN6gRFSs7aM1u6IwBCBSLeAPjN/NkZ+PuGLd9IJtYYr
fS00Zf4DJgitcf2QQLqJqRa7rrhgRYfkUwKnEOzLpPZrO9QettXgTqfUcLnhzUeg
rzQZOSWJpp6M49UEIR7y7kfa20WrXJytWeLfmwbYyVqwhhAC9iG3d7T1j5BGH20o
raywmu3LGzHwMauSvXjbybuQ0fi/u+v8ui7DjReiaHL1yMWmZq8obq6UE9ay1eNt
oj2pURRZVceyub3T97D+nJYav+rQPl/EEav6X/0XUCzlSFPzgC8l3hT92DWw5TNv
RfzSjpFaJFOFfHn2uXB+6rqQIpWUVSTFqMfHd9qZG5ZpnwPB0/XBnmWA3G79oSIt
6WKE/p3IfkmkklhfMOcbi+B8m1U4/ts6RT/ut0ZL7ZW03DbU5kgoZdCHp0lwDHRM
ASIH+hErRGBYzFOWJ8wlBZzWgz53plBwzdeazPWuGaqZyDIz6ttaAK0KmYvOSkv1
Et0wKX/Sai5MpSu7uBCyB4TyEvWhRJY5zaBI1K3rkYRFBKdA9Y7G+dkbO8yAU7Yd
VqykN5Exh/jGnsOqpQyo/cEFfMC0NHtD5xOwFj1tYEsJIVehlLU8vwAU745cAw84
0UglbTqEVCtlKAGDJsfMLig4sW6yKfsMk+EeniGA4tvCzA9Ns0bxb/kTWeVBvqJ1
rPnDZU/XSptc5VgHr5Nq1liJpvaER3SbyNrmW5FuDLsakdvWt6ssAwMO0J+amzkL
1KjmlASymSEhHOByoWpK1yl2Lr7oEO7ZOhAeIMlT5bdStEa4QfHiM5aD4+sWbKlb
wfQolTL/tciIEnJagVHx+lHiPP9d856Mgq3nf2ZvrRUri2JCvx2T1DWTltVahIkF
4efaSbTOzNyieCMmzlRwiUetL+btHnIhRRli/1YXNVHdEYMpDYUlqXC9S3dhWjva
fuz+0KKdrro6R5vOWzhsyZN9vmDhM/gU28nl1Ie7TtQ8rqNT6u7bsrnzX6mKtZFp
miio0mudOG71lqHbAxyHNd3b9xbFXwXuIt1wTZkDHsgcKx5kIkUmonOBzVtMXKxq
ElLI+zMfAmGuOdpNaBzUL1fwlB+pEuUa1REbs67sufRjRdtqzhPc5js7YY/Z7//u
k89PtRAUEYU+nX4fKZ35RtjwOmg5plKTiYxVuJbAQHKSN8eX07V+5JOeK+E0xVVh
aOyttOteufed43S/aptf3mhQkhQBYBkCRsQIT/ffI0m9QhMZP3JUHrWJWZ3JImkn
Q6c+jKSIl+eXgFpKoMHNc5JKOapUzT1ztzz5JyiMo4287uljrfjw+4oR8K2M/an9
6ZjG2h2hlUTilpzvTWA4P89BfIeAadyRJvhFpKMjEquefMmvJ/GvotQT7LRveqpV
yKNAivhpqFBFgsgVfSmq9/tzMmUKDLjM0pxBt32V9ux0LcukckT+KAg0ZRhlZcgV
NB8O2RNUqjnEU/+5hrHL1zHo/BZJ8hD1NjA+2qYinGTfTm7hkw2UFYTl1YHABqzH
9TYBg4Og3UIow1FGds6tK3X9n4UfOLm9XkQzt9158RSLwmq+lpF28xYu/C6lmB0+
4ssig6fkD2scVO6cfAp4gxUvXV7a4a06yfDGwT56bXulsnVb+Ygxck44cenXgEzk
ISVijGzHV5tvX9L/Xubg3W4aXHzDWx527DBnjigOImA2d+ydLUjGEZ6LiIPane8V
jGQ2jhOlhE/buaHSFjV0KzO3Oc1o8HkCcbllNJJ6G2tWCEZQDO2tP7yeoqv3L0/h
tLErVEIggdfLVBFfnqf4YSoVJUkLfXr+SFiz3HKqFhVtJwmbjZ79kz1/FY2lyMUe
v960et5dM8jMfwMJOpPO8HfA0K/AhRtCsXXODS+ezczOVD6t0pk2qu5FqQQO579X
du2cE7XitrfqdQqRYA6GKJ37kazIJ5kshSbTlkpTwQpj0TR5Btq1fLTHTnZnp52w
SMme3/Ct41PBsG1Y787jfwi2Qhd0k4LfK96h3xVhTdXJOEDiSBkZ3Fs+X+0NXuPW
E/6MEKar4MCXOYT6O5fBrlvSVgyDbejQUwgCG0EPFOa7HTBYYBDH3k5q+VPKdYjc
jdTZmd3JUxlLFjgXXpTopxxrGGkxuN/kqd+A43Fnz8xpgtyVl61/g0sKpVWBMDyT
24tequahBA99TT3l7KiTwQe+6zfYC+ks/Y9Ok98ia3g5T7ak6me8r5xj9INKudgF
bpwzoXdYa3Rk43ee0lvVf6JCynKYvZDdjOzR48PWIaSAOzsNLvLCwoWgzG8n1vYH
QUUEU87A+LXiRM5HFzbQsIWeCxhhgXUPKY5xZgAC35wcQoYbS8+wZn18g3YTIHrN
hltbUxZcCtbfsVTmB2im7ybqUselpBZZf0bxrWCWvWvGwLdzK8UmZhBog/G8iWXu
bBtQ6k9toyNk+arIfd1imGFRXxOGDW6JpYedMe3tG22iozui/8rjImhxr9n8GS7r
N8ILJjpjPLWPlMqBizp5CaIdGxmXR6r56UNrY+jL0xGwLnYzNAZ0VrnokyPy8QHv
1IMvyjBZlLTGYf1NJVv1KGD8lHX2/q8/gM383wI6WirphhQHrrIGWGBytm8KJ5Oz
P0KsHhliD/uxX+rcMFf1QeaJa26ZrwZuQifR2EZxk07HsYVMW0OCn2if0rTn0mjo
FlOhaLiQSgJCcCFtV5TAhJHj22UPymIi4H2CCVxoIu4I77sliPD4z3Hu0SfmUiV6
6ovMAbHVIkRAlnGszNuwuoKl9+SDJ6soFh/hfsdK54RzbAgqQnli7JLY1j9lc9WB
r9SqySXLdbEch05XTGus92xyO9Dh9SHndUG4ZpUN4AZGq3bruQiugVrCpK6YkBM0
+osZYm8m0g/VAFNrLA+OVDhKquoILICRED2vqj5kMo8aH8nxbE3oXDa1j7Z8Bax3
IjeZnhQaiRlXSeOw7oNj6nR/Z7rvOF+6Kckuh3Fc2rTo3f7zMUpgmHFuHn3jZOpG
buvStPAr3Oj1RzmNBVZxspvE9J4kVgCkcKRlf+eeitXcN8LxRKLhGkVO/Z+35X8i
pLH6GMs02xoB9wWBnl4chrz8ykYkLQpesIVjyC5GS4Gfsv+gJgFamJ1wjBghaXJu
Y+yvftckTnnceSG5GL7trX2736gEUJASpMthxjjopoz/5ZsviM/khajXzXZGe5JU
5F5jWAqxQm+K3MA+1BA7V05+ZTOGQxY4q5ndFIFqjc+QXNvdVo5ywJxB0hL96fbZ
Q+KeXx5j6LRafl5/PHblfzrzm6b5C8uqnCsDfDRNMeQv791s2R6l4RwXP8nI8XQD
Eo3sgU1HGK0toOlXOtryw8KKparWPo1Mcl0G9ca+z3E9zoe6BSmEW2oOMpew+yDO
6MFNX6HBhgS+IN7xMtzKqAVLNF0yTqyhR6BR+5ems2fThW+KUfRGLzDvvi9nXswf
5jJTJenWSvS5aqvzEb3K5xHVfwaUhKS2QHpQaxVTHi9FBuMKP8hJ3EI/60lFyoTK
Ebcuwho2D5rIXlm/Jjj3W82xYku8bC0Yke+Fyqx/N5MHCq9jM45H8folmKOsizBN
qhMdJtrvAyhW/ZgIXUNfl6jNJy89pxGyegMDQPdjqbeQTA//n8pXKdOTlA9yWoIr
ipaXFBNIzZHjYQwkLfuf5fuL7XSlD5jtq8qUzFwUamMrnt3dSTd8MzuoCVVRjFok
jzcLgTGMDKsM6cUwZHYFCLdUqfMcHMZGPvjb2RPm7VDiUuJiDWNTdiAuxfJiIp2m
+ouaGJXbVkG13pSvoBfxCikcNd3GwLkWf73kArYKeXm1ZPjiP5lqd5cBcZjTpppy
3+bhRGF6Gkd1ZPekMSkplmMUUtP606S983FiRxSRlKpnYRb7Wq90hpOkKtYDdMR2
OlRR2xeWrVI2sGxzz3iWsezfiitUy2NG+QqDHdK1GBqbwFLlBRFnRdEhAsbl3heV
/kIY246smqdNXrjk2YHw98QWOjwvyqJSCwHBvx75s0q82w/bE8k8TV6mONYotLH1
F1PsOp1CqP9JD2yT6343jEYnZ6tuzKKeBzkV/jr3Fi4+crTg+hNjq80Pa2gs9RE2
UAem5qBr5Df+KwATqmnvYmOcjEJ3WM1WZDKS553pbPjq1xZVftxg8z8/i664gei1
sPf2LJ2PZizry4+scO/pJDT/AdjVFWrngH/XdD3Rb78tLVXJpFdtWt/zEOW0JcjS
TsrDh1ra+obzOjnJv+TAPHFdrDnuEmEmf621FJ1ih/A1sCk5rEYHOxdNNMD44nip
R0mrojgYevy7oGnpQ91p3vUU5Pi2NlaYf6YNcSbrwS7qb0oAlPQJTk3ylWju892K
Kz6Oj0xwerlVv3bNCd+kfAj8qu611WX3F7ZjgSqG+nAQjnbePHk7hfnd371eLn9z
b7e7GFo0NdwbMBml1ssNtHcGS2fWUgfVeNYXezOC3H5XYEn157+evtNsLMkSHCVR
BlqOUPp09eE3e7a+xBtK5Efn+5oh1GEBgQnATKR6mdBtp19DCYjudN6XPhT+Abnb
3KWmvUdoQRgqnPYCr/84NiZzeTpxiih2PQpzRH/IXhLA9EUefFfjCS5SALvSOXkv
DFhT2JOgXHTYGlPRXLRv983exL7e0fIpL0216fc446j98080GefG3LVtIRZCxZdL
j3DWypUtZ4QhjmwKlBuj4XKVvAjEOJp5nRYwTvSPyfVB31jtrsi10J2jNxefx4Bp
Wo/iyNGd/RW8ajk1tEdNde5Yz4iiRa9e8aoatomgFMXelNJwj7LLO0zo2jDZfhTN
LF8W+0E+37VE/4aXB1Ps/gK2HaYC20GHLD3JxnkJy1Ir+yP6OX0jXe0dUtLL0ngA
Ht/AO8369Fv0OTxiou/QGsDqXrJao2cjxQCil9TpTBfz33H5TV5EUZmJm+4C6rhV
myrPYQxRUSmjLsrSmzhFpjJd1UPbibwFYhEyCYV1VMSyGTDngIHG5DUpKdaozhAS
HeWV6k3Vs3Saj7IfEAuaQXgCU+tM76fErDFstDHfN2czouSFbboKZOcDaBmm6PqX
Uef4RpsTxhskRbSteTzDuOKN2L0SJLE9FZ42gUEMUalvUOQJDLc1Nh/vcc3MDQPe
jU+1RisDx3YYewdIKipMooQlmZqDvZINvUTAOmI06Nxl7+LaMYz2WgybEN90k5Zp
/VQfPTFsxywCb4z4v7HLPWPGckdl4Q4LPYOnAMEBtEIWmIOqAQT1y0MigphGPMs1
NuYARGDGQAE65cYHRyiL3ghA+PBnk27pQ7H/xNg1bytjOksfRQ2Em40JqMsD6cpX
XnSMy8imhE3GpF+j6mrRjSUL81cGBwPWXNtSdgDVfOLqIlx5D4PADJYlXrVBhTQg
rpufarINmlEb/UdWNSfoVQkaJL2n4+Vimvo5tB3Ooys6uVLBpusFWu5CmgYlZdxa
bh3NRwoqRGwfW3iGW7WCw6JboH3XHkn0wYsazLHuTtZTsgjgvAfKBxYDJoTYexHg
mduhzD1HjNyKcmPKCf/BBYbjzGhzOL6e7+E4tYewvYwzh+IHnEAcdqFbxaVqRMeM
OAk8Lsa+35xu4y2x6PuknicgbkCee7QnOCMq+mZt2JZKbhNroLtKlJ3htRtjiuUj
WQGGl5E+EXgXZW3o5L5A1gUclMorToLF2VcdPX1uKFdIanxI36hmdgqZ7A/IwU1R
uzkvjYy56cF5BX+KjEeZY2iPA51JdkRONbVkWL/ZC/fZ73I0DHWlj0o4YLkM+QVE
2ygpiKaC/HuJLFXBfSXxS+Xcr8MpWkX8ta/tj5lPyX0bZOz3chgve90T7OlAG0So
eFUdPZy55UaNa84S2ELN8KarEY13j2B+uMyjAlXaF7qQL4bh36YFRWFWjkX6WT6f
+DOuRL6y+dfegp7x6Rw5lq0a0Axs9i65oMKGuQGvJZSgd8ZiREl4Ewf4jEb045dw
fsy3Nk5YRk91ILbXI8LtoeorJAvcfkArIb+5XJa/gHJM8gtB+ly+ZbGSbkPmq0Nz
STzyTLNiEEirx7zWlZSgc9vN+y1UF083YWHWrm899BL3N8ILMjRneDZjOHu5PwyF
S8muUk4lL6Cj8f8dZMa/UmD6MLfr+GkeRTAP2A0+wB3pEhrAZM4sRaPVHwy6OpC7
Hnvfh9DhIu282DWUjympaWTHBm4g+YeEMSdNNQSslIDAtHHNCDBJVW7DKWyBnwyz
OWQgEIHm5TpP8p/FqhHwJqIEbMaJcVKP6r1MlZc6uCBtqxUrwZMuynJ+QSTbTOkB
vBTq/m3cZXgGAb0fDk6TN5BTZVokw/KkDZ1UIn7LAh9FvKoyV1sC3IcyJepcjNIS
u7VU7yyD0E/VUKfyVEqqTvToRKHFx2oCyYlC84i+wrv991lo4ksDc0pJfD4NNsoo
ZXeFp5X/vq1QDx/VrHoNNryg+IQAJGPXPoNAf+gDdX/ROBWn9UaUsgWakYZyL2W4
1yRWLUuHLPYqzM1wacwV5ixZbuIf7pkzKJYFwPKjpHJ2M0EaOpIP8TbfNPqqmabn
gxP2BC4wQyEI+v99R2o1tMvSQUUaL6+TYQZTIhpYOIIkEl2JtqEj2aTT/3jf9rlR
7ZpmmjsOx0/bv0wAF//4rBFmA42mBzSzBJhf+lnW5MieTimB0TgXyPKFHRo3e4dr
tfae95uep6PrOT0tNikpIZrQAw2p2uCYepuC5sgV7KEISTjveGr2Xv5tC34SYE31
rXWpwi4SUBGCHXTS7Fz4LzgkLTl9JtDA/5TJ5Ok9kS2m9LXA/bszUoiJr+Q1g9gc
o+pYXf3oA6JnknzHbxK3KHItdMWOebcRb/xGg01nFbKI/rKEVlGcQ6kk1+2yl2uB
sY4zlGOuaUXVmseudxxeEUu44PviV9HMf7ONTrk6NwJqmTv+m5LHCJMdZ/NgaFtR
mVy6B5Kf4j4ZyfVAF9G7bcZI6xjJhLv3YKFZ28Q6OWXpZoqWC2IvDZNwN0kolgIm
k6n5tbx/1LXH5fGXK6M+BCTzeIWrTaCBnpZ5qwmsxrJnAsjYlIUF2rmkBLVUFHzO
lserLlCPvVbxIfnKSaBFqOV2sMJk4iD0nBEC3g+YzOjtF9od3NV7vJVbz+sADTrQ
vDl+ywbcR6TF7LnhqKY7GFPzA736aB4AT2gWmPvA67Dpz2wycIyjP4RWDte8Ith4
6Io7a6PbH+1DYPZsPhiCTcu72jNeEsS7sELl72ahRYz8z46SV6F7703NQaHf+gai
ZOCChNaBdP4K49ZAuBr1Uh8JTBxhTOk1eAOtImICwN425t8vRRXDUDfCw3dYekT0
d2gP8m8hCuD1XW5Bf3oSJ/DdOpdkqpIO2Uoc14u4uW2j9kr0qbyE+8gFxdrFF+EM
HZEh78xSudamj9S0A+sQqX3XJGfPRImmGP56uXyF3h1QzH0ZIzgcaO7FwMgjvHL5
alr4ZnLxbXXMN+a4UhPRnjvNwrzujgOAbp1h7fTOyCdPnOBNOlNEVfOUM8P7KFl7
LO0DnS0Qw2GR90f74mwL8smSuSVwjqLir5LQQtYbbdGeOUAP8HWXdVVQEKDzGoBm
M5vBLzH4olDlguSz/KbVtF6K7Wr+Qh1lnSkgaLLkmrg+y7Kf4Qz0FImGCMl3oTt8
nhIGUlGMCnPfYNPieYKiQLOYbF1DW4h6M5terlIhSch3fXSNgB30qPgRcUjXWRZY
KM0gU06fls48FVInhhaWvwl3o9wcs0Wz5Qj9abT3PWVFu3oSg35Cr4ddW0SfVBPb
6f//cXG13kvx6ReqSUrKz2m1NAH1b/Q3TXlRJa7wX8PTze+mYg2AEQMIbPrDLkPZ
Ub/9szJj9Ifh4wWuw4poLKLx0jgOoYorp6e/0aODRX+VEw4xDGlAGVLHPzBLZtb7
EwWaLLqjttxf+JdtaRGuaGTOPQyjZ1tSfFJctrwGjJ6SqCeS1KcWA47MVNxmAl6L
aE4DUQpxi+U6tKGrOMJ9YhuVhcRtOKyngiXwvO+qgcg3Q80ynv25R5x9wGgl8+mz
kItrlZrqTrAX83zNELklUz7pPinBGlS4ctoWaAS27W21GMUtZPwfrBrFsRDPwIlx
j1z2LpspZYj3WzoErSJSjdW+l9gHi5b3Ofve/foD2kTVCwcmoZ100Tvwji+bbv6z
TjMjVa3y3Ajcm44py3iK5EzW9FLSHjsofMFvNNohqT3As1TECKqGnWTtAgk1FaZh
FMAfQyyMBgDdL+suE1G2P5TM4FtalnPd7ufY0od9FZK3bY0EpfwrvulFEM2iYMjb
tnvhWtxDIjYlTaQTTg/unSf+B05ZGXHrueD1fseoY4SJjAgPEWcEO4MbtjqHiUTE
bIz/CV9EUXnyTfk9dKCxptDsVYSuthbB+kpKGT9SdADNeltvtqA18eyY5guGKyyX
2QkKvHmNrVeo/DNwwDFuQXJaT3lFa+anBb32wJLFf77mrJqeLI41yO0N/Bt7m4bJ
OKWzo3+JU9prVVzgAt/tDKJbh0mETXlQCiRsWUUY8Nmlm6z7fxY93yImuulhHBYJ
mybgqh45m8Aj+OcKtT37rWcjE9vCVWiBAgAzdUGWPBeanluxXdKsHNLgajdIyXmr
InL8LLDYEqmPMyRF2IunFAhy3m03Up54t3u11ZyycucIjSOXcKLubNX4yccYlCyA
nwqRMVfGLJqV10apxYNG4BkFG+ZrYBGs5JAyZfkJQSb5ja1eLCLbefG9XW0xTbaS
hc0Sv3+FHdpZ0MhUJfBZNUweDW4ljipgvfjnL521vV+AiL/FMD3XQtVzdM+jJn95
uijM8ApkHUrWgsHjoYK3FqdI/enPNyYu8uvHzB8wkZT8lYcraBjK28V4nGZnety5
R5FPQbQNfC0+N0ozPFdSo4XKOsTILc1UXCU/Yw79IUAffyuVUCkDG6plpfbQdPnp
II9bbrZ8+eOPLIjlSj2yDXahCUMPixKFpKkbePsyZS8cEuIEZ+jQi44PpDLUcs9R
PTL7tnsYh8nWViQxmJDQlvHGfeQ7cw71Tj0encAXQj12sHVBU8OxtlZ3fePyMsRD
Tb75+cZybGhk0Cwn2Zd3ECSW0NsZC2NialAvD2/Ti5sJfql2DiLrlpEdsZd1xWEf
BdGygDGRtnWFZ4jds8opPpl4ldo8Ux3QBs/gi2DHNv1feKEWH2w9h1YK8db2VGNt
STs1N9UgNJHmT8JGU8aipKSERJXnL/CgQBk2wsx+FRs0wY/bF9cOaMscR6xArso3
hJe5+fhq/JhcgXmCmYgHKKw/G4p/MWyXw1KLPuMYmhubtclPLx6051lXbcvDcDu4
nvgbsS4MDRIBl7kpAp59knVe+wdA2qSxCJ7zye7CetAYExN5t5RHD2NUVureRotO
C5Si0Tp7x7LM/kku7QvsGWTTwuKPvqh4qiL6C1fdye2V9LKMFBvqv2Fy1JM1W7Dy
MiUgyctb1+pFwCFosDz2i5VaQOLlvsJLh4W+N55jFxkOak0z0aaG7h2Gi2OL5daU
1eufZd6CizbpLrDUUoSkRanHrbjKRCHU9zUmNyTizGOnFgcX52DNkzTooLQ2M1Os
CnjbBPshNLPN9f6sFoF8vMuv+CdBCDLxdtZ8+pWjg44mB4rP27GXbR0nzTvUq6IA
pr/+eISFV6IiAHfVPGnjeByhr5W4l7zlnXDtoeQm3vmkleOGKKBXEhex5ApeOO0Y
o/K3o3F0oPLkIqhte/Dww9MLPy+hCOd5qb5jq99WHtawsn0M2teVj/Wd2ecPkqNf
EQm2/Ksd9hUQTSh4nGdeQffWXggIgkgAsJTN967/QUtMSLyPLEdLzZ6lX1DbfGL2
xlgAwE5SBz2AM9tMl8L/GJ9zYogj42M5fptDG4ZH/ntHT1IEcnNmurQt+nP8Jt+i
YnPJoy5g+kw84HTfTg9iG7OpucUjNJPGd/hDzJHmqyt8kNAVo1lxfgWlmA9RtRhR
NkLLFzWz39azor5PPo9PL/5wi3Ni4BqgsDWv9VsLTlms2u3dmBgn/OtPg0m4deIZ
92n0dQ3HfUSKMIwocSlm+r8wNZPR2xXnUBW0iGURTL8G1Bdsfm4Avy4kDmKe5GmL
bm6v58sjF/payqQiYlkmyVlZsJ8xTIe+GjkKgqy26rPk8q74j2jo3W5ZxDFa/Abn
W4YjsR8ALh09f5hUF8X0p2YCPe+Esd8gRXzTuhAIS5kqdrKFmZpRnG2cSBrxuEYU
mYnX20HWwSyqlN1+PaV+JolKVMoovIrVxP+Pz4KfycQY/4NGXZuNcZMwL7jSq9Lt
iuRzNaM1Kc8W5QU2ln05roRzSAqbY1yDWTQ1VkcAxwUxYZsTrF884Bs0H2np3Ck0
dTQm3MIHKReq20wveMPdQ+bnaMnl+kdTFz75OrwWlonjYTIOS4HR3NTtyDqzjPjS
0pGkwlRAN5/eDlNQqPOHWgxas3C+eKBu6EtksgSR4Rjc8vzU8het3GggA1+cWhnv
piMW0JhOMns7IDo7in2vcRfE28N31NDSWnyakLPdLno/BNK7FlWBLZINuWxlGcYQ
e2UPdLMt6pvCdUAKO33F3P362bdzjsy1IbtoprxzU0dRcc/AoVac5e3cEh6DbMC5
ZS6K6N78rr26OoJ4mA8oppy7UAgK9jP5JyM1UhXKL2G/30A2q5g6lCfTs0h9G0QK
8vTRcXHn0Voq4JkzNB8vq7okNbkNy7O/3vQeyhlM4hnDVAXjcH/ZyTmUPqxexpS+
tEKO8F7ltooqWusaSeHmCazejk2tA1cCEtjPFa69FDaQu59HEqiktU/6Vw0Xy2BI
5GzSHzt5fsFZQZCJ3YXnC9Vfs9zzH6mLeYEOkNnrxPWPKpfLbSPxuy0qaGE1kNce
/dTAj4JAcqUkvnpGksvhdwu020xwXyg3t6uFCiUVHHe8CpNFbiqNKlz5Hsm1D/Jd
djz/O+EdL8ItcXs0shbVoV/Y3aB314f/XAf9nwded5u/aEE5wqxEePsWADPA8qeB
FRpOs31Guqi2q3N2iQ3OhOVoLDy9kwzwYXVcmt4VuchHBKRhaU/OBxF3GTh9MqlH
VFYaxYJnsFWIqbx1yYe+5XPkv6nkVALxcz48VN3MqbVNmjJs114FVjCk1Ua/PbZU
lFyf2JZAMmYtB0XrHAcoNr2fUSa3J15RQgqZ7mmMbdgkPYmhBdvpyd5Y2wmc8fBr
r2U6Ir1xWCeXDUljgL9cpW2+jkT0/BmsYz9uR9PtueKOGoke6VYg2kOClAos7BD6
jEuLKESJC0M8H2CUWnlEuC/0xiRb5y1maxRf0HmkdpBrIDcjVuov2+IWNXNyWeTj
AlT2rhX25awwVCmRjGRjVuCBNU58H7ZffVkkAX9uTc9z+hGnd/2rfVcqVyr5gXPQ
41fwa/YEqhLWwwi1bDI5v7dpJcByZo84QPA73EHurMBsoB4SIzNKgr02hkko6NTi
VwX9QOsVxWTqDlQqjTfxsaLt8L3jcdlZFVbBeSU1ZHX4YFAV05pu9qbmTZb/kRUX
LaVoGuxyxuvKM6cKDvM4srrfPyQ7Ivhfb1BbWaY+TksmOLX2Sep+lkpYNHob3eeE
fU1oaQymARgWULWRGBxWz9Qetyj4sS4L67lSICQhCq0WVy9TjZoXIFux5Omc/T/m
B/XHCBamfHB+HnfgkrZN3D9WvQlCCaC11XFWCGe0YJD8c0SIyhrUJaQfB4YAtoZG
KasO6qGBu6RLXypjy9yArIxSxPNGCvG06l/eSf/AibzU5ISvNL5aVm8cAucn5+2f
GLnwlEIlUiGmPNqida1+9Sb9UUDPzhNb4xFc7+Ql0bqO+rYE1RUX6AijOgVNqy2/
KJhemUJ91kAhZhpfhESVrfVzoPw95ip2JRzgjJtCNt7V6VBorEDslwUoXqgFh0dh
d69hseDmf7vqc8b277obo4WFkd+9j2lwyjS2WxP0ooCRTW+1Ee8zhK0fSwnoPXfJ
sRj6eZPgtpJoT1tQyiB7vOg2k5gmgjkYOVwSxTeXTjurhOirn+pOumU30t2LZHTi
unVuEoNSvf+VpseWtfsOy6vMOwqHszjByRdARcGOkqgp5dH/yi0UGi5erCH+bfdr
lC3KUxCl6/UEOKp3qjcI3GCVyozapTAxUTCSAEWtGw+UbFeS3Infk1uo93aAP+cL
26rzFTNi00LOrttA6dzaIsYS1qhCamCeAmhd/vi8w2Y25Tipwwv2Ferw4MnbNAXt
pjz3/FZ84WUTNMwVaZx08m+KB+6ZgYRwbelwDOw4BErkO2PBd+7Ry6zxNus5vcGM
RJuBtwPa3dHVljK9B0MKoKBdCXeADlJ06aZh1Rjs8un5VTd18RYYwsqKLpmv5dnv
b1H9PoMb+s03cGwbSQQ+xfjAsbV9FwZH5egkRv9LOGAR3Ks3+016vacBjlAWe47z
f7wt5QEU/AwiPpaWr/T9/2P5MzDzj9aGOAmQaxOf6PElH+/5bMgP+BvYa9zj6BEy
YDSFeTngFimZs3MOI1UJicyUAqbS3Kl7/plBOqFQTM6lKr0OawgoK56aTg+ND9m6
32egwEKtS3li1CV1pCuwKhSI6KS2YaJOKt7vu5ectYIkN1OyIAvkCkJS5BY/jNcS
WlovP9FKvJP1sLBWKj/BbaW6evWMSjzelRlpirBw0O6jmh2ptzqL1fUDOxtxXmbm
710aFiVl6p+bJAB6xlmQADu9t90/6wYs43qRgXkuqFILPye0Vr69Qj+ermvef5FA
qdHjW9gtYfcQ8UsUale8VFjdLb3OMQRnCeDAyv6bUCvI0Q0kfK4V7/NnJLH45OnV
GYWjskJ6FdCVFVJfO/ks4t4iqJ342ll5Szn0rcLS3e7r5i/BMAw9y1M3EQaXt0L/
lH4GNzzurBb7VqDXQVmY3RkSQaeHt//gi+TGLsIDDy7fG08QdJZVJav46PE1ckI1
Rmes5iqDTHNsjivIuqn3yqqCltg+Uf3U5Vppmqpqtd5RraG8MA7m2CrmE/pOjdRz
zYoCYi7y7NFK+kIDrKSeZq9eesvYoyzjCaQ+gqgrqkyB/jQKQlStyp5Bxi8SyJmz
94mpUQ+pSOUNqg1akn+Flsh3oGN7Lf1t68qIpgbxvXTmFBdx+7ePbRpWRJV+EibP
aObmyMM77UvJxPhugQ3oA8ykWreYS4/X3tqom2JhN8DJUfe06mSzmUD788tLb/RZ
h1d0cP5/0733tkyJSpRgEGzMpGkL+0h4NMmtPso906RB+3NOVA2axcYksci3f7dG
cJPNIXroQ32zW+j2eIsB7ftzh/dinyBpRZbjSyXkGvzTMBZaSr+1M3DKs8bDXfKp
nHqW/yZoOLSTrGN0dxYO77pYbPWVyxHBvstHhbPPBshFMbQxJm07JB1QMBr1fdnf
dLKRrnLnXtLsaHvpgkT5XFA5u4jIN8VfO7Ayrawm3/RukKyQ+2EZwG6To3Q8JXy+
L9rBxRigouDqA1a4b7u/KqwOOvw2wq9LznIlGGVuaUL/bInqWSexyGoQyaA9cVlz
9g4kP2/j7BrxnFe9gyTTim9IywszFJoQc7Jo9mSE0YyLpY6xaA7rMhR50RNGuf19
YFq4b9qhY5K+bg+88ynoAUIAnnMWZZErh2jIcX5t+XHuymtUBsybktrVZY0BXx3c
Jbzvi7iMBwLIXxvrRJP7Kp60Pl7bHZzQQFXYVFvw3nMw3FBhL6b8o6JWBNvP7n4p
uLtkcbHlBKrihE5AY6u2uzr/o26PkGTv/Vsa+gO+zxZgA5nyP3jqlBFi8fBq51V1
Aj4cdvVJHVl3bKIf4+m4z9wix/hzw0wA2xdV3E9kGMEz8jowLMWxOzMYrylsvN6g
WPZNObV09E44kY9hLOC9nQc4IclfTD6JshF7k7NJu6ioFlPK2vemZNjl9/o9MmT9
4GOqX3yKWhAd91C1svX6ENvoiBoQUPVSTOmDnLYgjyMz8yfKFG2N9rR6ODoBQeK2
99J9rZQCM4HCBd1pa/lOEJPZ3ZdojRLKeL4rdk//pmX4i4QIYLpymwSRclTamBgS
3tHOx0haD9OFK10hpVXDMDrMURHRwrVWu3aK6ZCrfDVLKzOsAQ4h7KWTISaZjCWK
qowKC/69ZoKEHRKJVQkLkHJJc56Iot2wmhvHwQj/u0AcUvL/n/eqNlds8S/M97NT
nMrglibVNzpbqcUCmceSeDCfpUvneUMGQnX+lwdrj1r2KAHz+jpfugO/XAgdxk+O
3KI61nX9xdoczOLmFdZ/Kmttj7kATzlHE1dgAyJ/VxMNzZ6vbxhDd450PnkVxS2b
O6t6aSmoWgR47AFTh3seMl12ewxZ1/jMzdInVH1mB/xCVJmNqN7laHlElyWU+5Xm
xH7Re+/DmXwkDzzX7AhwABqHPiTntj1iKsEi4MucdLzHwZ4lqn7b+Gn3sI3tdHxD
bYIHN1l6fN9X5geI69YvDzE2K31xYIF5eUdiNsZimPCAYUiCrMAq0jKXCnu6pAIV
w9cdbGBGzQHgILWRzIb7GtWysxGp0+SNzIA7VWv1DVcAdXqCWmJ4DR+Ra2Ap+6hX
wBJuo5gnR3ZomnqzLIRSx4W0GzQVJNDTzL5wNYtgRrIeRL42j6TbhvPCqB5lm7qV
QyKAzUPspRbxBP9B5RiH0upwjuNrue4QIeTVsXODOCx7cjZ3C+AqfFsDpHO9+WMo
wfRSc7JMFAE/Akdvi65eLN5cTn09K9lBpHMAvZPr9lniou/wINRviHaDpHiGn6D4
Audw3v9V+12wB61mZWKRtJZIyaBs6GSlMPqraM5tnBSCDmWLubnx2KkY1iCrX4gj
8cnILHbTkKTptxEB/3zbSi1da7PV/vEk49zBl+3Z2JXtNi/6zei8aDfOpUBbB/+B
2glNHnj/BESCc68TPVk5dy2GiTxAYjx/Di0qLogEyEq8V4/Y2Kkrk++pJit1KSDZ
LoI0FQuKe+C7neKJ3Hvb4lFkX1oo/RjNJBUurlsa6vsgQRXJkhAW43ki1O+fAz+3
QRVTLNgJxR7r4Rasq0EQ03u8SNOS5thUMKlAZtWQHkfBfp2kXEkcBJFqSOiwkr+X
xEFp6Jb45icyUTa+8MAHUY7Axv0E2wJ94qSmBYkSOPKiV0S/ZTmJIvTd2EkQMyGM
ZuDBs6Nk8CMc5vHnmyPrr0gsBk0dhTiKk6ix5FWrzrLGI5ZTVcVHZFDGe7UOkDl7
svgCkjXubBsZJj6i5FjX2lKeJDLScYXvEFhrZKAPES4dtNjLtaBzHyRxa4hlc55s
GVfYhoXWmactZF+m6l7aYrOustIHM1L5l1jBvh/SQzUBC2dEdee7/7IgpMpSdBdT
umb1MgQkLm4vesBN5k1luGmSN7dao7+G5/N5z8jGV7YX7/seT8+rDbUh0RqRURdX
jVzjKipwT3gjIDA9L35tCfNqBxqH97tWiJ5lkQzvqCwth+5PU2/3nUqV7BH6RH55
deCct9XbZ6DhcwbVY50QScNApPW+uYAM0BmFFI1hC6anCtA5qpbOHVUS/gPyEq4h
l/5N1cc4TGbiixIVOEi+yZDrDy/5sGN1GtW8DabQjOPsmudBYSPs/7uqpUP2HWjX
hr2u2qx0n322pLeC/YEyn9Z0+RGOeAsfWQOsH6IQgO3RlvV9lXJ7ipmZjebapCI1
BIPUcFWnSacOGdscXorAyLjereP7zpWvDtmEnA6JCfT4T66jqBH88uWYzczRZLaz
0DvIEmOPnC2Q/ikdo99/FBIvux2u8+bWjg3zzDLMbDIFqRYsLYBDTLmnKBI08Mcj
MVoccFs7fDHjV9oNgnyD9wLa5PTnkGZFNvlygsaUm7HGFQAW+4ihT+FfO6cnGpSt
4q+kar5N3U3FY5WvK7sqltU/TTaURE4hhTy4I9fsPCEqs/DeJLAIW+aKQw4rWEnx
xDw6TGyLJbLw6IMa26J1LfrrqtC1j2Ats3t17M9XxSOaG4wi5ArZ3ikloLxvrULO
dnz6rzLKW4pup7LzscLZLXkAv7JC9Grxv/4FIhDJQBqtVKFPOW7mynQs+X+Kr1iA
VTHN75gClZ1QCMzxXPhj6Vj4K6Vd+/WV3nLO/VXuPBarV+cWJyzx8YyhOAZj6QWw
GnBVFJm2VoW1Oj06noikUrM2Sr22RtBi5aYNBCG11gdOBXHzHJgC8DxbPftcO6PN
ajIDuHFuWEtuBiVOesKLV3qtueq7KEl0ngOerBfVgrVnHZmRb/KBiRD6lpN/bzj0
DSexeQ3MYD4qJnKHpJq5+ga1XgfgZqhp1QnFvQIqEJo4cLTy5R2ai9STGUdfEGnM
4q8VWACgJyzCn5G5tEOCOfb2xdRmDbPBouEQgWLbQzY2GxgOPEnOSoCsdIESV7sm
MIpqJB6xisGokJMIGVzswX3KRR/s03Cwax9TZD7+QWiu7HdMU39xr4/Ebf1Y2nEp
/DG8QtKxe/Lnfq2+qZN6eST6p9M7iD+1WFZ6ZxZPiX6EjY11trhPVSbCKgclVwcx
evRkPBEqw+jE7tSXspIKUBXrW8z1wdGHl55FZ57fAo6e1EkmO/v+arByhd6ZzBL1
KlBphnq/FGD9ahqpKBsqTZ6zToiFlum7JkqFoAs/CsIVGC3i/e2asXA98pdEi6XR
vYnMXvxmQVF+khgl0LWkDmdLetAOW5qlmQ8OP2evuZuqjgbc8SqTPT+/qsrGoJXR
OkxNT+O2FZWv5+oxqeo7idBgyDLcwBO3JADP85R34pmVcCwTBiIXQNuHankgf3XR
rlOOoEXcP4ftC64K8nq535Ex5sNfk+SLGuS39On3vsCfGZEXhBljdXdwgwQlaAcW
oXPoN0waMNGPa13ay91iqREsnx7O9il8XzLMR3kP/3zH8v+3O2dBA3cisehUJoYr
JhQZ0r0qG+DgSk/k/oMc9TdfiQWjZ9siOw4t9eGm7UOpC8cC902KYuRtUesPBkVu
qo/Y+nYidwhb/CTXpeZ3DZU61xtSI8AXkHwivRCmKSkyV4uDJ/2n0x01FLpWwyKr
+gUl1PsVF6Eqji6CeN4OWarChKi1wveog1ZWJcOhvCPmdyslIbt06eJGtsfw8cbn
2LrcLmneTC4vnge1I55Xn38GlLHEvtwBIUZUhCylzaHjB0ZlLa7un1Jpk5b7978h
oMTQDFmbzguJtTcc4Rr4LFECY70ohYlUwWGZhTwDJsYxexdGf/s8ufRd6SEknt02
mTV974hz7GR6ih5whKn83NEX3La4gg/wOidXWvsWi7qxEzDXIpy/41VYQg1v3XOL
UHKmPgz1S+RKo80aY5BGUHm3ZFEjCrk4gz2FFJOLSDADhTfdluqanpAgum2IxWJq
6/cK0mrnZH5Plj9xlFihBwNNMB2E5cL+07i8kNgfPrb05YGBlHfri4iMlEI3F+Vb
LzlrHAKp89ND+QwAzNQDy/muEHn0ByEa14S2hlMDR+WA1IkTklAsz+nnJ1EOImVP
iYiLaYsGyYU86Z7BxmLFt3+4zXfE90ChonE7CmQ1hOh4yBKgX2KI0tY3mlaYWE36
+/XRqhTJl/HqUtGMpm6hz4ut2/6mrFu80qQ/sNIPHAnz+WAof/QCxziOsvrrxfxA
dyWaMESFRsp1adCYoCWOPNV9OPqHpjzv0iVcJ3DFhnn7eKEaYeTlm2x0v5Y4HAo8
l/1Tn8pbnSf18Nb2caLEjhPB9pTXQpdjC20Gv9oYmaIc26D0nRM7O3uWrPWEW0l2
11RaxP3fF61C+7Jd3FY4TRB6zowX9u8pKkZButiFAiSpFHzOXHloeJEgxRrX3CiU
txn6siKaWMgN1SZ/FBS6sfdcZ77AIyleqNBk9yA9QORtgMSc+xeG6eKsz3/HliG+
INR1LzLUwQXFXBFmO6Th6rxWVWao8mCfYxUYg9k8wSCA7VY5ENtkn7AEE3wjkJ1F
JiOGEuEu+CN4OmjR1i8Rox2BTT1FIeGkUo2sbQBgGACzC57mdJ/cyQ2Bqu40UC3y
JU8VBtCY/WLm4p0Gs5mCWv6i9rqG5jp+oCiOn/+NJihflp1W9I7DG9Frchr5nml1
HG9tjJDd1C2eQdm5x5fpbFHhoaS9F+FwPwEF5UcC8GQEinTBwP69QFoyCDoJJtx3
PkT/NMVTCG04G7e+BQ0+bFxWc9iQ1We7+9fp9BPHpxWYmR7sj1QuUk9vnXnspUwX
7Y+FDx5h8hREpJqKCP8fy+XbPX7Z8oT7cVlEVrFzLXyKwdgSSEnqIlCBZjXTQ5KS
TIL+vx2OAck8bZswhQZgXic/i+aZlMGBkdVyrVRbQEQfG9/IIi5XcQTa8Fjbqr63
cnFdHieZDbgcRxR+UOSAbHEB78UE2KxLzNVI7gZ84ZGYCMINaKWHFcqwRdwfZ+U5
Of8/t95LqF/07QeV76+4Qz7Sr2p4dZiHyHAViJpJKREHETfnltQj8Wyp1G3D4oHg
gRLVlKxP4Yaz/m8rbtBEpHKicYrSb7C1UpXLEnWcK0GeCBJDGHcJRggcExi4Kbfl
AVQPSSSAVE2yCNLB0UBuuMikVP57A2ZDKQCugMq/LweX2nKtYULEb82ZFQSCzHoZ
tnr164YDvu8iIgeMbcVRvgOwM65u0aisJgEq00u8T6RBSUZDO5ihXqu+sNFgz4b2
6ti3FP3PFlY83kBtGsjkpvENP2FjImnrGe7fqcveZQoMwmEKgPtSG++BXzUIDL8B
tvBoYP3s6K5yRV9UEv9KcmVaPIkdD4TFLgujXNmaxeiymbyE/V1Erm3MCaashBEc
+xZAOEfZATT5XicpkYYOcsDt4SrN9eOlgBhKWRZbZbhQy59/0JLcKg8RJrHgz5Ur
QdeqAchlJWvVdB4ohICqTTiXMLFJGBtk2KfDdODS7yoqgnfSMjzq/NPEErjaMXd5
xu5bIzCcZOLaQqyBsCkkksECm1K/VpM2376HYHkRKAlXh3JBb2NVoTThM+8K+HbV
nfgjVJPz/xISk60rLx8Qn6Q45c0H7RPF9Ywc9U90OBowfJ9vzqqL4hY863HWekpB
vLr+4z6J2HFmw/1brd2CCWc24GnK2nbTMpyDQV4JzFbV+MZk8kcEU8Qd+dYVEgLT
+mJ3ZQxT9clxRevIFJJbqQ73vTiW8aHj3/VGLM+ret7AvHHzCYWaVb8Q78YK6ry5
eoT4BSiklV0wZSc+mLRlKRJcvyuKJLhVyCSTCBwxX9B2D8a97Y717cv0LWORypCn
YjvsRv/1jg0IlzUtSnpTnsM01MuIKYYcpAsQfUC/CuOne6HQoVnMWzyGlTDhESaK
u6Y5zK9G3jmN/RlzmJPRsaZ5I2JVQBR9rEcHgfLH76JfZIi33r0lI/QiW43HJrrK
0jQ6TYndSxUYKtXo/z9w9V/JFTXKupcPHTCF/8NjA6Okqa2IV9yqjYYmeLAC5prH
QlIJwAB6KPiUuayWEVpGx7r3e/s9m88u5S/NHNRbxnQtGlRGZKp1D0s4KKPx1tuX
B4DXnx31Vlbd3VDxQ6l4L2Iutfx4vQeRgAGmZotZeMF0uEvRrijY/m5AM36Ueq2y
F5809E7Jzhn33o+tP4PMRUGKgMtm+g+dAu1456gn95LVb1rumJ+HiEFXaeN3+m9o
Dgjdodpl2tFuIwZ0P60g3ZP44Ok+2xdzhOQWphGTADrdv7HQYNu/XjjOU55cj9Mn
CiX4R1k4223niGux0DQMMESBPTv0IgNB1mQkCa7nL9LX3UkvqYN+FQ0IyDh7aJad
C0Rl7x5gDP79EIBtiU/R0d0WJ5jV5MIu51ve2ck9LkLI0I6WG1LcTSD0PJEmWJVl
iaU0UyGDv6QoKO48/vpuxU2GbdA093WwDbC6Nn4Z9UPI4gpbv1i3mPGELjjNKQD2
OtrUxXMbf+UT1EtYAfykjnPM+VNhkLhJUFC26nahxXBjCmXPxMBAN3D1K8cjas8N
LBIno/BEjfBIOIbULxS9h2CYMpfs/XKxTD7PI/aa9E628AbCLUeeb0gfidKoCYMP
dCjqIFqRh5avjAdUDmgRbVuW/TQwBRuRgitmP+C6BTFk1/KhcCvgWWQTDQfYyc59
M9vNT4sX/NKwP1THWM1H5g4zzTSAOupG1iiuRuw/yhSiObweRaTJOQUyyPsK5sfz
qPWFIPZQy1RhVYu5sZQLfr/0lD1P9r0naOzCR+ACZrgjgHLJU3If5x/RxO3Dv7+V
+1b6Cp2giF51GWsIi5DypxoSV3d6RU40e8l0AReffDF5SPbGjKFoTYtipGFk/eu4
acphiNro3keBmyeoINLhvd+bVjwGhoQ0u1RAOFziPjbcw1a/Lln0jkhX46S3FRQN
8xhvkleprButcVLb581tJgexBUXX4S1R5mq12iL5yg2oYLynbXpvLsRRFt41b8Tk
mVDtpF4Q0OXdxE1kFIpFwhFRMUZIBRtNMHmMr9JzDCXSIxoFPzGCp9MfaZ5ib7T6
sJ3PP1SyF5agSFlocmtwkL1eCvf9gwOKqiO17ze7FIOXzxB3EUgSnG+rfDJxBEkj
h1mJivTuXjthlW0ERQK3qQcpLqzFB3TtDWDXPFNmOgkch9MwdYQibNPsHqBfjskn
GSdXnYee1acfeU/La9F96MBuod0ZQA6+CcGBdEKiUGycEZhLYP+uvefl1xgA/7zx
mLDxLvU3/vQJSILBcSvUDg5U1+TOHRh6lftIDtN9xjMu9eIsbM3jzpaqcSNEq9d/
V/LN35qD1eqLDySVsiSATOXHysO9o3/PLfv9rnSg/2bgfqIqTDKfh84XXgxXaSJw
A6VQ+W11aRlAmpBoevwssOpXLvG8gkT/cuW6Gzo4D4zCcm8MAivGLeThN0JSq9uK
7IrlOpUxo+P4ayEcPdZedluZm8+cp23TrNC5B+n7iVSzOt7iVgTC9tZLRWQGF3ft
2DSa5fyFIkSYQn6QLaFHiiXNZZJRvPSwgAhp2zL6u79gYhwwbD46sEa9KMS3Oc8O
aZ0on+IpKDxHEPp5xAdjw2Nxhg8EIbxwpe7dxJeo3hqcz8N0oMDpCrbl4I2iEw2R
0nhKB775znqNtutFfb+OoCZQ3fxbpJXawA2Uj0HUR7FUESrga2JJL/gfR/efUaEI
wOxTEzGvY+DPag6Qv9faWl1j8dnAcLzQNWoIEpVM9jFMEpCsNRxXfNGUaBhH/F7/
55Uq9NGHxAtI72H+64JfAlkzP3hjIHw3ncPhpf1KpOMAFNllOpW0jYK9EjGvTFal
2+6UPo7NNcYqVSSIh3Jv8nNXgwNuZvbWUavRnLrNuOyW0jrnoqVcstMV6mGQ0BS+
Ldnj2CQseobnmyBfbOZNwIBSyluDTBVcP8VlMgWP+a5o55T1gQh/eMcJ8Q+8elB3
bL4hZ986K+8tErWJJHdxTpeITRWhq1GvTJZlVNnSedZiIAfMPQnKou+PiSlQa4lb
GQqtHp62sNUgJiIvIJRn6BShukVyn2uI9s7Xk4I8nGrkw5uL+L2QpO1FqT8ehFcU
Ek3d6etrVf1qOgDOlUWjYEPtjGRp7IBMv2DPjj6Vwf8qGEGeHo7nJeNwonj0U9RH
qpzDvnlHpNhrtg0sl9h19oHbFirQG8KRDTuthZLD0OA4uKpwxrqlJ46/Kq01XlY9
VcVuBcKUp05DdZYnJhtSv+xH+CZjWvfdWcexIGBaUFU2QGnBP8rhWMoub7wT6DzT
tFDRUybEijaA+ycV/3LOPqsaPsbWzsPvrityUDjuiCPbuNBSFgPpbOa8574kJibs
ebIx008rjQLgHwitk+6xx7ZL6qtK2IH6J+D6dma3ZKg2GmVhME/zred4rGzNmuSd
SrTldr+taO4YKih1SeYFt3BTQ0MO4REu4+P0JVOPg0raVVIJR70Y1S46coLw1+UT
LAnBEU2WiDHA76VzjcA/QpTQA0MBt+/YUzDOU0/XFcMiQygu8OrnB2Vpd0mRCcx5
5bn2PTj53vkdmJG3nQq4twFOnbThjMNQgxGJpG+6HwA6kL41b5lDQYcYerT6DpK3
Wog4NxQXntBy1ecoyqYHW7q/vGVk286KjovGziRnql+ZipfSoLLNmwdlTyNrE2ym
smglgg9+TCg+DweAGAKaIEgCxkpSjHts6r83ppE7WrK16EKuDFvk3mRpeLnbMSfv
LXSNcPDjl5+6VgZYN0hHCBZjkqrksXeId+r8lRU/2uA5E34nxC59PZmt3WVlXDlJ
Rawv+DvFu66iTkSul15YyFJsAKveMA02MsrpcCRU61ViBh8DwhGRh7nOAohZ1Lbn
9dyDX2soP64pYO5RfiE2Kf63m0MU4PiYex5j1pEhRooQGVqKYHp6Ax8unvJR6dvb
0r6F0SR2dphwVcU30CqtQamGOJr0qIdnrkTEA+QZUjKc5pnIoSnl++CWw+O8IuMD
s7jNcz7oLAUdClBxz22IxSnW22Ei+M1WocUsFxSmFQF/GoseNpXoCQtWcxC1Z0U9
Uxj7OGTecFMKscA0JZdgH547p1MBGCGqIcst1MsPL2eD1IzoOqBvlm+SMXf0rGA8
WJReFi35PC0rG+U8H/ketDZH6Q/X96CW1tfh+aplPhpM9EQzM7/lID+JhqVDn1Uf
9jbHkqe57w3y1F5Mcc/+Vlamwzwxm4qfN884I1jHTQ7LJestMI8bB+RkIpacVh4B
7krP6sMq9rUdJY/1tNCLlOlwc6tzVeR04ZshuSxR9emsxWa2u2wm3+vmYR8s9Ucw
VeFGM4znwzEXAiF6eHQEP/3PR1L//Mx5h2MfyNK8lYKooO0kVHqlzFDWy17eIY0B
8WN2w15f91nETRxgXwBqceyX4ldtTJ14+7sSfplds/0WayXsK0/2WjWfZN6GwTtO
q+ioz32GgfDYLkkKEZSSgqbvF6xzx3OA4Q5v1QfT3qyUrrWTYqg6DSoQUXSQepxg
Lc0f7FVMqLtWxU18z7xqX2B5UfSZ6IWvDA/AoyH+HzHQxD7AhZTqGaklFzuWzUNt
PxbJ070ztAgni5KztJZOkCbJcoI9/OcoJae5MfVoSKyCRxiV4g8iKQaa13vehMQD
4Fl/WayEWdpoNMQqlsgG0XD0tGuiCFoyScSmeZp6o7XaBRL2K2P4I+CXcVGufduL
NdlJzwJQNQ6pDy7ykbCy97XuTBEAphkWt2m6TuHctDVqhxt9ab2WSREhZZqwYHSC
vV8WR6S4Qym6Ot4/4JMCgzBkjF1MDzjsswyJJ3VjLlaN5XRXBs9tUdKdpPzxatNj
tShMS8CNudQg2ahgkvY0Z6wLKLopaKkomE16wCAIYxLBAuWr0por4VVUl2OrERTi
hWjObz77pEhWTzEGLnlZg0tTJivcKfrGzMsX637AVRjTK7mZ5l45V7H9DhSgRpAw
CQM9KJntZFWds892XPrIep0tO+s7HHylzQjC5Fr/85WmJaHS4QYKKcro5tvxn6Ob
VfRjBWIBRankFG3IGirWTdGt/2sxJWbNi4BXCUw4ErJoniT4rwrc2t0D4azvnWLr
Po4ofjwi9SC/DbHPVlIX4D2yW3M4711PfW0lFXrzooaUm7yPRP7T9g9Y2v3pEqW+
mWzELCy/c6MlKv4GF+ez8Uv3j5DTQ3aLsjXTvzIuE2YOJQOJI7UaHP1pUI1ZMOln
wOS3KLwMihzhOALGieSO5w9rOI2SMtsQKWaOrnGoj30qh4gO2k94Af/UVUtGQAyA
Zk1+u5nQpYjz9LUSeCiqIjZ+mKqxsi7UnKHMCr6UFvu1a5YYTZBGe/Bq3kXxfUG7
nASTQQnjQKX/Z+LY0teJs6mjK72o04ksxG2As6i2S9p1aLSH0vZyPeUT4u5FCXPN
2BGEBckiyHbRIPVp7ZPuWNrSZIZNTTN3pXiegZn+SMMPv0L2R1dXDQKuZlRmOHVZ
xVDmWbPrFrMxRlRPpNoTgenbpr0T0TldlBXMe9c8ONEdU5DonnhG9kvqPA5vyc98
RsgS76zv05Hh3f2F2iWA3eBt/DZsyQOqEFAxVxnlZvwEaDm+qoWBHJ4qohGesCqB
LJKWC/55k1DY7Wuxu3PsZ2XklaTya7C/FLBum1Jo8apOE60EjN+ouEC1fiYJ0leB
BXVu74Rh8kksQMShTGSEoTEeYa1aS9XPA1P1mJT7my202tY67JJPEXdrzit8FkJM
9lk1zYDxtylqG1MQD1AAIXX0EWQzajls8u/37pfIyvCer/X02/QZa+sr6rLQdKQq
ozBbL5ODZoJRxZkxnn/kxZH+Cc6gRBHxNvxLrMijAkhuTj+FYnzeonxeAzOGJ8EB
2IKWqIxwkwdPAiPG7h70soKvOjDG3TDBPbQhvSyWhMHf3WqI/d16vuCiLvXqk84r
W/sV5kizAUMH415NZbXpbnWO53VY73G907ANvZGiffVuJVIQxBBXWZ5Nd5Zd6h42
LeSB90MaExz2UfXxiAxVy2TWDOoG0W7WKFtSYoo6QnS0mnyJMpsGyC8YF5Dnl2gw
wuIq3G49c+zSdRamE0Rd+2jKf13iYDeFTXqtZcJSese/xzg8y05W6zdaDr71WO5n
0BYp84P6MJ26Z3mPAeNtp5/qwqPUBNyviDhD+U646IxctzDpyD1Byb8VoGZmp4xK
Q+uUEHT6SuxnvdCzIX4SNVGuJvDNnh6UUVSq7h/XIB0KEpVhERSQ/rO0w80M1WCB
XT9s9qUYcK6Uei+TRMTAcUCeq4aOnZ1KerCBwxlQVIg7k5fc1ts50g/xRFd1lZUI
nREYWv5lKa3AEV5t0iND73fYCOTXAtDOZs+NHtiYLN1lLl0Cb0H8XpxTYts4MUYI
OVfg/nK7XDHixGVMaZ9l5/G1jt+1p5E0gYzG9DpKllqMq3iXff37u04E3lYBfxoS
hPIDYPAV6+D5f9wXF/qfF74rBZTfDs0L102uaetz3R75WgwKzaECYTGJ3McSiHcd
zBBRvQ3kU+F2lEK4lZhNWfwgoGuhfCgMECae2ml8zG4OsidOozl/cNiP6XxCAUv2
qmozEEpKazzqBSdJsrBDcT+lM/GOtrQuoAvLOgupb11tleWJhaXDAVWooPaA0P/g
iM/yOdSGq7IPQvDi4BY26R3pUwpvqEL7tTmaOkkAEsE+/0f5f4RhIZF5BtVWX+vz
HKvVbyK1SCyCx9TbykyCvFU/W0EL7Bwge5Klx8JJC2F1UVS7GTGYwo76NVrsRmAY
WIS/4PQ2IdccMJP4k3c+wMDR8GLhc0tpNz1a86zSZ/WJmRZbyqfKD6sEGqSe7PqV
A/1Ualq+Mb+fdYllCoGJTA4ilbRbTdz1bEt9tdHl9w8vgphY56qcP5lE7Clq7YW9
++UuCRJwdn6pmLnoMNaNXnsgPtcUk4xYuieZx0AjXZPkiqqf2lRIBEg4jbJpGwnV
i2scWnGGB8U7N1HV8g6B7lb+kBDXd8mx3XypBMPV0waJKXCOLJ1QxWKUJNledX7m
XpRJYkuboODn8yQFNyEFWMXbG/EM7DnSPRVCrtEWK+rD+IufDRNM6Vpg/BaXTLII
gliTVttbMzIaLfc3rIlY6k/k/gIQ08kxL2eQzGzJKNw+l57VmGlkXm6bQ5hea2kr
FWGIp9Be5VaMFM22+n2wMhbybJGlMpjyw+VApTcq3mtMaA0LDMo0aLWyTgIXGj0H
amk7mnlTlTXOxXJUbMXWlsEGxRfPkBuPnngxmh4ouzhL61SNhQskl9oS9haTC6pN
KAUguLyxoiFpJMS7buJR/QNVD08/7Rl+6Fr47LkFB4o2BLzzvew3U6t50ND4q+KN
hjT8ijooFLM7pRVJhwhnyLHfWLGWSvFjHNzXRLYNA53chrtq2HKbT7HWpCrYAqMF
7NkKY0pq81EEubAt/pAIAzWhFMYUsyIHIZolNHqHxn45gkh2I00qTY0BOg4hRc+c
KnThBdFiZXAB/NatuxK3uQZxhJmtIkC/K2QXyWS3IbWU4F8PDiI/4qJ51yUnzwjJ
59W2UehYtWR5WsP2lIk6wHcQTSk++OL7pUK817Zdq/MCa8+KK7H+B2/gv42EyJiz
svDexVIsASd90nDc5CDG8sj/diXF6hPZwOFSKoBdhXnaeptQ6G5YKg2sj2hvepTH
dhcXk08hCDsfbYfSLhP7gMxHYhIP0FdwyrAwk4s1qmyq7I95L27DjC0SPEwQQ+Mq
0aneCxCwz5u1OgH2tKmdgCMMonja3+d32GmuQodomBvYVQXIsg42NRqXyOeUvr6v
FWF8NB2X3rNDW+19VWV8HyDa0JAM2vQPULGPxBIqsxZG9g78ND3g+StHNH97h/zk
kRgeCkGoqIqi1KBb4KDpmBI/VKLaZ7pKuO/0B/pIgggPojP2usmq15LbOD0EH0rg
m/Uqikta0FiSxHSpUCKTnIbDEToQiDDaClnyW0rLvQfGrSXuEw37R9nahX4dXRY+
09icn5+vT3FFHUIJb8YBDJJ3jfrlXGPnAdChV+3mbztStIS3v4ZGFq0xBp/gwr9O
ygDzvY9hQR6zvQXpxkc4EI49RcDVoEdU9d17X+mzYsFFdkIEnpPv+NbBeH1+PtzX
kfyGoVPXlazbYvTh9oNDizz1ISAuADFfHc/kbUJGDlPstejd7vnf6XnWLZUAMDHD
ZE+7Cb2a97WB71qriPxD0tpbi7o33AhndIpeluCxIMg7Nm3G09yP2lHn22VIcmek
+EpUMfpTMwvxt2rdVqB2trnw+8gKqQRMJKkNnvlU0KdnW60DXXPwAPsjpPbTdlUs
eWda7Rsbv7Iw9XpcpcX+6ZWK6oAEQ7sjc972At1Q9/UWlEx0t4GXtaRzPIro9Ncs
ngvG4rLQqiFYhTu7K1dt/UZHurU/4qs9avkoIO4odRl3/yJKck4WmYNxw3XwLEuM
4RH0jkIb6ZsKML+DkD540cPsUuSRVxmVfjWgbGZ3pLZg3MNP8a/0kFrIsWUS/SFQ
Pl469HcSXGlfbpwO3jwTz/gn04pMv8otxwXQIF3Iu8UhTfZWMoCgu99cnEzv4wUO
wm2rEaPrnGCfM9doK+BQ5UhFrc/OHOnTYjTBle3mjgpE0vkjbdtQUHMkAUSm6rck
RixTh04fM6KkPfwOGAFzUnA9qbxm4jJV92Dp74VOIsx6B8nPkyjNqsViop1UsGfZ
ZG6iyT5NCeMN2rnOVX1rJHLOYK16sVQJF3xsG8eUwNKeNRL0inlDYOQ/5JBWm+Tk
Cyg4+pfB7ShmPGNPv9dDQPA3rRFdp1nyeks3iEoEULJNy1/m0nqGLEClL9Kke0S/
UI++3nmtFNo6elqhJe7kdyups8gCROE5ApHEBrmCiJh0Pk4HvesdAgyETinNeRYL
Zij0BT2kH1siQRVCUj2B0WnR5XKVKH5yFBTUqbFcOeL3ypDZg7HvBjW5oFLyRLH4
6lz2W0gIZT0DcJMTOIQSR2dIn2w0Pf3HmFPratxCqTxMtqtsO8xkJo0mGoMt9HjA
mPkwoPbW3/b6mTLcmwsD9aEUcg3ZenGpeW6r/Wq/nzWWZ4MrQxsAouF2Ymqmy7sc
4LOjiUjqn1pxddhJnRRtlNEQfVCzQT8lh+R/aiXC3Uy3J6fS/BupK25IBoUIqOyW
hQUF0aXyAh0w9hLbwoo6W92SOYG7RL4LnKJs0QRQ9xRJNSbgNdFalIpivrjn9dRc
la+8ZoOl/vPv4ZQAm77XbetfLLbkKn8pjt0r9yN0cLv6tCnUWK4BKM9I5EMk1S5/
/zCYey1NWYM6QA9iY1CBy9E75Dwike/GAr8AJiGycEMHOXpL7CjNI3T5WS/GnzZz
5BAz9W5+8zItNKARN+Q6p+H60fU2U1yAKBZn/pOyhKG7Y6jK12+TO+HzCVEXdH1s
9W4G7VqIzYiGUx4dZPcQbiDKLUkWLnhaWeMRsu2iLO9SRTQ4n/kKxK1hvIXsewJy
QUTDebMsf89zMrsvPX6KG/YxClAoKeli6ixGJsEr6Qn/xBBLwQe1I5B+Tu19/GLV
dqic7NNIbqRWhFoT58cRowZDlmq4REvOpFfXUfaRZNxN3OqZ/XlwgBu3LadaB54T
14eQc4TyQ3TsUtDR7/35b5z8uADAFW4Br/4yaqYvpp2k0FHtjBa1UiqyQjFj6Wc/
yslct23p+BjYUOHXR54W2//bfdREYnIYMOL1tcM025Ts2Wl5Li3cCo/rVlRJIIPs
MixT0G2rToXH8a598EyQk1MHNjac4JX7rl+BbYrJLY8L6WTnE1sITPw9PmkLbFFD
5KD2fp2DfQsCwKsUKjvkbDnG94JoWB+qFL3SDPkrCLiDV2tSw4EgnY9VXVRP4Ifs
/2ZR/yZNeFls5KIuO5P6RGePEAfQ8u97cLai5yCauwZdDSYqAyVWB9P5GHzf3BBi
LRMVcmx3uUfl5TArAy822s0fSiv6PJ4PTFyOls3xKBVuZ7XUaUL7lyr9B5PrZ/p2
BUMUhTJvFLAFangxSuWH6u7TNWtUk+cpBpzdoTPGqupelvSOTdinWpiMjy598Scg
cK4gZkjrNjYz5bT2YjSK/efabu5Ogrn5D+dQSngHymn+/sbRAyFNAL/sAcVwkluX
enTbX8l8R+f5qXwjHvU1O4czxpouBRfnckTgKNEzOSikkS43t6utj+i9rGFbYKVV
1a0vjguJPD9lLHY2Zv2EdJS4CqOz+HdWoMiEDtOEcYhu396e58tF0ro/S/gWYizt
L6jec8y+wpGA7PeOY0mE0Czj6f20eJ8N3WBWvsylQ8NU/eF+kddujhtBvskHw8rn
2osoJCDX3BKGHYEJmae/spGte9tm6D1CKifp9fzXdgx9NS4JNr4bEoXkI6jusBzX
9bKfn8FKTUFg6JBaW8YtwiYOCPPvpJspW6v2DQhhV42cvUtuXaonxyFLl5ewrxz4
cWb1+tCc8SA4FxqHMFVIfbNgPnGsBdVr13Z5SpvtVV1Zo0pl2QvKm7wbQVIhdR+o
JLH/LRVrbp9YC5f32/ag/VMIoxmhCJs+KZsPjRW7xeGqwnBQEKB5PjHwwNnvifqJ
eLIX3xma+WGvguqNlECHyceMHjcspcXatmH2XxVEskz1+i1mN9kKigG8O6xh0TGs
pIRIKnpcNcXkHf+3sQPZ7wqm1BUz5A9fVgRLq+Khlun0dvFwZWsDp4Gfk8975FmS
ZM1UdrJLLud7c7lnqIAvR60aoddjsFMtJlu9Ecr/5zNum3gFGdsznj6myMi689h3
QptVvo1iw7grHPrHhqpmjlUuc35HFiRAUhUakWgtEwREoTnF72Dn+sLZmTQjO9mZ
Aws5FqnDixHdxTvFQrv25AYQnuXpOSOL6BxLK2ytf79Xpm7JyvQARAKHIOSU0xJJ
iP7UhsVPSo3/NVlXkGic6IVrIvQddB4hE+VF0WBgr1/fD9/ljd89jzR6JDp5lAkD
M4Dqq4RbrjlrrhEJJWMGErd0ANX4oegQfj5dBbiSnhWcAB9VsOZPj04ytH2c3DIG
bZcbAgrQPftP0T4FXfoevsSjhi5LwUq+/0uyJpDj8v1ZZtaZoM7IJmAVR0f6chbi
UQefZCj6uZYe4eZxC5dJa9OJoAkM/b+w4hNcdXr10o8SUzxHPNFKN5GIYUtvAdBx
wN3u7R1vfym0CBkM2bQWzSg0rrH9+KRTMtK6L7Bax07gOXO6Q6zC0foZJ6cN+Q0G
npr0HG2ahanv3MwsdLbbPqkx/HbE3yoMv+g1L0Ckh7qXkk5mTez7K6dnPEt/SW+c
K3210WxRoG9TOsCZzl/1BCWDGyNo2YHNgNuqVTZvaoC42T6dLjCXOLjrl5PLVKIv
6DEzpgufXxrcBYldlRZYWkzGGlbWcBC2rfCRSZxGSU700Vu7lovGxqJZUXxbUwzq
WIewQ3548dW1YYCm49UTzWuvoumN4O3uhTzGcYjBRU7qMq8o2u4y5u5vQ3tOUOje
HlXT0VGgZdUo+DX1IzKrn1d912DVqIyAvNDAb5JnHYxMeqbWl1zqMzsujBC9PBRP
X6XUd+qkSGxHL4XoxpqJoARHwhoOejGa/KqsXtJsdJLUnjWbYvkO4zSo24I4QQfC
nZEYRtv8CI6NBy8J17RToAlNUqT+rE7taSZ4mPEekaZ2sACmFqiHlcTy7thz2fV9
qt7p//4ZNtmlxA9c1YyodFJk9xjd4SbnB3argmWhPY4Yokdlxj25J4EsgaNagQ93
V9Z28k+j0ZgtJIQF8VHe2SR6k9+3wWNaDEBE5vXAR4/xEOM8737Q0I/xtibkB0k5
AqB+br3973kGX4VfSQy2o8uCcO8772lelvXI8K+FsjfA55h9EixaMn3W57ZOea/W
srvyqyMAwZMhPgv+GNw8SfK1FEtNtEalSVF6/Ge7wqK4/VeCg1A672U6mbLgrOzs
EaoHS7W+nuAxcRngI7S+TPaKtkjFoivekiAnfSycuTJxMcmIAafzC3bvnPPOzjdc
uD1l5y9UE+7Ub+RWqAegHYpr2NB8h/RnQbpVI9GQi4706905KlID6jSLPVjKwpi5
nCMhL/jfHT2BvUwvhCRk4kCvF33JqGiqroy601aOsQ+MzP+ckbG9XysjpZJYPL6Y
yXDckCbKI+Hcr8oAIm4nR+Ic+UYrok5jS8caHGGrT3+8CpS6cH1ayRICQVde+fZH
pySckm9UfBlBjX+6U91wHviN4GsYrYna8PS2Y6tyunYFEYG1HiMCmjQtFoNa6dWH
c6gJjEVWNG36VKNrsyeWA2R8eJiKAShn+G55KTATKAveZ0JsJ/bqwc971/WAppqH
7x+t58gIqYLMF6Y3OczAvQ4WdtzB+/sryfBppVl+QGVG7wd+625x/lHCI1dUFV84
TjVxUl+wivcGFRQ/JXtQfH5s+3eXoEWcGvqESN6wM8Xj8zdEk3yv/6Q6lT4JkYwd
HDHMrzbVOsIAk8ltLZ8ujClD3YW42oYfQajPdhzShRIC2/kvX4dRa8NDOUeopahz
6j0BtR2yNxKl1kkpr7bVxWHJGjMWk0Bx2HE+qc/fucH8O+uY0FjGTG39ZcIvd26A
qUgelaGzgEKF0EkJMXPU3nDaJmVs7P81HZFd1BnJw9AeEZmRemJ6BdBMnRgx+ML9
VctlyfD21cq1ETJJ+QilMhf8bh7Ozxnt5+kAXzU+g2ZCUFiwHqNIzQmYq45N7k8U
zJtyLE6qvac1h45HwxMLaNgon4ONrK/WmvwBIOi2R7OrUL/JUjaeIPbNuGudj9J+
J7z/JRHcfVmAe+DTVhqbLRAPZjvGxl1GI9u/sH6m0FXCs3z80ksXDulW4cVQeeqA
yz8e1F9+75Pox9w2l/3h/YEuEexknzmbEexlKZQy32kSKfHrgQ83mcjYVCio6UHC
5ijVJNp9+1kgJ0zBdOE6nKnTJkYaXD82TacWaVjsdeqoTB56s158Ha0oAjCO2jAl
hJoEKyHy6xQnVuHhNFNeCgPcb+w/PIRGzKUJt1LjPvwgbRLtNTwb7oQ7VN2UnyXR
RVvptpCW8ZB8S6A3ikY7+OFuF1idwPoACB/x+x4bThYkUtqFHkJsBV7T1vfnRWbt
N6Uc5BVdjGxPPdYsd0i0Led7UeoGdTps/8zO3ezykIelkk1TJNGaEf9IlQKQy7fU
n/nHaaOAgvrkJymSTPiCPRO5zhaXPGT2LTjTEI5UBLV16RWyrb4k1tldd8SKHAI+
lNn78T1EPjPC1PblGr18jlHwRUZwA7fH77ZklAmJgOG4jGrmDfIRqrkWFZYxV4Be
+QkKfAocUoBzX9wSgd04lRwrBkfGAFKevuZzLySGDtmtKTAWaB7tFOE4y0P2O601
N/mTvi2sWEIMR9dpIYYqpzz6S/dqb3Fm0JBwFZyLZJoUKUXgFQUkwqAsDUByhDFo
TALPKez1AYG/AS0HZ+cmado3So5lIVUiUI217SOuWQFAZpYjFjaTrkXj+bPxRXPu
/EiQnQOiBJLccRuv0UAfins9cWIg3AO0P5CB+dq/ETCNvSmRFyJ7P/BusK0SpSaj
x2fqVxgBiRx3575fCGNWdJvx9TO9I09krTl+oa1r8Vqw7E8mx+sP6djmgtYFvPok
jmn+PL0adLTvT7SxKjFRY046cujAinp6Ra5dhVWADwDhriWilXwUfxK4AFzwvA1b
uRBMLhSKiEqwMOhfgig/9baHKsW9IaDMxMgcFWlEgRE5MVerNr1w/1d7zm0o5R3C
/RZn/ZP0zZSXHx4srruw97oX2le0f6J2HbYyof1lUpk0Ex9Z5AQid6o1siCK8fdB
rRpDgHz1ryKJv4cdopj4XCQ1IsMJTYjAaV6JRL6FfCMXOPnMeoQC7JC1ZLvwPHlv
K5SPhJKDIM/hGiAIn284abx9/ongeE1M/ov3fruUTmGCT/+CP+hGv3kSq1X14fnk
osKoLep/gV1RaT4hQrgDTTGveNuwO/lMkH30uMxfE7lOjTHP3drM6XTM4tZ95Drp
UboG3ieSLkqrDriltjmKyd5DHZbxNu3lqtPWdIg+Dsgg5Pd5MM4Yzj/K89GQFnGk
ueyByl2J5Pmkb+qZ5nqc9hpxKZhAsNWx0EnT3z5ikIGZDME1KsH+EkHW3pQTuQYu
lfi0RObNQmUnVZvTg7sxHazKQrPClmzZlZA0lMULfrQEnXVHb9yfpzos/3sPCXpD
MviCJo4SkbBRRZ2yUuCA5pFyaxOptkK4+dgH4sGcJKJIlEkr0+8uw5C5cXLD9eJB
d9XiSk0+RZCMtbfjH/VLJnpVtqm8TVlWocOTXqKsxfPoP92G/hMhLk4XIa2ZhYG9
7WF3t+JykdI5EU05/VzGop/H4SYES9jAugewHtTic9KJj/JffLVo6iXE9FaocQ75
bsqg+r1Lm27XWneMtCFnG2+cCklF06L6ekE1r/+w/Ogn4ihvNiLEvr+2LFKYWIlj
l+paKTpFvkODVTXlSRm7xMkWfDK2kgA5+23S9YyAHpTbx1VET5dqDdc8VArDlOd6
UwrHWc+4UcSLyYV1jEzX1Ky5UzRMDHR39SiJLC2aV0Wse1VUY8Vqka3QW9qN4KW5
V8vLY9CRGu5WGTTFgFxxjAekRMY2RAglaT2hT7E28S9FXIoxbiO+e2zMuc0csgjb
BoyUp4a8sXlV/5uOxQRNVyyWB0ypRZ88NJs5TSGpQSD69pjskzNsWbOgQpQRF/Ta
R3FjFVrtxOf26b8N3146HZP85rLlpyHkpSfg7RKcWOvsxM/nF2XIW6/ymglndU8k
zG0CN15bDES2el5NsjLnbq5H9goxDzfP5saoqfEwLGIASMZ0yiiF0W+DVUBLAozf
7iupKT9upyvPvZbUAocCiUSkhLHtXqO0MK7qmq66Ne5qLodkxH4Bet/4XOpBBAHs
tdwAt1GxBNCXIntQTOu8md/SWWKeiKX2LqFUwAaWCzlbjo4TBsN7jdmvHb7CaMIA
6+F7xcBCirKr+QJriWKP0r+z6JZmGsWKxxP+IpRA5MUwQ4PFjih/rOCcXl7vnICK
2EwRoKRcGfnZt9TQwc2cd+kMgFfENn7jPho2ZGdJf4PPtABCaedwA4PdiVQXVgDw
q6xB7pd+xF0VOMZO1Duh9vlhcp+aPn6qQTGxT+Xcq2TwsKufbGID1agRglSJqiEU
bhihlu6u/o5bItNG8c1yLu52KGhPEtJlbFDXt8W3FNZ5I6TdAuGihgxajFpkkFBF
jlilcpcxsI8EZIp1UEGcDnpzzpomH+gxZgo1fbNRVkDZYvFSqfxLQrY+TkaMlkdN
blB8u0ltVnDTu8ELkQiSauYXSB/Wsjy5ngLbVQcgrnpoZx/RKkiP5rbdOWWEqHgO
0yMH2zmdm6j/r+Za0nUCjKhqWfD/G5s/HUbFk4OaOqBXUJ+c5Kjo9q6q/87eyw8i
7NuyARuJcqh9+AkU2hU7mzBDFIQtn8WVj7iRmrdyPPyQ9B5x9PtP9Hx/JT+GK11+
owwcA+67DNVDPe6k/tgLt2Ebs6cWheXO+HsscfSDWe90sz+0HEAC71D82ghJpOYO
5sik+h9H8vQGVQrdqhDDzr1uZyicRvjGy7ik3H4dhzeIxYZYDox1IVm1I/+5FY1W
bzE8kcWtLOQHtmZvqEsYnSwc/T16Z8K8stQ8IZkC3i5raqUivuf8PTSk2Sw5GrLb
6FlYTRc6elAnGw7oDbwwJnihEaLzw8u9yUH6vbvETR5VLGAYxs5dKMAQt1RO/NUg
+fjWPimOKiY606E+BUyiIG1Htn8wMS1hMVpP+ZyPT5IiTtdgw4/m+PjWECXAinRQ
eO/def4ZsFFyMCfCk6HL85g9pi3MLdatNtMux+aFkRkf2pvBnHZi45wGKoM9F+FO
EKGHsGY+sDjMINXDQ4KVwg56JxUos9xHfxuqkRI7DjCaZEJLpd5pgie1/K0nuVAC
ZFYtBKSrPO2JVpC5AQ825m4EYRikdmKPVpZCbRxr5WfUcp4hgmnopEi+xbk0mGUy
F9ItzbKSHqd4KpvcvbjyMlAGhScE50BtJxwlED2Z7xusyPr0lCLj+Vh0eMmA7yz1
Zbp9oC2yaQkYoR3i4Mr5Cpx7mVVG5Ko4csIfctUxPtI8EHl5mrS7qi9e8hsLMeeo
jkkQUI62fzAnEeGqxwHoifqZiw9Z95qhsGpQSo7oepqs4NiugSqKTyspK9UMZo75
SfwvL/U3lV/lxUJ0uB9AhIlT/TRUps5I5Z5okxbz4TPRi16QjCnQym6tIg026LNc
oWnlzSwziNZTBEdqm3nlpusXSGxN7gy5IYOZntgiIYGrb+nt8Xl9AZtos2cHd/RT
aeNG7yriuJnEsZK17m416HQadk+Qd77gDrIiLch0UnDTQdhdx34XQFcuiW5oPj0H
aLr6E7rNdFS1aM73yIf4xmgryS8alMVCb/ZIMah8jZckpIqjbirPWQfgryjbCJhZ
GhH77daAVgdJEjoH5V6iykqBWaMfU/MYWF3B+cMhJvlqAmCpV3UYgZRDM2DRK5+a
VoCqmugCT+1rVIvYYKrKzjvlOpX+wmFR9Pc1R+fM3RpUBTX4hIXFjTWrNYMwCPIJ
xP1ULUkW/I+ROe64+3Rt42JGhSs+sukn/mOqvUEkWnkR1JDlDS6YGjA2cMH0s8jT
JDyZiwxzI8g9nuDemql/SspXamDglrJVEH/VnibHNyIhyyQk4/HmUV0IlyBKqACL
5gvIxLOQY87suaUq01lhjbfgEm3VmmYNUPqugqDA9VN2x2inde0modUSWWj9IXRS
p6uiGE5aUqmd4UEfbEI74clceugNOPRLDKkwPbUB+X6PuPJmx9ROmX1qHVcpIqHU
tqm5neHdGbkYgMeXN3wUH6s7O4QYjGM15AqP4AvEWrS/cpNWfliwFCWd+eai9+Wp
oU/wFEmNdO4d9pssPr/0oz/rV5VnFnjYqkNpa5O8hZt6F3ekYmjodP/sIFMBpTkd
6Que6m/qktDdo0Z4C4F89wv4MSSA0nSQKM9Rw/VkJui46JyjIzEyFjqsQwP6s00j
fRwiAR8JvEGytlbhsmIM1AYMJExNqwILEiRZpcazN3DvV/BNh7fnG/FLYJrvS0GP
5CvkiQFdrHI1stI+SbCeuangGP5it/nt0+mhRPQMMpf5CryUrb2pscWgkSrFMXOX
t4eWNLnS1qDxlvV0k1MCadrzZ+TlnP57xj6xug8NK7y8RWrv/o3YBT4trm28GmEn
E5vxGJywuAvqEdhdjJqRDf3OLsOaRpE1BsAEZsZ+xkJjMvXw5F0HO9SPDA4/mr52
p8i5ZukRK6dozC09zfj331yUM7ZVY2zlbsesRZElcF7C8tczXd6IwC9s6IEQx9Kr
csp5WtdBD2TIWvVZsmzV2wF01Dvi3FeR29Z7kuEVWOTxrcDbafdkSoO7e1YeCIbU
OLVrde8cjGP+hTbckDUbxQRuWp8Eb6khcrEm20oVcQovD187+kZEXRLsTGjJ+v6W
Ho3fUbScxWkzFqQo9ZtDzZ2Xs7E2UYb2K23ZglUgg5aDTp9EI5eOT/9/2MpIuFxq
kvBwSoFNuriI9DOM33xzcNiAXhtqKGRTzWFOLuBJtwtVRBhTKKg6bQqzRb+Wln0U
51g557Amnp6fMBRcA7EMNuB3M0KAgmLszZA3JW42LEG1JEY1s7Ji/Ki88A/ZVmeN
aBS+ffjEdv/JZzqcKHjq5TifobQPoXdf188E26P6msVDAbRdxEHO/I6lV0qiouA4
8VYxELDA9VyAtDfLDJnym6xd8AfT6uUOl1jUwCuzICK5/77o5Pb5sPruSX08Dfqo
VQCv2g0eWtfGM5wqskVHM4wgg+disqdXRYkrNcMSMibL9kzEywnbZiFtJ19246AV
+y0m1O7lm+6LEcEJPpx72wPaYJ8dZvhnL5tpraDpmb/TxYhd7PK9+ae7n6usu/xY
2QstbZwwGe8lypPvoOJoXowTfrVQ0I0EKP3GuCNPY0JyBE9Q40PxUNgXBmq4nBJe
+RTkixLFidNA0GMzQtA1KtQ1GQxlxwrFkfYXBlZW/Bcrf/jD1Oq3aslIwY94+akb
0tDtS21+2pgbKzA4rZUGugwGGu1NuJsNPOCOywqGiGLNLgShDEPy81UgXZbgKFAa
xXjZdkjPfi6t+pL/OtK/3Cq5A/kJ6bdHerAkjwsJqIytm3RGsKhzZ4nGlrSCt1dM
vMLBsc4jxqxRSHIaIszMCpRAN9ZssNWFYqjrjvOyuOfPrRAE8nI8GZTBQ9DmZbzG
SdoU/XUl6TPDyFEJ7tcnNZQ8P6MsAwBQvnxTlxlOt6KcX7pkjsTF66FksyKgEahO
bawD0YNi7eOg/Q9T1Za4RsdRZ5gYMWuifUPQ+FSQSMm8Y+NXXK8TZbMB/O8Ec7X1
VjeqBWkUdP89yggMOAaUEbZLu3NSooaqpyF+PX+upBpAX/gT+hHfNzujbn8igdkb
/KECoKf9PvDZkTWGiPBBzPE1+ZCBTyMVhODSl2/G7lv8F+ZW7oD8wNfVNCTTWLru
aSNT3TnDK0esrrJH4aVv1Mqc58P68jbehYQJOO1Fq7d7NNmV7tSPT5GNtgjDvGm1
3gthl9Zk0Bvlzk2aYW4ySdmwiSUyMVBi1h55iT1Dz/LSqahLeIgWKPq5yVAzvdk4
JuixPaswmFHBP7nQxvq1ALEEWXxnENSswjOEpcw+0XTcl7OE0GW6ORm6KMv+sZwN
lCiP84N2uH+Avls6P9wHm3BET42/F/OEaaoBw8R//Oo=
`pragma protect end_protected
