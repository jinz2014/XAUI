// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
I3zpowSyiHD+ikvR95AnOVPIitpVt1pKmu3v3Mv/p0m5ycubbHIfxztppDNuxwR4
V/2fbZ0pBV7doqIgbQm96g+H6E9Vs2vL5j5d/i04j9hLuCnRfx0ReTJPaVSyRWFV
OqfkdZcV8RuRTBUMmG/AuLpopKMmHhXTPOORkFE4bkg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
oiO14rC0xWYm4+6GBpdK5I1JXZa/iBxrKyarIe3aizg297a8Qj/X7F5NlSM+7UKg
01GEa+wyOIkC1hX81sZPa0FYB2ezWp1X+v+DpNWaXIiCiETblp+vDvSWe66xecRN
Knjg4ElO6vNb+H9edRL/M0WWTsTir1TIitdVSmv2VgnBdac0UubM0tWdskvoG9Xc
wN+m/ZrUKTbbwKNkNSuZtlbr7gukLzjnlYt87gL1B0/HsmPBy+nF5EaVm98MyQxc
7DIRdznNVGLb0RUD/73jrySxCLtLY82Dwp1dq5fNmu/ZZGoEvVaDRXWeNNEwJYre
pv6WO31ftQPJpWAKqup9h6TWhvW43rWJdFZ/Uhdz12NoyPe0uqqOEuSvlxRdNcx5
OIpsqmo03vVOdsWsS8zBKJTrSnFUXcfI5Pvg2G/2eoyxc5n0Aob97thTJ5VmrdYM
nE8kzqA8sjQHbMb97s7pS74omD6t9MjCRRkCl0IuyjXrmQAqqHmJdaZ/0530LfDf
9F6jl2LkwEsnDr8fEbMIa5a4WAMhhRMQ3FHRCkIRbwoNb8uU9wgIZIr8j70V4UG+
aQgRUOCOUZ6itVaC6nOqCJZJ05FqOwa1HehTEKj/LEDvbmwJqj/UHmSARKXiviwC
xqCp7BGr/wi+MMn8jLqFBb6qAXqlPIQQobAqXaMo3voQlpeIjWK46g8crIFTTKak
JrTT6gCKPzUC+QUqI5bbjmd7ZkB6NivL35D0eMjffMXF7XvWCKAXwwv42CLogPfp
Dx/urbsL9m7Lqj3UbtV7zgMkCsQtW2qVvzXXPuFTkfVq3fmF7dZp7ayhBuVsL+Mg
O9B3GI8Dm6AT+HtnSdb3mgpVes1R2rLXx1BXVnfAxru+jBruNvWEgdjBAqvwSt4v
SqxaDaUY/5a97wQsExfoAcy7b9OD8qXl/FNiK4XxcBZLwC6oBgkeoeCQZfDDrfwC
U9w+SRZPvycr7byhUsahgLEsWto7Cxs4dV0+z82ski4rqzjOSOOrl66u7YG4rTf3
TWWaymlrOi4BzisSw/o3ADy8WyfI8rnAlVYdIt8SkTu5UzUdM0cq82pZw41vaNuN
4hepz2nt2VYyMMb7SmiNsUeB0Yw2Z1zhNqgdvd9ntX2T3xCIqV2W3wpybXi1OYQC
3eJdoPHDTLmyIZifnB8uUKB1EmoFuqKS0cV+We5yBwaUTQ/0vrRBmlaf4RaUSNcy
lLvTPTmw9pRRNQzfgjFq/TyMQKu0K5OhdSY3hIgiHnDXt6/+GLN6KXiTCbpvQnos
gNUGrTfvhdauDG9eKPPN8zliVCSCMG3+e3F6nNuWvBwXHRLh2BcbmmU5bjWqTmBA
p0rPgDlRA0FLUDXyDzlPU4G9Ka2sRtvuG/n+QkWF3wtnY4sRvL6J/oDO/gm3uxwC
st1FsWTpNNhP8G9cSqO+MyEUvZsEDrUXiC7nT9g+hZrYewhKuzKirCzDe48m+we8
OO6c3Ga2ocqZwXptIP1SYNAzSa2tGlgOovEGbENoCMGHeOkwnFWW6gQcRdCnLl6r
rdI1O9MnL3ceTFA+uqeEDASp8JVicJUOKT5W/BGqSLIZh2EILJIWw3UKZuMqPtrO
Hj7r+w+iuDnKK6ccQhOllyvGa6roFXTKaX/mtUKrz4JyOKjifVFyUpVnjr6LR6eB
kKg6tUTxIA31uMYkJrfjTwOO1xWR2uTEbBP4xqJl1kkdwyY7Tuq8rhDb0R+7MCde
SQZ1iRM6YNNW+hX9+fi7L8Fon52sNPkax87aK+I1g4QEQIo2G3nDRhn/3/rhq4kh
7RL/SQr5VkOVXGTmkSofrZHIkYU0SBnZpTGrT4GXEbyJFCx0cVA1x7CuKah1jPmR
2dmzQx1BjBLxTeDBbiFr0seyx6TErujo/u+tDaawClvedjv01VuRq5FvZQcXXI7p
zA0rN73Oj+2XYcaG5TmEdw7eBiE1UL/wUzXygMjoOCCHTkbl3QxVC7rIote6rBT8
EO32M4Z2nN/sfy0DTNQUAQ4oVO88E9I2W5egCcQ0rlOw0V2hTaq+krBGCyzvj25+
CQCzh8Syz/5+lJr++qXilsT6OPjjmm7JszMqtMLCVhZ7acPvJS2L8WRXP5wAHV7y
0IJPIaq/uC3B/fBjjWEZB6mQ/wzD0eYLzOFytZ98DbbEwfdpUkXIlPG5mHtduAgY
C20Bf9ABZv21gIpgt4p2i7pS4ny7rq5zKLZkUQGRFmZP9NktTjzqhgdhokZFNZ1Q
SlU8EFjp29wOTOb05W4nzH6SVpUnakpeqZcNrTNrkHNifviXRyydt8ibZG162eP3
lzyAH5LfiRf9fiNEeGBV9nWbRoP5NKmSfgPagrMsGlPKsbef7Cc4zP1aoobn27k6
Wn/RfOxOvUZVAReFpcWRIjfA4dQQILHwXCMp3lKAjGw/Oon7eElR8qsej0RIFGEI
CJFZOyqhYHLa6iRKzvudn9LJnO+M3pk24VwupEWoknFSOZDcjyBbqvd3m05byEfA
U4WYpoWXjEaBEYXbrQujmMf7KikrIaxHb76uvjj0YUxUOx3OjEtpGNYrIVCVOAEV
jgPBjBf7c8mv6wWYXdxE7JvTEm3xVAo6D6/mPyEu0jboxRghkz9o+QgmhRnIMxTF
0K4YVwNrg1qp0UA4cGKL+3eTF8xhTGklX1bDvEnX2VZ/lRasklwZbaz6tTTdUDd/
EwRkrWSuUnQdDlqP0W7NdfgUKwW1/OGpAWfM8NLPP7ggqDcEsQRy649Q52Tc8Y2F
UlwZ23j4rAdQgJzIrT9m7oEqZvlMtPDqbnwxA8Vg0P626BZYDcI4SD6GreCeOJD4
Z3p1MSBLST14mznE6jtM1p4GUxnUvBXcUUDCMXn9owxJBchdl9p2uCVI6W//jZ7U
2WHTXrhsBFH9jOWYNVSE6CtwtKP+Qvfj2eaoAkmXcY2NalHOWGbT1JA/k1pMpP3t
YLBWMKnl8gA6MFxJblACwJlvNjMrbsNLo53BjYnLJ05udkNH7uIeMR+M0Y9NTzEH
mGR9l5JdJQVVtbEud4ujDWeTY6vV8VcsfBlPVH/FLfWDGlochBZWuuAwtmyfJ4F9
kYiN7E8fHZOoXieLjXKMrOE3UaI6cWoY4DMM4p8DKeRqAdfgi+LAUWlANtnvehYE
Bqi8kS7l/U4SYjkG/i2q/7CTJ4r5YBsGlSbLNwAJE7cSmWO7CJmZL/6W/WCZosON
Amj5iYe2Iay3QG8K/Y10dAeEbZF2PrWHDjOzWgZAPM+Hl4tSVNn40JDClnKeVqOr
+aIhhYHKceUejcwIKjzR7lDoBKhNKmMwJ8VL54fIjZ0Mnk5I+2l2HchOKgprOprR
h6fcYCjkwBqUUHajKLgSpQAiZDBPeZXzuwnFu2yST79JDKvroKwUnTdTvm+0Xk5m
SyzbXHAIoG+w0u9XQT/hwDHLrESROTE7aksBHuu8l5bu78mQ0esqyONb6gi+ZRzW
T/WbgRPSAhPUraICpRhk9/imjne2Ss9uOXQvozCjgwvJ4imh3+rCr7CiM8zYBpdw
cgCtIP1Y+iJHkAxxmUe/EdH/YDWQOYkOeOI9v6YhCmf2osOPNPc3r8Gs7qc0jgBz
LXLi+XNaPlwubI+mlVqqEtNnwiE/fsJ6DYwKRVKl2LSk+vQlZr9un16IfxzZXAaR
uUTFkA9oVzaOHuf46ZBGb3LQdM3G8HHlezt6rA9yrEYfOqi3u/jASVyLbtVIkKHn
KZMXQ1Du2FN0ssqgzGB38iiDVdwk8ThO3caPpKlYk1K45Mujg4qC62c9l7t64TvU
qFtJNXofeLXtR8tUOyzeEJe3WJ6ppjHsCucQ1kX42wQRAVRr6zGvkSt4XIsDdIdb
mt9ZEgcNLBFOioi8cosOKhPJz/Jue+dbkyhpf6JqqO0OApJCv//b7wrP/XIWA36l
K/YVCPYJlReoI+qKXvGS4fwUd046O4b415PoFjJ2YYgL7y7vGTzWmZpZsfYpYUkV
qPEjQ6rhx8oXMgW+kwNCz6+Y+drx+O1z1724/1R3FOYwacet8NYK0M8k98RpHISS
aEAZQDVqncDADx58/LRRE6F7OENfIs/WbI+nBlwP6SaHwUUHgR+lT/I1dpi7W+2k
vKnUYpr63y0XAXceOq3WJ9LBrspTHNFG0kynhQVt0OZ50aIoLs9lYaeVbDHZChc0
arSLNMCl/+IumSAVs9VtpXaGF5QYYw7aIk9CSJgyTwBRl5yl5p9QBrjkVIcVOh++
72bSLqZ/m4oJH0jb5E6Z/Vkp7k60eEKQZTgrj8R3QBmNb5p/T5z98YlxR52Tf3Hv
wf7Ehi1s9yS4voZmUCeMyuQzvhPjvVfg4rUyg93wv6nlC1h+hWx9HE7l9OM5N7iT
2U7i/i7pZFw/mFoEfd3x1XgkscO8qQVYfTqoi29RRMD6Ry0vQDi0N6doxmdUXYno
OUWme1bRokNSRdgQ+cYwcDEZXafF717ocEbySU827tUBwiV+Y3CaF84D5CjGXoGL
LI+ihpgPAMxCs9QJ9cUWitE+yBu6bjuD2JJqDtG9K8iUBRfxJi4rDfpSZqUu+Jd2
tOS8AbFz+w0xwhH57hamLDNCNengLMZ/yfrnfVRCF+2qFijuzxb1AsVOxxmDPjB/
/g1aVehffQgY8E+aljULMxeHJjN02R1CtefLkQELlboU+k/hpK7qbatG43FNi+Yi
kuI3AD+roZUL3HwGok9DD0asZ+yVC314Zlml80EQwvaj0xnXhxYDRrL7flXVfqxq
lqAeTYaPlwi2YDlLlyKuGMURBq2DXhzY7FEK/uEkTHr6YrQRYz2b+Y2/CqtQ0MFW
0Imq43MD8wzAqYLIGtxptPWV+MnJ7UlX8JAMkfDCSjOb7YjfY8h6yOuC5FIn+30I
ocZ41B2KXdkX1EfLM9vEADDXaUWslzqwmrjQwuo047EuSE9sAE/u6h/YQ0ij+lH/
biRcdnIkJftSD1ZqQajyFJNNMDtcowvsVa9cH1H/QGBBTo9Y9B50DugIkls4cUXS
HrW/1OqxWhQWEEEp57WIL751AAyDvIDQdDRRQVElgNhIqEEPfYLcyrFoREpSFfIT
SZKxZGZcpjfF2hJyFz4g3tFQV096DaW0aD3cl9LvN0S+kTJmgrUAZ3u8PL5XHTSQ
GEEPuTUGsYYM6MpGDPCFzM95Kfxop5wqH4p6jBGt/tbT8Ak3hX3uQQJqJepP0vjx
6VX60jNtSqWplLCyIxPhkBNv07zUUEQew/iSXsVxD0n+fkZossW1VbKzkGFuIX5l
U0PFUYgIXDAp+KgprCQ2+TF/EcGYKPsLS1wTtS4yK9StKjTbL1K9WLhL1MhpgAxm
6umTlnhMfWSshjHgP8mxoZng7vtZ0t+IRal424MYxsu/lxNN7QPEG/FOCa2rxnVc
z05RFrKzcmSzwxSF/U7OeuJU6knAP2Q/GGwDQT5JXgnA6ocd1c2WbsbukR02XXNX
sbXk1Sj07x7q8HkEULHTpekEqP4oUj3vl4FSErY/QbvZEc5lu/jYq5kdR/RcQnPF
sGHBQH1n4mpbqmxgO+LE95A+tpoPD5OtNVmuJw6ugAtW7ufkhIAqTQ7d6vh76OUk
JVUmk4tzflP9CO7HSz2gRsG75y+ug2WHvZYkMGr0ywPnQRHzyFCnrlofknqkZAYt
rAJAuFyiBFUxs3Pj44HD4SZJvhAmB/C1ORVrO6jH7arWaAED1yW+5DyyHtQS2L7g
oTfPN48OIcHby4Yqy9e6+g1MYpYjxtREpKrZK39JL9b1tXk0+iptLcM9mnt3t7kR
aFj2tUfUWdPDlCcFeXACAkWLM/L1CJTrJ0aaGno4oXWnAyktY9Ydi8/7cfsXETn1
7tPgmSHex8Om2YZqt6WP3MT4xxld2Is8dVIjq5VGp7+RFk9yXzgIQfq1NI9CCj7d
I8GqK9caIFjwmAPK/AY64Dtndz4fLfC6j99AV6N0U4lgPn5UjJ3m3GMX+Rv2KaFE
0a/sW4oaCIItObNExA6uTAfDxBdbmr2rJSBXgaYbTOaJwHRgEJQeed7BnBCHI4vi
Y8kOZ1/5rLqFLXcpXhgTIsnSpRjzozmfyr6h+sbvmYlqVTLvUxh3CG/sftdJPtSU
ZaDEtfGeu/y72NIk4LcX5luN+1EHuIHW/rFviR4jBqyrZsD6VEzp/du+sPdeibUl
0bQdF73/pR6/+bdSefZ79vCvs9JuAxToHfUfBTfO2GZcy9oPu/ZT10SSXKv7sDSs
azEGKXNktdBd0irisOQfhsO0oB+8yFry1DgOa+OURKSVYBV72Pv6WzsrTwf7fuT3
ZHkwi3TiKNRyR6GJPLXFtuBdQg9ilyOSKMDGuZBLIlEo6rAMY9RASF5809ZvIcum
Lwp+AUeedpBMqlFr93h0Syqwy/lGUBn6RKzWNNS4L6tUCBleHuLxIrbBeYF8CL0B
NEIBxHt+lWWSvu3FCd0A0EbXuchOzPHUq2wfTeXpWj+GLm2piv/Bp5tRE4DSON/H
1bBsL5/2fuXbScqyv60tKT2gL3RxlB4ZSzLkfAAgxA1sse5UWuJVFo//ek+pRRZZ
VpcJbYyhYVq8sSzDJ1Iup7sjuuwEwiHTQi79AJmnv1dl77PrU1UIc8CBd9HZo3Ne
inPhuBxnLke5GMWco9xqOXmIjDEvwJX2Rwg3XnaHVoblDFL4fWCDaL72XzApsLkN
OBDFowldwihErmPTNQWNs0/HH7zOE3pU9LUzPsaoFD4JPrn5N+D/rkCBjwfgqODn
61dm+cttbWUTsheF3vdWJoAiBhwXGf5JXxVbQn+53ob1/C2X5g1Y5536pn735vjp
rnlAgsP83XO5+L4RcxVqQwomjNRl1INTuvqQYymG7dt3dJ7tVkmBVh7hd0Mto23p
50B6KvCCA6NjS7hPVPCcgPYs/Q0+M6uZmHMbmhLftWviPkj598B4whYKJ0+BdL1t
Jj9tIGYuw2vS3GnOiOveF1tmP/dJiAzmEjfpBDb+TG8vSd1YGZ9E0IEVl8hK6j7e
3buO8FW9DWpeK7UpGPR5Ro8QrLM/i7YkLjlAPfYro1IT/BBShUhRfxiax9PaV5LX
OdpjHAxYOOX3Og/y7o6nVCtDi9qFeOojnz9mlsdaIpcu5AhghY7iKTXH7fjGNpmf
+/bBj9tyEIcnsrszKmGxdIKVFa/Z1XY9AA9C6sigj+x52IrHnycQ6ceKihmSoW++
0+yPZlixW1paSZSRCyfkCYOgePo2HXj0I3ZocH9R7c+SYiYI9ljk5y/NtgWko7mC
Fbz0c+aim9GNktFmiiWBPqnHwkYR/wakRjXSRMoQLwePoIN5dp+skDRiH7FzfoLT
XzWk4ciubxGsc3ydgEkB8vMAjKCk/4hETn/ZAj4J1kbuec/2VID9CFq7FSNYwD9D
BB1e4tk78PzERfWhLkC2R8zpFz7PFFf2Kawa11NiVI8hITb5XyGHvdGG3PEDKjeh
tVgS2MDfHrGp0fOxI6CSLpPEwRwwppYqY5oE3ijgyoUtGp8UfbD4+T+gsjSpDq+G
mCbnb+WeFPIWAZNoPgLksjUXcm/IIPzNysk0OHKPre824Imswz31kt4hcutIVZA7
mZKSKwYS5lOMk4gKHKAEnp6i62DbXkG2dcbLbrOIGdijF1XbZeNnNiO03Mr+3Hdb
yMmycUhNp+i11g8sL0apB+l6sG4pdcyS9EqVO9swsvbVSaGQlbqPaYLdE/SW2Kya
0SamKB2XJqR50s3N47IiHfrHI+RFbvghkJ7cmoeV3X7HxuR9g/WMjxm/geoNiQ6r
gJhcl9JNvi1X0VH7Msucli/xffXjo3Babiuu0+BtR+whHZNn7AH04Ovp7B18gYYq
+sdKu2h8r5SlRq0siJsoHDKJOy3i0FkYAo533g/H0DfS57TFyWEuLhzSjPwdzRRG
fBq/uUEYPUYDA87FHkxqP0exDiNFNnzoss5gPhwixHwSyQSjBfZBmWOudeyBBC6B
UklA+49YPzAYJijGOBocO9U38VWWKOXu8dYhH9fQJdiS1daAMMYc38QM8EEM3m7/
DS/DRJkxMmXsU4Ozd1DTwKT5R26r/wtuWKXad16sWr47CEkmVQVTSrYU0b+6hIbv
DWjF2BOSr1mwgln8wvdZ9RdDOVR5Qqtxi9fJS1lvl2pTnO1AlxWCGpo5GDS7gB71
fNlOBEJp5u7mu87TYIugJPK+SpN1Ep66ilNcGaY6GXyib912RwRkxoH4v+Nnq0wx
bOdE/TB5UYQQClFGfrlzuqflSsnNl8/63tkjq9r4bQj8EC2RImqJ/wg/d/1okh4u
lBm3FESPAPvtziWYbMMy03a9JUkFERtkUEXNnP7MkXolBZ1IOGYVG04F4txL7xgZ
ryeSeN50tTnTd2d0vJKurSZGnWEEjY/H6GCYkdTfSQwIf4D+Esu+5XSbHEHLYjea
5SA99zKDtXv/zkt6DNfXGrCN8T5xSzzc5WzLX/taJFc5zvcSe5JjysgsgfKSKZdq
/bvJCHMQeU6hR2y8oAU28W99vEt13QKa3gdYoncJ9oLZ/AA3ooLb5LZMGwmCdYQq
rtC43ZCJjCx85mBsxtnvrrbdlEtkycaMhTt265/RT9UdovR2nlwQZ3BKYthMYhuA
H/gLDqpKEltLh4DtZj6DwpfDaRhr6CzaAFwiwcBMIb//vuaFy59rYXOIYmbB0Rih
08msaPUfTb9Gey52e24d8vPLJHth+prpCOfJG3r0yG0I69xzv/SBqBJQW9UisEId
L/2cDwg5MPYixE0Cd2ExZY9KTbSIyHDgGN7+bWMbhlBTh33xO1G1EhKZEtiC3hMs
tEq2mDkDDnpbXQeDTSjlgRCTzvy/jTIQjIrsSITgQNmsRxaT753eZxit8inBrGNt
j2PBHNOok3V4RASYp9b5dU8S0i03RP0pQRu+em4L4jvVzS8WtpiqiZj/Wz9ep6q4
/5bC68KbY+uLQ21eXgzZSbkO3YcRG+nttvV7s8CCfCBQzrZVPq1kVWI7fwBqPOjH
b+tnbOC7n6uleyjs41uC1T2TEhpFp5btIPsyQlo2MTqnR8TRiXiZtJ9N5SIb9eQO
irFXnsHfyRLWYl3HorLT/IqlEcn5F+NMxCGoCV/zjy/o/pNJEssdDeph8r4BlJn+
8ocIVjWCHFc9kT8i34QD1ELwvdbbv3DabhdzS+vH0gXPBrmWQvBwy6eCb9CjHYsP
CAq0spbm4Ip/ziVU0XSo6JIsIom9jYkmbG2N8B2V42+6/JmOwWu2Z7wPcdRTWUcw
0CawbXzpLgP8tG1vQK2q6U0DMqsWLo01EgmueWyIXTK8mYuAP2oOO/Wy0W1HEk1S
U5UesbB+IxYAmayix3HQVRfPwzBsrmqybsrmXVy/oRa4mDxPHAXWsWGhvKppT4ul
ZA6DQg6/hxfdvvw5AJk/tPSDCO5ykOKpttX0A1rLEMxI297M1wT81nB0w/0P5d0c
HtEIRFfVNsrUSqQ5Q4eaOAlubxVtCpy2Fmf6v3Bi3upwYQZLrQy23IqaJmEHu/bQ
cWwPdM3POhAbcQkm5BIwSEEuC/v86K4GpUdp5eZphfJ/4k0kzuEW+ZOudmi+79r3
s/qr8Lj+ZZ+zhEDHGKTEdxHL1ZBMRzqAXDTTRaJgpSpnko1AVpr+pFs24xxJ6ImD
uh9Z7vYCknEqo1OiW+QFf/eDj9NuOlfzut2LYnfXQXF2481QFPyek5eXDBq+HQqy
pXrqBvHO7B5f8CejU35tIvZm4KsSIFtRgRzN01UsbsKuyVlDF9zFKz8KS3c8t8yY
Mq5FXz8moeCCkiSqyhxGnujuSDsYL3nT+8TMrTChPn1I4x1IrwEbgTvZl34CdU+a
tzafkuK3gaYP86cJ08pybwqxe4x3ca2ogw8e+j7wBa5c0NC9lfgg7VTguS31/p83
GlsQtVcQ2s1QYWFbjgTsZgnwsdBhzTSvxaZvYH7WRTBS1nwIUAHh8iHEIZ11HjL/
KwwJnVjMMYaZIfTJrLdUe9mbcLLHTSJMvZ3rpxMBMCldWnqANGjXC8qWNDGVIQyG
2PMMu98P+rxWdZEqFah0ANkjnBI5YvFmnQpT7bOCLDyDND8LwTc9mOtoFmJr+QAZ
HviThMRHngDsqIegNYpa/IP6yMK59AqYdB72aUMsnNeuxygbdQYFxpgjbg3t3et6
BSEVfDdVoCMfdd8/5IhdmXCttdSVcxBLzgBxZEDCGox1sJm83EyJbgiamSBjyYSH
jRZrOxngxDZWnjqaswvBnjSMs4GZosJ3Ph/0m8PLKtEGGFBMA6fOLUchl6kVycjm
xNuyeMyH6SQ6XfNjW61V7njkNvUWi+93MkNIUBiV5/VOVuQbYNpmJ/eySAUfcmVw
NGzlQ/5uoxRztFUu98RYz1xkuW0Ex1YS0hNDb4ogYRS6Gvi+YwHz6l1FCqz86NBd
LbD+0Z0aUk8Ox3sds1gnHvJOt6xe7j8OL49Tx3uSwLNyX2bzUI+1SeqQDDQT4atH
dCxmfCphTL/WdGlwXPiWOXtrN/lc63S/gPkhhbsic6ja0t75VG7LpFp4oiFYOL7H
D42S5wpPcyXa6iRgiJ2Wn55SBKHQWPubgJifFdBCsFICSH/6ofq+e+mAjiLBQyHU
Vvb+p9od88DP3ngPVyrGXZ2+UwT87z9w0D6WlE28DxZzFggaoljcgXMqPoIdkaIp
e8o56QYIoV9VjkK9PRmqjGXc9lTIT93oOPNgyysYXR3oSzQKHWh/Ou7T5awfsHjn
AyXJ1bx/YNqT9YzjB+lC0ySp1V0ZArjO5T9p/21NQ0vEb74dlCdGVBvTziM0C5Kn
oSSBmo+7CT2Kx+kqA1gYAP7vhaCgCzrWIrLHUdns5wz1rUKgsx/74bw2awVIiFkq
7/ASqrSnPqRbX3IFiS40Q1YX16NFYBWwM4p+x9TQ968CyXeQqAQA5Wo+0hv86zM8
MiP5bZCcZa3W0x9nr9SR0mKZJwTylgZpxMQegT2tOl3hOBu3oNexbGz3tLofwlAJ
ejZSlMh/sCauMUcjdaJyBETUBwhS/wodMP6VqpvZxMJHIvL9HZvxqsNRKyTc0vNY
HANLVTKSoDz2be6uvqV4Tw==
`pragma protect end_protected
