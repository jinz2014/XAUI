// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cAd6KoBN7V7a2i5LnYAMHY9OV29W7HnhQfWGsGHiXdLDDgjW62KIfwOZ+Ti8VkgN
ShmP5AB+rPjJeCrT9qvfgjZvdNFIxXbzBoRU0hH8FWeoulUZA6tXgRuC76lWbl5k
EgRsLRMeTUHp1G3cWg6LVGRPU9wlpA/lRk6kFxUc3og=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28320)
Ce31SeUGwLI2O2aZA8AoWsWw/jnQv7fgvoQVgcu+t3o14I5Lo1WvIv2NjTrsvjcE
s6P/q6blppOekj6aT2l/Np6KC3cdz+GuNj3r41Rv1ee0j1bDHvnG7Yb9dOoO9ulB
n11vVZDbB0iDhCVUhCUJRZQiJatJE+fa3kV2pX7zHlmNrvxabS1Lcru3FlmSWt1t
g2IO0B8i0u00n/9iikS03x58q0OA8XWtjWM1S7f5b+iqeesuHh2YJluRBxA03yFG
ySz98iTgmwoKDqJYFWiwVQmLJTzjGWybcY4+/qymjzjUgrYBQ5OXGBlH6JI/lzt2
w///Qv2bMOTo6Xx7QgSUcN12YFVpR4ZyocJEAsEnsz9p0QWg6FMLMhyBoL75g7l2
D5tGBM+wXzrmVn9JhVBsM4ogHRD2t6HCJRQxMl42I2YzFq1avwbbsse8JZMoiD4O
9ks8Ou+RmY0e7t6Ev2tExGGkuOa8UfXvVMivL2WgaEjMwdg97pm0QQuPaS8PRLG+
/o7z5ZAkO/q84y570YLQsqOGKy5N8Wr0vZQP/14ZTFrHySow6OUkNQ3HHqNwB8lZ
gFs7Ap/qQLIr94Abb1X2K95Qh07vOQ80NcrRg4nywGT2ZEjp6Pdli0gIK4+T+IN2
EbSjfAMxPTFQGqtO50Js2fnDkcDVgFV56R8wBxqebe4+zB76WlNrbZF9oJup+pCm
JzJMXYq+FsfbA6wcRqynWSgvP3f9sNVqjnri8JsCHm9E7R/bDByKDSJWDaLAS8Qs
qcfJ9vHuHvHQyWl4tYibkz3ekesrWDpr4ev+qFAnyrteF5wnLX/dtlNGjRdoKjeu
1LWkK76CIqU+yvksVtz3gsGJ7DTsGSX28xtpZiTj2dRptc39ler5LY2CGgXF59AW
8mx5E+c86qgjqbV2oG0lu3Qi4EPPCepRbgnl8KodYxrGEUoqvgDjfLAyWOuFlnac
r1SvHRfSDMgJAihX73KxBEwZacJD+tw+oztOgbZhz76rZyk9jBm6ZblGBK55qC7r
Y1CAQmtAvzaIdBTFT71YKRU7ctiRGyDnW2iUyW1M8XOHyKz/Rxhw+LbV0+IDJkyQ
QHKbBLtwiGaFIesk4fM9wlCrSAE/S8QmMPqlGPdfisyCv5rOXwht1OYF5vMieA0Y
nPgg1UF4Iz6K1B1kHqNxuU/I2XTma/UkLYOCvcnV6nIq+g7cXshLOh2/82T1z1PJ
ZzlhbKTIDXLkpHzNdWorDoBxo2H0HR4SHpH4ewnFEY2adcm50xV5boUoTVme6eMA
MSW3QFtHV7HnSsP15/c4209xGjdd4exZ4TXzf4NmbMM3ATwbJ/TSHtiKgTt3E7Ll
hMstHrY5uoW7JcjnFn6XzyYLuQs59dN2r9pV/u6kzPHsXpS4GSJ9koabGMzIp4BZ
KX1jA1dhQRywMSdrFVgq8rN7rKJMxX8aqdwjeDQYArwv2LqCX+8P9KxTjSCeb4ff
mzKX/pd92qmr+fppiFdI3iZyiZoHYiQbl86Y4yh4DkVCeRo9LetBKXdHTVgRYMhx
n5YC4ZU6upzlWO3qmbAgMU8/2TSIOsF/w7WAO5R5MLS3bs0Xj4NfgXoyNXkxkyAK
KQpXfK3XZGGrgxIX7FAX/N254Mkp4fQjMYqtK/Wj3pwG6Ceu7j1K9uct8icbom1R
OInsJxeH7y8+uG9s9JIhiRP81b5BcdKeRP+kT4vvOK10PLwgNmWda9pYwvDrJna5
all3Qfe3zW1wB8CpUmLtZrb3/XagJooMDsKYaRlTDBDihLLlZ4VrfpRujveWeeRx
MzPNKqNBnUXcL9ISGdTnhLOYtgp/OroeyJKaHv6+X/LeDYPXRvpVwogUppfumWwm
OfIIvkAGyh6ESLGSnpF7HVXdyhco9eoe97oebQHMhGmmnhU5A8zgp/I7FEPolKbq
62RxB2Xz5JNWJpC61bPTtfKI08dRx21tUlTHerwI2wLOAlXHYrD3pmRGJq9A4W5D
f4PsVwefvQX1rbTi4Rk7rGMU0spio0joofjVZPS5hYIPIiOZDUol5ANL9xv1xoXn
ThJxzU8GKyQvnrj7TGf6J7ZGiKxRrh6irgSSnOexxFMW1XMDOavjACyCOSGbeHKB
WVRDSb1B7C+9qOeG/eSnvEQnTi1dXo0JikmYS3KfQGAvwvUjd+RPZv5ZQB2TN/bh
qtlpGmc0ySpyH85MQPqB4Bv3khmPV+ivmYS9B5Z3sfRCQvEChx9C1moFn3Do3iyX
3VxlCA2B6+OrZJvlb5cdsKCf2wO3lhf5V0RCAKCB5jN/1Yea2eRavqEYx0xkvKtW
O3NAPeKUJ0AO1lSDYnAWfiHZGjyvzqT6ltThBQX44IT9WOdWFz+sONUeJnh6rZUF
1P3SYWWfEEVDl5D4QVwhoLmEE/LL0voEyxBhmv2LfXacfuRbNdb7FrQpLCfiKJot
u4j7HIciQEt8zNn9y48uZtsy7ZBIhTJfQSIhUaqtBlIX7MgN1SFtY/Hyo1Y1+XSq
qI+hnWOpu/55elX3PnmOqhhAtb/BPk36vDggfDuxtHYiVu2TqLw1KoQ2G1ksrlFQ
VrYTQ6ZXQYh37nFKqxiuUPnE6RE9Wubb0P5ex0qKvvhIzVO0lx2mbWW4VuHn15Wx
ne+FzT+khx1OK9T+5CNYSajD3srZt61KVyafFMLmO22soBFJ4DIx+C3HLKGPqc0i
yaN5bXzEtC3jfzfK+qGtMJa6V6oDIXCHQTN1EJ/iMGlKEBy4LIzkZmNEZrlzmk/r
htE/ZBwCl0vMuNgTuooOgK4Fp3WM1xeXP1q/8YY/55QujP+6sLJDJhGheFJi8Izp
+Cy6dQylh4f611+DwR9nmxDoFZ3sG2nRQxsEHrlyXaNmTkBY7iqGEFFCOAQBse3e
xvcSHyyGve9+smBasPWa2cV/Bs+bgygFYMHG7COc0t6u5ga+YDdCbXt7A2prdhbh
2em9lARyTUXg7+HzMnOfc4aQnEiS0hTgRa1QrVG+A9DSUknG3uPnKKiwqSu3Mld0
waHSURygeXrqYV9h0tbMzdB8RkKI5U/1oZk0/uIrCvUMu34ee1D7kgUpEEPoSslr
pdRI4zNEPm38HWunAB9nJmDu2aeyZOBRA4O/o/YxYla9BrGQYz6IPe9acjisGwjV
rxCdd8BI92Iq0kKgdzh3YSI2jvFmfXXlvX9XTljTrzp95W7TGVDT2PEf12dDfG7/
Dw9ZSlW5zf2Ah3JuUwVY+Wqxe3UvYgPkyILHLY+fVzswEDxZX7Gh7LB1dgxUU+lP
X6vhwwPLlTvUmAq6aDWdjRFS/uMmcaBaLHmtePY8gvojNMlrwFOtbIlJWF7Gc0Xp
fjA+Eht5FMJxkl3YpGuqhU9pOs0ZzdEC9NYtjENqj4d81lCHOh/TBbyb58oGEjbS
a1gqAzzYZLoSLLQlQa4IJ5BEINB01ZyPp/GctaEMS7hGs43xvPhluEFpMm9cETS+
BnH5DHkXsggTDXvrBK+W6Nd3jdzxyZXWOV4IMZnrLEUQrbi+pDrf0igFaPManJh2
psmhyZ9pj0iWvlO0FVOcMpTZsSM7qIi8FL0TGJAJW+ZUUuFXvq1u5Op7oS9MXe0G
NhC9RmK20BoFCin/Pj6bUC1MtT1oMtikhAQzIDQaUL5QykpHKFX7MBvBdbuVjex5
Y7+noO5X5LjjnWZyjamKRfUeudFtXRoEoGqdAZbFIPOse2O3S9vF0R6uDdVIyJkC
yVTGVCUpAdm65aN/oH2x+lg9OOLXTJC6EZF4lIi9m1cM5vrotqyp4XBBGv2YZQu6
0G4a6aOZ8BQipxAONqV4UCWu4pTYqW0NG/0xAqM1xCfs8/69PgXjtwwzJzzskmPp
v6y6Zrjyzr+2lQXedxFODLTtpHdm29QKNPLLpvgLMZ+3l8MPqG65svqFVFH8Fp8x
GzviZeEZ2q8iI/EvVIy0uvCX+DZsQPmX5W4Q9kEgzAIDbWUJ5SUA9N8Z+XIER5IL
Str1+LZUxtaJmPYzfXyrVo7H/k/z+nRPwm4YFTkfGN5xuSy6/luZ3p+Vkb7mmvTD
Tmoq6KZGGgzR+HJPouBgO8BpkzOZn5yfSrGWFrl3TH3jwo1WWodFI0zA7nFgnLlg
DS6FFG17XaQIZhfd9jcpTVb0KE0zgIjW5u2RVUP6sWBrSpPZ2CZIut8A56bXTzIk
r9aREvq0FnXWmrIXsc/NwDoNSMvUPc9HCrOJ+MYIo0nvw6qqQEvRAsCSyasvS5gn
Kji5pLKyQ0orQTPGFxDDbre4kMPIg6/ZJLORLIjjwDnmFQRfuD2c0lQzWyBzDW0S
Dq/uBJ0NZo6rll08qATV6xK++UbrTMA3alajOvUgcqy2pr2fnGf+ed66hfIfTshz
Umtc+t6/Hizxft+EMTP9M5TDBG+upUIaqm8sEqFAddtaFK8dZjgLVzjrP9zzpoeA
/UhO7LRn2Ui70yZsDUOk0eEdae5YOHni9xcTfk04VN4VBaO8eefFyhdsRnHn3bGG
8VRivCcJRx+DaKlcr301ug/iR6eHkGLYKn64RXeVBrM/sgY9htWy4TT2tb/CjPpf
Q0Ix67OO6SpEMWHNMGKH5+w+PHCW656Rvv8+kspAH+zX3L44PR0qubME4vWyy45R
4ljszEClmtx1IWKYrthIwAlm0AaxRlGjwRkkGogtTikwky6R8jPS5WHYypfAP+ov
DWZzGRl38qv/Rhqv5OQFegx+tO79YxnYJy9buYURNYSfzCnnTVgGQsBYdC9QuySs
FUfc1kkBhwUtPTSTMskS0u9zIKR8VF9GjxZO015aXdnXZFa8pCY1f5DT+ZWeqfbf
OG1xWWaanhcx3rm9gRd/wT6rVJ83X/dSqRIcSQIYU6LK2gRiCfVnsWBAOhmOF5PJ
EdxVWmuk2O+8qL9ZEBJy2iCuInr81lwxIJr4pMOov930zKqC6M/dYrTwqLERLMPv
Y9Dd7GB+DfpLJUzHKzrt64mXJG4v2+DcwSayGVOcU0+D4bQGt7cAqnyYRf/VgG60
OSwrKtjGq4fx2g3Xb8YvWzB+cVWvyqUf4CzINtwAUimkLArU6IjwsR7vhKuQu3jt
vkyxYJHiKBTpWYGV0NL5/wMM9TeJLwKUm8MTbW4B14vyI7xPzhM9ipy8/pqVUmIF
5KhhFo5IDLP2g0pmxS2N4K4G7ndl3eyi11dupKVbK3fgVOBgWFXWf5dODKHpZ4xT
9+6zyb/ep1Em012PR6X9JuuO5L3cig0+vvv/pX8Bl6/LqZi7xHXbgl+J3boKSldz
+mW/X+pzkc+acs11b7i2o4Vv5twxoKO2OkqMXiHfmTZU9IvV2IyqZd3LAS8DQbnV
G9UuN/XG4CyX6/KwJNfRe3Oo32MBqe5rVD9TbQUCjYOzbEAjuwi3RAVXdPpw45Ff
6gGymlHapH/F9UcR3HfxP8IZQjCp/nCwHmO/iFme5n6v71r+YyO2z/+cNqPJCEwJ
2HLSdFpwLva0Cfl4nhiMHCe0JTB8hJ1m8WkusPsypfvzbmy16COpV5OeEXEZxv3j
Z6QmC8QnAvOJOtBH/mqhd/MEGHhuwFRuNhMhIgNBCzWULB04Fh3RTOInk94wli7S
/b9SZToxG5m4kseUqXCsK2COspT8wWq1BAHDGV7ZbxbFzfikqSJFL4SI4LoUtrIR
OH6w60d7LHKaAvQwQj+63R6bKhuYJwzp+txKlDlMA8eejtqv9uTndd+GbHd2Xh96
eTeLMWywwcsmTQHGL/XhNzK/m66uXp2g0INThYyX87EcSQ+XgOg4zVPbPy9o+FNT
Mj38DIVDgI4PeV6gwtPFj2DTf0g/g1v+YQTbttLUEI07MUSTq1gfBr1aKu6MVu3T
PfKv4TScImphwfz0mtOyjuUAYuc5tNIIKDcyXTUodvS1/unFDjy85M2nH0xkH6jB
xCziUXhc66ojyr5kLu/Re+WxcGSkHhNBZN0ZEw0P1MB+ncWhZIIygeLy8kA8JFDs
niUJZFZFyi8YnmeYtfm9IAGvRHumUDT+0yZGuZmHoDfttGC+IeDH74M20ku3egF6
4bv/AOQQV8gwaSLyOuY0+d9zHs0eCfcixs3aEI0j77L6V9SlpVl71jH9RR+zJdWf
aSprvn3QVjh1uQ5dzy8q39K4D4viyq0Lrid57nmQm9it0agMNJpDwZ+M4vl87HKh
CatMpi2TGy6CdbckNF4L+5B1/A/R2PCm672JGmkY9Mg3wbBfO3yAHfxCGGszj6qV
JoOz+NHRVW9rPxOvQgpp2vrdS45Qc6Phd3I9nNVKCale2eC1pHesOlLCN7cmEU2l
XYmZK/D71M6xRmZOEL6oSjQuwG1O/RluJJNFNrOpvDkWnFYz4WIDWLzebCqKDIZ2
+2ut9mOz8P2wcIvlVAH5AXhTgEf5xWnEJxa+ZObUHF5jyjoBGVwPkQg1eborPbF2
RvDq45+MLF0zY5eMXLqFBuE4OfWZTEBzZoLw6O80SmxiUrLLSV6MBviNe6ODapRE
KQKu9X7keL6IkdIWd0GsFM83IL2ZaMA19ktIbeANild/zL0M3dA9F2fJHct6Z6ym
/eH65gDee5rp504UgFjxqY1A+cqQdKf94pLfcsky1/KAuavwPSKfjZFZH5G/mztN
bI/ZIX0IKhd+uGxrjmzuNZovIiW5PIKaH+tRue+KJDi1jnsTo5pSydcpRNzTBbpv
+zqqhFCQOH79H9Pm1UxjtJF8GBcQRJ6POsMgaF9GvQfZACo81aCPhlVT5dTUQL3H
pzwp/MDwweyZyB9OKa/BHTqEfYQyYhV64d8MxXvDkcRiwXlZPBGmVqnvEcA30BER
9j8PGbCmoFh0utQfq7DTEU7V2e4RLaCB6uUVw7o0Qy8d/ffOwl0wSSpVV6M1+3T2
n+dd04ES3oZEgAjiYDIvymKrBhwjo3dQ3mWRrTbN31gOfFsV+oadSXyXePto2J5i
9m0/senpbGLpxfEMYrhx+3jJL6NMxhlFJFLWCva2GVFA44Ex6DaGf1pm0uQYvZJv
QyfgT8t59++qFXHQchQyqPyNiq+VZQJsfsog0/lbNSbGn9i3G6Yv789jI9BBhc6o
/FIhYa8SawHLiIb/F/GdfH+jSUhew0l4+0P58hTy9BcEElq7bOeRXt9NiLP6vmTV
sHiX2E4A2tRQE9+J3rjziMSSdGYIqAW7MCD8ogjPwhl3QSVGmnw08LPlwvMQ0iDV
NJAkKVhj08pNHIYixm47JvCDAfleNiZrbRb6EEmPdd3dWr6tzsZ4M591Bron11qp
Njuf+tGwH5oOE3DHrcqS57XLvofbN7xAueZEGtXQhMO1KupEs51sK5pgep27l6PG
OH06aLBsnXYH7P9cyBg0d7MNxSqViaB/Kkpb+fl6c4dItdTkpm6mspNYDt86Ja5b
vuBZenwjgC8SSV7QiVe8sNlNCKFhcXyXnx9MFDy/m01TTTEF+HwVtd1XUgWa0g/4
9kr+4xKGuvUUXIcoqsKWxfbCl65iQ00yixO5Yi29KzhF9Eylr6Yu7XgD5FCV76sX
ZSzAX71S58hLL9/jWQWohtWZ7ujZT3CM+vTNY7kBWgdmANLnx50xhOb2j37kjRAu
3sUK1j5kXWyWbgwcbR/NBOuCHWUhO25e1+gCLYoUe0rij1GgBEfpKjZujgyxZf/z
cUaQxkQK5ppIEP/IJ6TK1gcODI6yzfyz8+6W6ukXC9R2WMGVwHEhN1o2ObDTt1AU
YWwLmybChrA0ZqUflhADyGvTV2DOHZVlys+kQC9OAbT1q1Bj4O32SYtUr/XTlFGY
z+xRoIRXBkwQTCFciw8iTepv2xX/VvwQQeKuX4mk59NDaaMTlRMlp0UOCjJJfETn
JiZuZPW2bqqnKRonk3aWBJYXnjYi0RxapqEJ0ZUfDz2FrV3bxhci3TONSIJx9ulC
ZuovZaAsmWf2rKRv5pEzhiQf08vSo562/Lp/UXlrKhHBc4OHhboT7JVhQbH9v5ij
ZEwbIXrV0Cku0Z6LaRUTpMV4Dp66wUPSem3RfelApvXchN3Kq5kMocS+6F4DfPfr
Mria5XT5pEa30V6QZtgTJ1kGR94Zfz0F9/49BGmShePXwxbJTVkrellbAzejZUjg
ix4Xcsu3drJzbQ8hNzRhoqjZ7fhOVwA1L7i7QYudvI+W4l5BNaymYlphN7FfsYwD
KNirsNLIZn4hUwiQkwfHFRZnV+uKe03bMnTRwyq0ED6sV2ntMi2lQjrmrbM2DuYj
y1f5AiLcg3mqvjKKWpKza5KbBss0+h+4myaSzd+vCQJUjHuAj0z8qAb0DvJ6MH5i
i4+QLGHxF1Rwfvebd8ttWA5TyBcTQQchs/J+qkpM5Pb0XKhyZpe9NPHfVdnhcrxT
lIuHLbfFOSeA4eihFF5AyAdHr5/Zcokc21/7/6HHqc/LOEg5cHK1kyF4sF/8FKiU
s4HOx1H+x+AwVJtuOcpnyi/SNHfQMJ29WORXuBhm8vykGqyZWs5XzrLaKsXl+CrB
A3cdHxAZzARht9katiYeI8UUiEAckNgLmaeKIi9Nfl2zhixS/7CpNJfnabRRbNVy
bz3DvpzToFGBQrOljXjk6beMuGBxl4jmy3jrCNooPo+BC9ZBrbpLBHWUwlf8vrk5
8FVYnNKS+a54ViyjPt+Jk/Xp8csLKn8GfN1flYetVsQg1DggUJUbKRhLimWeaYPz
B5I/WcKMKFrzVYGOt7h/v7rdVYQzVrR2x9eZ4R+STp3Zt32bk+9xmNJZOSVdf9BN
3obsNLbx2ZKqSVQ87xwVbxxlso7FDedz6eHWIwiZNUoL3p/vMj6cHj2XSNTV9AOo
eCznMmWKoPukyZHy5BowzpTvl/SIwVEAU4rv5dYhfOL+DabEjy91xnYtVLWT4hiJ
T9GpnzUpLJbTho1jMMhjp7qrpMpquD1It0FUTnJs1ZRL0o8EQAL7Ua3QALiasT1a
fR/JmoXockflrf7NSkUCwh9jKhX7J5amHGfsnqjdkvgBiUtbcfyqNgBBUuZnyriZ
sLLAEC+hGREdGX3DRtsksmh1vonLp3WJwf8E1T3GSsMEkyNUNUFhdq2O11mVKWtJ
K2FpjUl77c6fHtKKyjh5DGMGZQKZLOSLGESCaornO1MWazJa7jJ8t0U28xbBI4XT
7wonk6gE9igfJjOJqfr43nci6O0umjSmi5R+Bka7QiSmEBLjiDrZPlk6qWAJJ3tV
vQ3dU23v8RA51dw+BJFo/EL3FCEuC8m+SXvAKymqKhZn79C2/FzwEsrmg/a/m3Jx
zO5qUrzbKml5i1xIMumlhIyhyU9mdxxzxmrTtS4ro6UdsO7Z3qgoerqyzse6/jbc
TmiXTeQsPVkmOHsGAbJ1S0rBIt/KbATd3qJ7WaMyDM6vkhPsSkCV63vRBE0IZlYr
6U6/8f6m0dEOGICtPo/dOY1S64zZ1A/JQpfN3BLqDlA2ibUbb0CwSbH+PmOI9Ibm
hMb+Ne9jV2hZnc9BxYjXSm6SCjcNSc5JdnyP8706p/rQ/jHhqZKILzKe8XQU6U1J
8wp/FRCxWAbyStJ93IhXFZv8pXjKLyVkUZ6KQbTfpFuMtvgaY1D0G2Bk6KwLFktd
GZ53H/HXJj5S06Obtw9cEgjZ/4W7tFcO6yHFvw6v5VdXscQp7cMmR5UletJ9iho+
dg7jDhvUh7R2FRyOq1hjtXUsoD2vLjxzfg8sOyCbS/CAKdzQ6B7fvlLJqGmaFEsW
qsz1NwbHoXtJofbSRxHS8tKsfiTvC8qThwC3B4KNT8L5fVrOnFr8pVeDM/5NRD51
0F1Mc+Tw0N+plTNlYul96PIW7rJWsb0z0Odt2dKhwPildroxiJl961mGTXqlIi/R
DAMbWzxvGJFhxxM/eLYFRt5bZW9QOlHeekBZnwzJWxJSe/9PN2Mx3RcUuLVVSa50
xMiic3OWosWyoZgsf4z89qAuOg60BswbzZKyLpu79+qTvW7GCNQcWf3xoEWrbB8U
3E1UvPKy50VPjjTWnvetiYzUuOnxN58AryXmtyTbel5d4eFuG6f44dBzFFaRzN43
f2YZKAQ2ex6xCmR+HY6OwFJ4w5UkeSl2GQXfEpCOyHUxqaL1kyA8uIOv8LwC5kMr
8x2a6/2/iyTbPiRg83APZgQqgAFN56fT2/LeLX9pAlMNXXcLkBWioh5wfLYCVJVf
RIFPUgG7/KWKIH3k59OwfpeuSKQ7ngAtLbQ9corGj/eNsoGnoIW6H0ZWGg7SXNhj
EBTMwZYjtXh3LdbQ2W6gz20/c44LRwQJYf3ejxLfgkeBMb1pjeEPB67C3fyKwUUa
cLQUWqHvj5cOVzjyyqyrazcl06ic8whqzjePyzJ1P5/0ppk5/kIQtlfLiJuF1ilI
r+Ku/1rOlU5bjSEIL6pU2DIOWj5bMoIZ8KcTyMUwjbANrHvPiouvoS/7Gz3TMALN
nHXQpbf0/H9XzYEPAJhyCEboPPYBx84a6qIxA6BPvwKECdUDLA7bOP4cbKtuviq4
o4FtD6vM8XjYHEfPbGN4cJPli7JgBJkFFI8BaTdcFeka07EAAG07qpWAPkO+lz1u
8lkLxHnN69/zhw7316siIFgVqPlWA6XLf06On8l7PFixKw1HoGJRIWx620qX12/I
0+n8Ux7mOSAySksOj6KOFodZwvnzKeG6U3rpJHETkFPqU83qmrNj5XI22nU///tb
m+AbJooKAwIwyxIXcY2RS5sfgi+5waURHDwU0c9d1H2M8qfKXX7dc8pT/ZaGIA+t
ZNqxR13cTL4mOsj+bxUWjTcaN1oo6FAk0rksE+szJU+hWCvTCn/r7txXsYVFQAxX
MsXdLeW3/ErO5ZV4w0IN/NTQAqtnzR8WQj4dIqZh5wMu30P8mm3DnGrUA12wHxvI
M6Ts0wV3Gi8UI4eSvKOqlx+mveBgCiIiK1Y7nsCXIr8qgVDXRYDOYBdL2yYCE2+J
XrtbLFz0cgD7vwr7zG9UKy3Z8dftg7Eu64wFRlYUe6QDneWvVntHHA5+vJ6woyv+
iFu1y56cMNGjQ3gM4qExF19TFSsk0H3XgdvSiq3VcvuzXM0qCTftR2HWiy1tZTvl
RWjHXiLFKjO7G3WtCL1cdYAqany35NDtaQjMHuwuXh1Jd2Ez6G2ROni3R9UzGnt0
vVAQQcm+J094xBaykl0WrueIet8Llv/4vvTobFBgUx/b61p8sgTtr7vz3ayRlTOL
M7VtiveOqDTuvRxvQxQzN33oDoAI9H6W30SgpxIji9k1aKrR27E3OxLSVK7Apx20
lpmqn3BuKo8PTxL2rfApcd1aXI76w1r3zJqH1Tq2x+jjVNVofq1UyKS3vCvmOv5J
JiOcIStwyOXcnszfzjc9UVJ6bt61aauKKHuHXJpkr8MPbE9WBxN/3z5v2L5Y1+dz
tEYBNNCkfJr2+blB326F5uY7t7dCy9Jlb4MKks2LRu1Hc9ipFMppTt1wW90RCn6L
AxQJfOJY1QZb4Lw9BVCuDUobi/fRAOVPAhhHjnQOYAETFnpQrRnNo8raVTVMBXxL
39RAYxDX9KnYCq5bHHPl4RX5QsLrwI+RyxxYz6534XFwRv1cFmy72/nkgEjVM6lo
gI08kY62EL2gVjYHSdKRy3ayBRGEtoSdBfXctITUpLFv+/ktyJ2Atb5wTl25Cla0
3QSwdJPM5queZ5as6qrdq1PxbAlXp3T68qUCjId4rMR4PrWRIy2Bt4lx/pMdJ+d8
CZlAya6XAR09i3XDXTfvupuPTxQftrsK5nKgAJUyeQIkkj+1RBgCkTbNCPfXqHWu
FruwK9yk9GBaX0iXF3MA/uXmubH0AFKOrvzbKQOgIYP2hj1vrY+C2+kYGXQrs0l7
uF9KaOHpY6DOYh0Zk1atYK+B1uPzL1tmXMWkx/opUqhnas/Q0bzx2mbCwf94N6ET
7/vOKoj3pFqb75qGMzorMSPWt2uQ/UDwCjAF/YAHqHQ+RMnnAunQEfLcAdTzXhu/
+q2lJ6LKoJ4JqSQO2OhxoH56YSl8W1Sa7dZdp7NT3BVpu9TZXx9rujDOEBz2b4PV
w25RQZcBkJ98OPJdo2BQ3jYfdBiaqpmXMNerNG24/DFKAUTJO13nHlxXa4yYYkLs
kgiNvX+wMXFXr7aiZi4ay9W3KxVJFflWDD5HojbEBGUPFU33pHx7bFaROrhvgEDi
4eEgH2eTJULvBJ52Cz5pgiKbm+RYXZYs2AmSOj8BjP9zPI1nHeFOtxpwUJYK1BTq
fjq8tRlHvynf7t78kyIV1CJvgsxMjne+EQQNsPuNZRbRaKsMnIKuzKphfJgf1Rm4
e6PNCCv9ZJDWG9WxTQjkXRoxWkAPX9jHa/wLBoLlNK5EMd7Bd3SY+qNvt717F753
cLyORro0lCwc5OiQ7JNz0gMkvs3ctl3bCPWuaA2NNxh4B3gGple9IfRLZy9HzFMp
CpbApYRd/9qQNLDOzlGvxFJ4Ecl4EmJoHePD/qjupMvOickiBYYeNs7AAPeqyLZH
PuQMP/F9E6OT89Z15xM/oz/EC/rVZB3jW7I9HFRxR8NC6V8+qrBYIJ7XNY8gb96f
0Yq0u+YirPqzzOJfUEU7nFKi8z82g46PrJe43dYq0cjBufopSERQNEnQUYKh6EOt
hcioaSa9SPU4kNQba8xPpYA55yDsnJX2MQh4wJHzirX8r5u8lj8mFO1kZ3/2mAGG
DcWy6Bgr+U84dUGZ4P1Ahsvx4iSECNrxVkv9tLVcgNAbPaG6UdQSCtYFokdd0mpG
9RQoA7lRBKj6A74kCreZK56xRrW/r0OA1kIaRCOMYTPFLd8P8S5XM66BLYaYMPIX
EV5LjITpbSS8rVZo+xG25mYiZYdutBfMBhK7DTTKQcDUS/tbpaJ0HuWELtPgSXqX
KQ8Jty5WIEL2sSZmEv1tLx5za0RphmM+rFdm7e6hJu+Hgnoc4guiV0BRr5v5zXOV
A1rSpsJgwVBs28veMTh3LIOd4eXwIE2kzm3kPqovqvqfR+RPhHeAOiLQpZ7YjFEa
BLgvlr4gaU6iepm/OZs/Xr2Ntx4l35mQ9ZpRsao820R4g329bKnLmdzPFYQrHy5G
DF0SVpBG3+tw9GX670Lve4cWNBZ9ZvGjh67gPenlbfZmxrsYfabTMc9c2W2wW8EP
JcYpch/mgR7CxwH6KfdLseXYBGozyJuT2L8VdHEzMQkaFJcBS1o36AVI5tdWM+ec
UAP8LJO/6/8GF1LeNy5y+zO3ZxnVldirvnoQke8Udq61Exw1dBVEfOJIoht/oY0v
spge+N0KfufZouDZyXnrR2GUvZ37hkAdoTXKiv3KYPHrHcd2NhdX1WAZ7UYRZ28z
4wYxPNpXAvcP1XrHptpFOxzTWUvxwoAg/phaSm+X0Vjx3J+JF1Iu6ktJBKvoo3RC
GMbqn+p62FddApGw06eo5oCp6nxomWUB+HaRw42ajQn7HFDtpeUEMxoHh9BXSXTx
7s6C5M+DiIPtu0iGHgvDhzs9GTVLk/EM1z+Uhr+kARPihErC20/OcsFCWOYJrtsV
9GdXV81aFoAHjq9zPG8F7HpForVtDJhbLgwa96axKP/3f8dX/EiZBO/wyn2C1IqH
F+gmaiK6tzNFZnS75uonE4jZIVa9Qz7cFkLjwMmgJe6h9YHAa5/02m9qDdHixRwY
xa1Vr12OJGtw705o04j07jde/DUiJL1Jc23YUqcEh3jcf3fqUDzkUlGFNgiLwTao
b7sliXFPe8Om1qvOyO5+cpKIKa1suYZ2N20jxXQpkRzg54+vBbazLdMvqTIgPDWk
EEvxEx+LfvDFyi8lvQC9m1iGq8soyxsgh69+20QAovler7R2nGhQua9qTDvshUwz
Hr15GlLu9+oMbp0+m0fus9nE1vickPnyxs7rqTiXNRi1KU2lFb8cjVWVTqhv6Pcm
WBa45ydHa8KiPkm+X3/uA9oqmz3qeLSgoZYHjtqdIVheVw8rdyDdcM1T9RUGJwWN
U+mgEogfKGt8WX6PN2rYfZ8bh3dT0C+SIeq94iYAUUZyI6rbCWbPpHWcRbxSWfmD
pnoDr1iPjkcfaKnTRf7/8sIkcM0RUWAGiO+4MgLpvKJsjTJXVK8Ed2DV8Zg3MFBQ
Ur4ft8pIp/PJ+/6RiNjnbR4HH1FRx5M3v6hYAMWjeCQHAU4bRsGmP2fTQD2xlmb5
Hpyl359QgnWx3quAlF+RwvtKNL8TzPt+RGz4ziw/RFXuchTb1zMQrB0unrnVJJrh
0l7UQ2G37QWq9APjkwv+EuBV27pXE8P5X8GBZ4nSNiV2GcVit/FIyz4rUxj/6q2o
YrvUO375GMmKIX+XEK391/ZQhlGL5gkqZfNrIZGr94yjI7Iu8jq3PYwfrONJy1A5
n3QzOIeXFq0qUFZTAetXSMcS594nFm8bHnihUNcJ9XgbaNpLop/J6B89Nmyn7opj
3IyLxe43g/OpR05VPtB79OCJ4h+l7qPVGNgxdE7GTA98uYsFXgTlSQ7K/EykmPWz
luNqSphJoqKjwug1qGMteIUw6MkZpmd8l3gh7+50GWWz3UZofJ4Es78B/H/uhtgb
nHC2piE1RaY1fb7bdzm8S3fiy4qOtmXUuwsxvfj9KwHvFqenuiwXT1N1CRhqZ2hz
DN9sm2ZTRKHUc4CQoQF2dDJlIgoBhooX8eINiIx/F02/v8/xqD5iVF/yW0nSN3Fh
bXVsf3LuGJl3EcuibsZKb3W2Gf98zD2NeXn1PkaiyavRI9hE1A+gORssH0IsykvP
/Wv4T+egiEb1gXkmAF4P9+nh41kbCuz84hF6ylAdQXqCmD6cMWyru6j32Il9Eliv
2enb1q8iDYr7mGS+OFJT159QEKVKGmfHsVn34rtYR5w4CuApknBz0/xcDFBofE6a
4IWwxnbbh6jAoeY+LTGHxq7mEWObNyoZSyjW4oJEbKVZdP0HfS7U3Jr23YlhhzyY
KoT2pSEVm8woQun5Lk4z1W926G8eirv51ov61iJLdbk8swcOz3o4vFUM83RlvYeI
0YA9Any8xLwkRNYXyOecGFf3wuxibYLkJSKv933xgE+5u2vU0VOJ5oEYiK/8FGFJ
EVcCy7eg08VGuFbWf2A7Lb4mPmAjeNheAvOEY9aHoWE0jtgWSljd1HvcSV3H8KJ1
sZf4TYl5yYukXn3Ghc2JG5O55TQfFvmV3KtIK8TXeHuvItA24oD7Y9k98/+ZFkos
rrU+2g2TgQzsd76uCO5o0sgTLAo8UJBqm2HrWsjBDHiG4i6U+NzGQWcMyh7egy4b
lGnapsJbKRaY6j5v+3RM32hk48TYoK+uZ52wPoPQnuwB9BN0KaNo5Rt0nbUuuRKq
aeTxTznXvlDrKh+zricEI6y+y1wctAg58GReNYT99kjJvH6xLD2PLb3Ng0+pmrP7
xBA0tyQz4000mWdC7IYE7XJmMl69KGPq0ux2/vLGgdJaGor3m53Cr4/TxLwFbqGW
mTjkoxwqvkscIXCuCeOiAvXJxebBOMDyEP49sLKWvniLneS+CRtEtTSfTv/h8nyX
j4i39kXh3kvYEsjklJqR4gQ1X4AAl4LzTkSYYIyAkez6f2rPeksc31NvKole0O1G
q23/wek02Iz9iOLBZOeP5tixfSOwhCnqUOCZlZbhJJVWp0zT81JJMBjziiVjVWq3
My1VB6Te7KGOtdChBzJWz8EzeOVV0WQNJU/MFJ0SlVdlPx1yWBhv+L4nZWLk3KFV
/ii5zz81cNHXQJT7xU3+R2N0cxoqL/umniz/uuRk+apveI3viGSXujV2rTxNV+Mt
1hx2v7pGeteWk1ctLOApLgUgWiBLkhvHXByvjic04ztc+2wrglYEJ98uG06qoSWO
/aMdbmAEVMh1Zx1f9g9/nosHWkx6/CPRShviUVnBxp0/uVJhne+uCzg6R+imREYp
4OBKgpWILjBLPEOJlNm4WocU/zyaVJEQnp89Qaw7GfXPZkhGt+NgazJ+rPh8pmuO
H3C9LoHJDwmCzp9Zo5O6NEc71/GiiFioXQEY6kmhG1yufYpZ926CdE4no99A8Gis
eBJDIxXsVrJ4K12AOW08waxl+g8M+KnitfxHwV+JTi6GduneUzCdkCrDqm+dieeG
HNfvRsZn4FQfU07kioMB0SQTKPKKkjm2O/Q9o41xSejEGk8ob6HYR0BD25fTs4Bj
4ljEFj/esdlHT+ddK0hjD6VYNbz8c1XjE43VicWbcu3Pqbl92tJ/OkNE2uHTzhoX
HnFxBETVD43XczZ2fAsICY6kWxntx9UOX61FJaROf2Cp2ACEAhs/votTTmlP5qle
7b2mgL/HF68/fWdCgWZg2w3GfrdM9gHKtQOqgDcTBigOGFF8aChHMx4Dp1lmZj0b
QsFclkZUZIQQJdYMEJS6oEX0+vscerODUxeYkkx2riz3NUTkwithTFUqf70hPpB2
aa/X10Ml58aE6WmwmZ4YtIGPWyuTKuCPyw2tMr4uW0n/4zBHNq+uOXrz0rIHQ+cE
GPsFkAknzGjEXhc5hKOoqB+fzghIYbaIpvtxeuvCRLip3GAnGd0l+2EQnJp+1k1X
0nJy8dZVOMfPcHQ20QWYgcZ85aziWN5vrrCNKUTDxXSBcs+pIFa1wea+IdOfNQru
beWnPhgrCWj2SMn6nBM07PLC8Y7bxtihl63YfmzzbmpHn7aJnieIyGqPCkPv4Mz8
D6zjAaIsIghoJYL02Ms0lDIz2m58dA2aWmWPwy6LlgNfSZmS96s8780jP8IgnP7c
1bHR4m2jwawCOVqaSgpIgZUGfZtWgL6wgsSOaiXhUkq7QaLW91dnz4RmvATDR+xQ
tZXaUz8BxV76HBzojxN28g2IZAp2PJHVCooH5D97GK8HsfuqJQIqSfOTlJI3Yigx
lftMv3xPbyyriJOO6UvCIbQL/CUxtj3cfFgpjaytHuog5s2D+2wCxsVExyOOzf6+
YBTohb574I95Kk+T2WEr4H14Uad94baSScdbc4172pCgS2Uo8IgXWHBLNWjbHxeT
Pf6Ec12xbRaVFDthmRmn+FbOAAJkoAEHAyFXAvbzk0AonWPhqQLYotakkiTykfzL
D3N/CUTmKjwpahw02yh6D1QbpByApNBkFJxvu+ByfUXZhW/Chbyvn/1WvFgUmAyn
MQ2fCwt+YtHFd6njWFOqmXVpihES7BziOUbNSNQiVFJyeLwWzIs6bPDWnZeyfsTl
O0WJVG8hf4bqO4/VfeeNgzj0y/CixpF8lPFQaGv0XSAIlcRVMvYkGGytFlOB60EQ
Hwn0RxL7Sr6MBobHv180C1ZPKEtM709XyshFAMr3F4MFDFrIEpL2QwbfCOMlohuC
8e/YjwrGOF8eau3E/IG+b0gWpf36B7tb1V26fOouUWg9m0/O/7dNa23d8BboY9TR
Iza+dG2ACTKgN5yhEhVSbDe4XHSPkmRdUGMVAVvDXEimbypl2RMhdA7ghknZyijk
i/7ufY/qEgCo1s0jHAUXLv0hB8FeiuBz5VMHdGSXZa/xEJYJf1ZpZARAlCAfa5I5
39Pbb/xTtvdS4vlecdliad4/IjsKuTFsazal49kSlICmHqoxyjylIOh2NctZAPcY
yCHXvp+tPRn1ZdBYEiQkMtvT6ysKI/ZdMvSTRcbhIG8eFMeu/1ox0Ab2Y4FKmfD2
mnHyWtcuD36jf0sFXNFM2bmhGNZzhaBLpmXCvxexaXyUTl+RcBAHRPDot53XtSUX
04BTeG6/7w/FI4xp/aeoryq16PyhXawYr3osyYTba0AyEhLy9c1QAJt3w5MwITdY
eyVsim6GR+eS1/q8N0nNhrkfB60mLd78yIlpCogEydSppBuR8ry38a9RHg97DbVC
o8dcn+MwhA7Jau8tSvhvRfVaA4Jqy6UmRuKMArcxWRzY+zB5X7Y/8Z2s/iGm/gei
fybJJm37F1shw+NiZg0HfZpjAVDS4t2s2MXEzUBHvtC4ZN4j6pbvajWCVM8LhX2K
6t5NHcbLi8kJQ03jK1fttF7JF3iisoGbDSjHLbqQfS7tF8wdOJV/4M+Y58I9rwg6
7rpPcmvkNm0yNp4iR3bRE9TRY+EykC1jba5Ka8qqwql/5Gtx7FlMvNaTZ27gf+Yo
ITqtkzb9XkiCVEyc0gUjJYXEx2bVTTyIZs3HC9AED2eZNEIVD2kDT/yHUz3080N1
NpW5M3jsj6Z/sZHs3vEcN9zggkEd0Ha5sSyWfo5jIqQZoG73ngM5BNy4mNavhuDd
NvuDtbW1fs5jOR5i0aQ72+5tVYG86OB84d3MqiSED6OrB7pd56lAcC4mtSfrAgcT
h6MCy9UIzVEjaG6L5bS/FEel2f21J6Ib+3sZ4tOS9iEecjxpRTgwuFCLZmqSj9dd
F3j5eWws8X4No2W6zgPK13FC/lE+YLrIQJVE1w11WTuNNFyQ8LgH7mdz7aN4DJNB
kbD8ezmI5P0Wl5MPNpWM5Xf3+dwKNbnmgQyTdLpP+EOShbn4PwFUfwbEhAfNlrYz
QVKYZkQirdB2xIW7/tb8kYbqgHMMm2USW+LGCn2R7VtCeFZLROmzzNGjSaowyDIy
Hmv/GA1xu5hgnkcSK6BiO7+9wl5O+m6mZUXMMRWuHGQsmuBJKwzeFmHSSkB6H6bg
lnnNJuN6eGhuA/E9DmUp1zgsewWJo6Rl3MyiMNSuiAtKlbndFvktnsmjkC5RHYD6
rVIlgcGVhD/IXVauYU8ynT22fF5bNE727f6l3VgM6+clUM3JpcL7/4LmIm4SFrIa
80vm/AW97a6sSdNmpzXsk72VKZWLXBm91IAk8O4VG17M3Y5UvtcM6/hQLg5J4tiC
jPtYcakutuOfns2+1ZQJsiAAwGHL8Mf0r5ujoNgXOCOA8WF/SazIO4T1SYzF7iO3
J5Xr7yX6x9yqcBsmvhPF9teMiTdPkaxPvmMvou3fbutFG9x4orvfVVHucbLJCxEM
HV5+vA1jIClTcry9W8TNIvNjiWL5481r1aLwhZ0Syf5DJEtMLjdiEYwbyajF3fdd
EwBgTJLOHosmoA3IiQNr+cHEhBw53u++idA2XNoi0P6u3MQRxey9OWlLi7lI8evQ
2rYmBr0h8NHBDvnryEoFRGqpSw4lhDSt5v/4PRqpUI7MhsLqr62EhHsv3Xzk1Upb
JJ14OlBBD1mstfZ0rKsgk2+q7yYzcxcN67b4fwVDrxCtHi9G+xIZz/3xH700h4c9
v9TX+mFQCLN32EVlDKRjbM+5kiAW5zhcy4Z17CtIOoxrhkYrPeEhNV15Wyqfhda5
T4SCz1ZHLh7i0BKsHyiRESrQtb4y0n45el71oMOqFhK0QRJfZVPM4cduanGpiVTJ
J4f1BuoLiqmBqIcsgj+fe4fBfIGMfmDOvbvX3thittbmqnpB1ryWawk9Mo5o0PAm
MC83e+b1orCh3INuMjq7WvpQBEA2k0slxDSRrdRJ6JoQwc4BhFnzO750ZStcwzS9
kLqhGQN1B1dJN18PHtt42Qavf1NZbR3eH6SD1DocQSu6ZGThX+/a6noPcDyqVRSb
Ze8PFWtU8TqfkfEic/4Uk8yTBFm69JDWMWRTCj0kz1iEL3Foa8ufXa2Qaa+GE3XW
CBLu+IoMQkwxiMrCs/us87tSoepGIiJ9xpR6qoHEKDW7Rye9ku/VBQudZWWzY/gP
jkcn39AeK7lhQurnn16EoxypAKPr5XRmW3GvEumKzHfYBxuIXrUzvCan0hp/6DKg
1Hce3wCMh8jwBxJ+UgA4MOg/rIBP6JydxsdArRMowUfltyzrjLuPSqsElyIx432D
Rw11TrLYumdr5VyHnkDnxttL2DzcG6s6UuAduISwPYfIiX1ydmBEAJSpjWnEmkN+
r6CO2dCCF/iGKieBig+inF9Ajnz3bSGs7Fu1+DEQwk2Kb3+iNc9eBLFwglYQK5eQ
GvNgnCkZJJ7tea0avdWmiqjiUMohZ4rn46qEx6XmG2RPiX+fev0evrZZoj9PPAd/
5UO3Q2xZbLYAwjH012J2G7SauFsc7Sy3ECVhy7iWDe+QmNt0A0gqAn7q2D8kmnAI
2RXnmkTU3BOeXyWT6PihFL6fvHjIAof8YtqT4IqLXErOGcqRDhutTFoduj0T6X9M
wUqmo1GxNGmotXzbQRMZJHlvhzy7OqmZTh/W3Iq3FKjYuObaM8/ayoIcifMWZoNt
i4C0BAAfsE/XLhskVA2+dPCibsfAUpVkvI+7l4lEYBLT3wCCKywEqtjUYJlJPgQz
bPfxydFPmz4l2mM3DqjdcPwkhBaLjG0sF6Cl+A4XdxJZZzO1hU4OfNRZsTKu8y1W
Xc+RdUS7CJfvJRSVBNDvsNma8yNjsT+LCuLiUfDUGAU8arPCYKwH37JCno3bN0ca
BiMAhgI7MCWkjVsNyLxoEosVWdU1FCvL45oLOdlamZi0PsuzlNQRo5QRXiTZIiCp
5ZjeW5UJI2Q2wYFo6upHQ8kUcDwjdfjjBrYYORAzylevblchczcE1kJHk9mY5QDA
CpPpfer7SAVi9u5GsS9RIui2yVXnfkl5xrStmWB0cq2y1pb/tV9IaTui/2ipaw+Y
EwNmyy4+6KLP+RfdnIvN645Zg9VAPZEaLGXAFq9WoZesbJ+zaLYyGVqqEtFgBoDT
wqeeTmaP8sWE9xyvIiYR3gxvoHXkoRHxnKMWE44qAVJggtQmS+IhZEW8z42fu5p0
bnOJx5fCmzPggCv1UsdLDBNfGXdwWqsY5LLLdwzrQ/BrBJrycPuxulEb8gIu4jkP
85gxx8eeVDYc0Bx1GUF4iWWi9t9tkmO8o+z8OKx8EMZ7PjKZa6KzJKxI3/AOi7CD
o5DVUKAN/wpvuDARWRsOw+XLBjcQD3FqG0GXaTFSDX2RZgRVCaXZAYY1AiFieIM7
33SZyQSYkPIKsCZwKxF35EqkqHBNjEWkmVKtW9xkbRx0QtN9zfZolyCS9Aj0/MRo
U9eB40vSP972l82DdcgtmGCsJXDpz78JhCWGxA1WbISdXwiuEEKVYsR0Q8xGllyz
eeLbXmUSAOFWmOyPhohJ3VijvFaT69g9/zly3XGuJKnywFA4gFGsa54kdRSpJogp
dJT5TZfI3e/4oAUTwY0Mx45cNeMAaJWI6jV7fNFLpkxp0Iwc/i1MOvK1LUpVRABU
m/0vGD84mp393O8QfiIOwHzMSe4PKhrbtWZjaKcVIAlimyqrvo8sIkZ6TEHh7QUf
DLM+1wiIEAc2lRwewDgRmOhIHVVQqJY5SLRosQulh0CgE1VXQDfezhcTdPc84pgS
OK9bvrINUK7mPqx0XVI/BxvKodChhYXcubcUJIpD4u82vJK/Xl8dIxkqyfbe1KZ8
z3FAs9/3GWD96UtPhVWXD7FHBIt30KlrtfYPHonGuA/4oooRXd0N86exVTxU8NQ+
6zp4IOZoPZ6ToTuhfD0iuV4u8rEkvM/gzIZYlK8VjvH5XJy2guQ/7uEaQFts5v14
mYSauck8R68h3YBlQURohXuZOIb5Zg5JjzS30NnHHxKJjMHp7j6P/ohGL9K/uOr1
hs6M7bOjVQBvKPll6AsKQFtCeBtS1Jw+iZehmJJLN3P7kUiWWUO1UG2pjE5rRRhC
CYXG9ap9F4Tme5B1ydqfJsF12cC97r5rDKJg4OSnQ9PfCJygEvlxeuk1IRmmNNTe
bHtg8/Mu2Ue6W+WcCn3L9zY1fQKqKA+JJ5Di7Rabkih8UAPWzj2QKGbH5nHbglsN
GthcptQLHbFHyFVumug3hRMKE6B+6B27n+kE9wpiVZ10kgZDpyWHeSJeh+pyLmgJ
PCae1ate1ioYGxzG9NlpKNqsfe6/KZ4iXDKHtMF6pnPIUEbkiIlAHm4Mwo1OuN8p
j+dlP1dvanYa0xGeEyU77fXKiKwH5duY/M0rqr4RwpXDwkFdQJsBpLZuw/oyZuTo
cY/ES0cxcx3PqJQZ9IHAY5bBhl9F8X6lf+755/f+rj/Dc2T/7FiRWhHJwj/srFhF
ySPA7DQ+LUiERngZAUBU6koHI9kOzDJJ8lOw7kDav+n/tOsw7hjIKEGVTpeF5G/n
qCymtcKg5cCaCWdHRG5wO2I7iRZ2s9I0/hIMwWNoHry9gIHjWZLP88pd0pVMXCAA
52rz/R+e2imL6Pso1GobCwaG2vi0w16Q+r4//kjdmviK9h0ACIlwxtkZ/S+wdqoY
pbBjqFP8xNKHixQ9F9fq+OHtBjC1aupzNJyQTAJzMS5E2MEwxGz2qrQ+uSpegEKx
T/FoZb1n+9vFOQPglyGmywL14ufvIzJb7RjUsymoCcf3XlIRb5vtozYHIkVfAlPS
w2sHBYCOXQff7X7H6VbQA5j2dKG5JuK1I8s6N11GcOnFKnYQTJh2aAVbAZfyVWus
ZYNHeCL2qGjLYBi1BhhCA1e4vPqhL0HATs27LJOPltgqXp2ncfCV5qTGMuNwsCPU
vfSTBakP9DKkngUy6Erj149fqkfyme27o9peX2iuqVBRDPFMpoC/3lS0h1+nxk2p
XsNdrwQrHy9bKOBZTtPYz3LK/PaIT9JYRh1NxyGIGQGGB3PU0IYUbRyRkGnyP1C+
Ese+Rz05NMcyPsQQlT2PK6WsqxsMwRxYZ0qgc0ELNjihMOXfRUiwIhjC/anTSWC8
hUnlZq1p52Rfvf9W2+ZOMbqtR+CeZaiG0p3UEXW5AMB+TBuYsLjJV86KMFx7ZcQW
9nnV8zmNBjGIGtkDP37l7IDBhYSTHDstWnUfI7PruFCHre9YFcm3UM08wZ8+CiJ4
1bcJDFGXKgbKtPSaSuFC6wdDPUlHJkyTuCxwss5gZDdZinTa95QW27sBmZO8pNpr
eI1ivmD+y5gFK2qv6b+QZDDp1wZ3zJKuu1qKl5o1lppIP4LcKkVeWZD1B4nzJiX0
xgGR78yoLRjAfA3cgPy8bT9BpPiJLIdT0r/jF78PvGh+qKs93YCbUbezRAFNeido
0UC+gKLXE0JZneYWqJeoZGWApk7R+T2+V4MtJlF5Fi+DJVbAg9/E6iDK6t/1KwFP
t2aSWC3QRBnWjkiiWowDto5xze0NcXgRy+jdn0opFGXhGuzQvFIpRAIDktxSZwH/
NC2GxORB0IzxmA+ucnuJ/izrLqPC/mEJfU3j+CjR/TElNouWWrr5K7x7MOFVO2bq
ydFHkuPFfaOAffCluvw/Qqqv23aEuihwf3KWBA42arlXf0dbNJg9jMvpQuBgnZO4
ZCwsoAr9NkhXVQY7CV+sqmXujSnUn8u8MHif5Kr9El1PVSV0ZNQY1TKttT6fuZuM
2O6sGRMi4klDuuwMHTBqQVbnuc3xeHX7w5r8kQ6LMN3XeiBq/8Lp3T9tL7vtJwFT
RVKUPUt+CZkKL4yDB3TcqEvGdC8uttfKcWSf61tcQFxWe6unDU9d/Uai+W1TPrl5
dJAo8Lu9T32TBkK3WN4eWhdrt6NSYSY3rdcnaNfdle2+GvVG99R+Pf2C1lVvmMO7
5oNpT+sPzBZtIeUHLMQO+ry5Y9+uBeDSll6177JMf4RSI3IgJm0t+d0+CNttD0PV
Zsd7jyMlzgxg5nYULAfQI1lOCHINsjf5xBcThePYY16fFIUD7RLWjv3Lqg0CZFC3
PcSkNwa0OJw3BRO3OxXjBDeKHM9p+NSzOXsgri/kw5cTwkCwvfKLz57ULasBRj6K
glpUQRaeTfz9qb+15WS08yzoKPDq9IvUspk895ptWaS5PKFUh13XNrZT3In/+TqU
OqExuybSClq8u7yvUsGKxc505M1Ee8c6Z9LRPm9NanR6g2rqzFXEn4ejkyTy8Dll
Ipv0wzPdcK+mnHkNKvjWJl+fZ4wuhdBK/YNC3lhXTKNTrtKW0l55VCznALO0o0J5
p+wFNfDj7FcgK99AsOye8yNoU7xWzIhf20UnIihWZdTYykuPJeLJ8rQA/LqSYLvv
ixKSJ2ebp5x+41Od64QZR06aU+Wnn/sw2JAgqeuMprRddJcEe0PI+KOiTkbjUH/p
oV4MxMXxri6kq0dHZlR5d0DpNofprXWyCrbt2m+ldJOgBPleK5XWuyi1mj1fW8ug
zWkrdMX0IRImZJWqbFYAO19cn42C6anlafkcBS6NsyFBssRw2uFjqYCdNytTOLU0
ugtOGSqFw8d1ETltQOyEWjm6t9GU4wp7mjMy7oET/VVBO800GpFWHl/SNcEorOpQ
VJgCWJZlWS2ZjAAjRQADrseReg+S2TRDRlzqjBNnxxW+r7m4dgQu5o/0JMvW/1rE
wxvMKOOG5I4CBovC+wCkMY9eGi4pyOYMRfKupS/3+yhHsWnWWO1T4dFcVJ0c+uiU
buZo4O/P67HQvygXdrxK0fnV6pnxw5crhDk550kYjAMhU6G1PS7T3ViZWyt1lVLX
GGWnQEHMSgyLak/34507n3s0f7zlLKAjcNarfUfKUo/iLFsVCHbvkl4GRoQo7ja4
0+wPFsxqnT2ZwXY5V8KkOdqaEdERSx9ksQNlCKDPmH96f0O0NkYN0INOmv0BCUcH
lz59NNrc+G0OM0H1ESE9/vUfExN0KEUW3gkQR0kCOFEsTaQ0o9mbVrzgNNcwTR14
H4b4ugW2tNYZmadLR7RoR/w9M/XnPENDh8fFpaRtTi7Ylt3FW/7vB4/oXbi52Hne
q4X2jtc1QOYlTyLLVkUyJI08iB/UGWIUxUirkSkAfGsLwkyER6waOyO1NYzoV05N
NHoqaIga3tr8UDBo8YFedSgX7LMF64LCWSKrFfgFsiDPeuNM1Jq+h7WVIgVSVHIE
dCX6XPAiGrwteRrxkHwR0F6Hc1C+pFVkOUIrJQzI24SD7vP8+SvLTPD7cA1b0bKi
U5RQwHSQPJq1disbfoso/4cCL7302+TqBXTCnrnsHpd10meo/PixyVKW/hl2OuRZ
2I7s2Gz44xsuVJaqZPyvlRJimF7xwQT5M5lwLYIDzaC2S0yd6TcL7K7WhOPVQtS+
Uwn4EQ4Uxhj13htJS8xMPXemKMwx0jLbXVR272BGg1ChKG05/CzNCNkCVIoFEdTd
bl7n2h4ipYVwRMHiaLDWHCuzjH43n5/gpcST/ZFortOfXcX/9x/4eJvtK+gfu7sW
kY3ODvGY35HY2JqVyyFaowpJVAvLcVUwihHzSuw7V3sWqSgrv79BhRPaJuhNGvj2
LeTdiEetLqUoMZSUXqUBwByk04kYyWfV1eE7O9/HR4mkD06DlExWclHSaQRPu8XM
YSyY7keg+0eAcbr7zjKervESqyVUMe/znPJnF4bOo0trcJiZYUfDGp3vzWTnCfwQ
nvxqPvH+FGgz6/aucJSSbAccG4jx6byvWI37xu2wa48MJf1gldYx3+UKvs7/KonL
1YkoFOOtOEIchVS1Thr/o3IryKm6PsgmcwUkTCS9l7IjsK6DEe6ra3c6KsUFT8Nt
ayzC+IRe+ikw7hqggv8RAVxoZJ0P+S08mfyfX4hE0RiafbldcmlOs+3jKPAWp0d1
ACV5KCCi2GSmnO9Vl89ezNdUjPMZDSoU3/KN5LxlxaQCRM6TJyxU1yCXbj6F4QL/
ya+N+K8KLE/J/LzYhrM5jTbV1dX1bVy7f1T6OMcAzZmxQ02Jk6ZX4d6GpWSk3tP2
ZWdBBvbLRvM5L39KGFsDrL/CgXJHLUrg4Nf5XrA8AHtlnxOwHCDkqdppbeytBSpZ
LL4T3MH9sa3FjZ+7lWcunhkoC5eipLPn8KflpkWuGJmANCMsgOpnOJvwrOA4/ALB
37HbWUjw/8h2g2Htv+tUXiW0K+2OMB9ZSSOvU0zI6SCUoHKFtCOFrLMUd6zjPY8z
Cfd+hIMpJ2Y3Hg5MpaNm2gscXfq2tFohkPcfgGz+SGQgNYderIIurro7zosYHiCy
5Y8X1Js1RcsX7HxnpaquOtGLKoTB7Y6ekzmH8qu+DPTK0fYWib+4t7vEJ562A01q
1DLBywC+ortuxHynVftS7zm0PnVSZxrMcJthoxoiNg+hg1ErqU87oKbWDFEf2ClF
LCFjueAFlMUKnV9OYoUNoUOMk0eELWaecEKUuol8EjPrTgsjyT8TAZUgnNJEgfZk
+tqTuffsheev10vl9TbHQV+SX53MO8yE6qw86AO9jy2KoQinYTbisMyDs+UN3VSX
6I/X5Jxh6bKKylOtHV+a7fY17RH08ZSrzWRj+RmvV35a9TS8Wl94P9kNaRYW1ppk
obHihEHa3A3ppoacC5MHNcECUE0JxXcnNuDiRdc/iuSHTWz5bLAlZ5RP9OSzBFFK
u2eSDU/Qyco9W2kvdJVVoToy/fDG2XnOh0u0qqcuEZrTNjFhfTfBXC7p7pqet1sh
jqQu/pEKwwggCgHXEeqEiUMZhcHhThBIaBLq/IpkmpzfmSWXpOS4jKnNc8YOy2gv
XP1S8IEAZoQe5SgBe8q/rnCyw5AMXp4O1D8Wjg5dk62obHoc0FNsGLfa0JZljrMu
Re+IFSCinGbLwIideCUsonhWr90atMU+B73ZnyOUR0QkcRtEVduDoknmqKAiGJRr
OltH9aublMv+eUuf1mHt1kHXGp666vCSR5VBx5clTaOLdFE1DZnAPrw0zXgsm9GQ
r0bHqnuQ5HhvMZZtNW9pd3Q6Onj/PAaJKkf2PrtI5+hwl1XlE0xfJ51FhPsx6WJH
i2HGs4rpAGI1QOmnN32LOCib1+ggH5Rj/JH2sdFAOmS7TELANDUxV65+WYpLI20a
sZQxbAQ7XLS4NGvJqN5vWn+qQIBlOzoirs9iADpe6ucPje3vrTXqC/8QdRzuGei7
LSoqqU1sUSLxHU5Qq80y5wkfNHDWv7mnejoq73M3vu+ti9MyBR5UdWDf/j5ZhpLQ
wNiZjVltKsCJGLvy7O7fTWoURQHeVBgxEtW0v1PRIzjWI4YMyZM2vqgjBmW79WU+
n5bfylwCNeFTDHHTVBpAdxwR1lcWU7E/1TmAe1HF1Ha+SX5jS5ShWU5oaIq4dKsC
Qi6g7gusk13xymy0x3FtROAlqbCJbcXJU33zC3xOlV0zVyI5glYXLF/sPjViFo1E
PO0UD3Frv6z6Y0cBYuZx/cSl8jYQLu04UNHf+mW/Loui9fuNpeaUZSQiEJ3F2Lbt
Kzqw9ZfA41h8uZ+cL+KmGbU4PF67bEG+26FGuPOrrGpGiEBOo0gWPCsiIIZYUVVD
kQbNdPnet9dOsL0CBSUyrfAfwNPEEacOE7vHX1aZlKdnX5X1013rzM3Er5B0RhEV
l7xEiaptjqJYL2MKUajg05DlZf6EYcD6NLAoaiQLUNqmwHrMBDIN5di7Tok/bW2v
YxgvepWzfF+wxawznosJWEudPHgIdqClG/BfyMLrE6Jq7vfMDa3CLKp1K4cdAYjG
VEt/S6CcebR3zqCJA5z4Xy8OttCOOL22bQSDjytePWnDEywfttQL4a1Ax2ssjIYF
Ghsjft7wbnj4Aw38qOTSqW616SKLBCRbicAiP3xCnLNqY+irle8SwDNf3+ElgKKy
djf8AmwHAqB17R0x9YwCfPpoIcZDwEkiPgF/nS0SUUdrbzwkrPW0ffuiN4zrMeXc
O3CFWlkN2Mkpd6jNW4LoO4G9kQQZUvbgIq3HO4DWJAq2VYBR4uCT8PWL0DEugzuU
qQk8SM5nQJn5/bC+xT3urlwrA+D+9V1sL1lcOVF4s7PXv+/klRuFifexfvuP0iAT
svDK45226PYPW888D6SpziFZiQ00/l1nL0eT/Lu5AbUvKD2evxka4RVsGjthGBYc
B7/LZ9nIiJ18d09WkjnpH7E6SQMOKrjnlK4mhz80b7cs0WZrpAe1C2MviD8q9v0F
jFzzmuOl4FMlaXdqzzX8K8nn2IHaO6ZUJTv1dfdml7qhoiqPsO0jd0lfB69YosYZ
2k6A6P50VA+BSaIBJdJWHg5/DokmmSrW5r3KsQ5e2B3mOnQvBSREtHQB6+EmF1e5
gIMUmFYvHW7ye6ysM/jlhfEBK45UWgpDZSTxzuWup82nsg25aNNvSAaLPqxZ6cY2
hZK8iVEr6RrhTg4E+RNqtHRMoeHcItC3Lb1s3h4TEpCDwh7nQ2IWIGoo1ZXtvSzz
UNrlWgkxtdI9p1P7rs5ym9QuPJPBzIl1BqL0DeIMrY6ZeQrcmvoZjHst22/HAVLI
YyB9tF13E1Pft/TInZDG/dWeOANzx7o4L0tXa0wnoxIddap+Icv4WhhJwstNoCPc
v5XpyFEvSQOOaoufQHyh62sUY3k25SKHeksYqkZR/bknzhT/FIyyZi3qR/G6UELC
S3o5S63H0R1MbHry2z3c1WizMb/duwhcugvfpBe2uPVVeICGJGS+/aeR0JHCVBqB
6X2qvL5cO6FpEL2VYTq8IN67nIlp4oyMxKQxDzErNE4xL60H3IG61g1nm0NL9sL2
8UzeoTeEeNaJBi+GvpwKzozc1JkYh8fweW7hGv/6RM7Brcmy3VNCwvTi1AljmA1e
zGUvWDkENsULfo/wcBydM2/VdT9xZ5h3eO4EH3Jy62kGzvIbVbxg+B+1UnyWwFfz
pyzfavtcjGBC23cayd/thFQhtAC43T8qvS4p73rEVsWssONNB60v+dyg+M3BGwOt
InquctxjpXwfhezKhr6cXmXPLAOEwmrX2V7MHfH7AYdfIGSQn29+ZBuzLotVJsnN
6BiLHRC5SNyVW8T0qsJOG4n0LJtSs4be7xugdTBnqeiYqz6rJ5vRon17Mr9FZxnM
U4ayGMLQUB661YUpkwwOmCceBt/KOEPlk7q++m3slEjqX4w6igGDyeZur7iNgtM1
l8zXzdpQUnBBZP7wCGjW20oftXjrVYTkzG6UE7QI4xN4Pj3m3hDHs3sRuJqdGTOr
88ZUahBMTsUONXyJQE2Y9HMFWGVMpLiclvd9jBWZxYb5lxkYgLENHnzJBTezMbdL
l+nzuEaoR30qwh3F8rxujU1feUEttBkdplhP0OyKGWXJid5IT0IEEA8AsprEcz+M
uy6koJ4jycd4CVz3uHJaHqkelSIJC0kiJs1ju32bTle2ohTyQDlcO7Py+O6TpOOY
LV4OPEjdTxs5pQ5i+iz0ZBGLDnZ1DaQ6PKQdRiMjvUijO2ESPMMUU8h9oh5o9psP
z/dWRpUBYOJgF7uQyYJS5N+e6RCWCAKqeKlNhxrjESOkk88OOI3016G/ZE57Miy4
akcd11QRYDHP+YZbs9OXdLptwyURr3vAq16xlEbXlV6KA8FXCmDtS3Y21YmhbHmU
z3vwcRx6XKF0Ocfb6MOiDc6B9Q0P/h4xy0yhBG9kTW9aU8J0N3U+FyBy44xDogz7
W1kelTH6w8084J0BvHT7qbTwvgsVgRalJf2RR/sZGKReeXQFB/ntFvb/ZXC1riJ4
n9tOf4rtTNIN1415Qv3sEVI5urW//HLho2iVHJCKgVRpKph8EkpUUGw/e6u3+8H/
yco2U00Wpbj0cH36psFxOvIEAdHbxJQ2TSnBirtEN13inbtuMTgzINRsq5a/YuH9
Bwb8+/jnKU3dWosEUpltGZ8gC3cK5azD/6KcsZtNSXIw3nx0aPLePMdS88lVlgrV
tLtpqXwOQu6P1WyhLtT0Sx458YYNDhZ8xerkiO/UzUJmFelm7cLs3+z8FQ3DA9xq
qBBODDICMh8UBbFYU5q463wneRH0Bh8/8SKPwa32fAJ0erlSGS/2fpahCkBHTvru
AI7N2FdHfyqnmroT41sB2XUnS0ImhuvBng5wEUEG/H+kjDTrjgo+CYfCpxDbnVze
P3kb5tBiK6rWa32w6NJj/GD+Y6km1ASOGsgoBGB6OgRCyoqXLEsKE8v59bHn0QFe
TWOUUkqHsB3aTqp+zb125rGzeK8v43ORT0oL7NioLPUPJ88bfb/ciENJ99Hx7UJj
r8at414j74a9NxO1mVtlJn2qRo8wkThsvvHpPyvGueIRX9VFIU4Dde6CPm88XTXm
/H3VBE8idd9EvtmV8OoTUyAbmumx82hdkBJnylWHdJgJByow19vkqpo2ex7atlzG
9bUpU7uqj0FR8sKy6tscH7ckJ1lzmenstL0wBIUKiYemTOb1wJKXQyVWRdk1sJMf
Q3IeE45FHceBcVKiumFG7ae/XtfhwazeiI8o3jTCunK/6OAQKKLB+GJcya/z4W+o
WpUUBYZUeQZ44CSZpmpnL4xc/hHA7FSgy03VhHAGcc/g/I8dPUI5SIQiFtpxaPdO
YjDxRgfCBjWpLcyyB8DNc+BL4BUr625rB1nWvsTeeJ+TiQ6eaauXzw4z93rNP+R7
MfRVjcGvgWjDAuU4CDPgoORPJa62NXw/soaivwdoQlmdYU5t44uWb2Jo7Yj93R9f
hBnIVIqeubZd1atqeaLX3omhLxKQmnCHA2t5FvXzGgm66TRLpr3VZRXJK7bn8dpa
44sRisw+ZgJUSHEQqjqVQYJylcyg1Z7NNX6L6rD3rsxr9dE5k6d7Vfaf8/cW/pLN
Q8sT+qPCGkm5MDaXc9+BdWC/8AMoVbDRptNx1sMcVmkOevnQiazLPlvKWMWZg7bQ
ukGzZV1WnRAD5q7c0ztwxNxKPVl8uCZ9llUbyY1GVNXNuGmc7RIQFhPXvm1GXFax
7EWO7FXcDOVJIIFmNonsfS1PMSAgtTQoLKcB30dd8kgpP/cO3ABMx+ryUrjn3cht
uah892b2IgJDtekfw/w+5tzdK7542Y76HKp8r93FFE18TA4U4+Em8ib9KK7o+E1Q
oyAPW7nRNm3dbDL7rsUE8fuR0shFBhoSjn5+8esPlRebvLdcRHaPFv4j/TTqMz72
HJZTriLEib2qvdKdDQC1zcQxSBkfZsLzsw9fBwGkHKiMK99RljdhANoih7S3qGOI
sgc6BIcakFQZbmDcW7LVMddeRR5N88sl3enMHEvxPoJlY6SVYOPfTrjEIA5FnJpU
qlYy5zkcQbjYTlTrj7pIbyMs4DfvBqyqhVlUWd8yH6UgiOSe1KMiWGAjnI6JPOUA
1Xr2wzyKcMu/y1VIWAdNR7DRxN4wOky1DhkDti0OEoWHG+6J1MQQgv9fN++FVufZ
/poEhk3y29O/Nn3sLEl8nhBN4/sHYieRCpAKMycJbLFVd+g6XDpFZsGVvpVsz6ry
kHJuqkM70ABUdND7O3o73AAu0agu5nu9tY45q0ouC/iJdSg9d10rFre9XZRXV9Se
IIp2MR20WPPvuIcknL3AlNFdmBP6L9nu/i3/xqngJk0bd3O8/SMN4z8UjOgEp2Fs
dy8XxB2RCGRmtJGKTEYK0oq8lquUYjHmi/rhgr/N7Z6ul26rFtr0NJD2tq/X0ykp
eOkkK4BIil/YGDfct3Gp6ku4J0Wm4oRaUR4svA7kyIzZ7vuTPMp1+83nzFkPTvIa
6bTDNDVbw4geDmGAdtbjXga+y32yFS49ik4HRscyp8UYWmwtNO4FHp+OF7oDxRs/
oSxewhiFL/pQ/l4XLgE0cMQDs9YjHmFFc+HrllZO9Ue9GVxLRY/AeNxWDt6JFB3Q
oIs3sP3jP1f0UUrjbF/2m6EQUReHSnsMo1P7a+PiilGm4fR+2eVUYwR0lCicf0yQ
g2KQy14raAcmaEqNYjFP8R8InvrcTWb+bAl/NVqP6D85BF4ndjh6Ox4boh5Nxnyo
M3XiJAFcmzwJ7kI4SYqb4EkCmVoUB3/4uoferaqdy4glIbPNkbaiL7M24cQDaggL
t0k8XtIzQOmc7380LGlyqzV88CrgWqrxfCKs0CEdwmzNmB3RJuORojI0w8p2Z2m0
UoysXbjdu+eZuLM1p1pBIFgz6xW+pTZaPprYR3UcgtOTiPbB9AL1K1D6tWrKBqu3
oUq3RvKbOPB/gBIf9HhLS7yAuvjHyNsjBm/+ks4kPZlcKBGumx52wrTkpYHPjbw0
ZpRqivWC3gjItI5TyhJmiZbiDrmuu+31G0in3DGSYroPbrLsssrgGSdQadcBDE/Z
BdaoTt59TdvAsueZIP5vbhjz8YS7SIYGyCCJI0CEbiZnahvx9npPvl2cqTIs3xBc
AzpjiiYJ3tKiiydImXTEKjEPvBo8FhLoCGchXtrla1Fa9/7Z0bhHDslD3XaYQWrH
2v+UEIQeRNrWYvebwB3Oa9nePAHRHIkmyJwM9ZbdTzUSnuqfZO+vQe1DaJLqQnFe
Xd+ixFMrey4ZBVXmPkOLBicXxTsrjM3V/j4h78RWHqHpbcStOaPZCDILuqy4RCNx
pvLbeET2WTM0HoGTQjJ7jwlaYmm08RXq5aAs5/0zUn2jQVMveVkbhX4jHDPf0HP5
SPiGZ4BDFp+bo85jya0AURF9060sWXde+f2zW6P5JPgG4lZFTmruz6WmTD3hWwIb
cTVjTHt7zMejWJFZujZI8fkN6eBGhUmRZaY0Ln6Nz12sBslhu2pTK6EgT+Ho5uAD
7IR7ug2nVTzbrnTBb0TMUlBWfrzaUKDp6vTaP9jo2IXtfEiFHDria+GOzEz7ZSKC
S3bJGcr+FwZ4Z9LkDNDwt0zd4T835yGJbhDTe55L0DyJ0KFPMLo6hnSrT8KzzVv8
Hdk4idozE0L+iIj4mbCSkz1JjSSlCKcWLyoCSPlc2b9tY+gfrVaZzrpuqM0Q+ejr
3pucZWsmy7OC4Xa6a0obFjNmQQgXPVxJQAIGFYDiLmG1WUm7gwQ9pZTf+vwX5hBA
glVvaJyZ+FJEV1iqgIWHnWO5BUeXPLA3Drsv6+odTlzEb0F2ipxKa9BxWl2XVq0y
VgnyQ6pYx2GrvuxwvFCedyLPJmmPek4gFfuyve9BUZU7J3tBHGZ5SViz2y07wTdK
muEj8Fk7cZ/SS03G9R42NQ6+7R7L1PB/iHRiw+zwW6JxCiP41Z5GA+OKoNc0uqg+
gEUCI0fBvJ6/nY0chkeQYQFIuIzhA/C5cn5aCUxQdtmyO8bHq2BkVasDQNMw/naO
V+BbIanrkYk5YXE+dT+HK6ZOlinxRAxwDPib0phyCPfFEmcp2ys5DgSSd0jtIoeZ
C06A1p4rxxR9Sfk/xSTLjgGxF3ECF4+NhAA9mTWYSM42WFtmR7Y/qj0VxLIJbhHB
3k/6K8Pb3OJ7WqSkeVPDhrjWoNY1W3XTKTM+liEfiY3b10sJOUCRGDRGuoFdCkVP
AVX3H2GosmIvSKP/zOm6DlVuMLIxU589Hiqxsh8TQvgwQ9zgY7enafpf64LkEFDG
YsB+lB4k+L+y+a86tf45bVRVpueVe8KlJm8X0AFQ1kRcYtyeCJ2yU2GEeDbkww5K
DB94jizNBZO7WA8i3zmpULRt5hGYW0/+HWXyJx4RvgXidOltPZMoHqidHjVOA+BW
/F6+Yc39eCSE3b1y79lKNWL0q9F1U7q75v3YGXx66anY3/NjMtZZ+OJxRPSSCDhy
O2kYa82TRNO1uqO4wzNcS68W0JTPf5PHWE2fICg+Ooofbg3rVjNrpEXmDXa4exF7
4KYq4zy2VrO4LmV1WC+bsQnSij8bq94coKebeqIXtyCDpZRmFl8QA9GwncXqwHYf
7brpXkHojk/ZSjkedEmzI68uIOOTCwDanzSccT0JF1NWgJ0oC/6gLPvzPr1qkGYC
k9GQ3vWuDQl9aa7XDZB/cFAN7NwJys+Rvl1fWoE+zsMZBIgOc5Q7DIaB9JbCYWq+
hs+DRoHsshxhy/XqB0XCv5W9W+XdUoH8+P7LB90O6P7vHL66r/26ZN+RMXHUKpTC
HSpNVv9GkmQ7OOcVCofEYkbjxjmnEVwea/op6d5XbheWJZpHABWrPTXCb3jvHYfh
2fA36ogD+p1+r/rOSEcHlJgqAfS9JrTOfE/vP1bCYeIC9zSY82hxD65KD1sciemt
1kMVI6EtaRjjEVDBtJbUzoAF7ynVvlw6+pxvQIyX582kTUCRtyXso0tlXASvLj+E
NnvIgsAUg+S9HBEHuOPTQ37LfSxtam7ybkA8dZt02YIAXAhtTfU8KJQx63y/WPeS
Qww78bunONxaoojq6Hj6e4b5UGWJ9jlHcoWfxrogYhfe2wf3ZqMy26ApQPogqzOp
AkNklKJ56uWmmvvkVzXhim731+iWicbBKjbDTD4ksGtg+HcZ/xuqq3qN2CVBKuXh
uYPHUGSMgNih2mvvupETAqOjeFfqGQynOTo8J5nkUodVbzjOx3sTf6QpsNvPUqQU
ehixAeh+pR6ZVI/U9X9o2pEplr6fscQfcMctSOzhD5w0DmP2dVOy9VnFfvBvnUIj
Xt8ZLZrHbAUWt9K0ef74Pp2OvIIMeWwnpRbKShsqoz6i5kpfqTMGCqECqlfmwcQ1
MFJYtRmCXRKq2jWDQFcN+U+9nAUblFQ7KBd7KC/fJq7HiAe2Bm+VrVKsaHlVWvrI
J/lDKVWBWd3LrL67vtZsgWwzFKLDO444a2rocCevRuq29p6HQJRKNjojTjRNxqNg
Oaa9X6ElCM+3y1qa29fPokJYm/p1KYGxqAm3+rEhAL8Y9/JnotDOHaJNDKXIR87I
ruJ0zOu3SBfWhrUvr5yzsDIzLoAo6ISVB6MfMCbMPbjVeBYHyn9EVpO4drWbb6Bv
p2yDlN9+7QXhInHi07kmUMh5RgAGquINjh394O1saywwYzRxKjbE5GryFrB0rA12
Wl0UF4HuzbvB9SB/g5s2XmUVDVIN+RScjHrZLx3p+mDkFl04vi3DcxxiB4j172IJ
uSZRZtv41lhp1wqdfSrVXNRVmF4ubseKeOQHEjnHNepOec2KewmcEwjGwHUJzwwR
xkDdKhDe1i0XzBkCgvDm8oL9pUSU7T/zBnpWS1oAToe4Mx9SOrOsGAXo35t0eS3G
rr9k5IdxPvqnn2nbeLnsFzkCOOFF358ytqdSmXXHfHyU+9RO0cSCMHVfbFC55QZj
9zOTNvkCD5hHq7Mcou1mh5XyCbclaagHL7HLN1LgkaSLHdCoAVtnAyHC2oqX/kGq
cUjAdPpYnVVbBprRHUtL2RFDYwhhOm2qSupliaYbW4U0J6wx5/Lkz3gy33dJb1+M
OVTmF9SXQSrpR9stT9Lr/w34GO48UNTfAuhBDW/jFpzbFMabaV3fCgvNuaZMoFGL
aaA6ErWNv7EanPPK3bn9mdTm+Rf5FVpKN82k84lxO2TtNEI+5xI7+lIzKbcc1M1T
jM9ZKx0i7PAXPiqkeQUKwJdwacCh1/BCq1376fswflC/1E/ege49giJpLESVudeB
ZiRMnyhEKYasvhl835qvAWGPXae3VdEIlLfE8GrIfCQ06B/Twc/Wa/qZS0K6z8l5
G3eadPMe2hccD34Leb0u4lgt5ffYNu8s/gRKTQkTIb0MvmCzNkyFMOe349Gnopoj
nEYKv+kaqycplatTjJ3lHPSqtmoj3aKaGFTEboCYT/E/2PH7lfII08fVmFOu5TDu
axk5q/XxsCq6vf1DquSko8BKUrF6X4qu+yUYAR+QtPTeN2qw+l921qlE5VcG85Fw
BhncDU2R2qEcOYqrKHn2zR8qQcEh5h9WdTcK5dqbH0Lzb3gk7voXzdGvbYqF1Pe6
uqyPfGfcrAXhso9Z4CaJPIW7o2Karnh4bHjqBR/Qj/g/mN/jIiMi60oDl3mN60Ri
wmpLw58CZK52TBmaC4IPtJGDMQtVfUoKBwgkZguLMW5hzpHbnCYy3jJKhUIMKkUo
UDEpbmaYM1rUGKjXJ6GWgR/zebXBtOnirBIt1CkPq6BBSkIxcZTCw85ybG5oui0M
mZxyLAbp+5+fDvf9KczNRZtfonirr+cViZ8JpQUSZdzvqYxk97C+1pUSbL7LZbeo
3fOAvWnQSGY8GRVaK/z5gOXHPL7by0lnMUEip4uw8bein5dL34BcZacsXkdnwFr2
2/XKS/xovq6Wd1ci+a+zmgQB/aM7LgAq+DPMawKUStwHYfIe0t0ymZOdlFVCfq0Y
vQu2EE0sRzM9YKPiGrnyN3xCeFubId3IXpAHCHUZ/DxwSXym0V14cVn9Jwi6STcQ
wogTrbbl21pGHoKzAbS2steS+YssIKbEUVC6Qv+yaLdJk7azPozyPvmys06uQMlR
37G+q1M/otGwIFokJMzPWmXj9PdplEnaNRGnpY6h0U1VR8ZIpZJn90FZYyJvs6rM
7LsWyicTGB8LIxc3XoP+dSyMioSZoSznblqaNi/8BRkF5u8UsE79zIr/T2f4395x
nfy5o5ElGMAWN9a1EFQZ6xJ3Cr8bb70iSCdBpUnVOqOyVTCW79SA/WMMXiYKf7BO
HldZXaqtPZsxPj718QCniptEUa2Q7WVQbdj8vYc1qID3nYKFZke4iISh0iOjTssa
AlVmr2Mx11PYLh9AHoehmbK/xGDsUY8d9vbYVSbnoF4qz5gZJ6QJn3xK6y8jx8GH
wCm4V00/f5M+0hIPdwlvEc9VJHf3Q1kRs09wwAGDF7D6vqVxjCz2CcFbuvaKJO1N
rTFEcUf6YggTTt1HUk5/KSn0fLYxrihiEGvxQTsGNokgEoaStmLK8MydP9KL1nRv
hqpRBo9Nw3KymloSVELonA+qoZ5nhcmSXqvPco+MPsHY/LIWcTVmNR/0K/qywVCA
2xoiqBCFiZMd+0XauLXnY0ScPRITI30Au/RfGsbcB+Q+DJ5lKxgIpDqVNbZazUJg
eapQAW3Jis0Npav1Nx0x1aF/VtfZVGe8ikJtgeXCYnqX6rdAMB/OUDd1et7GFNbu
8HdUsUptKzqudyUitv6HS4QacPPzhTqSXRpr1W2LQsZ1yMqHjt+VN8P2pCnAdUYa
9zhn7vQw/oj/hI14bEosbfCf9eZ0s9f73lCL/0hDK/h64/eM4gskOVsHBc3mX7yu
dv59M30wmBio5mO1UjK0gV4xtEa6NID4i1/p9PjGrMmMDiwTWTR+kjzrZxUTSn7e
GA1HLRj6bE4OBRiaHr+Qb7S7/riIR6GPsRCEIYO7mR825IV6g/YKT/dEUWayyL4x
WmstGoaarMpCrnoberslUsShqU9LyIk03j5pB8JzpNfQOUwIX3NLRLj7Lv7rzmj/
+eAVYnowdsgZriUKr+NlFRVsFSIsj9fi8vzIj0VJdbGw5K+Gl7v+SNSUFR95m4Lm
xgjtLGL4EKKeO1w2j+jBaE4nFZ7xjE3W8bYZ/lnI6lbQRSLSrIYBNOIChE6tFViD
xpQoGUgR/c1f2MNdqx7djapLRL37IJmQeGZybgDIvAtL0XLMgzpRP+sL8IMc9p3i
0T1XWdXfrN828BP52EgnMWOvi5+D2OwOhyXn82Pq/SfgFGU0dPA5k/EoZ84Ihml5
wVvNf1ChDCMmj4dy+Q/n/77ZSHaomLb4IX/KtT1v++3/3IANBBAer6zBDSwL2bGA
e2aF9G1uV+1Lb6aEnT0ew3cNhcExo7VBfrGNGaYww7nfMHNnUW3McUbcU3Hz1uU2
/ycB43C4KPZbyksIh6gyFBCiUkET+Xg26dRZ850vhG8bjnPKnv1DFRgV1HLOETea
8wUbVT1R41sygjjhs8UYMwyRw2YpUoUyqFF8CQZupvpxJtkNl2gp1Nrscj3tJLQs
RJRZniRgWBJDU6nt0iROmEQ9zVQYzt8F5hSuZESAKr24okOHm/5j2xh4ee1SWyME
mtj1eKIjPWJsb4jH1Kkez9+B2nK5NEa24A0FCoS2EOWEqLgItRvDWWSDOQL9CVV5
F+RgWhb6FyT1BlauNy3i4bQIYNXl7NdVP2PtXLxOOIiyXLt7/qdYnRRs0EiSZmBZ
GU5RvlEVGqJjX9wlD5BCUoKAfx6wUBCFv22BYR2FDiH2euV1uGdLgo+5grXj4SgG
VzzJ/90k/4mzBXLwA7qKiuTJpnBZe1rGDz//1LkHS50UzOCUzRwipiP9muMolBkq
h+EDQ+3X5FgyGLqwR55SduwffXYlNiQpA5u6D6xeXreaEccuBcK5SAZQx7xzerpd
T0ZTiglggwUiW9C19yAMHuI3pIrM4X2gW9tmKQtQ6QZKFFdh540rWVkLR1lOGTHT
KmXCgNVgHMnX2udGlOl46mJtJCuYUvJEs2IlyHod3sp1i724MlYuw/Pl/i3uLVMS
JKlDv5wRPzZ6qAKewLQF+NF6H0kV0f+u/olAtIEGu+TEKay9PZuV4xZIGPvjVRXh
`pragma protect end_protected
