// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JZw4wiDbTYu6yzykGgP9tmsaZ5vA516c6VBhoxWA2WHZMzzs4pgmS9w3OHgMPQde
L63wQE8Szt99c7fWxqTiyGrrt5WTPenRUT9s0IEMCaneq4HDNCFm8HrL+xo0PoLt
CFus8knC2wr1t6ltMjC3RZlc/tvv1wKJWKg5hsqL7K0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 91392)
B+7Ju93e648AH6eBrPDOzpmdgAvPLQffbcJ72lmcApywCRnuFx2mW7wTly77wpeq
XCQagoeNfOyWD8/qhhm18lXv0pVbFEqYC2gASgtCCoZw0Ra4WmCtSXiN0ORPKrVL
c/OvXBPMfNE/lDFmZwpY0V2iAvEYl3x+WxQpRg0IYoQpE4yJC4YpqBuktTWEL6Hc
KtBzNRRnH9iP0dapM45HWS3wJnakqU2RtxKspqIc7MZIF3yeUw3bkEhZwz2vAF9h
LTr66d+yC3jl/lLIdwfj1MABgocj7UW8ElP+CvhF4HfP7k2/30IBt3cpzjRj1Osk
rTBpD6aEP7hMqwDt9bj5HeTD+fHw+CpjrkyI0oYXlhXU5ximvXVJ+oHdeqlS3SgP
eKcuZ7lGk3Up1WD8zU+yUfXeMrzIGpHPI352ZhEPMG14k+5ASUsxFHXvvUajLOXz
jDRPJkaxwx8DSTyYww3SQ+IK7mbqC1laxYPu+vG7glvnW1USgBrJ9fRrZIqz8kU0
F33+QloJlbBF0nRSQi3YBtGZgxYhnJhQcy5NIgaIVHAR3f+fS7/hZjA9ec+M3Kbu
ZuXEAGBSb1RZnRyUJNqTQNvZncXD/DUNGL+3XiVg3L7IXNITUjfjNhb91Y/tYFHJ
EageFooRMW9/dKdLJOktpjPjjon5013mz/Dh8v0FKuqufeyc4o6mgnQgFgPeRb/i
uJUo9n9gXtTqHBPd5UCffaK0ys7cxn8K7Oz5AfZ90a2klD4jD4Tda9xp+hZzfWGB
IcsUL+2Nnj27+rowGnsmVrLLliWZ4CDXUDC5lN3c628g/wM9ahmblRQFpi8ZRWsH
omlP04mvY/zTqY93u5Amkdugus8BgbHKubbGe2j0930C4PJjy2UQxoURuFisHQlT
hFIxQH1Mrrgl+iau17MlzJM8uatrRWNqDii8ZcVCCNxK/6yinLCjzahupfBD2wqC
Pn/mWzDNt9fPnKjQ8mIr6vewWdzYIYxVUxXlS7ZU+NHOKVO4TYvZDZ7Gf/ShiVyc
WhjbPvZntVBc0crnjql2D9j0Dzzh6Gp95KGEtUf5XPd8/AYrW9Wf43f45Rzo2gfQ
8ZR3Z0qKNxtX/0LDuHziGRfzQwR9M+p8BbyTrmkKbB0cXBS+8IF/rMm7naGobV5P
O7kBhkBbXuJadAFOWbIrOmGOtQnfh6dAkfkTx45fZuEE2MH6b1f2ddjgS9CRbFD0
owM3cEbTRd9f/ZSIEdTCl/LVlsGWjVEzzToQkRiM6FaDua/5bSi1zMyb45iMZy9C
2kxoW8mDh3omm7sElKK5oXiz4oZSHL0Q+OsAqACCY7dhS76uLyxvP/ogfi8MnlRr
7EhnmusmqgjLkz6IX2L8FMJAHjwQzPIsQ5Lhd4LlXkrogYBpPgTRVOsQMcQ6Oqfk
3Ye/2YqZOyYiijHb7Gt4WuP1izTQ9kd7r923kqNTRB5bwDO35JawaMorjzh185Hs
jbGMDE+l7HtRzIvyLEoRpE33LA/S8aodxNGVFKKfJx+ygJroGf3ToWW0ytHkzPVu
3HmQbvJM2tG6uCva3QYsl5lK0uPLnSz7bp9ZUc+VO7Y927zYmXgS/DiJHJYfyIYs
UrU61deD3KmPxQKGuvj0rR9mb1oI4kcmqU+3Sek4jaNWvRyMRjUL/wXVEZ2SMX9I
GROFyg8ASjNlRXrkjCy6STjEHxFEyTS+URitgeagTPVHyKfb0C3k7kmI4/R6ZLA2
bxZBoN54mKxh+cuDriKA+acTXQo7w+s6YCSTeQDgEkKWjZXEGbWDjU1l5oqM8HBb
MLloLEb9Q/T1Wx243ROO1JMfJl+tofRiqECe8bfw7Wb9lGtNuJLScmL6CcxihbnD
67LYk8JpFjnvt62fQdK/uXcG5IMHDzSo9Sbh9et5t+pBkJTnxLqAKpdnizVJ0GId
09bFey9OH4Skf5pDyBvHUsb0vXlxpkFO6a9n6ES/BZXoDNXh4oGCpqcTu5NUVQi3
WO3F1oX6l/yjPsFUqyFsw1nD8FUXzMASQlmR0gSMaqBOg7AmZHIyal/F4Ie39YCN
Y9YQIgIAhK+Xhh1E293q/xZGZNjw4Jv08Vt+0yHHKYzD2nRC9yaCo/xFY9oIkt0f
xMnorZjHCoYSwliJZfdUIYH4QUU064LS7SLkCifoBryxQnFwpkOhHWAsIJnYDCwU
79yBFJtu4gb1fCy25tj5dJG71ISgoav50CglLY9HnTXFp4xpPev+Zte7kkRBIhiH
ujz/abTocFYeNvChGBEx7xCogJnKBbyrnDq4/Sv/npiEiRfZLyTEpIR8H8ZhBIr5
8OhAtVj1hSGBp0aLUyDPYrz2JFRUJC4RrWh82GRGn/he9WMZrnQ/xpSUUzQ/l3Kd
ZOZVedmQebazdABMkmGD4cyIzUIrXb9Kt7nHH6tpBrhETZfvolD4OyFFvCLX9ZFF
P3c85TgmpxwfYHf+0RU2V2rLW+k+GKTbxfSS6Zdzd9aQIa2/M9z5Q9YHvFM5KOMB
VsPaV2Whf/iKHubbkPUzbtHlon2TMvSA4Wr7kWQ1JteZRFVq2JVCWeUD5eDQ/UJ0
WtswManFG+XKiDZIQzOfWH2F/mWUePtPCopq9XnY3C/Og8XPV9cBb8sNMgxHeyQT
KGB2q3v67Kps8OpNoWwtmcGjNG9AHVThX4g3luDHE1UzqqtolJsxfVLd9Aif8FEg
duixYOsOMUOho+0Nq1Sw81XNdWW3J0xDfsyJMXRdmq5qR4mokEPL/4UdGBhwQ7IU
C8IHtTRQE+Ojne+PNPIApkMb2owQaMLJBkhznQMYhBNGEDYX6+tGnFUTYgp3UsIc
DwsxPdgVS8aSgFh/AKTce/DjWJTgsTabOEZ7wFc01IaOR7eAqnhlz1I5GkJqmg43
1YlFcS2sTDbLnwKb4rFJLlymTxeWPbTbJ8p4yqg9s/xJHaqL20G5SPEavEKqc5rj
XIABxXbMlCsY4zjxVOoUTTSfi4scELdBcDUrAdRe/V6du6/b6YIERDiP9NztPQIG
UqqR4fvoKEsDYWr4txWJ4lD9l30xlLmTLW7gXtaavDtdoAU+pcLEjWhc7UqMjBdW
7e0QIYBgZBEilXGP63iqV7GH8/kVlrKAn7PSxx7X4ZWjUDGSJ15NwzYwq+RDoHEI
7/EM4Yt2BxWK2oqII3n1LGC+gpCncabfythpaBwqEmz6o7NJ4nc9DOp3CkKawd+j
FL6OkvWc6+7bzcoB5yE5VScFmJoKOwzb7DqXOF6JPeJR5pOfYCZSHNgYfVJ/mNKw
Yo6wluFyot/mx4+jfi2HSwJYhocAwGLp4ouAvW9JvptM2q9H9KWK87XdwNcXXbLm
XHqbf8twp2X9QxPoKMHiH9nYRHY5Cf4/SEjTS49t+oFb7oeo+ndQESFHN95KA9qY
OqOj3oCrwtmAwklweBW8A8tDl93ORiQpD8/mK+4V2ocn73WiE0rKFpKnDmD72jI4
p+1cq96SxAakzhj2KBU+1Jr1fLrAHdMcOphFkwVK9gLO+RlWnVzrmwQ9/9ny/XLI
kAOb6PBpEg0OeK9RnzCiMZx7JJaCUfSTc4XgIgHTdqjb08TkAl81g6NU4KFK6WDO
g8nUYso+Pc9ramGF8ayyICURLvbqCgMgxrGbzioeB5NwARK28iEikhEtQPqLZn3e
zf1jw6AKArzAGtBiQIoshvDLqf15vvTbeP7nnoxAJlQdyMwkbJBR9ei9Fcr3rsET
oFV6DZ8Fuc5TNSn7Fq9i4OJhiGut/mozA3MSXSmcff9HIJep9jAmWwP+rhqJKasS
TvR5DNBPmlnohyTqA0Fta1dYM/2MFSEerYUENovl2YyIICA9SnxtEbksGr1BRy0i
/dsk/9gyXg6V70vdnQfRUvigfz5G1DdLe+sOjQGiPEZJFBWx7m4QpplRhM20Y3bD
gnqb73zu08PtnLNofwjYIxrklfl92YJf2GydkL+yaE29A1J/z7FzZV44D8Xjz9xY
P5tsCPUw/Yc+V0r6Wbm3F2n9FW6T2eIK0GbR1VceAC/WsVPBAdf+Zr6xzLw9LYjS
ngbeGrw+LpSQab2KXdExo15JRECGr+1G/XlioQ6VUDtZ/GmW7NBSaAXqSSvnb/my
qiVy+x9Nct4H5xd49jqaXubTagbse/h2F4CkeIAm0W0fCeKkRZJvMl5MEf9WMnBC
mNhQudt+soKkb6cXTHKq4j+Sy2HJTWegsxQ1//T5wymoUT60QOYut7t3VQvyCmqe
Uczzr8mZQBkhxvL944Zqp0tcR713HzNlspbaLpJq1gWvLZlquHySQgIOgomYAzHr
orXYrqLQcUl5tXBjMRjLOCIhxCfDTF7LMHBdFJBvBQbe01dOsSNo623KrogFU/5u
FPtMDrHrfh5xxvK8rh+Q7gvJoq/H2URPktBwDpG1ZpR+Y3eMGweMxfzlFXUwSopR
NDv39/EKTCG8KEEwlD10sZetVJXx2/QGelHiBQCAvmL/DY9eyzfoYgjjbGiKX50z
yVFdg9p821Ipe3SivvCF63a4PGJHXECeY2i4euK4MtR1vaSjnu8m/OoDC0FQ7tC5
gEVAEkH1+/U0VTwbVcRAxbzKAnPGW7Y0eLIRm0KpArEmKd62hL4yRIo1rePAZE90
BJ8HncpdLh/FaGKYrsR1CY9qa9PjgZMsXLI389Ng5OaVycWUk5+WyoDlMGUioh/S
qHI1md4DMlyJoBruwnSbc3zSdDVEO2frNcOOqqHezvlU+eHfOnQ9ralueyscMKxm
0v1aER9Oavl6MrSG5nJpXcK+zVor9ylwNSBxdzCwyRAACy8l1fDGddxgfLMKW/0P
dstbBrnj45i2tTahUfEoZ9+KMY8w3M/d+iK2WpFWMupAwLKKssp/EpYNRHkoS7lq
TetK/529J6gCydZ1ZekU9EB5Y0vfK1qfF4nrhABlaUF3wLTC1B2bKp8a0EN72ek5
Bdn/PMbtmlKw2wqxadcszPAelNlpT+U08JpSYOvuN9DWXIrexELdQkOIHtqrGejj
bawekynQ87T4sXrxRWWpbXm8FlLtiEkAzgRKck4aoQRImWjJvcDC8UzOYaT0AmFI
3m1q1F94BVzVbO6j0ZYo0ufcGKe9L2tBPrQ1VYhnGOwO934T0yC+gq9rnB+4xRG1
L8cmBCedO9k0kwevuQ6dFnnRANyvxn4x+Jp8tG8nENX97l9jDeihYYQqzwsEfOIS
JA4u1UDF0i/c0KhweaY3grfNYoh6W9aZFC5FF76TZibT4senLPIJDp4sBgy9xVa+
SX+FL8P0LEj3FBxweRA2iuX7Iz69A4mZgZNvawiBWjix+/+BlkCThuZiH4Nd660s
NbivMKayR0arwe/RGi545fQ1eReFjHyCaJt7d6ERkyzngFTwci89o/xIaU97ce4s
l0WScc6esa283KbOx84xBVHQGkRJYGFqX1Q7eYP/V/FDeJ7wBdVTS/AiJCdNdRT3
ysVoFDDRQ96nOYCNH24/e7xCxxxD7IckhEU/ZbQov/BDnFLPZU9jIZDo+mhMTneS
+cMM0s7nVwBiHsQFV51Ob7WTFOfplH8uHFR2Fir6OUnqxwFWF3e3AhdtCgKXRor3
pprRhgfZZCSS/fFAI6fw1V7vdosp7BEo0+cZOIXNOcqxTf/KxpTNdWq5xAVL43or
iPogPuRHIKgM13Bp6xeYyQOUc+xVWNVlokkFXSEwKB0XYYfUMxONbV0FXripewKX
JiohtIaawRWlKNmoXzxfoxVbqAQ0+c3xYoiMU9cy1OieLnDn34IRpTpoJMONdgp6
1hfkvlEIJ8KIfbxKRhF+YZx73QKR5HzGhDbzll+kdHKRyiG5+nS5R8u3X8AZ4/C4
Vp/elOKUmjGhiYpJ95+pBupwMmquNYvUnSBwJF860jevXDYDe7DANM6wvrda35VJ
qw6GYBz/8TWKn3H2xTwva57AIx3Gg8HTDOg1Buq95caZx4A2y5KgIkFB2bqSN92j
al4nb0IKoWbaYQ9C8y4vWdHoLVrvjqvZhcZ74XV2WN1Rq09uney4FSLh2+0MClP1
x+NPK2TkuwsxrhGfo1+Q4D052oEuDr1Kv741w/RJiNR0XLz5XCKJ2aFh3lB37WZV
6NjT4lcRYfZMZ98dhYrp9x0asWfW5SlW58GdlHeAUpZDKt7x5d8pwcYEpDhnF03P
slaZw3RaLvbXCtya6wDTul2VFFY0XLFosl2ysb4BLOaQhNWwozLHCHnVLWnMGjGR
0N6s98K2gWcp2vCVxA3COuXNg6L8bIHgX5v6di4+hgSlCQqTJ1fD45E5yxuPpYQH
LuuTzTGlcEXYdcLf70XH+9vzbV5u+e/RnwZf/wscr6YFKj72Gtkj0Na8oKvGyeg1
b2glk4R5nFjQwqHSRr1Eu4qZCWhYNX87ViwyQJgXR6GOttxA5KPugcoKNFzlNjv+
cyqG3Hjlq3htborDlV/mO79N0X4IA0tAk2tSt5BmWsIwXVvwG5J040K+5pC0iFqs
w0HvDmYLrYPfUtQ6wA2mrJKcF4mw+Sdi+4pv7wG6ehfLOx+F3y3sOhRl7RLanfVV
iSybpmpuI3iPH7da/pPNUFPWjF4xAIWfDyM9o5nFgyf1cehcUwS1UueLllqprUwD
/OQuAnMgZkyr5OFv77lb++3H2VgulSZLovObOG6xouHZFrXr+c5Mo6VGo6MWbZ3F
ijdT1kJfz7ohwRNb49VKNzYaFDM6uFelkIUtIO8JEbq1CDvI758mSgY/vIIHO5qf
VteOyDIZEJ03rlcBnjvqQme5gmlvbrEn6h9d9/WCQoXBMuv9U6gnzLKULWdnDk9x
NkVWLvpuShUbvEyHNG6Bjewqqwh+pZBAN3v9QhOXntpl0MdC5pttLANn4/r+hZOy
taK3+Y/OfFa0UZochUm9GaJD1BsU+gX6vu12bHPkB+57RHTV0CwmwgWfauRLk9ic
dLRIKjmMsrES8LzAcA+Vb11Akd6G87IDjHZfjwXeKxMpZhuWbfYFEHHlaczX4swS
F8PLe45UWD0M5VIjpUducPwRXUtBuz/5SkKP0TDCR4oFNNX8oENgNDFoGK3PBHmk
/WMPB0oOBzn8+Dr/TqEbeUf3LSaNDEJyBANVPhtADHowvXUrffiYzDvtOLpUIfCY
IiWMx4G4DhWP3bmiqMOPQXzBY3Fie74Ytxy+jg+1+f2RzGOe6psvpn9nGjSX+NaT
6aOqSrZx7JNi+ZQdO9aRPRyXQzkT5doLlG8X6qzYqODDyKS6ZFlVcRtAPwmbhXpt
wL3lZ88ekx11KIln71XZosUpGh3sWd8BICmNoTKLD8L0hgpYFWuhCD4gsZprX0MC
f2XAZjVj1soRctBqEXNLRMX8sN57q0IbxnOValH+BVXDnyrV+n4H5zr38eBSJcsp
R6bMPnoUVKwYhwmY4f3Uh/3GaxrRRVSxbcweYxLQhZJ0UaBM06HHWeXqFaAPlWhA
/UcPHEQWgXR+BnjNyNtIBAOrXAgb4D6ejh9F0/wctC/PD5YUY+Rid0+oJwW98W9f
91D3Vtu7LFxmOxdvUrhfT1glLiTgh5azTAw0Y/4SLHo+I8Ufudinb+0xe1pAA7TJ
XbQ4Hp3jD9Dek6d3S75OrE2HPflGlmEFAPs04prTOeVZvQlrrW682nDucb7p9qVg
xZFFcF5id+OM2G+MBhdNhhPxpB00f+VzPqYW+fW7OIb8IFLHSgPHDL87tNfbzIQt
6fEntmJmELLLupmYYhRtWwdYx0rqW7v9zff5vvkT9B8LT60YOw7MIGF0uVAST1pQ
Crd/eAtsoS5XB1uzIcsgBOewg9NYiqktBVyGczHoRQWFFBC+LgR3TQVHzclpQQVV
VKxbdjjnAFKisA3IS2mrFh3i/mhA9FZW4DrAAzSa43srY/ggUIiZ57vO8RAtQIdK
z4B4mZpTX9eFiXJT59qpHeIsQy9D2sUhzN5+N+8kvU1PX20vIsXxYHNg8rtVuKV+
cenT1zPxiMHqHzhiAWUqqSCIUv6cXTcXAmEsm/IsrBDOQ0fwoZ8LDcU2lL2Ewzg8
3MpoAHfFJ28OaNZcoH/UzLAQAmoUxLOZOkhOFq4LAJRLD6HaeHxWQwOpfBV6daJ/
qWzAiBQOtACnig0Dn31c6uTxLgA4ZFDYmbLKLgvR3Z8mVVTeYF2XQ8zwLyFHZtqI
CRgrQixyeyzXNSrXsqGdrPoa19JYFwtl86EvcXHpm56OI/2/gDO+ZFFECVbuAjtN
OlJ3Se8nZ4ajFNFgIYbNwvoKGQr5ilrtduC4WpbJLsp8rfXtttdfGPel4zNoHSWa
ZvrmTYGQPIO4F383UhaJ0S3WFkBM+sAs86T0iNVm6maag+/SgQc9rD6qRzlXM0UT
EKREEEJIUM4QNkumZ1Ls9D5foz2hsh6fjmaLNhMl6nVCH3ITfXSWa+ToRp2+H1Rq
7FBnYhXJ6GbgDUhO9e5LSIqfYtYmu9Zj21FfNdAuD92nt8c4WYynTolFFuqz36UV
4TFGguWzOdeghk3H/e5bw4qoUmLMwi0KNc6vHzux69uF8ofAps8wHVeruhfrjh3z
YZukc2/oMEXgUrVmB/soPMW8ugdAR9M+oEjKhu5FWZvHqDKIIvNyww3Q4UxhTElM
rAR3jlwQJdg5TSKgiyUpghPwSTxGWuatzrPZYyWX/1zpG49lEmlja/SRwTNxiXCj
3Dz+VSAmn8h+dFDZvLqcvHtnpgMeQiLKe3DlEfUEYMvviehBTq17abz/hOT7HDn9
e59Dga0IHc+df8tUPMkSGoFXGo281vHlMVwnDus6be/jcnM8dlR2pQ9slXcHsO2c
3CFylK39a/jUivhC/apZk7LT3Q5mA2KAYzK60hAZxMT2eAyB+fJiQWI9oGdI50od
X5bEqEWHc0zF/0sFzGi8drboFyL83yUK82qeFSr7vwv2YV1RPPVE6MLYEZUG1Gl1
c5cHPPhVPiM0WVchbF+0owk6ugfSt6rGQg18Ej04XXyGeY4ULuu1ZjvwnPXK9rUM
2lUoETJyMkBjHDTAclBfSmtWl2tLml5uKwg9TtQelb2+I6znKUWGhIlfy0BpwPCN
40oCse8n6mEMclyiEjEjZS1kfRFKzl+pANjS4njSDOiyHfiDb3d0Z62k+INL4e4u
Ho2DViIsqMFxqJjT0Ia6HDRN+sSmd0nQXlI2DBwHjOKqst9ej+IOWc6ivMEoMLEU
38DzHiXsPwGGvgX/Jr6VnVqI/hcQpTMhZ0GR9mk5ecg7dvPRw5c02iAhB4v2lZsU
V+XBMB+FfeEZesuKoDLrv7dPt95Gicix12vwhl+/9Ze65tZhrxscGlXJtDYSCVxn
F/FrBLP/maMkBUGdoGiWwNY5a9+ZApnRzhfKR4+78ANMZPqzO68pc5T1UObeSD0q
Fo80wzD5eczwka3l79beUsnoknWAf2488pHKanZa0VPHRSBR4Crhm5pt7quoEpV9
05WrpRjFrTAiSMXWoh5/c/aWGVgxIBEZZ8uDIeD609cfCVzo2n3nrwaehZMjIYOP
NEvds3raCAOpCRC+SLyafIna26RHK1iifTw9gYAxVwL+MENkRyDxylqjqXGGXWdu
/w4iM8bnc4H8HF0DIJkAAfzcjnSaDJNpmR99uarqJoc2A1JO1b+bodo7PCdM5LQq
DPJvOBjCh/PuiuYjgVqRyW4AkMah20s+Bb0IZl97TcxgOrvi0O3Rgk5vj1PbOkFV
TbOpq7ReeoalgJbgGliU7alw7dNUfrmpRuqLtnWhsKEBIZuJGa04rpr6zY+yqkbM
f0Gn4Tk3u0NPQu6/+LhDty/LNbkH4qf08y1oZ8ZA/GxxQGlu9m4PG908bvxN0hwg
fBPKpU1pUfx3OVXc0GmYSZgN5cmGlD7QlrAzWaaBlwVi4SBc7monQRgD1lS1mikq
M8HdMf4qBNz5r/b14MDKZqnS7nEteLsTQuaAfCGeFbhKUhQWTlSphjpTbyXRznjm
ZayyTVwEkeI3T1q74MClsk6VQgRzDvkXef8vnw5a3sZFAaBQGMt3SA9fINTk9Fcn
vmM/Z9MFVdidhmlXsh11qd/FRdVz4yA++vlf41w+mi4NG4EVZ+oCVlw1vINIJ8Pl
hLW98a2NM9wNZ5zmb7/8CY9w6LuVa4G1kfi0FFlR2L5jhlOHGZn6oTfxp3/c/xvp
lmgGWbum2kcqwlTbfty94RkRS4s6kECuyGmMwzujqIWi4oYCb+JrddYFgnL690Ka
U1ContCXOKoS0KSV21eUcbaVLTLKBuQ4ShQkBybCWlYy9WMbsgxajGF9cKnuAx8L
oQ1wU2nXWIGEYL3/KXFfjaYsK7IrcqIDh1zGjhiELVgRydKVS6pRJTUITXFMFtyz
dUqLVZJ+qd8dLnHnC1yCoD6STirX4SCQMDNUfQJQpm0lzPsaHTeEcygLe+Yonszw
BnpEu/7y734xxH1SJi7bNyAl5+4luuJM91heDN3m0SkT1EQ66QQZ1dsV0lY8jbsl
v5ncnjBFjpGh2EnSPK7y81bOZqRjTM29KoQDgoIZ8vA65kjEroyoIcD3XPV4urS0
mOtD3nuFfFtcLld1VtDpjGo73v3ReRiSa6rH3OPmYJGCF8bU80+tANQADDfOLqrN
Rocy6GJ3pmE/OyMOGwKar/b6ex6Rb+kU/202MfMc3urnGERS1P/BoPrWMSbzxTc6
gSsEwfGVJdpmQr/EnuFAwXI1uvN48FY9wR0OSSpw5AoG/6fcfgrkD4FPOokROsaM
3/85J4M+pbpo/T7cwdbXxhBmcW807khL9FTS7ECIW9AMbRSTAHHuYsgFp9oN78NN
4T8MX3KxsIL1CCZN6/+8oVTLOc1b4bIfb0TNJr7xBSe23dUJ8LQRiiCTVt9RU5Tn
S+sTw5+ZgJgVs/Nc/a2TXwmnOw3PMEx3tGtXRvlvFWoJIqGerSpkFhmAEUfKrdxq
kJhctxWVwqwGVa5b4sYx/iypbVRiuzJ/Vry4PPkHufe7mFY9ttrz+hCXd/giEqgU
7L3dPcgq+aPSKVtrpqsDC0r4Zh3jSb9fF3LWtGnL3UEz/A0nCeJGJDwiY5NcBVmR
AzxgdH/ESUYjCcuzDxgUUqfHX4imWpuhmtIR90KGZ4Z1Z8Ns2Ok8m180LvJu4ObE
60Ca+/7qxuYm1rU5EkwUiwmyu7j4+APZGxATA746GPCDBOZvh9fowTa7jm0CXIe/
BJ17YDVO3RWtBkCfi2TTaRSRs9pPzbfFyU4llvxku6f8hbBIsRJi1A8BEKcIgPjw
M8VqGBeshVkfA/H73ZNGEuwlI87pDGGgUwPPfKfUxzZzWwCvuKi9D4sa34BHghZO
PvtqtEl0HFauiKEUfKZwYM6bEIc6TdacxsSMZqRe+2vgbD5Lci+rZioqIRi9n0WR
USfmYFrvtCrYpJH7juBBelhmC9sKusg/2GMgcM1pvdPRn2EyujZHJea9GQwRbAQN
U8tXpCEX7A6324Cyj2oEHuyKhEA8BuVyD+4w+/nW60+HFzf86LCUSwILmKPk5pVJ
nsANYhxbpq9IZi2zIsQrx0Xke6j1Peuu3+h9wDKWfTLxVjcDBHGtrbW1nJVjOeyC
kgpApeL12W5G+ZRfbC7ef01sI1r4zDiG4X7FO2FESa6vDEvfyoWpLRdQUNewNcEX
XcwoGAUi+d2G3woTklpA2Ou+JUyhVYvx0VYLscrmlE6bw903F4rFFisLSIm66JuG
AeiBjTwvwcdO9BxGpViTaXjrF/afEqi/inIFvX5sabo817svfFdDvUddAaRvyyZF
Q3sDycSwWvM3DlsqJPZXkl4pyeDHWXu1Z4rQO8HsWjvK25pCTxYr5lW0G8qlapc6
jYHUPZdVnOQG1af9RnVI67MuisoOwsto+TVO7tplyY9qmy4iHNHOLds34RrnekIo
F3g9RhjV2ocfIgoL7nIczXSW1I/JVPvq138C/h1cAMTFow4KHTtrnHkRW2OdW2oD
924ox1wA6jaDKad0+/SfaKD/0Ed5Dxh/S4TBEBQOw57JhMgMjR7HlpC2luD2S/2z
A/xuFNZBWF5y0dZ5GI9QBFMbB8s7V47vizqTYWifmF8jsqz6Wt3qZZ6wW/ymcfMk
WJqkXLrBIePVZBdaWZpA4DCpeXIL+u4eVtATiGtPTb0ojU/kW68OdL8Sd9ijlyuW
ytlLlbijDSLgEy+SOcTAOFUS7ftH+SPqb78Duu0aSG9Mt37++blILMvC9fdzcDFg
jENxh/v2mJDEw0T+EdHdbQ6+qK+SMamqEfYb2GDBLcImv58Eh9eIbMuC9uSXfIIl
vM0WUoEFumHdGB0RbCSbUjDE9h8LpiB/kO94U4/wHnLNKqVz9+4UYyvWRfOmIZZW
CUDJnSRaCvUx5hYqSikWfxibZy4Y4Fc20nBGCKluYZ6dIExI4hQFM6bS9IaE69tg
6f2tY5NSbqiwnKSlWkB1XwQwZkRJhu+WfurC6jfrVEsgIkmCGQ0vpWs6JpGb0BIt
24mOJQ2aebeefQZMviys6JDmKyFEhT0waRZNpc2fjFaWEb+E7pSu6ujbzEjIZHeR
0peb2e5tAE1tcqVT7swP6LcUreLKpLoVialJ4JWniSpU7TTao3MYs0xmqNa4lq2L
II4A2CuSDvOzyy2spWxr4BtoG/R7ateV+MHLWyZ8JCmNDo6RQh8Ec+I/ABYsCkyG
7tH2jk7w5Ndk+pcTlxoW0tkFM6qfXJTOPje9NjZQiY6KsG2sasKjMFQCsbwLHEf0
KlqHfUtUpguTpE+/9gJcxD4NqFWHc8+1BqMXRAIGCXc1NoC3jumt6IAiC3FEXeDz
8ovgkHhTAhBTctu8mrwmzbqDSG6MTEYUX2BCA4QBh+DWK50hWcQCbXfstieqPbBU
DnnY2HM5wW3i0lgzwgzlpnp56ekiieO3u15VNJbTY5V2hICJvKV1VVFe5OJhEL7M
241vLWr7dhjUU208CQJ8A4S1hkW6iByqD1D3l6vO/P5f+L+Skhfs2ZgQG+k1OqC7
OIqoSDJY8gy2W4slGUxNsDGlez5MSl71v9IieG+yiuXU7TIOQQ0yhmMdSJYWZKEx
x3GwygyZz4A8ax1GErWpO7HyE22HrK7mQ3PvZhUxrWjhfPQczol/mt3U3wMT4pXB
tFbCONtnIaCfwnQsmtOXpYwQd8SgPGauniPhyJ5lJ9VDCECvSj4tl9KyUPMpL047
3v2+N0/JXLLFM9Mqyi0gxHzNyOKnP81MJvEwIDlOp2yEg8YY80EwGpsd9BspOJ/T
9LqOul4Mv9Xp/kQgpope2LAALlAK2iR1o54gxKfykO+5JYtw05waBnjjz4nz5ZfF
GigyjIdSX554x6OwqlJpkRxbJl3X2GXI4spb/LTH7NTc343a1Mv77FTTvjnYI1im
qkYbdWkmUhmeGCnBoI79OPGM9raw2sS2/QnVaWMSDtNd0+r5Jd+m4dySOTaFftJp
gFrTyEXEEmLo+kqImH/3wFuvYIIgU70vRbXskn8z4sOVfbYCoYFg3kTl3WaicDeH
DIr0TqN3SSy5xd4K1DQbLAAVOekja362V/OgR6BvIDu+s/Iw2oaaWy5JowQmnT+J
qSHLNkHtoOxyKIbuVWhq9XdYYyznbnk1yqLBVTrvhEfIyCBnI7P45/aGBu9ePqiA
x+qTCg6qXGZvKHxvUsHevB7jiGv4qONEiF27MrnUkz7++lcWPfrQkctb8bOHm4L7
CL+N0eHfNCuLSzKepQ+1eoKkn6iDnSzYXO7tLU/ccsPEx2AUZBLIoaCIG1G1bMBM
UBbwvJj6P3RMfkqQeyQQST9m0UOOfFHHZAWDmyA5VkLFaMkZqjR+n+hCHIU2ZSJX
1LMTNn+3baKm/kgmiXZrqTsNGzxx5Pa+Ty6BotqbHW0PG0jv5avHck/ZuFzqOr5A
wTBx97iTd2EfmNwQNknd7ac8RSlB/KoOhhJoG4ROSSG34GpKsRme4a5YkhdbMyRf
sqJLyWoah2rpILirHLCu1J+V8UoebTTMXnxCCTibNwQoXOSLVqO6X1YnLoe8Tj3o
Bl6ytXaELwY05GUWQwTAw66NAjVPL+vbNzQuCyikPVyIzPHtwHq/p4kufpnZqLxt
DGBHwetJ1CWyL2ttLyVlvolidVxjsApm2Gn845J8aXV/x0o3e7sfvN1kWWzTH2hN
5h2DMSK3I/OWysuFkgoREihtQmpGo75dg6QoWckjoB0fGTluXo2uG9gzO9xqOHPU
6rQ/PUkpd/nlgJwlUdR+R4HOcc3DcqfoUYxY5Pc/WJmxyGVwTrXVqThh8sTo9zDn
WX81X1q+KI23qnicYy70enILKwsaoDnh1bscoNHwYtoNFRMSS5hEg/ohsTwxLiWy
9ysQUX9BohdmmTnsX24KZhT7w3Axjb4NNh9o/EQVmzkD8jn7pGdt05NVjiv9BfJ8
1S+cI+Rg5OVqZ0FCgKSdTmeBJgRN7T8hOd6t3Efw7e5vV3tVR5D8k3z07kBaAogj
B3vfMZ4nSKHl76nHcNq4mmEU72qyoKueV6czNgqmrJz0HEAavJ7x5Qx/Fe22J21D
f9yhUP0s+67kdHeP6JMNjallW23NvP1a0tWmB6NULm/GozXN6QawXUBlpFEnTJ9h
/tq4dpe1zW5mUa1uJTlRGm8PqZP3z24EG6tUPyv6CUyv8G5G4qJWLPWa2KkpMO+c
eRKAkgkD8lOVbdS/FukNCPGXqDj4nBP/6OIHujT0CYIpVPPLWyhKWbKHTorx8KCR
rZRSn0jB0kxLRKtPQg/UVHGVWBw+V9+YH5+tgd5anSrqHgLoGfiM4B88kYqWueJp
lHQhn9nswfI9fC2Hz4vxY4rbYKWsLQdn5ox7QZb+YyVLg00SbKeN7qYxzV9BusZS
pD0Ang5Thfdg4nY5JDvPyUIfuhFQNhHv+thUtfLHFt/Zpk2v2nnqY/BTSKLJC2Ck
Wuir5ktzT981CjX8lY1PwjUiankJBfJmyRbr+KsYJgrunTQV9a8gWKwRvXpVM8WJ
3wkRjPCJP9/8lc4m6YyyOb+i0s/6AlnE/JvfHSpKC9W5IRkOJaGBBw7euncmrs/r
Zre4eh+6a/0KFD5AJyDBl9al+Rbvc/zkq3mGiAY/OiyfSG0z9UBo+gAP2BRmtnAO
aJRHCSLf5sGPmRJyv0LzBBeXtNGjXV5rJpFOVl37x5pBF/wZzmcUHy3nRJpGZC/Y
9cGBOy3gsyoWdAEbX9iHM6DRfWWj/+iXiKGunf1c8Xdr/hAgtaf3yzpCbR7Y2d4W
jGJ4s4548xw3vBMDleiY8hfXA+pnzDoqiMs9IdGcI9bembyOnXUoBbf6IGbI+apR
tzdXDR/kFiwsxDrzTHdSFX+aGoqRtUqYZ+oe3L1LdMsKmG/uVQDi5rQ7/qxSvcTg
SLuvanoEuRo1hK759UQOuQjQNCCAmVcL9fgWT2h9YxDXbtxgx635wDwhPi71FdZT
VphOP8DEeloMBAAusiOybgmSj/nOtfWmhkZl1alxFxjrLv16OEOdBGEzVnE+/gLF
kdzoXTUegqQUbCw/rjHUm8e8zC/29UbjORlR1Gf+dQGH1y8mQ39UL2gYSTutoKmv
yr+grQeaAzPvEovAe5IpnAOOEqHwSMdZwdQIeVZHS5IA0egpVKNOzg3SKwp7By83
VwoeFpL7kUgbLre/wzdhFiJWgj6VnpFhDSNvbqgg5wcsLtZkbTK7TmrggU+VrKBy
ZjZXvRWh74IHm5pYIClO9Z1QJf+2k7wmbkPGa6gG2KfmsjTsziV92a83Up8hQ1/j
vYbLuun5feQEbstO9vbtIQDhOEHTA/SumGekdTNGcbDgIGhG0XngxoLUpafvFwC4
zQ1NnwfJ5CYZWCCvHqr4ahBFSwXeiH3fhYyaDoVSH/E6jBxO2AjzJZR2MeeA81mj
x8mrDwbX8raSrZi1Ix2ht2u2vHh2JPLtYo3IhRxIh+PLLv+Rt+S1Q6b5OQDtdtHs
i8SA7rMMWW9Bg1k1kf5tRWtbRToMlgDknkV9aBOwT6TbUcQQC5dVso1ODH1n4d1p
U7R9LnLU/xsVnLN04JXnlCwJIcmv7nWWYt4gbjgBRC8fwJd3ummuSgj95HhliEks
AJT/xSSMEsTDuenOpsM/fOxVH0/XEAqhMVyE8bWR//plwX0dEJDEHwjiKYaO8td8
2xn8tOWm0k7yB6n/Z8qCy6BmOFP+BABUPcXaiLJSRHO6PPaVyaM6MYTvzhSb8oUj
S9hOZflujVJTr4DEFWuy6KVy6o/QM0RT2yuVH0G6zJXGgxYfhibdFvtWdHU/zIK6
scZlKMoIW/Wy9FOQxTItMpCafoMjG1OzV7+0WjnhjuZnzXRV6mNsZ1K68COYG4hC
uMY7YmxX6NPA+r6JfUQUvbagbx/g7BYIu9vZG0M8CsVrIF3I/RXS2q/6PUAwaVV3
En2XgiJqQt750+U7tVFEhTYBckxrviQHSP+yNg2nsEVIXDEVDpDCVwzAc3MZ7+My
+Snqe8eTe7gY7XzevTM/Hg7RIVeBHJYZblOSt3u9/Jf6u3hcx+L1axM8YK+uRabf
M0c/RCFbZOa1jhdRByVNPjiyZfYe0zuKorpjRKQTnnprr9vD+Da9nqLUFDoPVM3P
hR+IfTEHr2m4E77pwefQESJgTisPv8J5NuIwADGv29vDIIKR4ZQhYaoyASjFz52e
fxfjNJtt/awTtSFCr0GiROacZEfs9FnuZ6Bi4GTE8dCnYqq2EmRyFw3KIrLHrI6e
CarB5F0k0lYfBRR3QxE/b2J7MegBY4G3Rqm8+L00auQeFIb1jRfQHRyq5HM/Y9TO
3Jj7SMXfixGDNkIMQ8OOjVlux01hbAGNrd77k68gAXZHVCBHy2lwlaC/U7szVswo
1mIIBiX3oLfBP0z2bLT5+iRaUXeAQ8kWNaMXCEqEWAszST3U5jnuE/bPeC9vpM5f
p6K3sxefhj39lqFA4ybtqCFVpSnZRLHVqRmZt8+SYc7ZSJOgTe1nBvcymQtoHo2a
cSoNigZ74cVsbsW+o/UwYVj4KlopuQ6n8I96OTfsV2hG89WvmRROcOyjUpqu/Qzx
r3hSV4vPdTrraGKfJJva6m0L3dLnaRlCoslVxFjBZ6oC9dRoFuc8hvjHcLknWCwh
sQ1fdTdx8C0vwkC9kQrmytMZQtEuNum1XL/PgaOotnelmbKCrC1TzjSb7q8r0eMA
I6iNxJhQbTeRLHP4KVP53M+zmSbE4SRQb11B7VEWsYqbmvgxyId9Y6nUUMUaXfUL
LfZ+qsHD73ya+ppwALP89xAphr713xQxKVQRY6RFLzfSh+wl++9QhDGjbUvl5EZU
l4LhcwcjJiZPIdwU/CxRsfm9ae44Cmhzg+Lz504b5O0RFaRbB+gnGbQw6BE88F6N
joS03xmxDAb3YRl8oI7a5/Ts531K/RCKK4LFDTkanR4W9gecQwAbw7Jkad70s3hI
H4vs3A0gpaGT5Xm9fVQDMMcADpYk5FpMjP+ZbPW0kPVF9cBwNLArWTSkxpLH2UrC
0M0CcQItmT2FI107/Y6ifgZsEFImTjIFOWBONqEwGR3HNZnZI2QClEGPlLiVj5ij
mTILOKNocDZXEcbbOdrJzrhwxQO66LbWzrcOcYFgoy4t7gOBGQzHGmERJZvV10FA
tXOe5y8u6/mwVWsIuGaklRsRcvt8scy8zgtQtzMnJTgU5QItNTkExX6Umln2fa1q
8AtIfYrJrKXCZHNgMiFeCSWqZDSquc+W5gTJn5wDlRWkr3bdAr7PbYs+8t6f0rb8
qTW3DmX1pm3lCiw/3FRCU0rkz0x8mcxXtupiz+r+J2rNW8hUxSSQFtHAU0ZCGjwk
Y7ee3h+xh7N8L5xJimm0vFN7auIMMW+tKL+AgVUZbwYF1Iv5LlDDbRDF1D7JI3S1
N57TX3kuXLwfgdK+kI1P9eMs4730PBMh2b7Fz7TSWlyztZtFiM7o19vwV1fUUINK
9hcHRI4uosBofVJOOcPkOLc05GBEaBgjK1ku5N14j9Xiw91BeNmEJbwes6TjuAuM
AALmbuNu5zjjRO5jCxqvXPMkXKr9cvu5FajmHsE0mKfY5fa+jZnEM7/fe4weO8Kv
y/KIf7q0yOOfCDAi1p+c0YRXl0nnu+0MT9fC0z+TkzrlIESKGhxmB1DlrMMVrlBh
xqjtxKlcYrIlKVY5/IWIZsQ3GQOKi5EJsvJK/LYR5Wj9FgLc2XO10UL7fgfCtwXJ
Z326Ll/5Mnk7V11aY0EkNsq33TV6j7UC9rrxP01nphndmYzkdFjWr5mLfvLm3c0W
yvB9N0U66s11O4W7SX57F1TlihvAt0LBFrirShvo5jBcGqS/TadB0Qsb+vWKnPZ9
7SV5QbImTEZ6FoSgWs3/mwQbzRja40392vbgBPSpGMn8dkEz0xstshUnRCiETKAg
87jdroK6uBp3vTBnOpyuyFh+nIufXqi3JOCHMrbOYq2kTWBaREv9VC0HYM194m8o
arR8s7cQFm3PueA6UB8OiaN8yPU+ILINXCk0lnXbTkULf6gl5OQFayvrmzZagGS0
Vgodi7002uZqk+wjUPT058lGzxrvhANjtCky5nyhqgxVrAC5Zb67fwTpzaky4wSx
enmVRZ8js/RWyZTmbMnFJASZh1eE9nf8Yun5Opay50vklV9upLhv8GHtqAcRfH3k
77ceXUzN7fsbx/Kx77kpuc6rHePPfMlHJmoKTfXjI/2f630uBpNXp4P9Frtgvd8A
kKaFp3QoOgcE0KwU7tL2bbOs4dZU81flYwD2ruJEBJQXvgy2m4psY6ZYqI3162dn
oP2hyJ+XQ6W/L4FRNqWQJBTTT3KWNhIJHaExjqOHWtk9EUo3rbVyqxloy842kZS0
eALzkuc3NgNSnGmb42ggCu21pRkVfw3kTcGpiVtLEIOl/XCowzB+steDkkRbHbaG
rtTezYf+7lPo2bfPSzDhMbN+L6BgzmAaXABFh2pvzfDv4Xvo0xv8QbhyT/O2WKS4
kotdHBn7uANitpdALpzd/ZTyT5JpJJ+aGi+vcByD0s8x6dS5iI1X+CN4nw3ckahM
eyUtC544YPvjuPvz0AtKaI/txjjDuFEapQsUyqe79emNJQTPcBGHJWyWfn9UNo7K
SBOuzGGskKTj4iV3ATV+ofA4geBQzo13TJFzahoghf6sLoNPUnx3nIxOFic02rAf
3C1/HaTBCzsTM9hJV8T2tU0qPzc7c5pIW44mvXM0p5xu0oMYqxPKeV3+L0/acF2d
LorQptWiWBDDQKdwcdQMJBMN79N3tj9BYR1OYlMwzvC5EgnWEW+fD2U24PqIZ7r3
Z/eiUFXe4cUFZ1Q0CejeLcSPg+HpIQHuM+5vEIDsi43qOc/8worPVU8aPZel0U1g
HBmj7XaJDbNW/OVVGuRqp/ETCpCgMuxfY2jbEJr3SfMq+AFMLdpu3mNdzeKoFIHp
ES2NeS9xvXfe0ENcyMoOaV0lqHLzx31YRKeBo7VOtI1Cmbs6Md30SAaJ03ccAPnI
Da51AsE7gnL9ZxW7umE7yFxpsa9ko3oXxN1UIGg658sbuG/b6KWRbLDf5EPY1RiM
rtEptnukvmc0KkbHt7Ss67uWatFzN6GbLlocOXwyqXSMD3jDPPH4SMFz2brUJeD4
B8WcuUU9ktsRPpC6pKKlgO7Oqv/1QAk6hC9GdhiT5Anr1VnZVGbyHfWYjtCHs/TF
Uo/1pA49qlFz/SYLRzSbvVo3ieXwviM+pxlvS6QicoKFuXLZkZAEYnUdPYUeo6pZ
nVoJ9QAAuh433AqY7Pm9IARawCqVZ0825YgmbVQjeeaXEJQDl1ib5dQP2D4248LZ
XW0mcFQYthp7YX7iSujsR6k7uHsLmDUqq4nmmYNYpW0d25I4S6nldQQCYx0qvdqO
ZEm1pV/eKY3OGKr3CeFpd4YkBm+UAE1zhnFDeUt6vYvLNmOdZ+7VmOr39a7lq3v/
vqyIL4NrrfoTFDndrLrmYniLRK4glnc0N5ubQXqc8bpvWFuFjs5jB3jyNmSfT3ZG
tbKI4499CjrMw4pxrAmDp4dIZrx/eamhglYgWt1Ten4pmXZaINQcykEH9qyZJ0f8
kZ8SfM0sv/L6daXkTq5wWqC9w6kND82xTW3oe4r+hurR1rnC78XIDzSvpXFF2Iwy
TKhEWww/zzC81jMT9ly4WWx5MCtwnUxIQgtr9JYlM6TOQVlUq+wUXLCWq/R/PEvx
VqwbcXoiztpRb28grs8wXJkFlUGIKRU8nDRy9u7L24QZX2hYcMThxEUz/+HRA/H9
XvGgGN4Kyg7rP+0+67Dxg+2/hkf2sMJulmO9s8yr37BZC9+gD3tXnEtGa74ax525
FH9R5HWrX0QZDsgLmXLLGZmaZyfy7tyq3bRv7AF3lL5nK63W55Xbo3mA4we/Ok88
kfoPa1+epBJuzpOGFW8kKcAMUvqoQZTUyOGbhas71h05zvuys40i754qR1o7EEeX
M+0C7rM5Alk1u1wGOddI252vMaTmhNZ1B2d9QHls2lH2aCuIZQrknw163isTqrJb
5StH1s18z8ukZOdBCH8jpJZjeHczX8JruMvHVqQ4Sh5UHftcT0sytiuR2jJFHTuY
QcAMVIOAgZQ+/Pb2hOhEZM1WKTeC3HGK5UV4KlkeOWaguUdykFNFLAhtbWd3uI/D
ESC/50vclm7FHaSNZyiomZQPVjG37fROQJc/AadHHF2ln1dy3GnOjEgrJZLc8Nmo
kR8ar+LR72vRzhHFR5lBPvpi8VUvIWD1r3LOiRQgGhAXCUvETQAPxSI7iiF6Hh9l
9IHFpf3Z3dEy94+kltGSinyLzL1Uu58ZAITyK+cyAJV2Jqqwaq/do1lmpyAhUN6c
r4JArjvzxHVLsDHQfI1IAtf4S3Qkk3cA1Nw/1UgF8RRFheqq0c2w8YzSK1iXWW+o
stWrQ9ZooAKzSQqX4hp+4ljcxL44o8DdjP219YiQWavs3XQY0/EZ1zxOuEtOax5t
NIVicIT7xBquyev/ApKPSWQiUUJNPvUzE8ErkplbdgetqrzEJDhAkQFXiRFGDAY9
w/PnVaj0jF+l67++wJwDI1PzXY7vJwxEfgi1FX6PJpD/m2MHpSrD0etGlzz98GVh
YqJkdwiPP798jvQny2KaQ5MDsjJYiHEGJBnkX9TbIdejG8uJp4Liv+doT3arFchU
hWQRqSNRReVzaU0MYG9Soz8yxlpY/PSAqf4x3CUDT+GHAQuxukg4gL+AUiHiXYR/
D4XqEE0Meaw/Vzib8MYajQQOemvLfTqjbadZWYDWFTpAw6AseXCcjumnXNlcIriW
C+/f0M5e1X2QdlfYxlPCTH/83CgfP2Yl+mLtWxAkUqGldmTtRRSpOBSqsZ2Dm/DO
iHwJk7/qwyzxZM6C+Nk95MoHMgqHEWggn1ySQOqY5fNcoW2GJyP4evhR9dARbXb7
2YVnPWk0BAEAwXAjGZtdutDDrYtlCtPzD7oUNXmT5Xyfj9hjtFZgniK/mWk7rzWT
K3rwBEZeMlCFuucgVA2v/DXbAQA+tiM+65WRCtcC2vjqgH4Quz3Huckg59rozR/K
w+xnO1ojTltqmEk8vFyTPYxXZSNj+eO3M5nSf4+itJ8iW4SeJF8EHYQzvQciwfW6
qJ22Wey+JfCQHOfFqA9cZ23oc7MMrz6zV2eK7I+XRd8388IKLD9rO8jAg1p2c6Pf
NUouVxzjI+im9zPtvb1CMZK4FFYV6CdjMppVmbMEgcUsVLLonpSSoWnjTkETrvUE
Bnakr/+MKXl6lIoRMMvw1K1oFG12gTu5kMzNZY18EHeu6UEyDQ8g2nbPPqh/8Cxv
XhSGOx3hZjTXRif7pZpn89Jedmur+IMjlLlqC4SEld3YtWapqMRupqXtm2sfoB3A
5H8igNDBdhq+IjI0RTtQzVu19lu18b6ilQ4UlAGyUU57gV6ym0aGamlvbh+dV8Uh
aXTMULOYVmgMoimlrTWfaSvcZtBpk/MtTCv3NgITj0hdClSVb872gQVxWEWAmyel
JZaxyOZYAWlYq+bBcIu534Ze14f7fnbHqnP3MNsdz9G3xBwC39i17sD8FMdNtMNk
j7lwNkRVqc8d5KAHqbrodOiHOUgZXetaZm+ImA69i39vC94PVwvzmCiwCLQxPhOD
3lHMY7GX6rqSfYY5whX74ZDGBKq9gT8yiA83V9LbbORT43OG79fbCPGdbb9BVsba
M/cia+Jigkvm3urIM5SHSmiKCRjiO07a9eLK8U4hA6DE7Aq+ZJmuIp0hHzSEElwR
14MhdzZi9zMG634bptKRUDOSvRGqvkgX7I8Cg7H+CvnnpGk2rjIfDjdfcO41bu1w
OwPfmsa60bFbPg8ZLVeXTywf1zgHtWKOrgqsjycnaqqHaEgu03lYdaqfFWheBND0
lXeIU1audp4cBkp2BKFT/Q7G0Lx+Pzusmd9TLH8kz96mKDXHdqdMY3LJyszVR8RE
aFmOMLhBdS/F1mbSlwwsvZ2wcBQjzQCaM3Zolo4oMAox9E2xksPI5TpGMWBZkRwO
uHF1SbA5bKl1tgdU2N9PsPmN3VE/uQAVjcjSvAqImNqRgwbnylzfGLtJ4lo5Mhel
OGRVz9PFELEg78JEWZvImjKtUiG8lQMs6YkL8pcVkhv5SV7PPnAZkatLuf9ej6t+
QxjlcJNXx/DcUPNbeLcHk0qd4dmzzT/rmgRvngNXGWNdjV376LljZRwXk9Hr2iQ0
aNdya+DBiYMWcLj+dxQxiGvhhb5WAhtnAfyPdEjkBLLpoy0Ahfbqi59/ajv9SYTY
iHJJaOuCFTagb4XhqQBxen0YVhRhlo0NuMwniOrvCAvyfSkOuwTbTrCr5mqubOk9
1KssbmVEKFOhLTWNJJMfwjb9KHpcyoHxUpxOjXw6kcGpv3AAWxZFtND7rWxu9nvZ
f+3QzycuT86X+VMIymGgIRcqREZ+eXcH7tTsFZAEX7FqkRIj0jlERaULjzzxut5L
hU4Fc6aW8yqhp1FEtHmcSFM4l9o68fML2+kUwCILGFD6h9OaHTCWh3hkvsXUpKSB
69BsoJTB41jUisHVy6vr1RNomz7ni6KzXqsuKwY/yverdEmNrorFN7nDYFGY36u5
7//OJv9WAkTz6huzJoV79ad4dcxUeGtF58g55bs9nWfN3le/ASpWOplm1UanYMny
w3oeeDRBlbF89eR3gaoxnBUEoKBZwvbRVUS5n6neA2uE+5kzv9E8KNf6PrsMb0yE
1clXQ0SyAZklZMMwQFFVXBBA+ZtWkAMm/XQgbnm416aUEOVpZOBW9z4UgTw6+mvG
NmsgEL4hmX90nvQqBJQS1ZbrlHawsDZF5kNq/NJFPjgVcyXCRFl4f70/nEk/6ehl
dgH3z0GatKiSBbKN3MuOkGHODDL3aEN8CZEM7a3MOAMS7GTONfdZVKs93kRjRwJo
2gudMZukG4lvnrEyLuH4nOBhvDe6co3YuL4Uo3jJccNGe1FgTq7ToQn3o3VnmE5l
SDQuW3Fud/1Tc5GbbmcP04OWEm+kAFlgKQpjXqeOK2iXrxoWREvALTSxQ+YOmnex
pFM7rtjnlTxB1r67Bmv+Wadxla4jri1CG1CHk3fejshQRhETuDyM/4BBx0LesOE5
AphQEpYv2EaU5q6Qww2Fg3lBu9e21bTC8cZlFBB7lWYFg81mfAD3vT1Skqby62/L
wFQo+F5epwOqGBZ2e9hxT5jhRSi1tamIOaGwoWlTTtHxtVp1M4VkugPOFy98du/e
GKZCduvKTfHMordaR1q5I6cmZY/VlI4l6ZA1C9zuC12d40c/D8l76dw3MERPi9cr
2HfpjuBJNYePj7pL61ro/dhklu0k1oOyFJQ0arzT5ItGHmRrSkpqMrHRp4D9cXgx
dCdgdfaI6wjrZ8dCGELivueDHMxRIO5CEa3PUnSqAlQSrNnonGoetjzvktmWlgXs
+q8YXNXmmlAKVMOsqqQowkIYMHqLoymiUwi+uTW21XQEylT0fuSWiISkh49ut7KX
7YiO7sRX32o5XaAOMTAtPszQYyzTwysiRlPL9j+xkotHrRZLOKc4mzf1cdyHUFau
7QH98JiwYoPIhJ5pN1omeyXw3qtUMEmcREqFbADSkFMAvyuAl/69bnU2wJrMm4E+
CXo92HfFQAX9YcoMKqPNK7uwQFFE4YqNpPr2h93GQRptOgrgMXtboDMcrwwNBnOf
MZYKiJoYjOHOd5xaD6Ai3kIbVu+pKknw6QKUH2MgOApbWptcTXlIUJW4IfR85oCF
s+C6JXVDrf47WZqrNgLTmafbSVQJga8V24YYfTiYxXpeG2qzCMrk1fIMq4MYikR1
dPGel+90QleZ+XSuoAAQjxg4hTCsjU4DsTRB0sPyL+HEoE72jwzG3bO+moAHQT7S
fFas91HKzXecGmFwQPBvsyp2+RE+LeyMJsF7lsl9LQ8JU1iACsWR4sNRYASXwYYb
2lQy8KVEUdR8izJLAnctGwk5cKjd12O2tWCfSgCD/700iRsfVfFvUpYNgg3ZsWkL
g4cJSBlC266SNpHYEUmCnyiQSa44LFcQ6esvecqZjTU6zX+zyfZDA2tWjYXFqlT3
91IV380K7QgPlk9R4lSpaEe3x0YSMIgvq8vE8JNqxNghzGajBf+X8wG5l/ELG7DR
X6XkBykS/r88BFjMGYHDEoAKefVrQZ61J27tiPFHMn3f9nvxUF7aL9jSw4hqltXD
WJaYPHty83tEuQpzfnvuhB2hkN6GgJqB3iLCYqORLxcfTm3PEAw8s95psnLuBIND
dYxkP9ikiF0/FFo5KDujd2NwrpqOrRxmEl3yyS1QaB6pSPd0B2Vp+omY8lX7D2od
7QNgu7O2y9973yxcSGJHnp1/9YdnH8s9thd/GXK1EPq0kLRcGkNCtKWc9v2aVinH
hiENDV4vpn7hfeFY/UAahtoEe6+vjOBB5I/EspS2D42YEdonqCYZfFsm4lVMpZ4j
FJSHWC+iUo/eMeSK4U4BC6PggxzRUZAKv5y4dkJVQrIVLCIpghuIwR6qYJ2jbCQt
LtqCgcSeViqOHXwXr9E9at80zbj7vfzTnZ9D5exr0wl7x390ciaILumN/gQ42Qtj
JjxUfyMMUzpdJV9BeF9EJpRINSM1BX/3C5z1oihamRN4lph80rNPhKJagfSYVCKe
DHRq3cXgthU88SNNgo0Vx9St9NIb1cH0jXBqTE0VQEAMH0+cXtQuFGN6encnPuKi
/66E4MhS9UJH1uci/HdN97CF0mi3CHCPW/e+rpTzw4gaEkGxj+F17/olpVzJ3QkQ
rSNeVTigf5HKfIxyygYz+nKUPdWCcNCCg/lQ9RlJ4LvkYyh1QN8hR+k6N3bA/F36
iUIrXKxRt8aUXk9WCShzYOpCpiBDfxBh9CPXkb2S3vb22URsWSwJC8JRVYVAZv89
+zvLkiF/g4d29JDvuWmxxz3KTIAa8eh2Y2psxwP0c/XfJ9WPDHJJkwxlP8CIbWM4
ULE0aeGmapScYkhTJfC/ifFQAe5an/W7J68yhS7kGp26cVaG0pjQ4URqRG5dPQo1
8hrokI/zza5o75/83W3W9q7M4pDjdlE5e1mhJ23pqckwaHTG2FO4MaWNDVcndGN1
eX0igShA+e0rok4q0hDM+vSfQ/bMShYrJMIr0R/zjKuJOQdHt6NTJTT2dhltZE6g
7EYQh0zAIp9vuJfmmPAzSL7niJVPhu+QB4/DKgS8epzf0ixc/aMAWChfrD7VLsmC
YusfcIt3jgvh3LOdA9ugLZVAzCDV2Jk/u+SSZ0E/q6ZDVuYzafVKIiPUl+ajdGcX
QKII0t/C0oG5naIhffqP4zv/eeCR2otNdQA5izq5VYsbX+4yNRBUK8D9br6nPUTi
+fPrGKjejWZr+92Q9tbPTEqd7ORgDEb7udPTswwvo3FnZ/yEGZ8alFl45bi232//
vfwr7+NFQOxHb0/9vNn5bSfmrZJyq2PCxg+oA3mLjBlGi5zzpf/QXkMmeXxt/B78
SnVlH6AwoZncyfrqOp9jKBiS4T/g5nqUQzLx+f5rBuu99/Jf0Hp4u0YtTDitTbqX
9ULRuSj2ObNwKTYBQxzZJry3JUaYFAkaKLZL0NdoaCeNjLk4ifr9YDR5z3QSdqkB
KFzxuRYc81vuA7knmH8uqoIDnwrqPaPZMvfydkyNLQppDJdiFHeYLXRs4tk8hFOW
ivnelfdzP+tnEnbKQc+eaMa2Imilfm0OEBtF80uhfj7raai/nr/V4yO9lE78/6eB
yD0719BfW+1TmxkG7Kl81DQ1hMJvCKON/JVo77svhsDc8kf55Hip6UxrMPPLqFT4
zGdwrTMwZ+XKcrGcLwN09LgClJwLgHc04oJCfxFv339wWl4r4ok9tHmyhwU1O/dj
lj9SW8lsPBN45y8jhgOlIBl3GEKMCUntsTn+jz/4LkjY0d1iqE8lovwoenJzN32+
+bjmbtBXtLew9vu3MCrjxku/m3y+dqOjpirCPBmOTQUHpdpoEvP6eB5pBdeEkl2O
ZgCnKKyAKIMGaplL88gAPkdU0aAt+cXFTOWHXsON9xMKBw/2OqjaxVM20aiexnQs
n7+SanLCCwyTTIwSoc7Wk3CetKgYenzUAigdgkIN8eGS9zhRC+/3Uh9wsLgHlqI3
9p58Y/UsevlWnuIAxMyUjhb7RelnpCG7npjEK73+VYR+3VWxsHcdJ5C4jAwS6vE4
S690+gbTVTprCoMbhNUOFgE8rq9ltIR/ux+O+DC73L9YICRgC1AFDa3Z0I1NHoHR
lHBYVKMvStcmh0fh6+1IG6U9KImbsaXTN7/tC7EgLY7ZKrqwKGVW0wJ3D7LWE9xh
m02/yjpNoA/5YIJkrdKe0Jb6pqQ0rJjoWAcjg0oAaey3Cn1hBSaaNpCpmzKOjSSc
yOfPO1LJQmVubz1WeLJ95frcsFrPCJn4QKbKG/8eo35Ro+o+Q1yPmyp71q3WcdiY
d2Bc3q27sCdOxOn+/PasSJVbQ/iILNlr0/Ppj8UK1biOn85daGatLQI/bXVo7k9R
hsPF+oT7fDKFqQUHQFPWIWawMUWIq92/e4quKacZkViAW3gJIgZwTgdR2iW075wt
JPVpA9Gf8VeR7xNm1tdnsCukb2VRVy6n5BkirUHEEz4R87bfsrnZztJpkGmorr9E
0mBJ6Emr4A4Cy1IEqPo2bbcsIrwS60Ey4b31tiDd4mGiJc3sUCsJEyi9tL2F2a+E
Hy/jfxg0ZIn5/bDY0D1i6k1SzWdTPjZotjLo85op/BAoO5OaOJn7DegetaSvBFII
H0ct7MsO0qSP+WjIwr3IXJWicxbEO4E2m+t6qrYKoVPOapIey/K1SHTLYB3ph45D
SRDSzVtRlliLqDemk0RyyDW5b8pUHi5eGlgmEf6BODsNwPg78jxOoto81J/z1w6v
y2UwfnWzhI7ie6yfQRA+WfC5UWbe4s4Zc5SuWzUq9uNDLibOnffQyUXLv/5JabD9
bFUFe51eVvkT5IG8DZtc1ci93zdedFp3Ztkm5CePM6YtzI8RbB5/NF7j2CIzK3Vh
ciwOPQ0E2HeLHaTZ2jjZvyvlU8oUX3aETq/BQPbueeWY0S3ea0tPFhXbWRbgwT/u
8HV9CS9yPJBrbKR4LEIpcI0/GUWu/XIPGsN82rsV1JB20DOQy9ZS9dXV7gI6/euY
DJrCe6SAV0Z64iR1uY4A1jDiUYQJqhzBr/2k75w/kyyYMlO+8xH8QT+V3eukVOIy
QnjdrEkoiFZP5QeYEiTcqBAQWhepHy/pGst2YtgVEw/kAjuTFYCXdd3RHnTHCyEs
+igb4f0NOInZuCENhzlWCH+ZOSpZNYFOWJYZxnTGradn4J5SuwdcXXMc0gFQDGjy
oLigKs7IwXBAxJRSNcugDXojFMDE0RFe63b+9X1Bldu+P0cBcLRESCVxlqgJIy6u
BF99mh8eEwzbSquFHLZk48uCStO3zup7L2j/kGdkcivNrYIoilJEe3USn1ngGUBY
WccofRu/Ypnr7/dMaZOZJwqyipitgsm1oRrA6EfQvDOZwKgNaImVepbg4QZs3vlE
pByXmhidGQOCeJThaFvayLpcjtmP7TpO3PN0hy71HOU8d1I8mxYt9Ng8R3LrAW5f
jHZSqQFiwLM2XMA+9XLUzjV5K4IUzULNkbTw7lcqAnxd0O9WJlN7Ab+3guRttEB7
JdW3Lk9eS3jswp3lvX8tIu4Fjs7epq2dj1giHG/QTetf8nw/shJ9C/8QjM3biX45
l080koYixhdYUOTaVctM/IwFgqW5+4do8gnEP2OSsXmKK2zqQctfqLScjF82nX3j
UNyLLdFppULyRuBMaW64IiLKKkybhwWhvwQpw0tSx4LAhibV4GcpLbvzpOQeOFP5
0fkaNONaTaPPeVnW50rgiLLVJXoR1+SPc8fsKjjYDuRw7zaA7icv2jyD1OxSnd2D
zsPmDCWsvPH+iRN/EPF0hJNvczuI6cshQCXP2U0YZ+vbQm9Q27diWLhZLWvnENCJ
/Q7ZYJ0bjwRiFYFqepIUUJqxoK7OthlFmcYzVYFgFEtSLFSxv1C2v1KcfzROqh6t
+4qMyfpAZ7OK0c/KK6Bti7wmnVLiQmwJ4uYP0XM/wOXz4aGtDAp6XtdTxZHI+J/J
SrspowkMb0Vhd9S1us+5XbGHXxEk2y49aspyAKaq2ID+ISEbBaSlXxGvkOkWezZi
3lPcS9dId1qO2r/PHcGvFYUtfo21p2qKBBjmQVpyV2Mv9CG3y8qoBS6RRqW7IcKl
Y84okdAO1qZ8mFwuhMGHXxla0YkPBHTz/LbB7sejOy08ghqYtJRQT3iDS2DbDiNE
vqjxOKokHZbNSz7olI8kKjlLUEtA+8BVIVzF4ZfRJBz/Wy745Kp0pV6opbs+XQ3U
X5uvjVnZ1tnLuKYxU7zA69vFUFan4TpJfyF8o2Y4ImiIe5+gicAooM3iSbbU0YDc
mPC955G0jhea7BohfOy3aFNJjyMOBfjAfOuzNcXKZuytNR6Snxs5fCQUAZSqszv4
BOQDWBx8LtgcUbbFRCu5fGglKvuttYuiGGRsvsoefjq0pH8UGL2cA6XXY0Mf40sl
Qk6kRy7gdUvnUT/O1F0/4w2UfXl+na3xsUNlLHPSuFZxq/pQ+8WQjDD4yZ8R4y3v
153e3t+G61j7vFYuH0vCKPuXCj0/4NmTZcens+T9Pllje0qzJBzFmmOe6XhMahzu
U+OUFxDH1kTIGA5N1qsITc6w0dImIDauH/D/3ZGEWbI/2jyjx6Ji7fmxHA4J7dE8
k0g7itXv6bySjhWGgHbET/ka/JHZnkwJ/2I+cKfI9hAlYSh7bt7AZ/DBRobg4W5G
cIA566HWs/O7MmeDLYjByN83AJqPdtWHFailmXOI/GZmqC20YjZh6Qm/S78f6MFW
QCXjmW2NQyAAC8s9Rv9jvDoZeKbQ5E+NoqPgpGmUctdclOtmg4XRwti0w573McNt
NvYJWL4AoJ7dN//nWh9DYlZPwjP3M5KFmOPNXUXGC1DUdTl1pNJ4SGnqtm1QDtiJ
BXFV+ERV6wwfAqAq+a0NWQSkLxEoUU8Zlkh31SjgJbBnKu6LiHizH4PxdsK6Fzr1
mHXNkH0Yu3vwLnUCaI85a0MjGgFUXxEr0WRhOvONH+YScLJ4fp56TgNuTZkdwWUO
ZNvv6u6cA1m98t7wuNrx8ktVP0ms3DgBE2UFvWRRDwHsEP+S1klnLLgoQx6TZ4ea
TfNApkSa97uTi16uMDEvAXO8GWoMAriG7W9XNcvAKa4bQQepHHnkNNhc1yHuufl+
guI3nN2D/CSoplxMag1AyCFKyqhLnyj+4FaEaspKs8tm63vPiwnOkNOXICpJOnM3
Ao7bnkygWbTqYIKhkugi4BQ3nvdw4bS1MmesWydAKMwa7E/oV3tvdCY9D+6JqwBv
dXGjQerAPhIdaQ0Fo8VE8zc0vSO29+W5n2wAbd+BlsL/6RC3sC7GAnaPgtevK99E
tOkf/f7zvtCAqGYuqvMO9QHzX5h5KteEX57Cb8qaNYE4etvSrjs9lQ+fXmZCrbEd
R9ZstVjdsEH3kxPb6sEC+DxQC3+OyyZ0a1zPUaScDs5DXdATs5fCG3NqDhbwccGY
uSxMrfd8aOmy9BwYspf8mym2ZV6rv8ex40viXTEphDGeikKZqPW91RaDegb+2GJx
qi8z2Hmmn1ol0j5TwqX/9Y3lUI0MTzWMxAdt71msyBWQygg0EIKpGEv/MjKPZCYU
6q2aivbY4DwSsom6BURDiEtlef1+z1wENwfJIfjx3HVTClFRlTdmSismh1fblx6X
MrFRuB3FG4iedccd0ogq5fJQ32JXXNlNs5Fb6VV55Y2/ElhG+I3x+fwYqXevjalW
tItjNjjwGdeRsOVzwAp7IaBuh7vrtDGjuTdk8uSc55mRnH26/inPgo3K7HN7dYID
tJi8Fp1ppKA1QLZpMlvPljjCWgZpvoLE/Z8y4JTMX+DJk2+m3caheelQRTJxnGdt
PgQrTH85L4csiBXc0TPuMjUbjQ42E383+T/yR73oH8I/ixAkLfqz0GASWeyVK1AL
5A3j+5HefSKAILf8oGDvOuf8Xd3iXy6Y0S4zl6Y2ub5ty+oEwMA4f668PC17Szce
v58faKjGySs6moruxSC1d+j4s24cz+5gkjZ8eLyXK6wMh3+yaG/EKBg3igbgnRUi
59CYuHThTGzqmkQ/FwVCE6qa23JevLm9TiON9C8xTy5oxj2ypnvMjQj9cmvZASHr
+jV/TBThtZE7sdVExo0mh8AE9EjmrFdslbXtgsf1BfAAquELebG97Qnbl0l3HBr9
pHgvk1vS3EaQNvEbs2pTpWXn46gjnUtok3/mvs5HptJw9i38wmwc8qyeaBJLeONZ
n6VwQMhy7ysKNc5xdgzVs4eSAfFsdbVN2epZnMfmcOSFQLJHRNQN684jzkowtSuU
ACQ5apf+gQz93zMKPl7p93pKGQI9ZEqcP2rTnsX6pOlVtzZKnyGiN4gy+OvTokqX
jdXo7LV5NGzzljqmNrjbrKBnsWdNoK0Y+sf5uPIJ3jFzJ/pFVtaExdoFoLMkgepx
NHUXh7d84pTy+UTPJ1OjEk1CssaGkvJC+/gE9Ymxc4j05TGj57nSnPOJaDm9tKim
QdA2hwPTFIfV8QLHKscXofMF+75dYj5iBaoRd3KNKRGkfD1Hfnv0J8MwHRQR+cl2
j/3XFdDS6fs2LbD5e5N9/+pB4RCIRwxJiNdr3SYKbqfERb+5zn1buXvo55u5GfxN
XMmagdPVHEIfsLWIzYPsHZsb0YF9CTGLLKuPRpSE/ThB4QVqTYxALtWRpWFOOTsu
SBY4M5b/MwvNF63uESoWv5YQRWPVpgg4r7i/XdCg1rN9SFp5/ppwDvKTvbDXyAob
xe1yg/UPB2mGlHli9Cou0XPCVw6cxSD7pSh+6awgay/PzKEJudpz1BUxCh1sv3Vj
2dSVajsC7GLL79arJivrWN70dqr1lcNxso7Ex9TaaMQfzyCyQ1eE4kD+ibJYdbyC
6x4g6vfA2dK8SsLi5P2vqTmtBmd87CMWq14VR0w5FUweJHH65KCbgrHBPlpoOH8n
UyLBXtQCP/GrScbC5ydUDv1OL6Jvz1G8TgTcOBpVwLT/aIo+/ExGi4nVYCCd/8A9
/aPdBCI/6m7efrufQTwEUUIcMx2k/p3kv9WpqV2ED2M9efzNYGdOwvrcp6z2DAxl
3fL5ItCdSbebCfRPuogtZp60MRzOnvzIf2ZG7sGxGOm4dR5dJKUfqn/XzePs9h89
bDOOOQsDHIRa5zpjyr+EXTxRhhd+6BPTKoGJ+bZ2kLkB7H96hzOymMAY6xrnp/mc
/3Fx9URWGEBnohOXGRkWCSFSUd7pvOCiYQ8U4EjlSWNu7lOy/pl1DBx41fO0Zktu
QCHcZrNF+pYTAuVBMo5siIN1gjzrGt8OR2x/S5DN1i/v3BFGpFh5g4PsB5p/DXMq
Tu5nORDtJ/R6MfpjMxpTi4jhzccq4EcqbjlRe0+KKSzHwJxzvv2/BiPLpe4+Nz+N
P/5twGBKd4W/FUuGfmCk9YE11DQbhsOnIP3FbQoPAPiV2VANXnNcj4SUD9K/5Qek
WtjryiIlnwIkRHVIdvskn+SoyfeFiSsPVsaTOharMqRQ4rHttufl1fF44CqW+3jT
uCEm5anOmz30i3wTOp7vVXCtSjGOPNcQHwpgdfFR1qqW7AHK0G65qQkRiuaWsl6o
8hN8R9UtKHiCq3a3GaZU0zbDcAf+QJY09Cqj5gdXXg6THx8m9j0xPGXe1xcIg/Ln
Mj7U67xOWke2KfMGATD+4p72xEk9AP4DROHfjwllt2N3rWfKY8GZ8YH1V7wiCYwv
+SIdcQxk2C4SV1mBkZy+zwI20eIyYks30LWZdzxPHmmj1rjelIag+vCjW8EmgM+3
68wA3w/+rc+F//6MIhBPCq+Y1PxB9Jy0ADKDM1fvIejvLhFfszY+nr2yp/d984GL
OEoX3rCB8Xxml1vNobzBC8RI9PkSTW5FNtEddLKqGgKbKTpkjW4AU/LflYUgCbzG
YKQJB6MSxKvKiLeqSxq6kOmPk9vDWBBqwUVagVszxKUIYk+yOHUoR9UYjjSvJ4RD
fQiCWEguQyac3C+Ejx1DIBYV6HtzRbwjMNAlnAFNrDgDxpsjczdJFuGweb5XDolw
bef/JN2RD4BbCkwFcTQeKhqU1QUX4Xjrlpe7gJKhcoP0mxY1yx4UUQvIp9S9SbD2
OnYuanfaf21ko9k36Vx46eOvqUpgtsWAFIFb4GAGvQrhkd9fe8JD38He5E5k6Rgw
0Xrqc0lPF7bQQ890aGxkclJNuOwKNF8Xd1pdWvyzyAKz4jqH2GNv21J86JdhE5Im
pxneFX+j5XSEwfPKjnd0Zgpqd/vGDd/N+gL6QuxvSkHl9A1OoAqohjhAGeU6+xQB
dR4VqzwMMxa91sZvqslY1pU6ip3yQSj+q4fzxgVloJJE/QRL2vC0ONGb/LPh4Oxl
e2eGDnfYCqiP/JvFObHErFkWL3JsfZNztu1KGzNlWuwEsSLG9Qs4hdW2CrWVuy3x
xcf/cxuMLRZmFofGO0OEPAuLbYEvETgCO1NUcckotkRUGRkQ1M29noGoRYIyxhOC
B13OYtUBv8tiNJSlLN9V4HE/aYSU/9mkKPiUJun8MymS+7dq41yXnTSlgdwwhfKB
1mJTegfBIzL12IF7aeZUTZU5Y73P83rChYjAob82acrSkKRh7XZvdJv/YX4R5mEj
/Us1ojfCshZLPvsGHUUj1moM2huFMFkKP9ALuH3yrNFjK/gteJAKMxtv/mv7kjNW
5Dqi5LCXtGIsP0dOiVUxZSdaYN6Tj2EGsLuMBJEgSejJaFMn5CjIfNXE/XQ/GzVt
AR/XYSRGlojDpH2k1j9TUTqonUFo8xeYD5vZBqaP2PXQt8/h9VmC191Prio5qHbz
CZqS47GVXuFobOoNYH+EEkmC2cdSRkaC9sQeYU6HmrkGM5hqHPikNSGcuFx8cDOg
sKrAebB4Tt2zlFLdGT8HQ6HVVjcOts61NNPEa+ugy4XwZAX1/w5eiH8SemJF5VHj
2sAN5h8BuJAKmtxA7Yq+iQlRBlROBAkXCgvQeUH+q+BL5iLiVTCPVua+E63BUa1t
Z/uYuNC0mlBnqki2I7IUXxWPmT2XUTTgUnj2u3zGLrvsBx2+2XPs7dDnBXBup+/K
IdGm71kRKNEOof1CzdYXH/KxOroY4M+eAUzrb+bEhZIxlgahnq4p1rLs1hbKBXeh
LG7vFk/VwBsGaonjmVl1yeAllASqLCOavP28v6bRJOZa9+bSMpDlENWSZ9HKM+2L
93gyzF+0pqSTdDTnL3E5hyND5Z9JBLvACJfeqnzTalmPgodazx0xpNBi5l8VM8v6
WkvSXVWDnYsSQr1yZUORtsr7AVcvMj3oj0LXKSDwxOHql2yV8MFYWaLfiK7Jmvd/
BWqNH8XOo2oLZhqRlWgCgB4c9lSo3C69gStdRKcHaCKNlDykAf/dURv4ycgjsazg
XLSQz2H/SQxq2ULI3scY8J1EIFwBaklO1RZzL8QcsXkh7deV/m6LXncKAkEE5B53
+H2tXQbs/K7fox9P/59S6UseJixlBwfvYw7s2bszKPolX4Q9edrcd8Rs938LuE+w
HR7sKULY6QNT9t4iRfNkcQE7sPeirbepaYIhbhhw5hiBhmooR26wfzDijt89m/NP
K+PIqUo1uBVZJZr+06r9LXVM2OVeiPx3ndXla0FtQS9rubz0c7SkqTksuqHtjfG9
/WicwQJze3JhLm/AWg4Q8sNnIIwULdDVVOAp7ZPLRsiEAM7VB/nXESgPF+zNwzgJ
2puDVOeD3yJpdFBVcnCe36YZKkt3AdI27Hr1+dFT5IeVMX+YL8MyoAM13yOFdlOn
xa+vCrgXVEqDPudRz2EZ7eTVXx8S1w8wKnXaijxV5YSqU4gDV4Hl0SR1jIK3l7yE
oF5AmEYzuLTcJPDzRIVkQG0dR8VMXlaf05yAPUhGLJM08JRw4uAElATQWljD5dW4
FgbYklVasbr03tioHVpwXZiolC7mBtkKhiWPLpsB2sOPOR7PwbLeVzMRWXa40VGm
DMFJuTYZZARo37NmCHv9edXNVT2j6qwT+vFX9utl9/xEm4t2n4IHWfcw16ItOw7J
CS86ii0HJcyCjJvygh4rK3YtlT/+U8JzM+RkjkV82hxxL/08HT2euzKVnYOLS507
YaF3RJsJmX05lcws7BBmlpWiUfy+KATUlQ9sAxDfguy1TrxUsFjyaCUajk6efOzh
DyQK0izqaMLZZXhJwjXnvRs19uo1M7K4aJxHUrPy8TVNv/B96vRzrvksD7zgMg2q
6abRLiQgpDFJKtKpK4eueG/bAWoY3qM+XNMq2cmnRmztpeG1g7IFD8icwOfIx5pc
MPCpkpE/ygeQJn6thWJIcqrK9sYmULr8Vor/1vjC6VE/6r+IRSQeIV2bjdHkChyz
nf5Rzvkw6WfBhUlxdnJp8Y5/gwBIZ0B1xa8SIbYaT1Gop+FL1ARBA+pgr1YLrESr
BdEpEz9rhTV7bkBgEVySHT5/03xIenWKqMZvd+ElFcDtR1hLE3dVrme21iFKAufl
Ztuo9bUkCrLe8GvCzS7JeqpXXknB2v5W8Q1LXcZ+0Ymg+MbtbvvTx270TtpLxrOK
S2T+VvB7FH/QY8v8TQ1fT4bIhIqvyUuseR5XtCuH//kuJUsZQk/RH8w2KrnyPptf
TCf1RNpSO7T52visnqVbFzOmEAxv6T/DaRtuPMTV21tMSzhps6Zy0puQvdHVBdma
E1CYrIUOVXij3MED2GUScknSJbadiWBey8VUDnu046lQQzhYwxtfBXOVajU69s6Y
aA6exaikQ9f+7F5zqnNWZw1wvbkpIe3lKmMhnWi9q9St2xv93Rr7mn4Cs0fRqmqI
aBWMjMILgP2rThtfeNP+ZzI9wW/EcylrYbG2ra9MSFRrHBCzIdID2sikkbcwezg+
vYU7Vq20sOhZu6pr4m9XPPYppMnpm0OGZFZnoYMPK64Myzrn/4mwS+3HHwdRX/2h
PaIa5wfqcfwUOqM65ZGMDOV7UkuOSwm6i/OCPnv2q5/JkLGygXvtLqKYtW7KrM+A
juLEpjIWx3AelZMyF6hZ2P7ueTmh8aGyMzczOCB61YX/hpH+srA2ZI7FFx2MZ62I
s3pEGe7uO++WhBVLb+piYmmWE4FZGFh7VEPqQTU5X0bOpvMAW6qLNnufcCPzQWAf
wpmbESns+qGCI+x6GrEgCkCr9JZQ7JNkvPvmDolt/uGFZSf2TUdgoc/eZ9482TT+
+jP9iM1WDKJUR8n2rwNORhBHAOkSJSKPpof8h/q9vrO9yAVv6xzn4AHxqzi3e6UQ
QcbCWTd4JPIW98f01aQG1czZD0jSumGWquYJJSvRH9AAsUo7QejUQWYL1q99mhfE
HLX/ljdWIQd4ywSL4ITjeNFuNga8JKFr9Rc/R8i1r+LYDvT1xF8Fp5Tm6j5oVpo1
YEQl8JVLydMNZaygYEFx/24OyCOskX8ZjQHSvjJzw1kl8HekKjc/CTiJxeaT6rrp
auABKnlU8mJZmVXrYburFdexxMlMqsu6KM0JCApNBVsSB+lAkw5fDa3G3KFtVitL
pfmNmRLA+Xw1Kfls+kFjediDX5r7W8YVhyNUvuQAA649okCLPkMT3A0jCJUgTQVX
7otO+gNX/F3d4VGXpAABmx2b7FUvvwtM6Guhp9L2blQNuafKXYyZQDFgo2gX6Vci
ubHc6dBdA8fPBgNtI8qsPEEThfN4MkVBHCs1MAcSFAkS8n7zMbi1XD20UbORI55I
pGz7z91ESfUXIwIbp+mFz+fs/1AQUyBeYhla2U6he8k+Ava2mA1PWiIrq/51dOQ+
rAXbUMHRbixWFJylKhH/Ewgq8tYckTL7gOkPnL/YvFUQU4Zxdt+b+7o3LcvTOvQV
39wajTGckVXgpAZ2ttQI5t+BCjPAJUndaJGqVWr4xbscPE3cropWDfdUCgtJ99oE
iW7AUx56hbOGPhPdjqrpRHJ89ufn4oyNu7iH1FUr6plD3vVgjz8nziGpfiMMpwG4
47Blg83Gtm1NvDzRJBVd7fhBwY+1hIopwOg2gpx+Z0xCHxuuSI3mmmreuX5UiRxP
wEra5Jxq6fhmqGOA4n/60CykrCah6CTCSH8zCgeLoO9L3yVgof31lkfITinbd29w
VWNHPoORjXmZcRjKBgpNFhmNNiwB563uH3B088PKA0K9e9mdgQIAwZbaUsnqgPMn
iztoeiK1bm+C3oDBohZKizypSd1P10gLTkldnQJ2tOzq7JJtmxG4JaZH9gAqvhIQ
ASx1VpVGvLPud4+EyEgenF010WaupKqNrtsBdieb1yVrt0nISMdLs3Ziz5d6P77I
y7PajPZmKneJQae19Jy6wOm8RUiz0v8m4PpoujuR/2hlhNy+o77Cos9lZMgitTXD
J42Ooutxu1WVrQFrj2gdG4jKrwymAI3NGqSNw30Kg17BxZRTLnbjhcJ7xCasUKNX
m0fV+1qvpH/bdDuZK1C3WHDtW1kBll0pasPlPjMQQdFEyWMkJkkOwUoMYkqW7UJb
ffHtwMayaB1EX8X5yg0wOdQP3eEvuJ3HeLcl3CTADLa4BPuc67VsP+SJVVCrVYyF
BJn0UZPCRP8revSLOuOjUAbvocBOs88ks1OHm/XxT/+eaAyVdpxBaRlcbNGCXa4L
aZas66FuTuv1bIfmbL/Am0Kf8/iSA2oju6zOXk8XUQRCFAdAiGdxdy8XOej/RbYK
xQiPSXCysc2As0vRHWSh1qTG/VBryKCJsOXFF1LeC2lJwglYaRWoE2sEooyMmjdo
H+hp2ntM109OXJypIOixeusj6DUEblhTwaBJ9Y3ZMi5ES8dtwaFZh06NbhgFNhYQ
XZ8tyRnaVyJf3sNfJ00kSSusjPmguZHASPva2e1TrExBH87mb7XGDOyqUPzQltOr
gMqWUS1THBEu/tWz3WDzYhwggLYqXP04iTGq6VEfwqakk9nqyJDBCtQQ6VA6+cU4
gHfQdf0FnZclVM9Tm0cw+pQhiLlQkis79yPbaWAlA1Iw2ZrMdc7jHflM/QLCL8rA
bqnPWXsCOW/IV9qdp736g1Jh7tY4SJxEbtewAdxOhNU6u/XV/GtmrcyWhsp8Jrs2
2tq8D4gMRHNWABIucGxiXwY1gQzLz7qYfc261YtZ/KdoOY5/E/GLjP8xDF6Ah+SD
IMvbhTxw0uwZ5lHB1+8jxGKaJ8rK3YV9sGqKV2APHeJg9ILFhUEUWnXV/OYUVu1k
LsZDJMWBsTtRuRfQ7ndxccrJRUEmn4owpZNULp7rc5p0iYnMV1aWgnfIamp2+YAl
E/R6l6h3KvL0sxSvMS1zLAr6K/pD0ltDnITyUQOm19at3iFDGdhAM5Aiuy1Vt+1L
Aw8gR7T2uURSbt6ArI4qJF55OymB2watr4lQnL/GkY8JvcZw5ZUzQZKH229qn9ud
XIKHqVBt0bYbg9K+HjPiXhAaPcSQkpXkEFFvcmQg9SLmd3pdUmqmfLjLsnEOmyNY
xkyvtfMlY1rSdFXOrSGglkrX6NIIZSFeDoRoxbiJa3HNiD+30raFXb26bDT/mZiD
tlvnBMT/W4sibpftOgOKsZAPgVZFYhkMlV9ys8iw2qrznyOEyrdYGFVBCfpYFX9B
PZXNWl3gN33DSqCj2LwXL1wingd73Kk4ENSkZipVxFwOgTuleTorn7TGbdt2BCCk
SYmMq/IKPOqmwR5NlS2PqMUFLJ4sfgx5fTda217TfucJJFSWPiItJdrUJnuvXXyE
ZLnlJmnZJx72IIPfxkmCGPMi8tjLEHennsIda9S5SRSUF+smh9qzykCzrvGtB5Iw
P62Vf45xeLtd0j1Y8jUCqa0DER0FXM57SP9aPHfNTvA5e5WMaCW/wFU1owOTtNCR
IUtiP4hotKq5inRJAnsjN4LyHp/EBUo3neXmM/4HNb60umjzCAFeg+KJkYoLNvX9
PtzwgsjxH2NISECgDN+8F3OaNK26/CR0e/cx5A1sltxRQRuv1Ls+YNLryeJ0Tq5D
5JuaxKBKJfsVTpf9g96pTeadP+swoxE9wD1Llolr+z8ldbok6EpOH/A9U5bmmLkt
sc37JNbkPor5VcKRB9mSWJYuxgqCZA6LhFGtDblY/1fQ68WnkSyUbW3T7erHlLAa
q8t2JT/sp2qlZjF8xwoJGMczUv8JKqNfgZv2iHhB3zHWIwdPcQuaJ+AmkEcqCBbs
jOxme1AbrfdjcchlWDqIIZtUsQxmVZNpreK14/aYMDLE0phCuAtzPVkNuHpKXpNU
8MXTvYeWqS2Xr76TcspTLcGJq6LGx4O6NrBSBY09UmcKHVnPpVvfEsJA/7lQOkYO
SIbX9QqV5rLCSfZb80nOpx1/OFgXa7bHqGbx3+mcRzgmTX3uPAbiTJTVJZY3c1PE
elEhDK8loLe1s58E6tfS3UJLRPRnO1ZGmPhAenIOQQZsGzRlBCLvkIYs5pRGVnXc
A/6GUVOuTdE7VogeNuZQ+dJ4PceEpF1NeWAfZFGOgfNWvDo6Kod4uVYiPkM5tAix
6QXfaqfkHOFzuOJQU2kB13m03BZNSooSYQbrbHYJGtoCIaaZRcnBa7bzwYIIh8d/
i2UYwx2LZMQYV8uarjQkWK9+kmPB5EnHlb1SdOA2Jpt40zuyRgQyc23ZdNy/h1OG
QM7kyqA+Z6FIx897WnIG54bEhBT4YoUyU+L4LJGyMqcbkRi1wDMBZ4lO++ku4UAU
n39Rp1D8PZlWkO8E0t7dUL5a/VhRk81AbzdhmPpU2JC77GOdktG+JRLqy84QWGog
sgzWSThTC0FTbf0R7cjSJcdganJVUFEzNKLYiOR6lwSGh8vOdZOcsXjrfFd8klT9
do1gTYdeQUaLy9UQDv1vlntpJDtuwlFhthcVfkI6draFHBzSLI0oQkj068OHGJRU
sEBDX5uxZuiYJzf7mRKXW5vVOHOPUdoAfJP0d2EmQkrDLedapmcthhQEzShSTWdG
lUB2pZAjn+TEX6YhIinS7d1GzfaZnvqXpaUYWx/oFlk+rgdefzDYG0Ug2NsmeMFe
ywC4wLgErGw3e3y8DbTnpHAKMFnJN7LjVcVcsM0QvTRL1M4ucFjWW3wcYtm5Jc93
qWMZ57fn2Apv5ZOTmsb5Ftxo8jOw4iqdzSlghg3ijhaKls0I5lP6c5SWuTg5KIfU
C6v7t0W85q++1V05djhW3lUf+3DwMqlsgyf96QFNBw3EIuC2RH50rUTkXyTX58Lu
TTo3crGp8VhTIFfH5wy43dWM5X3CxPuJuPUX7nNpspzGDJc9QBjru9ljowVS9b2d
sFiaxLyUQyZLUr1+x5LynJgWWND0r5gK7v9vhqAI20EKesnEoeLwmXbKvGTY8gvA
XodCiK5bKk3OCW3LSdfFjiX3syB0Kw8fmGXR85mx4GubKgcDzGBEDjQpo92D6cON
vxKkyWF+8vzfzrGMMAoiA/1+cDWWpEiVJE4jUq+xX0aE3HMqelWiS5z7KqLaKL7N
9L4mISRBEOhm2Vt8pZo/bOovd298nTlsuSWoybGGTERpwPriyXrfV44Gs35sNbd9
f1HOxEgu5DI1/PQXvNZOimtjkNFPrHXG0eMF3SfKf6nyRmZhvv2MBKwZBdf9W/2k
eEXD7qRDYakTvObIzlL3SwGKR0iIPqU7bWJZ0MmbshFQh0Z6T01UTfQenjVEb7Nh
7AQfTzBsrUr41G52YEMrB/gi9iVqlVj8+yGJbIH8wGL9hYnj35R3N/D/6EgtXzGc
5xcCh3i5aCooTqjER8dfNHuRLNjHsuMB0Xu9Nc0dcTHdA2YRa0k4WAaXDCcv2iYi
rBTFt1IYvPmpzsIk/lWBwMh3Pdb/Lfvt1e+JXCgtX1rJjSUF5o0GVJlNEUcD4KYT
z/oDbrsK8jnlmo2iDF4+mV2aRIzW+FgIG2c2CsUNgR5erIHGfFCgGY8Xn7V8sUmh
ZiSdc3ZlzuWxp7WilQgpzO0WtNvjkvc4ajOa0Khsy/noVTHhJlfvkmsSlbxf68GQ
5hl+rxTtb6C7Zs5w3ScLr8T2cGrtgfeO4wDImJMtCMGhkR3doF9Y8saH/iqYe0br
2cANA+dhSy0tyhBnrZES/IOAL7IzKBQPeCsag2pX71YjnqOezZRtPnB64X0A+G+h
/Ay7FLmmH+Xmct6Plrhpkqvy0F9tLnT48oM6pCKiay4/OdSeq39MbYxDzITMISh5
4FFhbk8NO3yWEyhWVVV+PKAJrVzELleIEgqMpssG1VeeYrAKLjfbVpYvUIGrnTlg
dEYG0A5tiyVVTfrrWjfU5yNZ3Gd9MFCsSKjMwip+2bRRnYXShcL10990bFJPtf3/
v1HDtStu4kVC0/snAxjg+5cCY4WDqSjAp40yUDyWhoVe+XhIAvWl0kPT0utNOS/l
Y/nUIHVQ8GjvaC3dBrNXWe1yaS/hal8aJDXRW/n4uD4XT2r8MhtMJ3fkSDehlJzn
2MUqZ62Ogg3IT3W9Q6TepQR5n1pgAEFhO/XyvOzDf+g9BBmfrXlc545tEE7GzOR4
+GhVbtjO8Lqi52dmDOp2dbVPBLjSDxsIApN0mTmJA+7BYq1VsEDKfKgmh1XDCv4J
u1WP74qceiMNPWW6itOd+EyczRQ1KCYHUcg+LYAib5cLxVuwLyVxtnl0M2J56u4p
kAFd4modMzlWyydc1TnhQY+IVFl9sVJQMpM5PE2F9gmcPlx5qhfIIi2UGgILcIvh
9SMGjMlnHH7Do7koI2se23P2+yHjWCO63iJ04RCABNzJ/sFRADqXkaxUzr+Q2sr7
CTgohzOYNxPzfi+vsNeCIXeJKPnKnFr7ULyPKv80Z5tnclL2h77rCh3OjuGAFI7A
khAOWlr0/JEHdye7kupc8SqrIwJEFfJKBSGTiKWRZXN9CeFTS+/c9exOB1pNzKXb
NLd9kSgPtdETEhQBr0ae6VMFq3wQsu97oSIMX2vQxfHYak2KfJ7BQbi6mBBoj2hM
aO49nuhJ67CdFh6hG3IkoWvkwma9sS8AMeQK7E3g16TSF4XKPN6Wn1wnYhIPR1RD
+OqXmLHIUrdR9NPNKFTiAsg/Ojj2f7mQ/VHdSRAea6VKsvffRTaHjKGTMGkumgZ9
jQCRl5aiD4i+blidfP5BiXosUCKxqcfIenB3qSerfcWhSEAst+4ExFrDngFPIVzd
bu6yCKpjZk7AiQqOjmZ7Ixu3UHmnIaw19jY94Ck5yMpIaV+SSciH+vnE6aKU/qej
SBrKhUL87WCqvIml6KMWNJcjsCCyIkNBeHvAbMmGagmffhUDy3OOLO2bSKKE2zBM
hfJh9u+1c8HGjGzhWPTBLskhsRYsgdp4WB7U60DGby8R8zVZUIzyVRR5AJsGf4Ra
lkURMB1JOSjOhaM2ZLe5KiXpONgtuyD56LIAuiqrgEs8WWRsrYKvDx3/PG1jfqd7
iCjEx5JBEoN13lM/YM440AwvmQf8y4K34jvDzLbMUSG4q1me9AUgCxiOegOFDwhb
yM9HNnAmepZJGZO+yrZoTxNMp/4wOzg7qYfFL4yLDxn1LpSAKH2CL2Wz+PUO4h3V
BAjACxu6UU3/TgnkZCmFbxcKJarbmdSyagMsk4KlKwj95qD5BiOzGIfThKDqFjZQ
deBfZO19AvlNEsq8Ci1cLZYfLmwD/TrTSRbvV0c/ufVseQfnU4vUFR9HqJN1BocK
njEohvlI4Vq/AZRkLZiRhKpLQITLUixSJHokFf4OckePA66ilLbVBZ3TwOHUlFmv
zR7DfCxkq/cdyAqTtBHRgh4QCnDlPS3XyEFVUOU/tE2NagxmH3b3imHLI6uzpDny
lDmisGwuFMBNoakAHNFiN2YXkFs1isnPLmYhh5z+xlO1Pl4CM3nZ1oO9TF22TJQ2
hjWlu7ufABEkAErZaxbniBS3cDfnNOSDtOENIS8SKCbCxPQd+8l72qHKX/eZ+ARh
CW8Jv1cFAZckV6faEfWDIrA6VLm/auQAnwipTIX3Kmb96NWqA8FNkpQdz2pHK0te
Ums8+W5fd8XOq6bO4M3dKJfFpFoC5TOSz/MuAElfRJwGLqu5rj3ia71aXwzwmFMl
qBHSGWpOCC0mCHoh3djJ11/0DN13aHdvgPGYFUhgFQCI+/6BhCTRax0+m1bqfDcE
nJyBdO2mjrJ4h8vaM8w02ND0UtMrIwgF1Md7mKJ5zTLB/eWeqbpDUH9HamRhNN/z
3oeDjdcEk1EVBfUWYhfyLR0KcFBYSYXcMahwJd9TJ8CP05u/wKmQoh+aI4qS4CL5
L1ms+mlRsNWnfBPSlvGh+rq6fcqCkkWZPouBmzu7C7fjGJJXE+MFy14Sf+vE8z9p
kcqhCMQddf+QzL3jOZ7TvfJHUdrFCxIhzJOEVCVIAt+NhZ7ZAIwnRkjtzhCeqxxm
y9vq3qZaD19//Ngx0oId+ZOU4HwHfbx785l6TVFUvmkNBd59Dk3y7dWFtfJezBaX
Pah8OAa6EGBQvH0s3K/IhbQh4fCXsh49afRvCh0pgtmN5YJYqcB69HiCpY1R4Ik+
tO/BfHGVxnuyFgi3j1nGgvuykLgyIyKbelbB0qij+Jlk/tgSa9LnJd6aljD7X+ak
ovBdE/3mfAD6Uv4Os/xuAZAOzYfgx1cq5hRmY2sLVkoVC3UAtuhoqETRDML6Cdtk
x6IYxz+ze/II7SuIqQZlRXk3X43mgpMiUq0hkIp2qR+/ej2CG0ptqJuA9/4MFGlb
otAW/MMg2W5JfFcBIFBIop7hJNAT4SlAI1pmKJuOeUf7xbcFHF4u3hbY6w/YSbMA
DKMHImDh36qVbHufYrgDBNXppRcPCtSb92Zii/hsa43pcvw+YVORCty7q+xUgTCA
g+k6C37kcIsIujzuL36Dyd3ttTowCOBOk5MfEb/N/B6xldf/F+EA9atbFVcQdoFR
mRBHI+n8sRMTmz8YvwRbkGCu5A6JvnXE1ANPb6ebCZdZdyjYS7H0BhyxbvmUwjtS
8oHn+dhUe+FYMb90VS8Vo08J2m48Kq7TZO/BcMK5RMhm5vCJbXZojFQN/u0IR95P
wklBInlDV8xK8+H22XCz8n8mRlSiF4TfbMxxszgyf8UFC6liubElfXIjnL1fT2Hw
C9DXrdBaXNXzu71snoWqAaPDtPFAJrqB6s7eUetA2gVaI/erZJvU5UYu5bh7FLhL
WMMIYliBHlPVbmy9w9LR39xyxYyanlUL4eztONTpSKgsN+PMw2fj/zvUAVz8dbbe
YFg7cJiGPmJfRN8rYqlQqebLCqD2Rmo4vzE3awNviWuvC0USaPknJFll0OV+Rsye
sj3lx8jcmJMStNkhlIh6e+47Wa1Wac6gRsY3eyOkEPtkG76aOx8yEb2/lZw0l2MY
Ansg4gnm/icLBxhgdFMGnCSC2a/sc4rW4KbJV48wlUt2xnynsffT8PLI1PxR+zo4
0Pi0sspT54D1IADIOdhxYrhdbkFJ/jHLvBG1/pUT+CZH5R7frvmqS3+/zjzq3szo
feB2otOYsrEJGs6kZpM2Y9KF03ZCop6bnJJpQ2KGdHOesGTdlwSfnuEfiGjo6IK1
If28ikWLIuCeLgBVX7kq6DeoEAPkGx9rWqlJJQ+ne8dS/0gKefSRCfMkb5eV8uTH
D+DlrCZwwe/SP50pmHhVDl6l+qIEvlH+tWhjmDnBgl5Vh8BsGXX2Z8Snj7AMPM9z
eSW3Kjw9VCSeqIEAQFjSSDAmWHtD58TwyOJbIx9aPRn1dj9IwfsbOeVsc+Ji31As
aifpU7poHcTT5qDHfszMDEc8qQo1UfGRMoxv0Bp5t/NKcAQ5TbhKkBb8a38LmRwq
S0tGzhnAIiVox/uNRGjFYz2kYmQTESDhf7rhLaqM5lJLdDn175RZ2M5VNKsqOoVh
EdqBoaaP0h2AblK9zSCEiLA/xteQJNFJUBiNdmytvFeMo4LHT5048GCHmcq6zJgd
MjsmPSuIvNhfroNaY3LrOBo57EeeKOotiKUp6L7J5NKPybrVRPkBBJ5qXxty6513
DplO5NPiA7DxqxG2VK2ojJkkSsl+6wUwlF6VgzSvMUNB/CZKX7nXaoKcBz96mrFO
gMBU12xruFSI8MQtg8o7WNoB12vK5RQ4vGeo9LTZQDHiYE37QN2y89xXvAohnCkp
er4m20nr2i3TYYisYS76AaNgY+BEXSmS19nJ6qWp/8pJIaXeRkWSQ8f05en7PxU8
nTc5cE8ZxG+yFwUZXyEx86BgxCHNrRrZ3AEVNUqDdN/eUCOr2B//LPvaUuUGfESN
oZ8RGWwR1ny2FyqaWyelccPk68rB4BwTG+ZFbPLPK4QwH0JX63GOOv5CW2YutEnk
jA4F9wt6ALGlL6nWIOjGg/RlfqkVRq0+c7IKtRLkSCo4E+EOcQNcswp448bHGlnO
NibhdGMpZG1HrBg7V2KBzT/GJzck79YU1yteEDgom2ZXHZvff5L9mLI281MfzNeF
23d/XIFIa/3+iUG7KU8NqV/ZdDbScGlvNHzRRO6HAebyEnNA9uOSHB6YOS/8HHmi
sHxckrOmRLxcOxF3qOUq+k9fRyD25CL+lLCY+0PRxxFhO23dlXi3jXvbvnuohRyG
BgG/S+l3Zn/ZzW6PD8MfK4SQ/46MY2vWG7ELH56s6fczDGBeDQ20xq7Hlz611qUu
nuG+TaSwQSskHKF6ZogwOlYkTHzYuKHVdDRj/ooTOBJK7lzPnw6ynaDLbkU4jRPQ
7QX6S0aXn21yYiGS623mAyS8Y1r3BrQIOR8++sZqbPo1C5pD6tgbp6xUAqmK/z7v
82yJDv+fMXzNBXgSGuaNDk4llN+E+AwB3g7rCm2WU5h1yiGzmQMAX5RfOannDW/q
e69inGjUsC1XC45dt5hkFgznOHHEedkfE233EHUXCRoACDuyNaX4FAT+D2aJZyxj
vrdnZvLcfYHzTrgELLU5hHTq5SX/iuVDpVEfmVOXX0n8kRA5b79OScJtwRons1d5
B8fO3vIuoH6Q9q+azSIL/5kjbmkUP+x7eNrzbiAE9cWv89o2WioCPKzoltoT0/M1
XsNPFs2WTxcmMsl1cvDEXLz8NUIJLfVIGr6WWumB0vnLMfJojvhtMiCiSiJhfquR
sWnnyoCH42l/TvoOF8mbOUeoXnroxjdF0blC/bILm8HfAJ7BH8q2m5NinnwJOTN9
nxevQKkNKHlGQ/Uyq/81PKW+jv/zP2FJu8bExWwmEOJJSMpfy0lOXSUzF59sUxrs
O5XCExFiaCxNo9IoigINt9K7O2Wz7fzA25wxflAfDEiQ8WaQIML8qJeHuq+U0aJQ
H8jvvd0R1Au7yLFAcLmlEgHh8mgmnjAqECNz7iJR6LCOArcXgarqLiAC4ZyWdiZc
TbfAqzPdiEXHQoluXTfH4lrWrldVZbPkGBO82XTxL7jnDMZYpjILbMuPdInzDCcU
RzobXbmesmkH2G4lygYJ/JsN1OSYm1Cifr9PsX5t9ZeuZmd2Wa2ECvRtgLklV+/Y
5crm/xMEhVxdiRmmmmZQX/jYlyvrDA2L/kVmdjqA66pBO+eImSJvL6uzF2KeYF28
CtmTUpqbFlbNsxECjbesh4F375FQzR58T8sGpxGmdeiB9Q5tlCVldY134Xopzncr
qcToLoXXruwWsSNBGzfqPxjIN8N1pJNe46nsY10qCdKvKkgWI5YLcxcfYPnZ6oTw
DEIdrOjZqw8jPKW2gikJwK8OEFh3RlDXaUsdYAarI25eADI7ALv/dYNZOHD3kBeJ
y0f2KLcJsqeiirFeBDqvLK6ozznZ/UULnPqndR7qm9jVlkxpgwFbBhtJUj7YJj2x
pd1+wpWN41NjfUaOykejCUjZ6ewPlQhOS9l0XbNTu+6ssbEp8hSZsQEphXuqxNrg
dAV2JdSslnrZDgoCJG8E5hf5r/gu6uJMKplEbaEnn7d8QK/Kg1J4/lD4w7JcY27i
PFJYIimdLpk4YvhHRfje0j5PXV1IkrojAAbuioEestiAaUtbF8+1kfIMQ4Gw5zds
P5LWjfA3VN7hwjs0a0xP7F0G8D8UVQblHvUZxJenaavr4AlsATVBqbH63bjAmTi3
0IxNB33CS9tNrzhlWFcPjnGzWfGogJ+bgdIawRj2B86hAN7511SzacWxQJy3Vxn3
J5FdCFL6tjdFuhOVwpR4FSOsL4pcm6SY7SFuR4emgD4lq5By8corsupbKUSb5PPq
AihGCeUEf8onHtxpb9/uCoxIQr1JiRIsbOnglOS2mnLQkYbApJN9EHkLFP8ec9EK
monJFHjmMa+bZ9lQ3v6khTR2iDw0HuM6vU3Mkn+Pc4e5ll1uTFb1V2oR5VmMSxQ3
x4rysTOOsaS8n+44Tgyv7WqK/1AR+83Tqy2pJ667MoW/IZsHV1+6bHmaeluZEiJO
fAMl7DezDuXIrGaoGlFuU4s/qBqC60Beb1/yVxUYosdC9E3ektasqn+xxzVbmF8W
mEQiXE4/E+8gFcS5hq9Z2YMXbGno3GVt5zGjAuBACwLW3nktELULI8nmfLm4mg65
Os0eknBBMMiSm0UURFUNJHh+v5vop9+RDqDwuS3vvOs+G3wpWkT6Y1x/YhJaELk7
Q0oVa42AndOJq3CH6zthPeVlYQnxz+Pjy94P055IQ1sbZgzhrWNqWCIwwMNPZOLZ
iC0Lux6x6uv1GZT+88VlrfnloSUYY9WPt0CtG8Y76cK92RULTyhoLeKfP2rc68l8
QCGrJqWWgXnGWorw6yHmIizbcbzKbUbNN/eQESQyTgJBKMqEzIxUI38rH3e09JXg
lbldxy1p+I4fM2xxt8nff5BmN/MHmBSmSJq+XnXUKQT2bTBBXY2sIPv9iydk2VZj
S7BMMPAZI6siokZuoZ2O0MgVSm7resFyuj1CkUdf9+cUezO5G1L2USDDK15UHxI/
iMJXuOFSV4MEcqWqqV1HW9GUUvyfzbvvqyml6PZdxIqCdkoCSpBFKpPtjYB9A6VJ
JWhAs3mbmSAlM9+wO7A7IFbne+xuSdc0/iueWj/X3hHpGRrypobkyX2dgnBjo8iz
ok7PVYuyrRt2JxKN5P5FobTorUQitFbrUWfVSkLnL7ompSMOPtGxPXFAdFztZsKZ
z4wk+KbnbQrtwUMGr4lH+2GJVnUOSXErxuToNMTjEyxBFu3Sn4PvYlAzHQa/qxYo
qeCdjzrRKVrf+ydHCIhBBPhsJvV3zdmPPIzRbhIwBENZwvzSHRggLyLgkVbr/nZ+
buMb35IZXhOTTkx0lQhVEKScwtowSo6D5CPBDAGXPkGL9hPCbYpUiSLVXP5C/Dh7
NH0aEc9L/2L+exDLXCKQIrb7XoGblXUn/xHwfVvmDVCBJJWq7ERPXVLoLMxR9Xkq
Wy4Bvfzv1JhOXUiTnCFWYT8DCXfWU54fROssWQz9e3rpzgZk7qlCgn35ixamU3Tl
nNX85f3Ka9k2QsQsEiGl9yMZ8TByamRxL7iNzPHQgHOrwy9IS3fFIfSocqOuTchE
ekcUnDiVVMogT82oc5f4Zg4aRnZgO+N5O6aB6KIj8YaA8mBQAFBP/nOp1ePNkylF
tir7540DD+3NT8JpP5qjSBikExpQL/DsiuANnPCZslEhUh5dSm0NuAhICHsLJMlR
67jWXVFbzRhw9Flp4ZwTNSyS9hNy8qwA9UWCHoQu542lPlxzqnliJIU28hprfzOU
s4BLBCpUEyDNYxgXwntsai5c3WLaf+LFyMxDTbhja/R4kwOCp1YhVzWPimbxeiEX
pz5I3dTRrUsJCl9SCDsRv8TLYSXKFhV0Qy4+Edu0OS6AJyUzed7pXSBmRmR0KR8q
0iUidaJtVcQMHVjKVcJMp2VpG+7eBHQ6eagy+T0EVStNxbdkqU4VOZSmgHy0ncms
7Uw0L252zFF9Kuk7RLqwBHkVU2Lky7tSJ232gPpUvjdmXW0cd5DnKp0R+ueOmFM1
4yCt4S/UH2houh1Mp9VHbzgFqF81Ivwx1CzsNZyuaRo4btYS8fq+bV/D6iIkyUE5
JSq39hTicAKVuYtb92XxALdonn/QuoblOclmEKMSHb4IKhc8Bj8KK1K+l3jLQNbF
K12YKzEguZUVDY+TcnhdzosPR+Ndc3Se+E7F0iX5ZrlHzAggLC/pGqncQyCPnynr
djoGrQGa8HHVzYivrhkrY0BWF5gxnXHFyFYwSSlQhozPN6CnI2J3anA8CQlTCZ1D
OzvrMVJuZoSYrS+TF1Q/RjfGfnENndnw/qCacbmfa4GGR9dWGjFbHu/ZnSnsOsGq
2FK1ryLBkOZW6QIW8+KgcbBN/wvNuGBvTsFucZF6rCUb7oAaXSTplkUuR3/FhoCl
PwY+krB7XRcRVKqGxa9Jtlj9QUbspSqWbOVzfJL2biK7NYiQpsxEP6G5W7I/oOfT
WWKM1UuYkIppOk+l3ux7Yo+pLoNQircISmqGzagV/kmQqT9aksXCuPc5Ca0SCifw
lkOnlKxVr/aZnhTtPsV/iBK2bX8gMLbP5cdEiOfpigLJJWpexUvvw7gaC2apaAeF
yvRcVBjts3sCSf9nahI1cqtDya7rnA/1/QFCgiXz6GrRB9jUm9pspl2mlzvbWBcG
lnGdK8NFghq6v7nzd7TzNwL7nSwAiFIcXmlwSyB5rNFtIL8l/vZMR9/vErNgl9hN
Qr5oCsZwJ/J2hABWNJ5Ilkd+86PTN5/+WLHDMRH+yeS3e7xpXvxZcOzSBjyT0HJr
/1+A9+jokEKQML0ATT+0BE0YOFkMCysnMSrqCYUjfkl4eqVhcID30Jc1aB4ZOxzN
RU9dzRW3wTN56C8dAUz54povjWbSOZgJrHLXYdqdR0jHy6UJ02KvmwMrzpHkPjLI
oBubZeGG6ty/LoFoIVaWX6KpZyPFdcIpN0eBy08S0GijwqzFrO16O0kBfF2lbaRN
vlquA2b6kkDoCTaUs8b1CfVx1VeQTDC8IfH/1VupNzszxudGcL/NdF23ZQ2RnOZd
K+kDtPN83j04Rr8MdD8scDlt9/lhVWajgkyfrXDI4D3iCMV9eoe1FQXMSznmQPzD
3/OuzlP/rr1MdxYSlRS6vH36tmf0Iv4Bpbm06j/Fs3qCPB5c3zibtQwStBARqOQy
IO4LhvMsAA5NrkVvSYgqfPRpsN3eLhEiTK8p7mD3q2FQnnfD/3CT+AzSvWcjLiGy
JZoQn4LhT7rOncfVjW4iW2ErsUKfIzy9nst0HCAwv+Ec4J+8eQLVxqYkmKQkYZYr
37NJiY9O5uDFXbmgDTgG0dJBtBGlVmxt+m6GUHviHc0BrLYikfeTqjm2c+AAuUwp
S6ZNSpAVZr8mTeRkU8aJ3LlGBaxNkULIuUO7Fvn/T3ulDKGW07RrE8zb/bAHxexw
vLpjumqf5+t2XTynkZ2y6tWJi9dKdOjyCXHvpTQAWeEDozRSX47SMDiKSA0CMFMO
h5LgPHWpbbmkhgLP0PGTH5y64IEZaK527fAVM3e13FANaZbBS/7LYHraLvpWhcfm
WJ31pu4he5HGxio+VljUxBcUnLnb6fhyItw/u7S8fVW3ADfd9uOzT8e4QcAD12Yq
maNjA5GFy6XXJDrzUFWgfekiK7Db+7k4hJKuuh+hFHajta9wk926liwnKotIfzZ+
HLOez4bDORks4tq4O3ZAa9iSVPcrg7RY/vxUqGf41oWQvQpSnwWv5Rh2ARl0F8eD
DFOnn+4mVrk+cH1Drkg6/v2Z1n4thEBnZY4moM2YHlVbfp+z+lA4gef7fF0RpbG5
x/4p7i5FP2sZCGPvwpae3Ts3TCIgHuRTBKYh4ARVfsM5peDDF+h+HiNSe81Ud624
ZB4wyg41YVz60QXbJvNQRY7KfqlxyVYA8qp/tNdPvZ3vdpjgeiVESHiBjCp7Sw8f
VYItLLefv+R27adZwrGuKm1Ghs9YkWzDpFGoz13rPAyQL/lPO3X7qQwwYkZ/GYnN
f5ZCqvcA5n58xBtvaHQ6b/r5hCib/rEaZNgaRnLKmjEcyBeW0AdWmNporJdRnkZK
YueCtokcOvOpQeXI8VOOk/keJNcBy0r7vcfiOYkbNWmwRirOOw8Qdjx+3PW6VTbA
Q9ldlpFLe4LSIQGv0NiZNdlJ/HxajhSm143BpAvXxJJC4oH/OzAf9bngfYBJwBib
esUbenmie4UxPpZijaPXOKWWuyxzWk3ZXNEwLJt04m/pfoWASK7kNJStDiz+0UG0
iw8PMDCIbRICVTvZCPuRo7nCrLDHKu3mM2Q/oDLPic6KZGcYiwYT+dVQRwBnfnLC
agBTpK/q0MBdhGFduzjJc3Y2cP28mwIvWXFBdmz7qTB/6XDUKO7oZZKPZPv+6zTI
atPmySwrbT3yOFyewZpUfMyvPiaWUGippWmoHkNWXhIiWcJRCZIH2IZm6ICa7L2e
aB1zBDHSn8gEWvcWtPIUwR8Z6LFRzvndqVtLug10MODFNs3cYscUXF8avfOLPPKx
+opr8morXdV+f9EcNCpFibIlllW7Wea8JbEzUO+P77DYGcM8/l8+mHVOExONg3J4
fvhV2PZVNS5R7ON99Pl8OZ54MHwrvPGIp5Fr79R9e+Rf4i1Djd40/4NGMN2GEXaR
+8LGVa8vNXUg8y/brjiePLjxzEA9yN+4EPZt6HVlNIAYOYHOIG0Eun9JK67rYdHH
BhDFWWa2oLgi0nyixY3GykvvRPCeKb/BxaohCbvmRD/WJZ1TsD8NpO0JrV6uK8zb
ls8cr5K530x0Hr0R4e42g0cWMpwZT7aC9kGwzJMqNou8KMb7hGHwyZPh0Yo27Yu/
ZIrIDPi2+CcI0ztwDE1vElWcMNGhJl9jyfpP7S3WrAgApU/uEuHBtoJv9d2IQwFL
uNvn0yYadrAI0qF9BrEc9MlECCUXIy6QPZ4OWji0pJMrBKVBw2HgpzOsWN/w6l3u
X+prpl32VxCaZpv9OhMmeCLLHbR+0mfyPuGELM3KO0N9ezbFdfM3PFJbgOjxgxFU
Dz5fmWDGVASIjXUcxfgBvJB0Yts6G0cHVWSGTBVfTk6Q4NPCOa4cJt0g59XGxPAr
aLAm78+yfrXHuChGybKtLW0upXRnOoGz62Z8qdXbPLl4ao/JDS0uNfBpqZD6Sjjp
x4jbhgDhPa3KPtHAH3XfsDDsTlZDhrtsgYD42SUs+WFllx6NOyXVF1ybfi3s/Q+W
f7R0sa79gH6UtE6K6bJrNk343SbApyZnXI1d052iMWVbJmnMt/kvTeo1JgRVbZvB
GGsW/wac+UKJEoyX0asXS9q3ZqtIEMumhJK3x0v0pv9Pz+Nd45Koe+kspmdB2efY
cAcGa2CTGH/P65GwcsMcAmlp6GKSXGMRhj/CLt0UfOYK1jgkSrLQ/9ltyT51eJjZ
/g4zn14m7aM5ZGRw8DzoJUnqstZGxplBmsA6u1gHmhekNzCJpvNkp7sb39lUenn2
jFPWH/Kfc34J04gKJq7KGZVWBw8y2f/2qjKon8duNaWyV/NBeLWF58BBQm7Y3Be2
10zQMEirUoc7alc8pmP9dpMqkXgFvYCsx4QNkWz2AQ8oSrxzGH7LKblG3J4ucuoT
dPrYqBUUQDoPRiNtbiwqNzRLrc7SMrn8uovGBc+Qhc5qVBFzkTexP3AJfpKuiBzX
td7S1hVi8V1SdWe4bJ+GkpBN3C/SGES/RirXDgUTVlZSyVwncuFLYWvzpZ/FLU5Y
ZVsGqSz1oRtXkwh8ehnjQuX40ITjP2awOv79uL41SURcXZlSBw9t2VrzqdW5FHIM
rTnDfkepQaw6IR5xgxo4YRQzRwWuIcVjXfUK4pLIqYry+FUwYwvyhetsjhhIuw4p
6Ox5GF4I9ixok7NWk39k1uW2z55IbRMy7TIHAExsou6Yvz7S93YpZtDQKnfJRXIv
QdjSBJ9+zlQjGCcJtr5NlPsVCDTuQqdhk79WiJd1RGX1OQM6eSKgoTtUCFWClH9T
3q/ErDuViaY0bKj8cvw5tfN+a2if5g56Sax3gVmfX6cvwKhAlHM2USt2F1gwKNGv
t6gTHsZ704tvfYchk9IUG2fE4TY99KBij4hTVM9TNeWx8JUq+3fzqR9s1uz9C+hN
KASTXT1oXyYLaE5iqsN6YDUZ5f0lX1n5pWkpxUQ5IlX1o19KREJeugdi1juAV4G6
a+2QF6LD9rAJBNiUZh4fVYurA7Z/XcSAYVrVtYdB1FZh2AIf3W2QViiz08lLU73L
YAE96M4awaI3adFdo2/njbBEJaCXoKFEQUae5nVxfKr1IGMRFY8tY2ikXbjDSvrS
ND5U8Q0OCECOCVmJyTsX+evT9e5qFTohO0+zCIWISjtMl8wN5ggaSFfO0qf5GZkD
2TrZ7GNNinxGvH0EqeLNdL1V1R7tAmk+IepW0XTq4EuwGQIiPGMbbzivU33dOIXq
GXK9Ib6lcg5b9m3b7g2ut47fFZB/W+KLSxLClZwbzqmneYsVabY8DK/c/qjLZ17c
txguqnKNNgE5lgWfW6ZrZvPHajMHsu5/9bkZQERhHrtAKyB9bGUUSNsNZQZV13DK
xFVp8MkaJI8X6NkxslyyHpVtFUZ7FxxQWutqrABiobBarWcstEVugzci3biVnA3G
QPt3gTJDCp+fzelhLb2+FlCxBs1fsMoFlcuz7fXXqVAclk1L1EwiB8Oh5/VC/3ze
akzmnxChDViWPuDjdWuEpCTzk9uRKILvt6oc1QF/10Q4NJ/jZX+VeYC5gtQ5M8ao
Kp45TVV2sf6+5WU8RCF2pDIUjRhep6hyQDkTvyvQ4578A++JUi80psZAkacknygo
C1E+155LL0QF4ZYK5kB8hqtCRQf/wp73Mqvl+rF17CkQgCo3stEvz1cL29ToigBz
A4CIlSWA+e6bVXoyDUD71/g0eLtMGJBhmnfVPrH0HQHJF/+q2y3Y9f9EP3YAUMgE
JkGdiU3jjy1URgGOb7lh51JVdNZELLAmnNKA16/UXSOKUikaf71dXpQ5RWp75k+Z
fK3VFZ+EfedS38pYvDzgz0Q49Mtd97BxAlGnAc87GgjeGtg6gypRyeB9S6G0s4BQ
9jxN8bQuvpFAje1h2sI4EkxguIhVyI/WocoogfymUTcgErL9HAnhSrhxrVbI3dPF
5K40F+fViNLab+c0R/5MHJkEqpgGEMO7yCQvb8PfqIfrNRVt6dMkOhi/Ws3eFSn3
Ejzb3N21F3jynYzeYtXFsSbBbzaKyv/Y7Obh485oYCzAS9XcA6gJYobYQOUf8BCZ
lkYXVQGPxpTb/ltu2t3T042zZHT43Oo0jlUG3zCdoEYcsmjy2Zr16WSxpSXeymBT
0fM2y5YGPw7+nfHl6AofCYdKxCW5UvhFOMAvvVtROigYwybuyPzLrPTFZcCEl0zn
5f6RUTmzpPduvrtLny+ESUScyUn6CZLFncNpDI2Ke9Ab9f2ii15wc24w1v+WJfqR
7gp+sfM3Lkwe08ZuAXMIv9Kc0j/x3TEX/eo9cr8vE182HY+eULMOLW9gOF23y4VE
itHdN6XGFrdQ8v7g0fLVhMZOPy1iHbMq34XrrfSixC4IYpwPY+xeAfuewJvTw+O5
9UdJnrjSnKvAFyQREvCLIKS6UepbmEdhOqjN9g9oivr1IMa2S7+CKr5lpznsedT6
2Znedb9KYtcFG1kMTj6Wk4dvYYPyhVKSsPPsPaPr9bnxwsqTrZcEQIapLQ+XXv1M
XSCZtyEifO0ZIJ4zjLYL8rTLOxWqEaeZzljt+kqtt3QqBkk2wu1snDX7eLqD281M
lNaiQYUCPQZp+nWUEUWcAUmgEoced/1Fki1CAheNgv5HuUVVdatwfESx0zvhi5ss
AiSagK+3rRlAziOKoO7Jlk26vEMayiCg0Iig88BqoEuZUpUX63f6EF2TkKcRFWeD
dHuLNCObBHVz0w+SJPey4DNQvyF5meR26UH4gW35jLsSb+8OZqVGqVh+9QUf6vWR
YBV3umTiBrJEs0VhN0IZ+rriXq3tpq02UksV1L21PBDvjrfoxgxAM9j6g19QdBfQ
d8qu6LFkeS+rNnWmba35+Prxt7uWZtJwBwjGqdzkhfVAgp9N3JsQGM+AA3P0D1Ij
IDkTdtx0f+24810smgR9nNfzIC0CCVpO4c9HZdF5mGk9sLn/SJb22oa6WUerguQU
pvtdE7/e1qBCoHitKKR/aPNP3yFcGjnAKW8c+cdHox04m8zT347xToys+BgrWVhx
/t7foi+a130FF7gx38izLsldPqUnHoIWYP/paw+SCkI2/x0rJEKK4AFLLZbTXD5a
WzpfghFdER6FTfvrHagwIEmWjX4rYgXqws1bb0403HPu9LXL/3erAjldwExL6iDs
ZmsUXBttctWSOt6xWWQP8vbpzLF5H5M3omP7cm4nLZDG6lgEUBL9tT0xEmLqKyYx
A6U5r9YBU2kXwI1b3l+GkDTBI2v3I19mXQ5QP+fyxOJPzET1nfldTKjk8ByQw2tO
duIXQzv1v2V2NSEZ3SETxBkkNKq8mRQls7kx3qMZS+tw++vuEEkDu//jRnKLDLs4
spbXgdF9qqxS/9nURI+tGV1j/w8OZa4+b0Kz0dGhLiJQS+fNfVz2eQXBzjJ+fm8J
ZTMG/HhR9tFhH1itt48nDCN35U9+RzAMuFowL5d3JfbElkk3mQOD2XPmbaf8djcZ
d9kY04FHnH4Oiix/uCjdsjkMM6mp9yNFYK71JZLkjrytw0jFqdhsUuC4g9tAdWwo
mfJJUQ4EjovuboV0vDFYQgA4C5Kzo6ZbZlXHCZslGu0QQ44AUkt9ExTMFwTn9W0w
sgn/MAKlHWOjOX4tcPbjDv9NrFHvwV4+uB5/Eqhh91PK8RELFwZmOtDGWPb2a85A
oc+V0nog+/ITKyLwcChHw8WY5mlQkOn4ox1A6y5klMavbHGYe5HqkFMUpGi7Zv7k
ulQ05JxxmpazaNdeVku1fBEXP3iK7b5paPjN9utG2+RL+fMNP/CCKGdlmixa+oq6
rfeAdi7lIgxL8WPT4+DUGKIzFPoRsMRqoBzJn6rUc/9h6WGpLdZ86JdbX9SKAzyQ
VvIYtSVNUx0iSsaFk6GnEkD3a4h0eUSwsyaKkQRGl+xeWC5Rf82TloOKRrlFkUD2
mocXU3I5P+4bPhB1kuqUj7OIQWNrYuu8MrPMtMyfcZRF3TSJkpAQAi5m/4rtcE78
4qce2jPYME5wjvyoWeUrJdUT3lgzWiQf6TRx716KVO95E/JGzBJjbvMQIp7gBUFr
aPuuW+XUwaAr9BId+hyWd/bFHbDXUV+X1VQTTLJj7P2BJk+Bo09eI9uDobQEmAez
Ml9cvHtMfXcnEV6pqgZ9r0Kpmt/d3DnwBER5phiqnz17pE2GkRO++zNX2RVBzF8Z
21oH2litZe0MB2h50bwBt2OzgqxvCEzK0hWglW90FNBT27iAuMpAbuSs1Hqr9gqj
+yqc8rQl677whz/GWzX3VxwAUmHG/aNdCI065RILc87HMSVbbpX68VeHIQCTfG8x
V2Pm7fJRzZgw3DGLfaCc4uVJQN7hlzRBsN7g/azHaRaNiaX+glXJxYjnBCqKSWB7
3BiwosOZgM/U9LJIid0JUrgdBsI4oD53Yfq1DeQ7SEguANKiSQ0rIqPq8krjOiZG
bgy8tjevZqDBiSpCNHcRQ9JNpJjofEV9UfOPAhf9Vh/iQJ62M+kvYNKWAcCHcPDy
UB4v8wKOqF28nO7lkMvVAuOzTP2ye2RnR6hbcMuCxquq+l1RousmMftqyk/2H2kV
aZ4d/S9uy8dMD24KCil4eQRT8wfvwa1lG3Qzs2/G6W/zre/qBjf84eVmGapGn4MH
QbvE64RlRi3vXGcWnufLJLWlt/iL73CP6Dj+pRQdEvwIgxtl5nNlJ8Md97KWICdj
Pz+ipG4nk4oO2tt80V66pkCmzH2ECRbKOTSctBIy+0sJZ8W62XvCbmSNmgRVAuN9
IrUcvCWpP4xv3u0dDuodlpUAwYJqZIS+RHQm2kpMmB4EC9OiiKaXCRt2qCmngnm9
/0G6ybGTIKya6Bg0iOcuYaXadEulhM6NuN+cc5ccvUE0uZK8GQ/aOqgl7J5Tw7Un
CxM6RxWn0q7KBYbTXdJN875H2zp++uw7EJTGimKHIxlzKZQMP/wT2F13Uo1nx32A
0AG9VDa9IBZ9sjIG2WK2RD4MOt8O3tc/h9lzR0oNwBuc4MBs5BXMG9BrOD30fp8j
YiOqAwG7LNgRnjYpcf0GqM26LAkmmGj9frlXvosaESJ7sEGOl8z2QnVdTaECh7Ip
21bV08+t9ihFJbdbW1HblA2ha1FqH2wMF75A3BD0V1Kyqkbi7BSEi5fMGhxcdG2j
mtl3FL18sGIb5NuQ0mFzOYoh6SeVMKPyet133p6RUDXlyCb3sOTDMcA3/jBuKg+9
UGw9uDQFANCl/qfssGegnA6FTWiA/tG6O5c1dpySCRO0xI7+v9xO772i/CVMZ/y+
jyNn1iriF+gPnIFPBqrSCPCgSAWZYlJzz3m0vNekFDoqFUOjdTFGUirj7PSFzFFg
keAHuIzNOkOt14ZGblWKUVOnF/ymUmYu8CP8LHueilqqvEUQ2ULhdQxAXP0ZanQp
R2lpeC2zNjjTaQmvYeeIvnxpmfifE0/TFANckLKn6zHligyNKkNv/ybkPusgXFYI
dd0ks1ZAVFqggii7eY89Iprq/J13KiEQHuG194L30lYvTY/nZ06Y+96YaYt9m60a
frVMVhaYYyiKG0b8nLr1gVjApFNGiFk2AeCWSRW1CnBFCJRsCgc0ekmvergA0lMy
jRrfVbeF38/wLyxyUStakP7DznQHT1sC3ISEq5U5ZtMze5dpYB2Y6fuc7V7rsV2M
YShlQuklwqXXMxHtWl162cP3NtqcmxcnTnmreaCAgQgVc0YWA+chuVCQOIiKYGgL
/9DdThXK9vEcmUSaTWiv7B+Eh4lv4X+U+Br03wmyE0wn9m2i+5cvLP1Zy6WRPgsL
wJXvLyam9Cq7aEB5WbjcJzQfqlLOXzYexucwEl78ZtpstlmlZQQSu0yLf97wl/qg
WU8W/AxAmP96+2G2kUrOtAV/cZAIrxJHo6ULffP2+m31UD9bVtMZX8br1s/dWzmq
okjIL+zsL4X43ETNiErwQWyUJEZIca+IqSAgYMGIolt+fmI51l13vvDOWmhXIWYZ
Sic3LVvXdt2+Xf7sCK2Bh7eEfZyNzeQPuFQvUZEH4bgTVWWP8wxNAO1ajU+HkpDo
G+ZGXUHT+762Wc16Ok4wgFtoNY8W/yNIlAMx2bhUkH5lSy7xMcaDvfZFdRMVgnyI
unKJxu1NhrFRlOPhdLtyMpFOcTCwRQn+XpdTEitt9vUucFB9HcjYaZy/AnSm4xab
w6oFS79GJK6eEWuE+ZMW0CUW/2LPdKjon72As2DWxqu/ki6R2cquoH3AoVTjkfoG
a10Dq3vAXZPRF5ZK6xwRIylewqKt+E8+USkgO/s2N4GoM40ZVDekkdLBc0SZ9Mvr
KO7gLd7UOdNUIj6wOPOJ2xHk+vRLnzN+CgijEcfx5qZithspP6dMP+ZB9sc1Ifov
G7c4G81cRBgIW4vty4pqDGzAfW0Jj1MdnPzTq6H3cso07ylBR/kgc1DL4mOGOzrI
JCEVGlwJk8GJwCYZOmur1WMC6BsU80tVEvwLG71T+4OqT4o1ANdySJYVVfkr/xR2
yctwz5UDxXR234yZbWsW776v8U7BolOuFoSQsSxCzH60CRaECUBu13LIlsHvxxdh
rTDAIWVFK4RsOCRnZI1PgNQ8ai9yXX9RdcfYr0DtDJ3SFn7W1+VsAWc8gryM+ZSQ
/AL3dueqfMNsEWKAVia9l4g8Iev2F7Y/S9QK0tC1Xz38kFOsFiBwN1kxjd+buPOZ
vlWwj9xv4T5p2tx62GAXVZ7A6Jmu5XjjRZhx8L4F69+dnd38/3i+uEe2iZwWAXcm
591rXYKtk/y80v4qMqHPsx6qeOUi6jIZ0Zercw6JCDPj08XFw5oPK4pdGRpRl9Tf
IhZnWs1TahtYVeSXquG+42JOqswLj1tShLW4mt1/tjUfjsGkI/2xUtzTw389CUzA
8SfSceB1Q037q1G4aFOwaTGEyNvr0JhMcLSktZdF5QsnEo34PoHOF/DCzqe4D5D7
r5OM7hc9nKolPF062zNM6SiZJ3gofgIuEiYxIekuNFI/93PhEHbOEKeoxkrgvjWd
CcGFLa8ePY8uXQGRHSo8d/MBjOn+PJrF//Mr/sGVBv9rD5TFfzJ49tYStpxjA0Sv
MAkdYcadQXYrwpMsK8xvoDDDb3/jvivcjjGOyBYz0FYkGtx8p3XnxgFabUu4xZVS
m1ku1Xz+7zLG1PwG7HXn0Kfssi7AArilG2ygPdjs0c0+HS6vo3FOj6Frm/EHJ4Fd
JEwcwXqdBEi/QgR88bsGfpKS3KkFPu0JAqhGzIevxzLyeYsRr4pebhLuccVvFvGl
CR2n9hxL3xk9nk/dz23quoNMLxzsbwnZfGiwN03f2jgc7GxjIWz/YiJJjktNxuLk
NborK/kg8D7RCyiZOROY7DaUFXytCdHKKwXKqecFEgRabfIJC1LUNv68tFhMlofT
j7x5pv3R/5V26hR7odb/mEJtMbBb0ONAaJdUACg0vZ6Yo2HZZQmTvdW9cr2/qjo+
Zov0X11AYHKyAAcRLc6UuHIrJwPuyw/u5x+wdicEDf+EBKUbAP9BeTnSfnv3nmkc
vBIzfev2fIlQhHYKcc/RUX2S0lMae6rwQSATFKPysn1uzcBBQzbzOqvK5aHzPa6b
9CiNTGAVo58TaelTDGj2rVEP1M05p83v2DtSTMaZ6aA5tT0s0I4ZxAvy3ngUeTIg
yifcaMTMHrXiBx9V7aFRImz1PZRj7UxETkKr1r17dfGaxv+ndLXQP0y23nycuQTG
BTESR2vbd+YpHzFRM57dynOE5sOzEnpj1ZN8DMKmnJWn29X26I1co/IGIowUv/qb
ptCJUFxOj6C2snkb0lHYup14fXmgYpWSSxOIJNn0ozeuWriqgsLGBaF/upFOgzch
oPyagXRNQckbYrXRsJbzKgkYofrcgJqDvkJkH1DVk+LuzDYMWCmAfooqH42J1ipD
8VejEr3lLcemgd0LKuACrGTi+apyWPyFj8MWPm8+hql4yX3cLkDCDLjV+GVFHn//
r5z2ujkGoeetWh50MSjC+WNkf43ZxdkhSl3769fec4snGK97DPnjvHBcP2JVD7NL
0a/tsUFl+eco74JV//04lHtv15wRcC0RB4joqTsKJVwVUd4JCeYrbtmfxe+V/htn
lzjuJOxkr9pONHvPZsAMSmuYbhJWupZaL7rdU6FLHUtWjfGroAE+I9X23Xo7A88p
cYWFd1kAV5DySKBbyK80OsBIXufsOqmCj2HuYPHmha0LdAoBsPL1biUtQPg7GDLg
QggygZRaM84avAtWS97+XTJkHSVIPRdk16RJeL/fTopHX55gemvK8nHmvk679C1C
/O3HXfYn9JPEb2WuDg1DK0FaWVjgdwRi9wJJUszEElsBPEI816Cd3iKZO7ye3iJE
cvIY9rrV9GcBNMkYC6N4YIc+t1IoxqUpRi+M4c2lixO4R7Jw66oe22oCGFvZHwgO
5pspEgCNpDAvP2DrVmH8Ls8k0xq7NLgqxFoF1k5By2zWIzsdj4+sQ9TtlLRVCjPM
MYwrA3DCcvpi+R445Z9FyvBN1aVjhpADuaZROHP44GmlH3GB/CxoLpE+ZxLXFUm4
Spfl0PhubQk9VuaeQftx/g7Na2eygsh5Icz3wW787BxNp7Ivao/6zhd5CBbpgEcC
mrHjux0hiuvD8JzdWaaU5Nb/lfdl539Ys3BVAWBf1YftPVgF7+fRF8JzX2zDGuqM
vMDXASGGTo1yIw/HJRe3asp98mdGqRHPI7jkLnWOvSVSmoZJEgzixs1/sEJQMaCQ
b4R4xk6poh1gaPj2avuSL/S5rxGSI4Lm7IrPtQQC2MzA/WDUwDfhQdoWkWcHxBhk
cC9qIUQTVLwHBrZ8QUVoRc9VIcviwYYWnjtRP7mCuagkhv/OQvSQzN5PtVE4fal7
/vGCuV1vOYJTUrdZyjnzBv+IR34/j2j2YpZLFJeDuCDxsPc0o1S8PK0xmq2Tvvx+
knkMXkFUFW+IEhtlV2sXMdg1zp/S6XnUkvyeONhWwu5s06sTmBKosGGGSnQfDyPw
8+AHXN9fwfxS9Zd1CTSztZq7tEVCw5kZ4MNf2XhSYEH1sleWYxyJn9HMUtW+2lM3
sSrDXUOeIF3hk9lJHTo83vnjztFEDlvCS/g7BruA4NXMWclORSmsnkuqvAs8vOMy
B3/gIFKNlHZskdk0JcfD8LxhCGhYbvFZB94IzQt5Bk7IJResMBbMD6QAqxmBQU4l
oSiCuky2MZgzaw7xGI+38eXQz/n3hUwINiFWg6yiOj1P6b4Y6pXxq1JrL9t6vRl4
DWOGWHK/g0GstnQXq5pXMGO3GPjLUyovq50EPVg4JO1ijObTfvKnFIUOMyIj3Jfa
cdKeye3jhD6gtDRFVOVFWPjaMub8LkOZnP0EqBpjasLUNrBe2hKUFtLFIpOcRNyJ
9I/OzOrfFVehZqJ2CFZ2/oBkB08PQRKL3eYP6uNEPcHBH5OrmuJjbgP8+OVI9sv0
FrBj0iR/L/U6h0KiqumElxU97HhBlWTViq+sn2fnfjth2JeFODFcexRuUyVrVpZ+
HM5y9SPP8QBnhuQTmYPEZgml2zHqczf5zjCutbHcSHEiVDiVsR3pcwdIWfhlvICD
MqY3xDRlrCyvK/NqX4Q+povBd0LUdfHpGu7h6Yu8be1ZwGjnisJoo+UvmTufiIHw
wnXqVaJnhmSSlwQh4T29pWmbfLvSj6B7BueCavx4/cfe6CUThaEbIig2n8r7mdmt
i9mw8D0aqVXMRG551KsOHHm0OeMNXUBSmcJjPw70qoNCbjswqL+U6E7OwRs82Lvo
ZqjOCFvUzp9f5eZCLUooCobgt6yTuaH1Z9Y/3ZztDvNhmXaM+1pzOP04YHX9zzXO
RmrKO3k99lH2CSM+tX1R3SJSkt4pFl+a+GhOTGZ+QQBEqz0XADXbx5+FrDkwH5V2
lV01TxqRsCaYnBtDy24djurMHklR6EHu8xLKzbi7Uz1fO8903jrfSJ/R4ZOF04c8
4488yFmaZoDh7JICoWr6hvrnZCKFAVlVEirWC/wInyTtulMfNcEzKKG2WDwMU+fT
A0Eso8zrQZbQ6nN1LxZZsVtflmUuUtGdVR9t59RG5Sr2tzDBwKjz9zAhBK9WgZU8
HPKgtajgCg/z8BNhkuE7zBM53iya0RKRqGWtk+qJrhFbUbBapyUpwlXdI6ZY+/Yl
D69BWNP7Y3M9sMBgLC6RVptT4dcx8VnM9AfW/R5SFFWWBaXkAK9IH26bmx4N9A4s
g9f/EPakcR/t+nxJnjBpZJ8rH8h52nOE2tJ5yXLMSqLyx0Avh9FNDylm3oayO3oZ
8FFriq9Fds9Op9UvtNJFCWncOvfHtW3FSw8nRHbazEhp2R1lWJhclbInPY1d2f+A
a1r/NFHysSY8mDcqx/8FoxAJFLNi7X1qPZwXd4rW4+NN3xovhuFMwGJ8pAlLpZDV
YTIa9ZpF5bGrGjv+JvoWKHQVMzkS111/ZW83KplvY8UIVt7m8jRLPMaG6lsyEKg+
aa1CZltqvSvDIcMcLyHtR9Xo/gB4TcDh1zDVMvxfmWJXHs7gI5JHa2CWXhI421il
dqgb5zF7uNpgGVvHFb+p+7Jh93ovHm2oID+dxRCwmyQlckRgdJqKpCYRJk8viXcJ
eXeNxgMoiVqXRa85KcXNBOuJ0luqlJKOjIMuq48Lg2f/FJfjqB5RdycDTGIZ174W
Oc3OZ6AM3IF4h0g8JyueZf9OM1DYvjEAJ06IS2xNHaXwmlcVY6iGVgVd5qJHxeWs
6O5EAhSzMmz06kRok1bD72oKDX6V8lvAPgREZllD5CIEOZ4QdqhE+P1JMe9fivo6
pgGcR+KN8lnhT+taODwQGGdZrhTENaIYFNsw9/Am3r9RTR+F3w59q9jG0bvegwpe
rLBkLTJESV/HCZtEYCuJ3OAyBYQZ/G5skWIm4i0ZB9NzDQ8zO11oxoE7lDi6aReg
O8lf/acV5/88/iOZwHQnKHoFLz9k1hZhVmlRHEX7h9ZlPCifLpC2I7+t8OZon7Gi
jFN7h507IoL6VrjUJRjbg4sl3azxIBf8j+vk3wuGNr6N3Rs25LbVjMxS4H9Z7kT0
GnMYyu0+xPhejFd6NVKpzgxITEnzAkLOhpp/J5IkGcpFQOpK8TmKD9sqBFIYO6zj
9wI5WCYfYOSg61AX40NMwK5RPJT7JeTuuY8hmcbH4MtHx0xyXFr+meEQn6SMOAjs
pThtlYP9Wvt5lff1n7OuvJC1Dk7pxqa05aQJ0cw/40NBChvusQVpzLiF2xNzV929
fm72bvnEQjvIOBA8IuF8PBDvr3h9CJ8/D9QR6dFuIUVd02RSRoj5MwcEsQ0Ek5Q7
dI9drGEZEU96z3t+hqRTPyOsOT6i6ZnJbMtCr2pFv/uRM+k1bDQIpaSxz5BOYt7v
ZX2HHzkLoyRDPswk3f/3lfXAfDILGmsB7Xx7FanTxyiXEsYC0lKEc+7K8U87Ja9Y
N+YEe9IuxxMpfut2aHBxImLMxBDsV8GFsqEMFSIAxBenIJwV/7J/zHD8qBTycJ6Y
8W5Lv9lCrSvfD5pFkVqFzYNxeS7hwFpAUwnwMlHbALfO2kyOvGk97t+nw+Mauuh+
K7PdnRY0aCsugfJ7MNqlGGMEAg7mr8FnDKYZ/aAlr0+Hh/lWAEWSJv/Q86WEewQb
jUiWwl9g0sFkhIZYuQV2F2WesmqQUEn32KD4Skeplh6flMpw12Kqet9mF+3jOcvO
AWvCmpa75WfjjqaCfuG8L8eLqP5VxQuyeXW/adqo354wvNObl1Obs7p0wlPaNlI7
lMWiQ3yYV96IKFE1ypCQrmBmJbsr2XHakPHoUNmFlgH/Ei/YwzQv2ETTKOJ204B/
l0bGYlWDu3hte8xQSrlTMpZHsvPfzplS57EXp5zqdlL/atbtkKc+PIEB9EExeYzP
d+aUcLFT5G9zCMEHSkTXnL2I0/AjpEyyhGcSZTUQPmdyMwP6ibHXLT0fJi97baqh
p7stYcTvtpSA2O2scq6a8WeebA3NxppiffPvc/rnO6p2QTh3UueR7TxNJFes4ILq
odUdtW93A0YFQoakhroHMUJeplW6p0e9b/pnkUVPkn7ri/qRPXWXQFitm1iJOeGi
iFAUPduPVAheVOcqXP2dAFQ55feti7fkAlKz+1tjKmEqrryC96XeDSFvZ0j8V/Z2
6dIgvnbkdVI5eZQQCW9LTGbopphbOk0QNZoxKwdAKpZxa44s6uhwFTlka7iH9fX/
FXLxilOWLr4ndUFDLE3bpk7waOi/rraKVtl00BMSqOkbv3z978iDwI2yiS3G7yYt
Pg6E8xoIP0ScMqu3L8FJXueStsiZv7SGDAb4Z1T8gqe3FAh/02iHLNMP5A8nYc0f
0a6H3svt3zuav4aaqzR7XPMh/B+hBTDFyi0IxPmWxFvYo26rGuCks0iFcMcuahp6
h8vHTGG86UcppGJx5rUyv8zo82/MOMAyoPJGoN02+UMPN4bi389K4gjj/L3ASZSD
/+zYQ8VFEn8zb4ejO8chSuN8N0OoqT9Fe23Tvhlg2pY/RbOu9fXceqNZJqi75PNb
RcXzI1Ba4qEblPKUJrt7NAFVlktRPqjnmvT1OwM4g0XOfcEVaD4DJ7KVNEfnTPHG
Qej/9YhRjy3B5mPpAHkhgvZttWwVxSWF1tFd+gYGwkSMap7xVU7nvlLSJH/nfLdc
zjAbZKCIvNGGsBUeSCETCJ4Fo8NI7yrN8MasXaEE1SHokxEJKpFOVgFW+ae6Og6u
f9HWzStnoCWe1es4p7o6rUmexB8VuZn79o8Xr29Nk5ydzp1nL3TNtHbNUm4I3kFK
2YYYfxaFRapHvXS2Sko0d9o8Dg/wTF1juJTYciP4c/p1CYuL/breakdvg0P28Mcy
4E0yxKDOMziL80CsLJ26DBF3YZONu8J7UbcpgeDCfl3vJHAgGDGL1BW+/hdKJINm
+tAfG1pTLvMW72lXWAvA3+I/FrQ9HZpGhB9/0czmBuJ96xJIIPlmOk+QlqPYJk2x
b1UW9se+FmdLibKKOsJ4+u/L8EDvhTa2tRePl4f3ZINGw6SBxi76RvBFANNyyPnr
sqxtyg5Z6kbgwvbmA5sc4ErgAjQVnsNHsLIQKF7muu5pf3qrFXyKU2Zj/bElzi2f
8jQ2O6FXDn+Ecx9Q8wNCWaA8znODJkdbswfLwo7clv1xpT/oY52mDYWnvJ+6YbYS
l6plKWeS+bS0fbFu4s8XouvtIoZaWG0BBglQ18J3rkqmV4Qe3ZCF+E3QmkWqIM6J
AXNYcFJfEvaC3mkeKiv/NHAdmyPyNfdnm2MTC9jks+LDzPyV0p6CY4Xhgxz94Qfx
lf896wTEhBa9u2lftDGCgmLnNfS7YA8kMGRZ5bgPeb1rzkAuqH7rU5tE7uLrlqBF
4nN7nNN5MEgWZpnTPpkFKSvABqQahAKSV0/Sz3xLzxs4wzuKRSPxncjrdNh8+uN3
9BzGg7MV1pnyatZB8o0RVZIbq2KwPeX+o7JeAV0DjFvpJ98/KbHfSR9ZWSTiEuNt
tE8Nt8cYvWq7Oawkju/8LB+ego8aapVlaX5RiTZxPf4KUJycClGMc4NMQkVPBiCP
YAjfD+u0oXiYLj5ipOVnDqdBpMgoUU/n6pgZM1g2VXwb/jmSv7PLU3aul0Pfwpmy
gKCQ4rRhWn5Dk+T+fFs5VMw6dmxdJ/55ekmyGtVfwcykPn+a/wyZdNSjXBLviaE7
HFV9xETDD+/7LdnTlTWDgw+Kta5I4wJRtXu1fWcimTsnM01cNadOfCrgb0iYHUzh
2a1KIaWU//Q4NdQZ3SvSYCzR+6EbbFtXKh1EnjRQD3iiUAKB4B4AKL2zDnHk5Fwy
bodl9KN0ldvWmQmKwrZCTsx3UMbmI2J8ar7BMnJ6+XEJu90oZ57CooDYWP8P/ikg
OvDkVAuJXwm8/waN22iRui+UzSVL6Sy1mj+H0NM3Uw/sTVsnTzv3bEoQnD7K3t1G
rPH9TsOy0Y2dNVPWEcBOaofTtegTHd24RbbXRI6pVD7iSqQHkcyzsbWe7bZEA+hP
A6qLJERx54sI+3P6tGm8E7tToM3gWGjSBHrXWSRlCHk0Ef2jydWlX9U0r0+PDNlD
E1tFt8csekkaO247gMJICpoE6wry+9J4n6FxEsh73nPdXgVmx91JQfpXUpujwY1k
3ZV+m+e+FU24rMkupcJKHge7JYQ++RQc5OeMTRc50FW+cGr/1E3B2faqEnxDuS0H
StOWQposyykMX9Mc3Y0Uax87iGUVbsEoCRdUBhoQq0YfeF4Lq0Oc61gupMcQWJe0
auXk6TKXRC8CXjVqVLIYRqkNmeiR/pYweTDmOkhvmIPHfW8t8qmyePKRAm2gVh29
s7qUDyCarpfUaP6gLx/AntLdhI85A6KAGU65PP0oI6SzlZBBOdnQ5tzSQ/uuIjzK
X0FeOwArfIn2x6qfk3DOz6FZkdyfpqfM+qsZtBWcQMiXB46fWhdgUofkCiKGnpz+
ExIuO5sq8AC7Ebc9ow+abZ7lF2ydzz9+B9OgE+fyDmvnsv5DcTfkT2qcjkS5pq8t
Etj5qzk+Fnwo23m24k/LYaULay/l3vBvsgSnkes9FQ1X/86YxyIXWPheufAxUbYb
TpxSvoNEJsiT59ZtWylxOIJjdlke6MgKC7KRgQgc3Y1wbmuSsoL8QRTXWQh/cfON
YqIeCNArT6jKMEcMqM9Wu/HMxYeDWoLBHGXhu37+3bUVO7vTtmH07HQZUtffbFRR
Am3pLFzElaeuJ17kGCz6ZM+lCWYDIC/NldD8l+FVYtEHWZMqth00GRoMgLn7ObdV
Olqiui114juQvSt25F5SWiBxA4qqeHyLg2JH4qi7xP1+NwonQSFNgRthSvEazUgH
6dOjnDZabUHpwKiJz3wn1bAeDi7WA86hVDMpNPOm8qAhmPTLr7bNkBanol4RkOEd
yAXZohMbhkoWLeMwK7nS7wJKQV04NXVzgES2UVbY/1hpQWTiQoEOyg4PS5zeqITK
3quJwfWHzFhnv5LqtFY0t8Ioowd71N50eunRaH5a2GkTZj86FYN9Oe6cg1yVo4U6
IB9roqjR34O36Z5PSxCPXCY4N2942a9D8iaI5QEukH4sMn9bunwe+KpFi7jDsonA
5Cp5syGpqxN1B0uOPEM9PJyTCqlmUN9fLqUBsSFhx9VxoJ1djvnievGEBv1pj9R9
8BhOjOmRS+ayNArRdFe7k5QVPG7uONuUK6m9MxHw+nYXclPBWo1OPkz+KIKD9cVa
0K7cKHWaakf5Otbqw0Woe/WxLzPt+qEmZkRSA2LV2G17TunRPohQzj2wgXdczpWU
IcGCAxFU/GxzeZRnNdppT2PqFb+LYLc4r5rbKzVetEbZX1gCpgMwlLEogDnQnd9T
W6vlopRKFQVKdQDeBsJ8KyUo9ex/UuFMnc3KOzgUOXhrDj5qgPtgKy7Uu3dFlZ3m
36ZvX531QqL1aYf172KoVNaqte1tle+qyicRXincA5ZKgxHhT9L1gDuT2Si1lMdu
uiP8qBtvFlGa6tEqCnW5nrNBadO5MVi7/IHYUQsazuBfIjPdtTVTJPWJdarTeUZy
Sxk5M9JHp3RMO/QI+1/bFE7guj3LysnuiE+MLQvpoPd962YByMvZpe/Ka8P23KUh
nQrT/dne+c6aoB3kvxu35z+PMtdPjRrYMRbekjXd/whHe+g+mlkXbFtDoy9swj6n
ag84ThmEMfaTBMYUHOJPuwPrzOfYMCQT9GTuxXYfoPloGaK+bxYjlNquS+R0HaDy
dMLav7X2Z2irLpnGMUEDn/OS6oSTofQDo47Z375yN1XdXKuB+LdNMnnUVfqvY8eI
4Kr1PjtspUZa41uvDj0Wk1wLgFWs8smUrxizFAKG78nQwEU3pgRAYhlI54pDqGnn
BMHspVj707GheAfQ0neHA+FIKlCXwld71uxiVRWms1DGBMag5I2S7deDYlkPvlBR
7prmnTcuMm0lYAeUYtbeaDbSj6UTekmMZo0GPpYYduPElz5Rsm4bLp6sG/UJNbfV
8wj/0KEYXuhArTgamnnc6FwXeSlBalLFF6wXkcktbqnaxw8NrxXHGLHu1ueUCIO2
YVtc5wRdC9zygof1DTvNNsS5iXwV3mPYDpJLPtd8AchH63jKaX4avE6N2p4WlOwF
EwBcg9ZfiAd+LgquvfKiwWHDUpLf8PISHtaCcOgQzQ4dF0n+2CRaRJqK9Y0PfT2x
32+dYpdIg/2PrcRxlRYPncahMygXpwoytl0caogRfXTqy5vcBM9q3ApUulNTDUxQ
eqRtLeIdTT9yFi78y32Hciq4isdmxIMFHqyTnhVZaaL5UqcZisLwrEL5I3zTbRzp
wN9s7CL0splyXfxpQs5cRk52xi2NMQD/9i2vGYmbZ5VT8foxOoOpTiZC4V5eChaJ
rJUZq1uc6AK/uI8MCF3tc0Fa5gyzC9F1ETCJE9SHMNBDJ8kkquNTHQOtHDC4XOgu
vS8Tgq5LVlqOMeYvJJVc9K9pVa8JTuCJKQiMYnHpwTrl5toZo7KiTlMDKmkBabES
z96Vk/+jEiWtgRLfo0CLhmPmu9uE5F03UaxHGmGpk33+tced0zT9KLbYZbNrEW3/
DdDvOE7xhSuHJz1Tj+PwExoGE/s9GzscanjyQbSOxbpaJ8KzQmivmlj3i/STR7Xm
CAkV5ok8NP99HFWfO+8bbnChJ+N+EzfyrVPuYGSYXOs4lquEAKa2FUCw0MaVv0Zr
pb5tiq4+ceZ9htQ/iOnxy9MXTnz3OuHB6u6xOTgnxLXzVzcDBhi7PEwjwX9Ix5rb
FSZlBMF6D8CJzOogEFRIRMqgbeFlxYZw4Fkxb5lb2ZNErQbC6IjIJysP9jUtBwTe
RKuhgli5c9IRRsPAs/gSC7lz7cLQHsLAjv/maHwOBBCGYFG631m89W1I/rITfVM4
zEWJLfCiETNPB2k25Wm9auJkwlhHao8Xk9iUoLl6uxn8GJVId8FKczqmrXVwUNM+
yn6zrnQAmMOstr6DQB6B+GiRv6IenZQjxJwmgBZYZDVeTcNTBW541fW/mlV4112k
PeyhsVObVNYdlt8oAJyrAlIwMSqqaI8NrLzOEzZxuLJdfEJUGt8p8hKZ+71pPvlf
vP5NvdWZgX1pP+6IPrg90Icn/H9sycJOOiOcxzsZF7BQNI/ECswbpbbV3j+Qx8Dy
lGEQBbjXgaX55X2OcIC7MwBonAZQr/aX8FB9+swOCBhNI/RA0bmcbRc4Jf1b/sh/
oqZxNNLrTztDOBMUaBkJ1U4U0+lVj1DHpjkakgV+EMIx3aU0gSZjUrrO4QSXclHd
OopHteT0XuhvO5133+t95jIN0+i5PPDPUtDjb9zp6OftiOcDE9oLaNkyp/C4PhGi
ITvSesMIMI+m4mgUS2PcPsirlH2jfcHrcmVgyGlcCeY6MCh8HqTY1Cw3pYLKR3cV
bwxXaMRKxrnPbp0notzm2vuhLCodZFm1suiiif9iWrzotOjoVfF5vPOxDDnjKcju
wKCi6VAzcBOtJUGQF4MbLBlvupjGE5twjpEqH4LpGTY6pdg0tA9kEO6rJrStiU8s
hfWsUNwOVgSrygRz9bNs1nUuvslhesLnvC2WVUO0SvHCH6fdPWVD3VGZkEZDqMZr
9oSMgkWvd/NZkmJ/SDk6ncKK57pQeK5VsqmKmSQGQnJQLUbsmWmTeaq0q/czVtPw
AOKtEZJCJLElqHZ4kOaP1NKupxTH1XUfbBkUkwArFVOvFJ+0GuiUBeX4QPWXgeiL
5OdPhvf7ssYxR3gybMF5ZSz4xxKp1dhSVLcDAcPZCrnREjFOTXFIhhjC4/2/tdpb
huiTW9OsYv2KyWRxFYts+JqkUxHxNNkCAWRlyCRg7oG/LMMost4SAPl0OMfrNFy1
YJfIzIaGFDU1nKuPcr3HtN0hVyoyYGrvqKrX6xGJXiJsRi7KiDFdxcSnE46u5s+0
O0TRWgoN5yLGT1svgo2OFIOA0rE4nXDTEFXoBIN/69R6dAxDHkZkTl3R38VtVj/S
NZwj0oBkWgJd/IJT7ww5pEuUPlqvs+frcHAyRTSjOMsVDpSBRsXWuwt+B9f+Kc8e
rn2Aa31opaCOc3xNsAj/llfiYyIfWCz90+lgvdGDYQwZABgDBDhpbVnLTtSJPj+C
97cAxBkCFofcnyB6CJV/7v5sA8iX+W+YG04h88iMQYs56+9qzuWjqvtv+7qxT3kC
ODn5GeyOLYF3ukvrSvGy+uq/MENoUTYP9nMM6eBTa1oduLG7VMl2MqLCGWiOr0dZ
9k83HiCtT4Y6PcsIc5E6jhLT9V+TmDYURpaeLE5RZQChBTGUpFCSAuYQxyK/Bpex
jKYzYBnyvrAkspYHKHvc1j4QnrBN6euOz38HbZ+1BHOmUisu9aoT6IQZEZOddwve
Nr4yLQGspXkmzzjHAz7AYcmD/aLS7xU1jVQKKoQEimTeZRRBhTesTR+hIwKHDHMg
EHHm/n0/o7tCbwZ6+dAPbdvZJWe0xal6nANApWqodRnyLgfGaanyX0YP3HZn7SaY
hbD2eejziq252QJ8jq7ruDVZLZZljDDgEwAsONipuxRzFr7r9zt8bSwQNeWLKh7R
r/ggr8scApk699L12SzB0mbgBu0krF+9zT6HZw+Gmacd/Nx9tH4muGZ2LejTAfh7
xaC16lRFw7QqDeFi4VxW4ZeA9OElOHhIUWUrkrAHkz0xL71KUYdrMlltjnPeaYHC
sjlRoGhdlJeVY4N7XGRUgdRzWR3ax8wsLz75DtC7lIaVodEC+rlDJE8wNak927S2
k52IElRQjUZZ9oHfNdi+8ko2clxXoMU8cGY5cqJk5eNSqW1V7lKEunwyQjdsSxmV
k27+xuJ7/d8+VacMtGXPK+RhVPzNfoTyXVFWdsI+Y/Hfy62i7xGyl/bC4X/7svMv
YXnmFrlbqybF+En6pUlR4zYyDRmZv4RlriTJydDNBURPj++fP221qIxJc16SdS98
FNT/UkbQxaO1/NZ9lQ4mPUVeZqkjGMQbgazfCz02qIMMzGNRCASJC9jN6diOkPdS
9DrgO3hwqHeLPFOK7dR1wf1Ii/BiGroUNYfy/TIisa8FflevtQbL9wQyz9Y7kMDc
2wlDs4RD3txNbydx8mgliHupv08X8BU9iCm/3o7SmjRySoeJEabIv5ioBdg2cFac
G7q56+GbQb6QbdMO8X+Ao1pxiutp1617x0PUhs5KTXPel3HKGrinNaKMrmPWn2JO
5mkMxQxoPoou6N29QrvkywRW8i6TLz0VRNevxvZUlW0neY1nY1jjsfPtF5rxy7aK
rgDt6lTNbIIpgmwm3IxWMT2C5H2dkUvIqjInCl9KWhjKrrOXBpAKlKycyH54x3aY
bvhnv3yBlM2waFkeN4yp1DmJsBm7qY4alD61Fe30cecSb+rZbzJ8SDQBznPQXFFh
/+JntYlLyaSMYMyOVXnL05j8tNz5MbMR59o87rIzQtznNBARvf69Ge9io65/AIWA
y9tNJmWPT3McjHVA+KqfscH2K6fMOltDEp5URYZT2H0frjMqKgoVyd4w3KEymLZ7
5e0Mtsjy7smIgDjrTSRzqlp4dByXqIc0Yd/IbvUnbngdeQ9xLxeIGlG1m2vJ5bgL
/K9SzGt2czpLf9bRljBBjCeYJLYSDAPrm6SwUc93jm6qkZY6rfOMd/J9Wyhsc8DT
lRYI+u0HbjlM5rSz/ADy7wHWOxswQMKAjLEmcTlCgz+rNGdSNzn2O7I68TfoAfWB
+QL6Y6ngw9uVFBwA2gq6p/Nub7/bNXTYjEmZb74/ttxNM7dqhaFtmNJ05qat8ped
paXUpTIfnX8cPcTTFYQax2frfnTIBEcHmuFOqgRnT/blJLbI1iPUfOdRVH85THsM
tKBSlWOuGRmrB51N3Pnfo4zKL74NC3UVV91v0PgwW+BK1iLqaPYApzB8VYQKizwd
KVby2B5YcyCNUX5g9UWb8dcgc7RbXaATveUmeZCcDt0g0MfT0HyoTELGsSMbTOTH
ZVaeB74CtKEnFYNcC+YGsEd2d3qIvz+c3+vNBuSJe5B822eBPUbqEOezTfzhi671
ltlQS5lDkMHOohunnrctZUgbZpOLuUa71bUxvRDFeqlJ/dzG86v1G9AMkgQy+5Lp
rNSG7iMaF017wBpdnDFq2/BYDoH0lXWFgSUYS7n8vY1QzLW0rZdUhzyYnuGPmXIa
/FHm92O2Gos8K1utUgKvB+bsRNYxjGNYT2D6r1zjIRBfkJ5ql/GpWcauN/OmCMAi
CcaRDm/cQ6CV6BT6swPvjocus5DrJKztBvdrQWYR2sOhOXBaYf3QdySwgetPzSYr
fxxipTkUQOX33wc6WvEUNaMkPbk18k1YtHTyHbp2JrrcwRHKcb0dWV0PFqA8lUzD
isbFtyqvV8BMBSl4ChoEgiTlPZrpUydgF/17BWlYcp+xXUSA9A1AaPEfCrnQNmtQ
2mC5TYaCDZQGzHz+MiDTS2kk5NBcpk5Uw4zWKb4d5oGDYNIxieYWc3l6nCgfMYTc
lTFYi+t/nRVBlXhzwd9wglaA5XiEj98Ne7AaFSWhIKUBCm3Q09kLxWO62CQIyquO
yIPkC6j1tvlKYwvho8VjkJJSR2MVRxWPVZs8WPpePVkhGEgBL4jVumZfLTkB3Kqf
38M+FjdD+mmZ6hs09tj418Aqq3JsP3We+lYI4/iVHQK+eBKYynmlv9RCi2efp2v3
FH6ujBDlIvD25s7u14Zg0i9LLDRh1CzeOUYVr1frUc5zLNQ1meitbPbQAJO7wclh
N2rwdPiZL/vlDqgMmQ1z0GlnMHuKa6Sx9f/fHSwE8A0ri0S2OxMiZkPw/udjfzgX
ZTZgHC6MznP/RmB4KC1gdf3ARTfdQw4+l0MY2zzrcZAKBzv/DSsmxGX5+Qmkf0h0
SRwY9inYKzrsMUKec5MwyELNZj+GhNCTeeisF7PQ1aXxnEMw39orBOOC4eYtCEbZ
6P4SQN/YQUfx+WpBpcXvGqtKALJPngsT96Za9sKmD48SX3ZZeHz2pcTyq7flsrwT
Pc8TgdAEFsJQtDVnm0mYOq5InF6PJt3Zf0agTi/7UZA8nCaPFF0pJYHmFEakdo5T
uJi9ssC1a39woiq1G0tL6JM6KsuhqL+xF131JcOh4fKFFJLOJbevq1tLYplVEN0w
KL//R1F504u2OGyhc1X/VcndWQqf0R8dwiOZJJ7Hrh3bZgcCK5hbGLZwAr6ELz81
OapU4AJHa5dVJblQHI4WH09nuBLyVlChyqkRvYm8k8g1fZoOh7EFTfIUtlAWvJmc
hOyIU1436+fAdO4szLQMJwwPCfjxq4ec+NSapmexSsxHTURjcMoVF1M8ZLW+U3ye
0evcHgTaXve0qMwksAEw9HkgMkZ5btbok4jMnovRIBf2mWrDiYjQuizWfZ/uLNBw
hq//SfyfqciCGRINA+1QfSk9ygCS2X7XvO1tAzYJzhcVuxs+klheV3Icn4qDiWeG
UgD4lZTWeWQ4xWlwTjtj/70wPvjzxYTYadKbl+nut1Ewn9neNji+gdrX4io8BR6y
sZKaa2ZJ/ZpfgARyB2zbvG1lRLWtp4AeRs71BGsB/EKKO+HXriTh72gUIKXzARJk
jOeUTNQS0UIRHMb/GgaZzeVpR3mvD9Qj0ICJK5+qEFl5C/8w/cdwlsmh6klrKxEk
UqvDCDGifI0LiE0mIeReaYUIzQMUwnu2Ap2IeOZ1Aq87LclaCj2lbw2L0MWtsmIX
Lr+CZJw+aSgI4XoqN6TFG6WwHFFscT2XlDlhlV06mvSr4zVEn5TJOs54WOa+jdD7
Au1Ztx0bwpwaMWy9GMNjXff9MlAEYvD0cssDGOvkPvuvlcq0R0cHqWrqc2rvLnh9
lJFDPCU6dEZuPNzaglUKcnSHudO/lDIC6f1fUj2qDFxdGU4EDH9dRy0ZfWOMpu45
CFVghVpla3AN3jc4ZjYk9GgtOr2ki+I/WejkYuvdkTlUYCfrl2PmEHkI/1Tt4Zv8
xU1vw9G9HgEUNtuw1nEWNiWThjMq8R4X9NG7JTDarApQYjyfttc+mN5zu3YPooW8
mw8UDf2aEjavBIKooPyM4j9xC2EpEBo2d8VdVUr7daJJ2tKw26XZ+ztiwUMeqO4r
/C/fHUMw+FlOij1FJIvIsK4G3A00I0/hRDhT3NzAbT4NzPPJ2IReg0Wh08/KuGTm
a2EKkgRfOl45Bw9LfHsC9yyIElkBzPNmUyH9otNCpASm0XLVmRPnmhjqyX1DGwaL
laWI6UF4e4vV0WEMTmUD7fphtRbpRNPbVqwyBz05Zl9ibjBQgwBmKaT8hss/USlW
CxCVvDQvGA2oG0pLpB1XkeqAVrl1PE+rUtZ9wcudXQnzg3dQr6DM8Sr1ZA2LlI7i
RnpNh2Zmv5rWSyEy0QNGgA6lkUC2z9k1GwKYQV/2UzeRb6+AvK15TKgGetsH7Hjl
1lZg3d0I4J8GoW5uW3C8Hd7XyOsRVt3Iil0eosfiNC4Sj6l5QKhxEq7IhqPGNDj6
vuXM6OOZZAubeg9r2shjHZfSXu1nUTcow8REbo19tiAIaOF7VPW/Gz6u2Aol2ZfD
7BQYgDliqvihRqJVZXqVtjXDwcIZjYRnJnBBE+zCVgSVoRxw93xG6CVhHBX0yI3p
2SELh2NWJEpYpE6cSzFs//ZVGsizyD9Jw0qjDdW+JBe+GPW5cMXb2NqAjPyHcGKg
B+DqVJEoWFrSvEzsTp39x7VW+dRnpzbgyLZHBNrrthubx/sxFa0oYG602BqKwmj+
A7gjae5VgoNrwBrCVPQnapNaRNc23OGWmc23rIk78whby6ghKghAZWWutY7D1rlF
2h5AQ0jgpivMTWyGjPjvtSTWnpNifhjtjco2NQA+nOLojZLBnJKwQCNyNMRI0+BX
OOnaPHp54fzOn8ne1WRraeJXbMcs7Ywb+J+uKNXANIOXPjGlx50+XbXZIEJikDYH
9+EvV6bsSvr1pS1cz9VHyOghrzooFBYrOkBhQLEvqIhtxLrbNVeaCkbL2b2MaRWt
cDIuo+Nwq0kdqwYnTQhgNBybAhm8k8aeC5gpDck3aKXaj9CTzqRJSgxkeQgcTUKC
hnGW/sd8Yyr08n2lQkF8hXxhBVzjzUgpqfClQEMJUg3llOg8rb7RMgVwxlAVRaL+
HuMQHBI4q5O0zlDPi3d/dNG5irbX//GAwpiwF6LpfNzhCw10EKGVoePCN1YSOGIW
1vfc1hBC6rGtFt50AsCP6n0Ls/j5z9Bl7LvfqsQ4M0uSTh6G+LioRFEQwrDtC+eH
qOFcty1RZNZNRerniaL5tTVJujNUcw2DVLX1Rf+qdtwdOYQ+awvwB0OsKkBO54zm
WFiLsOUvFI65qhwFA6h5oWF6c3FdKjizgigsw8LXb7jzTJnCpRODlZKe+UCX9AAU
gKw65w3SCI/yQTOixStdrYAcxy3n4orBJ55jjSvJY8zHKC6f66f7Iu+PCOajEJ6U
Eo/+YC8XhSALaqc7L8r8kwUlajcUKvpvmOYbcGm3wkBlfjYPZjx7z/MVqPrEpRKd
JlbMV5kwAXVLJxCqb59Gag7bT51sb2/knNwICOkMpTj/EFCJUlTE4b/AyKVs+XFC
+6iraX+0BI+vTZe47Yq5oSqSkSLFKgtqZVspF5rR8hwlJ7SV8nzmXHLM1KSN+bTg
N1tSnRQ1LMqiB1mShnwmB6Run9+EOI9c3TC6XMMK0r4uvAhsVyeh7wMx9OI7miAT
GbTvDzd8vYzGMQPktngPVkmmqe4VEBI84aw0ErJXdjniKq1xkjD7/iOchdDXGtT/
MZFshAurQUqvmrPI1y0JikGFpvc5sxpEX2M0ic+mQtwxq6MwtQIsJtr6+/7plY/r
YhtiFgbz0x6j95nFw0U/UwIqKxLNND0m0eRh9Hoy3xu309xnJyq3Mo/7bZQ0TFZh
f5NqPBrg1ENaSWt4MOUUp9Z3lm4x3VdgFTANHCHFePs1PggWdXcoS5hyDdazwVVU
TPTYqCdUgByLgcoE/cTle1y8WPWfCPgBLSvVNT//Mnov1sCsFdwx80rXbPtmZ5WZ
t3rRm9zKK+SzFzKGTmF5kv5FVRpXLob09FrzrecnJsObYIHNdK/9VAJB+Cwkq/9h
gqqkNpvxnXTami4FfE8p3G1hv3sfL+VRPw7mYAXgVRMWgeKhmjAvqmJTGY+BVCV1
WKNWcE6OroCyqKmz/Kp56fxl5VlLJLj4wxocKf9I1VpOniupK5hxm+vRpEYC6o+B
lNBcaxFMe+4J9/YvPUvC9apAuPwAd7UZy8bF3OjJ9qoRXlpzGrvJ9AX2OURoLwzC
IIRrplfAgHVVl+V4/EMZLpsl6aspimfKk8JoLUK5OCt5VH0K/nh4mkjaFF7TVB4b
7Z9iTxqTyzrFH3pPO+9Dogb8AlZOqsaT6+T7NsH99oQPo1WfPjHS15jxm3K08VYZ
/JAdeRcRpgUj53sKC6ajWeom6+R9VLiwpzysw/+5KeMrzw8yD0Tocl/5FkF7fXDU
XiFzSoiNMWOpZ6h97T76agwuG8f2PSZxbCyjNH2O+Ky0ch72Ut3UpY+DyptTTtKD
3St8iLc2+OBzrIt8ZBr37TX41XnXbsh9lZsha1Y3sTF3ZGi+bGmzfTJfRj5J0qhH
09hwmHFC671QJGt+S/9kUFGiVbr23izx1uSKEXXK0KarFFAP8MAMuW1nAKXDz0HN
4UWc3wgPu4yMtrBgBi7ujO31uPZO4vLtmBGshJ7ByYc36aEXylIUbBs2NXqpDc+R
Pk3ghF7KPZ+efUAOw7FVgctYYkWM8sUtIrWAUho/tTp0hcpqdPaPpMDu7lhtnId7
+UJ7L5vkA6l7lNHzv66LQxz60FyMyBDweq5rncTo0loTA3IC0bNaAPTWf1P1nn+x
YloFYhCsiV+wcMZ0a8FTeDVSiNo0dW6uTUV0Ah6u2aOHpSwc3l4i2YZuK8AV8x49
3c9SLS6ci1BvCie+8eI9L/zECjlo82OzAyvL8NV50/v1u7BHYD9AuuxId6zwX0IP
Wm13SONSEOkHxz3xsDaH6OT8vxENom5+db3F2CtAVv6lQWsrU5RhkYaTr0Dk/jog
RFdRadUhbVfU/hjpdVJXKgoZHb3pc7CLCyV8lv3MNXyjJWqBnUnN3yB37+yU49pv
uANqg6PStnKLeUa695kFDLjegQ6HzQ4qccrpsQaB7mP3nD48ZWI/RM0ICKczFA6G
SXQCnHxYqWzsCJNRFxWN3brRTii7aD80iToeAPFxKMyG41ysh6IZrTK/mBL3WhWg
c4yrnBNtj67h6dDcVJ5+Am1U+wGCeF56BE9brTlqgp0JGQ8wzPivcqSHAGgIDyB2
cTdQ0TWZah5HYMVy8x9kv//a0E3TbXRUlEhdtV4YFyDLOqt50zzrQafn1Ffow+5k
RQla+gxKaU9AJndbFl35ndXnTJkgj/LdpejH2rq/2NHzSd9pBwH9bPfv/pETISou
sJFcc9jU75OpKhVphaFIkFMu3tp8lNNGb2VL/vwuCXNsnVChU2ZCsu2lWqfnmk9O
w5W/AOrZ76Bjg8Q+NlvpglLZWGxu1T2sfXNOM3YJLmoWOvuHAHJ97h71dqctuyMY
YAwU2ULlbU4UJyE6unkckNK8OXaYMg/ezfZCw8ZzZWY6WkfPQc0A/j6u+CZ2U3n9
TrZcaG7sd8pVLP+0XAWJTt+Lb0Dm6JxYQMWp/r3pbmIMiaYfFIt4AaaOatF7WR1Y
I7LH+zEq2YMf/9ZGjaz3JqXk+sJAgHs6GDoTzmdncCc7wRsPTrMbwyrezeFtLka0
EsggqqRw0QrT1XJmkaQdz77ShW9Rc5n34Z7hkO7xIyOL4qZGu+C+eROwlMtdW3Xg
UE9uLgQDdQWWZ81wJQwe6Rbeb7ba7wV/Knb6vYuhofyrVfnUUdnMT+276We3Kdz0
S9yugEsPL0JRuwEqt/NGK2VnLpUWRo2BRrsU90scLUNX7isH7tU5sajDVJcNyn8Z
OuRaMp07eUZzkqNkRfY345NNc1ms6EJVmVuLAZ47jp4UAFMxxJsuULYMgBjE/IC8
2syvk9hWG4uAUN4n+Wcj01bBI54A19SyAltsy8hy2VZRAQve7DFktE4tDXnMns2H
luPxWfyyfgy3X+idBPjNf0ioubS+4h/SCp6gi11Q9bqC7D091FK01Xq+al1/IFUp
r3eWAdEr2tnK5KcBjoAAKb7C1UFQwDPCx7mv/ReKk5MHEJmvS/hwvGBB7KkrvYnz
7Z1dBb8efhRIhFHtjGlwz9pJALM5pFkygnwYyNfJ0DOm7WDr8jdhvxN5KzJTSAXp
T9oMQT/ROLaDDHsfM7LsnbDNe2DP7/YR+ScN8gNHxul/mVRA3eOolhUXUgAGe3yF
kS+Jzjsi/WYYphebYGYM3Nbjk64PSgncCO6vPjxZgnXsYpetF7bXTlDtToaKe22q
jsKGjUdcwwZmibWhQo/9wcm3O4SrkK2mU1Z4GgFKgG78BSTPw6kqNeBj87XeM3GG
fg2q2tEUxEGvcij2y7uNJtVD6m1frtejGH9qJoOdZp/hhSnXn9F/vNkcxeZR2oVV
c23xJR/BrHH/eV1D5+pZvcw4LLrBUcnEB2BXcK5vbhXbREBMXaIz3oEt73Sf/Kx5
QINkonKQK1mhtz2vwIC5g1GL8qfshYFIfubbrcs3aj6IklkyG4GDJ1k15k10PWQv
I52GOeOh6qm7kpdc5UZBPKaDN9Zdgcrk/5llnFqrz9W/0UdD3zk+1wwkFNNIpzFw
BKniFxK1F2/Z1l24KhLqT0gCUpwa2Eo8A5WnwJLOVBosQOlnhNyE723SKQgo3tYu
YATMgnmDkoBwi1KGSsmc92u3qGV9E2CSr4OeIkowz8RvDVY2RzJo8uWYW2CyZFkU
OVsom9cs8Q8eDqq+tmT0+WKTNrOqZh8hltdSZbv9Owmz2qFiPzzRP3XrsrO3ABkK
I1qHtb5DZrti82brzWpsX6oV8dy98/BmQ/apCkfEVKQT3Yw8myZWys637mrXTs2W
nUEVGACLH1iDF4d7G52Yo4x6xJBHWRdStuztFMHhPs67iABtsENH1rK33QijNnst
jjL59Ta31wVwkdNWK/sbOyIyHAwoGMAWvb4fYp6MhRT7VI4Q6QT3Lt6dqQ3bTPXy
MsKHeME1iaEOLjHadI1OKlzHyEFMBYPCNlaCvrn7v9UBChIpjzv/GqTeF53LZVfL
m2/w+ZlgVekOkFDQgSrak8e3boYDNVddiVu+TRUu/5+d48QgftgD+e/nUjyo2cnp
opX6aXv1SQc2wwAfGh3dag6U22JrdWxYCLkP+A+cZCgBJSpygivp7KasK3QigWJ9
nL41oyrnjka8r9gNKtEXAJcsFamADJPt5t6Ut4PKzjysMkgIAC7dfyAFi1DTj9tx
aHaB/SuxyPeynZ2KrnuQNwkP4x1tuq3aV4l9n/tqoETBGWO8hG8SyS+T/HL0mGcC
9Ce2O4ISNU5+W0gBttftI6C+sC2ws+z1XN1VnISvCpJNK8qnUn7kbjXQGcGWhN7q
Lm8tua/wNqTVkg5oUWGQRWV0CiDPwHJwk9qrf2pQfN73UgoWyXK7es+re+ylY612
p8lJaZP5NR1skjoKWBq8qOlKeDdEVxyHncdH104wjkYsodnLBp6sRiZFNa/je2KB
lRAlaetzcwqyHWOCXaWs8it1jEZzBm93AeL7uxLz+P/W4sGNF7ElBzQDVdQ3o8jt
iWQRgkPiDHPhhTyUkubOPYxicIWKmh4j9tinQatrXzlILsgnSz4Z96Q0Echu4N8X
y67RBR2xvBqePlVx8d+kCaEjGHiUEawaOg66gxlzZaa/OlxvNrKSy82axVlxxTLM
QJ5xUhzIOyFJSZSIyfFUz44VWCIARy7J6nIHVCr9c5kY3VsHhKhVBFQzo87vAEMp
BQAhmqRHCd8njZjagGUiiwRTrRFL7opk/UGdtwjoVXUc8QRg/VecYzGdk3HCohKC
j+zbaHDFqgOpC9vJ30t/JCiJOeD6UY/aCQTUvOlx4WcK91kwY5RlkE3kGr0llRJr
Mrn4nmyzwjfLPS1ubtSqdiGBuR0tW4xnNEfiRBoGVM2UaAEVwY4Np2ZgCZpJrg15
kd2miW8tRiHqNXCb+rgbnnLd7fba6OCOsflFhptqBNB5pkInQywpalmSy0aufEcu
uUxSUAZ9ZyibDZtC9mp3cBpl2MghnUk4KrCMk9UoPDMBAfKj6wkGhiBxpv1HP3cD
962B8W16zjVFERyYs47A05ob/mwAXu1tLQmXgnET/ASprdMggw6TeYcN1UhEdmI3
zydTbWnhKaB0OZCLBeuU9pm87aZs0N4L3XnkazRLEl7NXsawK2cQg+Z/uOYiANaB
+k9PXgk/N4w9fyVlXWkcsqOBnMBCqeSUsXxo1vofFl0gHfpI8Ct6f30si7F2Cxhq
LARALblkkWO7xvif/8IGRPU8NoZJiNxjdDWFUr1/4f/yDvXaWHqfRzy0pKRM6IZx
mxq1npTha6eWk2lz1RNjC5j/7qv47dzOPgQqD8HGVtdd8uJo6wzdn9nrQ7sLIRfh
24O6dDz6zXy8yGL3iN1JpJgStALeIVT01dRxZzz/qqc0eV1M/ZrjzSl7CQKhbDZt
DNTnxxHJXrYj7qYq8dEZeYawJbu0cnd/Njy++LUI2TP2cCk+Q77K/pamaFzpNnp3
MB7ITpysjg9zzPhbBAJkYz9PhLVF/VTEz7xX5OQeQ8RrUoz91iY1ysi91H7Y1Mtf
x8rMjYLUBee/7mMzVybmo9LfpdSsoi+mRVYw9Omcengg9YHnjw/xAvnCBy6GK2bv
mLACtqv2VeV2WBsmmafdPDc8gVIavvK1q7DiLJO6vIZuPzf5a5ygIaDtBc2wUnpJ
tELDIUXnbdU5qbIjnZ+JDf5DIV5i7qw12aVjcTCE38H6ZGH3ZhLBFMt+AHgpQJB6
bZNaJVCEurhvHl7SSCcV0rvGHp5QBu8h9PCPwZY55oGWZxEHifJBikJgs25TcDAG
05hn5AaagEYIaiYqpIsX+mu8VymLIfWPVDXRKa3EzwLGNVj9UNfX9gMMICNKpUdD
V34K0FDQA7ht7HJqTVcMjYU2QBJHUL8JT7WaryZB0hyymHodsfZKXQZ2mNYkmhBt
JKK37MSXVpVOWag4BsAD4kxqCnTQDEJVGIqa5nq91El6a0WHQdulU2bxw1BDmGVf
L+t6Kawx1+SowIHgbhXYW98UyXttb2UioLt7lcNdZt69V0N5JfEg7QoXeomjA+fr
YnJLJ4f7M5UPsE5Pg2Zv6sXv/C/8aBAPxNWQgWcSmKWMnFQ/qN85OdAwNooMODQf
NVffeDuGbRTdtnmRFADsrDk+E10BTMigIvtpogWu2gaH3OUT/5cPu6LIQDf/qkT4
ooFEVrHrxOp34AbUlCU50+AJP9kbgZgKMbjhb5HNdZsPz41Imi7uWd7z6B8zCGWl
TR0NpfbbzmcgZvPEi8XnzCNhF1vJtF2Fv/1Wm+TJ8rc35pykWhJJucAhzQUtLZVe
qooCohV1VDoa/qSFfX/pU4q/c6wVTrtZT4i6USXrghlb8ckB6jjxtAG2sy9wrhYq
eCcHAxK39n9rbPRcaszBiOE3XYxPSt7RcN6eqbOyWjMcbqL14cM+lpzwBeVXudDm
GQNnwwlbM2MuyMpkWi76ZMCMFwYJjTOebqffnrUXpwfTiBRMQg4bVgGaXvUIEJ3L
Ui5/Vx6ViGph4TnH02eK70DSppo9E0zSjm+ZnYte+KKLA1DAAkvvY82OGzj8zwVW
75IDMresGxVTRjtWmoOI25OFN+YQn4EmGYA7mi5S/PaZtuPHz7KVyRcieSCmCvTW
yrwWq2v0QJbaleOichr3chWq5Dip1Uw2ETKQz3svVN9ElU5+gotJdE46qqJMbV9e
9eAe8BL4UMvNaerJNMz6Elyx6VHn/A492JQKLasN3uiiZtYVHLlCd6CmUQpidu/W
cvEIjI5eFRnwhqycfcrRifakpXHq3Na/89680dI3iKwhYBO/2bdCTnaPlP8iUy34
ugrI98u3U5PBM5j6IDUxchf0aQ+3xiRzUm4ZOzLHYMObG5ZwQCJqK1ufyQDWK0lJ
kOxXCLFM4SJ8Cfx9ITVT0zkF2+Tt4671GQaXchhVCE3VXyRT2uKpInEZxnR3AyZY
yVRanbRHSFh4C2wscN3b28TBFPME54o6I0AzXWgu6/E5v1W/Jv+i9SFwjYEPwDuL
4Q2Udf7kqI/NoGYJAdORFU0DlfyVrJ7ycvxV4uVw+FhTx4+jRfhhtBb/KvLr82NQ
3jZOfdWruQoRNu/2hSJ+LHYftnejppdBEQLmI6wVeP3F1glonFNP9OvJ6Bs/eN7z
qubV+M2PPczr4UOqxmYzx2GpfpBQhe728w8U+M167/owsSzSv/PRbUIIo2+abZio
Oz1GNcW3kAVemevy1N91QR0CCIvdQW58r6hKgEHXTkpj/AYUWT1i7Nv0J9s+MAUM
EBUG8M+QXppiGyN3+L4l0nHEQIqFnE9oEMWcGJKYZ0w4wx4wxa2tXylQDNV25n/B
de4ZjLMU2rjSq5er7BFJeBwmnJTBnuy9K68GKS+8BBuvZHRgm2/c/6wU6+rC3TUd
rYstrSaznnI7fx1BlasioYbbgKzKVQn1zXtsIk2aBXF9lwGrMphfFBe7ZkcyV/db
F75wWF5B5I91XUNexSHjMCXUqb8EQvYbTnUdkNJ/SPFjB884UjOSPeDKXKvvt4Lk
tpW4eNwkb7jBJok8qhykbZGfeyQlfGUY3Au0vRCobkoaJVwBV1xAMke2z3peUBzh
rZAgWYdnr8KuzV37fkmk8cl82nXhNehqh0YkqN3RZkKwaF7Mgd4pUSk+PQwCH7U+
l4cXecd5GD2jX7f/LbDA1C0v+Grb7lf/oBKodWuoC06NaTX9qE2Nl5OZC3QL3ncx
E4UWScuH/ZBM3vsFfuHRdIaqNSA4K+k76grq7FF/mH+aXB6AnLu+nbkMwPxr95Zr
QyCqNhEyBPU9zv0C9Pg41stOctw3xnkDZNC4XKGnxKSKS2aOHR8SS4ckfOf7Vgub
bun39G5Ixcv5df6IZelLyPo2GvB8nljuE8iO0mwrRoC2c5kdz+SGRJ97xOzndCFo
ZKA0fZuEpLgifZz3WRRrtUIlF1VxEA5smtA9LW3Bhf59hmAqOVI/3l2ygeCDdRjp
m6Lr1ajN31Q+S5vm55Cm9IQ8m6fBo/YSi4DMxSsrW8yhHpfUHdQ+043WGQOcqgYi
7Eud4G4og6h5RgNCIx07ODHZad9eZdyVP+f/1WPMxvBS3OegBte2jJZqWOeenNxL
jYeuQp8qGJG4g0EXU7G2EyNa+shoToGHWVjYUmzGojveFdAA6lcT6y/DouUyCkKX
HJhN7mFePjldPa6xBvFTBT6CW6bKMmAWf616ZMWLVEP2LQo4lLntzgqYQ2Y5eDx+
YWYZvoqKesQ0qrStEkjbRzX8mTTADc0xmFeca/s/jhbh8OpupWAIra1OYW5Jp635
WUpUoj4bOUnuG0pusYT6C5GccTBo3GZDwX2yh3F+Desm3UsqwOYjc6w/DrxC33Qe
LkyNu67nqS1eXAT8lr6HTr1UKaJ9R2yrtEi/3EzESrkeZ6yHXHfX8RiQ0E9XMsvp
17PT2VDAswY1gkVbruh/pcl23pmgLjoEH0c42q6V1PXrUQwOcce01SCicHn2XXip
75N2B2/TgFC9LqILQOKklDKd2r3bk5Ng38bpWgFFGupQW1LDNC/4LkyrAaVRy1ha
81RVKt1cOuEMOMjHeNm6c+C6xLK5s+5DPIyb8GOB5Udl9ogl4rtsQrQE8NS8ld7z
ubutU59S10TQQhkKvHPdGzSTqvq0gFpRyQzOfKJSsH1HIF/y/DkA4SZVSuX7anLT
m5DkLghrMWLvUtk4tauivCa3b8X1j5Y9rDesXSotApzMYP02ZFkpYnTgeP6CW98S
phUXh7NELh0Bi/tdec1zLcysW691qZPciJQ1WnpLlJEuXuhFqxKiH+cEe5OuTSdk
CjQ7nUKZWbBAP49lzJ0NSUuFBR7N12/6cCvUIksbNa7I9NWdJSA3WxBXtS4fIlW3
cPawGQefotGYcrmJ8d02WmiM7tSHiHwFCmhmgCeguARRMhrdjvFNaYlaSnFsdgXv
wlw4VPN48+dmVAOvN4NRxm+t0L1LNCvsGY94KCqroMCnIVo9OdUkBAQkpPEepGxm
V8N9T5biuK+GA0wnhxHqeO7yN87BPPGO+qmcajK23KkTebcw8vZ2SqbqRCB1HVrW
Z1Lg4JMr7rF5vMCrdQJdbAT90LhQPCyL3WAGHAi9bHuB0dqW4uFOwqvuKbA/OgYw
rcnlqOk9ByZGY30Kh3LDM+7WnEOF/Q9NmM8VpCt09Cc/2VRRM0cZTS+v5g00Sp6o
NzR9FgDHiVE976lFLNp9djQxehKndW+2y2HYsG0UUzzb7+6VQThvKyMMRPtJlVv3
ZA8GVbrixnD53fNbKSGVCmTjq21BRd4BEF5KJixDWwjfuVS9NS8kATmd04/zjXWl
oCU1rsAiUwe1pQLXWdpiCHSUlDzhujmS1S37pocSKn/fQtQ4KvejoQo79o+YqAdr
oFhQaEkO5Iz+H8AVhTVFKl8R55MXpdlg5Ee3co/+w82gKsndRAkW9ZkgDzGrPfVt
/fmH/VStAkdrpO6JBT7VgmlLOYkVcZi8zZetB4rR3xElrHrQCrA6bN/HI3xPzNd6
dB6A1PKF/33v0u7Og1rU/p017yjg7vOy7apxsPr3oZLoFyyFmRTNphhq95xKiVbK
1PNGVABbNYdlNBo26gHmY+kNrAuennrosyqruu595ds9atVbY0eNpCgI8M8Z4yHc
UvZm/K4ZcZOGokw1K8TgHBOmN9xl3eJ4h+DnZWjQWPHvjOeYL9rzGtK23S5D+MdU
8wTsAYRtpONPdOqa8+N6JxYvWW2bwnfpPQ+H+wzrtmskeJ26TrKnOd3tvfqrnP3G
d+BN9nfXxMfZj+3EWkDDBzFSZtUkOYtltZrEI6yHe+67vUSdeEDTreVSVqBW1igi
VdnEGhTvzDfXODYljIsEMTgssg9aXvQtwMdPKpAlQCmnAYzsI28G+wwY+XjmEG2M
PiTJu6YGw71oJFekCYcGS8j5Wq75HWF5PXDLrNyFmB/dfoPRDOthspQGMHvgocd+
g2tl4ruZ6tCcQAzMx3aJGgpq80rJrxhvlGy7lKQrRfbdJKP5pMxf9np0gAzQuoOJ
wSzdiB5TN8XGq2dmaJg+wYCny0+xN196rTumw1U6isfVhINNP7ZO3gA63S7B09HW
FU/aBKBJc89eKMpRYghyTGNAnNy/cuU0/mc/jbggQ5W3Ckg1pCEImxTBrjjXwCBw
dPz//p2d0xsJqcfi8qNjEpJTzMEdjYUDbCQTNpcwFlX0zzzWnQp2QJep+7VjdZd+
iWJXL098mKtO0qKem9aEaT3JFq68nou2DClKiel2L+zWD9JPfkXOy5j4aKdhuArl
4qS5nX0ZuW9Odw23Y+Dq7GeT7s9NcQQKbqBV2AQUJzILQVhtxFooBD9+W+hJcBd4
WNLBmIF1zgIqd79ZwzIJNGHD7PtDBWrpVLeRslHijm/GfEbriJAOQGVzUdtLXl48
LJCWaeYiljSU18wycj0yK83AqVOWoaqSTarDn1pc35anaXqldzD5mo6CbDlaLatQ
+oMISCexbwGTvYc9u6MQzFjLCQo6DekuF9WTpvEVUtJxrf+5VEq+8VMiBj72rDwM
t520Lic6tJN8ghZ6dElHaf4ysKI6oKLuerzjlngkTR0/ZKgZTP1X5AKdc/Z4te9N
e7iH/ZD1SFNSnNUJvlWKGKNSRTmHCFbPdq/EYD1/NgQVtmlUKjI5/4+79MRhoyPK
fPbeIbkkhStADIbZ8fHypizEr0zYe2WKNnrihBZpriz+5gNJygFgijHc+qTl8D0W
d8K+/NY/3oPji378pIx6gh9EFOlQ8X5ijgDC4tbMS8hHGyp7l/sDJ/mgpFcptxpz
DIZIiX5x4GxuiiAPqldUYd3VP7CrRWbZp8HcQ4apReJ4a2P8np3hWYJVKmeLKOm1
CMq08X+rNADt2K7pp6glpxbKrTq857SnVmv4G/5gmJhqRGGM3xSg3PVGRgxg/5LT
P5T+nZbMaeZiotxGNgUXdS9d8+qBDIyKqKqGmmbZyuWhZ/KO0ZAbRKx+TR8aYO0z
O8/pSc7Ao341R3ZO+rNsAd/w/BEiKuzQ4R5xxlzodMA+uvFjfO4PAWGgAivcL1/c
Gv3InbctwGNZNtR4eDSWJ29Jcc98UTA2VpIqie+EPMSFIaDc8QYVziBm0eRyVLtq
+f+97wGXmaWO26GzcGjxIRSWxzK9L/6ZCZl5Uva/1crQCkBwiN3A0N45F0+Dr4pk
Z7Kpir5GweT5qWiXDbBbDcxcpAiMUUVHjWa7YMfszJ0LgbVlLjZthcoHjZqicKTF
ph7IgNOeXF0ZNyE9vIEJ1d/YPBruf1N+B4QYgSptxrnDqqFpbUaF89i3mjgjl2ms
lAQQk0cDfJhriI+tzGtpuj6gcmbqkUOvDcohxtn12SoJuyvI6s+A3R/mhOK3fMW1
HuHvaXYUI9/vS45f9YGKltOT7F/soKHH0QNs2s9V6XXaa3ciJf498yzWFy6H5c5q
D1X63bEZMUSyDWQ81FZi5hy5g/UCq9c10aETDLCSwClFnwJ1KKzXpW0Nvvjhd7W4
dFrpRkT2m1fKm4x6JnaSpqzpP4Bghkzg5NBWaxj1O/LHEcR+kOxST09DUJeW7TLE
GVE+9koMIiTy4MlTYAQrGuXdY2d3Dm6WBpYSbadq1MlihiQtLsQKyuJGqu8tdaWe
pLOGJWt9vWQTTIj/0sVmGuWclEWId3ZjVfQ9r1kScCQsbuxCm93UG0093l7VZ1K6
1Kp71Qlzn0XUvczpD0lPlQjfSEl5UamgWDBlsuVWUUUZTMhzhAQutkDk/g/b2wI5
W12PR55mqPMGY0GLTCo/N2UDy0SR9xMgUykLAXYcMiDfMY68TfQgIf3I5mTdhYPo
qh5z+Ca1nx95dtLDSBE/TnKeN5jCO3GDIAfby6qQ1gKgTHiiv5i64DQB/DkfguME
HrTLwEnbtqbuyfwQWJ+JhM0L2LLZXKCVQbCdYscrUGrsOn6/3Gdy5/LXwaInZhuB
df5HQfJR/cxJUhLO4pX4cTSMkhDyXrVpV38hjGm1ApTChGSZZJdrmpTacQl4OdeW
dvgBH00XSr56/GBFRITiqmxpC+slcsZhsHbvHhJJXy+0FtzCE/kgNJZ/1/fcMkLr
PrNr+AylUK2L6rY8rgh637D1lsNIDNVfabfDnQRQZXQhLKTahtRhtpPL26gRv+jh
hSLgC1AWnVZOSXN08lR8ZxqzZgrJRvFzBpfngRFESFIkoneX/cAARVD71gZ435i4
X4FiU02PKPI6Xfrqw/Y5oGJ8XlUSsRic3UbMKGba6OY1D0vaFIhcRiPCfNhDFvQ9
xgxQJSyhhoauEWmdex67s6aVNKXNOWVxowLnbeEPUmaMgu+yP8ko17E96rL7s48+
HHlm0mwunhhFt1Z8YtD44I2llY6slo8Ldvf+x9x/IoeLsk2KywA2Cj2c7yEYeb3T
cBWOaAqYfC1a63p++mfCJ53t+nzGUl80+X+y2H+HxJqKc0FqSJ5zoXMvuxTrr+va
0VkMEB2RyT6b13fNAdDUzBZcHzEmkxaicksLPZR8EkTu16/3SRJWhjhss1aMcbT2
4aaoCEYzYwn+ElFzOc6OsLrEOxElwMhd49O2G3qTEHxeUgIhEH0Wt693gj1J17eE
/Ri7pC35gPWGDXm0NEWYvCfHOr4llo69h0fuqcUGgaIoWzcKFu3iuyLKwTKHXM6d
ZjTcOWbpeztDSDYwMXAIQNrPhHGaVPWIxysdp3+U1TBwO16Xn4531A1IxspCIc3d
yBH0RFpinQTwlkH/O2gcS7Rm3u+/f6JlYmnfQoh6X76SMQMPeUd+iHqY8ygx3L2p
tJmY3w00kocG08YcDn5uKUtwBjqad/SKI670ZnKIj1Z93w96a42a3jy3xD2kEgGz
+3gdJ8Lq/buOkzDcpBZggGoiUi24pIOn0D4LrMAPoT0wgL/0gZPklk5Aml9sxWVb
JNi1yS5fe1cw8Vov/7Y0CKw4cvhWsj46jxNrMXe6Am/2lAiAk2dY4JB8ZAa3WDXt
fQ1CC7jmfgRF5dHaWxqgVaKrbBkP7Rm4XzSikWUkHFfut1I3EWPCN/Ma8JUUb3Mo
0lpsLadS22y0bjbyQUGti2dvHpc8nwmaf8HyLuYEneOU0rREnWyyy7yhUsPwTV5F
cNK7W0PXD4LMj/dI9jlAL7ntRFCFlS1X0p6kzZTfMf9K1sYMw9ZqFUw/jk4U6FXP
clKMhSLO/Molqj6tFDwWhnTl7bRVHK/uvSq0jZ2NCPJ+t3ubVn6P1FaHeeTCn0zj
engXOR77KdfWawdLIjMQoIuo5M1gjoH3+eOF2fMd/DSyxjYBNEuso57SnUmxqHc8
ORujhdEw0XoXyXElYCx8qy9aPDmzwlaa4fj9ISdhAty92VFwaoxDu/9kOMcL7nOt
5+LSNgF25U5rXqfXdG5oSncj+afnCZnuwxzHoYR9SvZv+WaacEMo0vWS7+3ZJ5qS
xvsAmEd3HtlTXcJPcoW4EphJbuZF1fe1S8rOhF0yFfwuTUx+IJIfIRIIMp0/zimc
xBXOPLMQ83JKZ74WpIDxrEUjlT3pV/7b2uK0/mWYPiFc55qllcutohdgmIMHcATo
3fuh83n/B/K9JJY3J9m2VdpwP5+icy3DGaxxPomnWMikQelASpkwxSUhEwkr7Qu0
1Qtylzu4+9pxd5u9LCdF8U+LG/tgld2PykIepJTv0TPmLg2z5NnqTNbf7KmGRFSI
BLDZHrovILLoVYPB53HtqdkHL+N0ViVCHQP8xylWCo2XJ71jIGk0W+YhleVdszun
vvSW4b/J1WrSS6of8e9wymBh5xtXwPkgeqNI4Qpvxi/WqsDqjzBR+39jzrPWchl4
Rbxm16JkKWzlyayudGui1F1mWt4UX9ZayLs4NQaeUGuWx+G+Wp3MJgOZhLvBzjMI
UqDqPiQrasK+vPjAVwVMfzaJFsagDkq2QxDinq8bFXGfzFDmSdtlHzngARLUVBg7
bPxhwMb+jolA3rrf0zOAdipATMA8TQMOCOUE2c8biK5Cp7hs4MoCYUBOLLuE5wMf
tsurwlFvMJFS9R98mW7fmkiuJLSGYzSdvob//sSbGGJyd2X1Sos8Uu0ummofxjSL
84KzWwJzXdwNjQ56UVqUkCnrDrBZsM++GCFp+KEDe5utg4NqarAaUrNQJe7Sdol5
mMNZ1Ge6FQsuj4JDly6j0R7Uzez1chsRHKxlHO4GkXFdALCVOp7VR+v+T51tb7wB
2m5aCRcMtAQf/yoLr2Et47UAI0gPPBlM0lWXAmIftEkbkzS7VOGf1wAVXKKTT95L
pvQ5WOQTbpfyECDpyk5ofY0TNKwsGxwh2OmO5WGexgyrh4uV+vAtBQRvBijKfJSj
d4abAavRV34sPiErC7sPFPdS9OgoB+Ga5Y/xrFqDFlOLbHT8ct0mHxnYwSJqNMnZ
DqCcmYrjgfC5l+SfOO8fuK3J7mqecXGI+70K1gGHa3hEuJb4ZlMWVVwfVz8nbl5i
3bc9YC4dAX80nj0zoXYyhEut00c+Bp97Vxm2JWpGWCEcUqPyrFf2Ih7UDidsLoaP
vcfL2bPI42cbgKf7qNVeXe9A6fyrFZ5Gm9+kftAJ7AtdrlOenixgJHDhDVxtB/tm
6Aos4E5P9F3p02dYpQ5SoR687j5veW4cQMufep9cJtZ3Jlu/SinCyjLXh+Q0ZYQN
Y1V2h120DE7Qz4B+2TCA1rGwVUUQEc415U6XPoK4i+k61hM2EDc5+oHokolkgL+5
Dzlu5ecK2gUJuxTj0jHhPu8T8O8108lg7UokRu9ae4uqMv7R0OSgeaFVJLPm5IRi
MhdgMK72xSMC+9eZ518kQf8/1ntaSSbMhZONqlL/M1AjyIxZEbwcWSOVA13YaBiq
gU2cEKxNLTgM/c5BjirT/EvBQKWyEdjAHISpvNsPB3SMzul6y/Jp4BkbynsN5Gag
Ygzg5NwBFd4UE2r1knJDb3qKpcM+qH6djOeqpzzmEZ7dhsBlg3yZ2vHv2NwhhxGs
690diy83Vc9qXIuHsABUgDsOl56ZPH3ZHUjRjteOwdOoPcr8Ztz/5MZSbq1SsAGc
gb7B/fVt+QR6HQPC7iHDv0F6wUP5dGnrFe2W7Fzz7cBNQpTmOqx7rE9OhCLYiee/
6pz2c36XX8VPMU2lW4YlKodCz27WRUNssgJe+51f3GkAq72T7Zb7LzUayI88nabp
BmITy2PdTI2Bn1/HodQ7NSCl+EbrDVBWZzmoPhxvZR2n1WDuo6MScvFSW2h4iK9+
fuJg4ncomrE8RQ/66u3Xu7PQpDwqUTZLN/7hH+Au5Uud8WtJVsMA+s992w8Q/3PT
dhT7+Pga6nXz8jyQEzja4W7/llJHw9aUDiYqqLUjbMAhz8j8bRStinB0qXQNsav5
sp7xSG2XEIn9HEUBUwdiV47Iw1bc5Llj7lAytqZ9Yb3j90gkxF1tuavAJoJgOXON
FdF53nYpG3+X9TDXhiRKBON7a2IruDA7gt1N7Mr87sP1Kanfaw4M24v8Bq2Bdfcf
GQg8ezDveXSWw4MqaXMxWctF1tuwG1MrK6+9/NaswB6pvBJiRsijMEjBYKCDDC+t
SaGMQngBRd3HCHnRAHjsSUWBmnTZxIInz3e5EaGGGVygXhxUJDRLeRaOXoF0i2XN
O73bWnADw/fA7nYjhDsOgpE8m/ah5HwYrehM8xK8YPQygL4mG9nS0K7XKA/byxHY
hkwSgsHB1i0yvikmBuULg2zXqxLslxVD7omaA2qIVKKKDCoWmu4gZ2w+fRXzCrKJ
y+PrjC0nxAihjSN0zclTzj2AhHJPN67Q8mFHIgfOh6WHAlIHYeiZP5MkFjoZhFjQ
ovDg2ZGWTaWUqeMQbVkS1CD4evIUh7GR3edVD3p7WhIBLZhuxTvgfeMTVtZwPKpC
I66NDYtUyJYZoPhq2X0kOCmM2CclMAqBSIsmkBRiV4P9hMrF2jCD62ySWzSoKnmC
/kuvdtl/RKkZYyb8u/w0g8gDBrNF5QjH4zVZl1l2kpp86tC1V/WuvnWNLvfZXRTZ
IWlMckHJFILzL6Kt4sN+cykRGSKTH/1jvTWnTjASBBgy9ukQYWO785lHJyYe6nZW
rLFDUNwhwb4L9eRE8e5FlDsASCF7QCyTTJrV3rNojD2+PbhPb6F93B6wQ9gSypY9
PyAbWEQ7YfyuvzaynYF8aKWGspTscbkfXjoOGe0pK04HJJaBkZfgJEhrLBMo1+Vi
S586hHC0IjA0r8KhEdbq1YeMuPUJ7fh9QPMf+y/p31HG7VqZVN5X1QcExVI8pvDv
VqYMcGZeSYX4iWhCo3Ep95k100zoplwGNYlCvcYkNCid7QXsPQx929mmIMMdMPUm
gkClKPfcIfkuJ+st6bwr493HTsoAmo/7FB23BwtEvIqXepRz0Bo2sBheIQB61NFB
hLZC7Y1HZrBcaPDA+Ixs8DqiVRR8Clsz+LeCkjqNMUHWePRo1ZzM7s+0A190HK7i
Y8LlbwX4rm0FcSAK7+MlxGam8cgyBYshbDnvRaehE1e8UrNblgUX3fMgcn56KY6L
5bFWn9ds0f/RUdBGpCyHh43Mj0D3bLOCpRYRu5etbJ+jQS4DHPYmJTuc1/M/P58V
4KWEgDezOyq/Y66ESIIefGRhTeGiqaxTXdPQFZc5xuW3OEyWNd4L/ZkY97c1wgIh
Y5WpgbkE0NL02yjgso7fme9yeMQQEN+ksnRAU8vF2X0pt88F0kAeAQOccL/7UiyR
k8DMNbaUOP6M+l+oJ/JIhuwryu0LMM68eGb/1bIj3CRF1aQHrhBXsyX+jLsEheA7
dEj9A7nAIrn4DnViXyJSjZo4+rZ04GZeCMSZjK9CxDgDRtSst0r4YlVT2rWKmqUW
0MKNVvsduthav+nLli80RE+vg2/CNyM6Y2mFgmkj1WWwleWOb/vV5OBOFGj2QcmP
lfNYqV3UHr0azyJNgDBHgXK+tQO+ksEHTJc1rDBPii8T/pa4W6oL1YM3f2nyrB5r
XZ3dfw/87hY20nrPTWA6345udRjEeQZZFFSZNwLIhMsMy3BxzyFq6KaoQfYdXMQw
mwuxA97E6C3xkW+a/FHdpyTVxg7Fm95KrUKvKJD2neYPUVve1o8cxPQTOVWKUoIB
FZvZ3XTesc9UlfR9vKmDCuQgdP652cEnybtmZA3kGqn2ya3MltggxZDadrJ0YrKU
U9MY6CwbP1rDVgqUkMzV5uXGsawTW1Me1gkn/LmPSG7yQqNOc/G0FD6ULExSprWq
PZFCkZzzIteZi6mJZgQ3YX3n6r1U37Y01yyV3IONPvdORBAhj+BZPC+OgVvX0CT6
GbA7GdsouRlCqhKyI6Qk5cgJuLCTikE+5Q7rMevkFu04Vlxb9vmy1qm2OYOi8Sfr
7PnlQ2l1rchmjeUTJ7i9UopY4zXp5YqfxlM5oB0gf1LU3JJHl6aFOCcrirvqfNXt
oUhSDqVirW9VQFka/BqG7nRQdZP1G3J0ED2yC5E7U/xZ5NNCLkT1p+xLgu2h86ps
aPRD4z50F6ZMrIf9YToqtsCzy7WBvc99ntTHNvR2M+OFp8QG0Vyw1NjFT6rSW/K/
75HjEvJlLQN2TJQNQpxNnlXImlYkbe4UXJ18GRkVR4rr5uTuVrTFssEylrtjaoC6
pW4vYdFFn95DcG9EpZLYeb2Ia0C3HGPpQ6MrRr72fxdhFNCYXkyRNeIVuYNsIH0U
DIArdSfnEHC1vUh2lKXMNRdD8HPQf/Q2yISU+zHlKTMTXXiK27QRFSiFne7VvUBy
SHvOq1M38TcpzTfAGT+cv3E3DBdmIQrE2es6R85oB/E3Obeaubn1YcY3On1y4YAh
z04yXdXYuW86pDaIHqykjlr2PbfPdEoS7VQFC2unmUk25J07rfoI9pupt/xrpQXY
QpOV+LnSX87n4+S4mDZylK3pgapzLmJAvzFooPpMHo20xzdwgOoRBpqSvJ4m+kzW
6Vqo2jWUqKoyxtqU55A+zWxIIbMGBs6cfkmH5sSmn5jA0AtDxLmwzqHmizz/o+nB
s867zAAePjLy75Tz24TMieNwgR2EUxtUlWP5yDS+T9xH5EPm/16vF9VAqM8MF74q
iDsKZ4tC9uIrlkKIVDCgCDIbB8hujHxTQqox3q6V09SNHWPNpzNdX4No6cqMl//3
i9NBc0X76Tcza9IEXXR7cvX8/nxPQ21TdfonUR6JzS/ihqS5KjJKgETEu3B1jvq0
4hFLsBIPpYvPcWja7xqdnj5mixMcYrNjIT4gJFjSKi2MvHOg+UIahW3qNvh4xFfo
yAdyAZc4ks8iQGQOwz52hkGNyoKaR6qJElv+oBBPX4d0EIiP1GI0n8JfhhRdwo0W
cqjobPeNsvipzkW40eUpR7NEEAtX9/wwOeOQltZu6dZ2PGrmvSvYG5Q/0enn53RG
V78zqId0ALvG/ChkqWfzAsriK0tELjwWmlQmsBvArjF6tq7PHhT7vAbJfJrI4iVf
udgtm64CleppFEt0phfW3uc0bKy+LGU+OzRmUxtBy7Y391ZIlYZJKEbwH0vRLXiA
qQySDOYQl9ENfOCwXKzgJKLZ29wpIVTBc5fGvXh7r93+uCLLtnMNbgILlBsIYA0S
xmcYIccY68J4dk+JfPoKG4CjEI7BfiR0YgiXiOG2appylXwZJygFeSL+zC0knncz
46ifJ++8D7kWEcGWrGHPFNhzf4K05fhMYxyNjNAaKYbd7TjIXWleGqstqvxiGO8L
5ROD0sgz8enm6+yf/I04BsSuz34k2fr14zZ0r/gJVkHumzELzobM4vIrff5C1jTN
IQlLWTQQCCZnzTUKPTM3Ccbeguc+choN52xIKbc4VpBp4a/e3AwnnTYv7bW4AiFC
5pVjOvqjxkJHK94Gk/cAELNcfXTxxthifbfaO4oDZJwC6iwRmMO5e1isxkD4+ViW
m0rWBL9NDPyDkP+/07/9nT3XEKbG4ulhvZdwQdRqKL13EWE9RXF/cDO+gRcqD8Ct
ygsKTr/yDFzNOnmUHIKyoZhQ5hBtYWQuMe7Oeg64HR++35J5cq2CiwBfeo0PF33o
M2HE43mW7rQR1m2didnEMnp70RnL62dyVVL8J4FIBxpy4yUyFtEyjR5Dy0Lpw9pv
ZCGQPem8gmfm2NvwNoUrFffNO+RSTNPFmGTjvKKvX/Rld7lN4CrZR9TTuwwzX80d
yCactJuoZ+9OsAB+3b3pC9ibuJJvxhfmDxuyZSFjRMtQL1hGmpluUq/6T2CX/zgY
b8mKqut4DFbT6rGrgaTxY5yAMHSisv6vdlznrdszBcqFnVaWR/yJGdy6nBbP3wG9
u+OoXCXtNqsZh6aQelynbAIOnNQG6IlELGiVvkca1USr5ee14nqPz3h64qN4+LCm
Phi/LUwRgbkW3QoAoYWOtfjEEI++iK9uWOzPTLhfAKmXAcoJb7g6t4w8/ZJatwBo
J9+dCE4TrAQwthl5N7nMS4f0E27DmGgr7DlgbeDQFKleUt3kHHAEEm4vsOSKWSzF
YzfSiEEKOO9bItBEILzJGaDBw161E5IRGPMtghJy1hM8DX2myOZP0/TcNJDIDwLD
KDisTaM4Mqjkpt6+Jb2XZ2CjINPu+tmXNdRG55b3oxikPV2fOKNOqkNK6wKUisgQ
zVx7lGMMY20u/tuZg6fTK/9fUsXKuunSbxhUTmSWraIZo9ErROcvM1hPD8o5eeZk
O2mg08vOGyPAwR1MbsbEQZyxasiJUDGNiE8PjjUzhGBexIR1qaLGde042xLHVY9h
RuAUA4bOueQF/dt8Fq77Jfih31IwbjClIIF4iQICqqvUXhdMwpED1junIQ4/nSk7
PSOBz0F/a/scgSl3bka1bAkP0tAg/N9h3ewSaMrdtzkPDr7uILQrbOX76CaqfLn6
XVwObOGMkZ5SD82SJToh2KIQY8kEdhmtpjxXqRS05OILLzpk3SZoFWolYvyqOVOE
rVCVUjPlQEVD+WfYnzOJoAo/X0iUJ9zPKBqf2jFQGRHrfc0Xic2NzWp1A6A5Z43H
et5C/POiL7fIcV6IThWOaGlZaMH53kgUxb0nUQwlwficWJ1vQjFvi9Jnd20bcoDp
qqcJ3RU4G1U9u/wExTCOS9OWgtfuIwHg1GVpVixEb+kpYoBnyQeT+lkNlzB1pgdG
rW4oWcP/BqmY04SlULp4HfhE6oizstCxn5Rg6hZZtn52aGecCZOfr0sA4Vpfy50n
T9xZflzNaNyveT6pZ9NN9byxHz60FiE5j2MzKWspK4xY4mJdQ8KHH0YzYDQpKAFx
4K0N8hwv6JqAHPi9eUtqP2mRV9KB03ijw6iNc/ReqE/FQlco+l92CG0xBgqS262F
jUpPOASTclE/si/EEX6BqajoMwIQd2PSQUCyRoUEzuVrzOo3FLRqHhp6OaRTRmDR
WRr0fEvJJxQpqKdM49eHYyulHRGcVB/18uBz5Re+GfGBzpfstL9ng9ZsQb1KjHj0
dculXSIFAO9CoU9BrtfajWTxmYd3veNLjoMtx3pOXpxcE6zugLe7m+9o+Zuet5tQ
/5qT6Zmknnndklz3bH/Iztxhw56dqrWqDeWI33hnBrEQwLtGJFJDLrsEWpm7mw/Q
Ktok0BxSsdgsLNkIHuTKVi/3IukCHXGxune0imhuX9+DTemBSpmQV2krb7ZOVfCY
K+MD+dBkMDe94s0abbX+1Tx7d2JH6oPJ+/SiOLUfQonLgMFR8ijdN9yfsEGzwiIH
1QMgAIKubsiUAnCYc6RgqYbK3Pf3rPigH13FFaNzJiPMWyZu42OLe1Er3RxheIUD
8DMWfU8jgKAPL2nLvQ7juHmaqOhx/q5Rp7aRT0xdoTuQmZWf++8Q1v0BXVjtH5/J
7Z0JanStqyv5aDwoUzLl1Z6dYE7CNQTSZ9B7Wyi7jenzp8jBZuKb13pn5K3FqJWE
7P1NVkJyT4Xa793tE+M/wz5kEFRncIdOi55c8GwBS5MttPcZTRVbRHjgJAka6Le7
tHNB61RYw9zzVyngzzbOLIbrTmh7VO5/JYsKXdh2Zyh+okjhy+wcY+dGPtSS9GpM
aqboNMP6qh07Sa218f3K7dmYD892pkbflkCiXKjC7Bk4DFkllB4t4NeLudfjYu4j
fxKWtBOwtHGe6aSI/1MBfg/A5yJO+VW/d+7yTSbIS+kinR+y8wAaBxkFGq80ThaD
amug3Ql2qYZjmlDFKOl0NAVWbFwX83XmDZGD0bGt2lyhbpolz8fvUlX9ecYPH2uW
7EeG9/Kpty7SprIfO8WYl2DsPA+aY11ndtkIl2UPIc6xxv2HPAAIUJ61arub8VtM
BgnuFmeo16gO1uBhL6aUbU66cnN9lOMcwfNuyeDfm2NtN4RwsEHC8nFtte4XuY3s
35u+rTSM5hwdClrpDJYJm08RcYWyjRTZC5d6s9RWK9rUSRmkV+M5iJ05bl6EB2bh
tOcKLunP7QIztVQaXxlLvIC6yYU8eNZSBSv4EznVX9m5reGWKJZynDkmCTRMCWe5
sH523qN7waWSL8WWO4WBq/mPL+eWki+qcag6MV9IQ85pn/UD2Gc3H4nhMpEvOKHI
miYjBmhf23XS95SjCN10LKGh/YjvygyAkq+8yIEo/OE1RrVqjAZLHlAtzL4zwxY+
8Mor6fvGtL1KWxT1tENgMyrrbiK8UD8IsXElc1qdvjE6bWmO3G6b3Dmu4ygKrRgi
6QI2Oh0PW9YxR9RBkISquwbJuxD/JQ/IzuOA+osG5F0BVVZuDRShqCkclGJtjxwj
nFYUV9uBfocq5+wcbPhMOWXbTS5+aobgriI2x1wsJG3cCWCHoegaY7jLIu6uOJGm
XSLoVqiirgXfiNYnVf0Su2sbH6EH7gHI/nbknRGgEQtbY6mW7B977Txj0R1ycg5F
l6G8AvACyetFxv/5QgJ4tUaZX2RUV9mUHSW4xbc9n/T7fzcQnxXdkWschr+r9NWc
V6WAUBvknv3rkE8eJuIwliSzfjKXKq2+LzOOgJADCLbclDzAoXtmfZoJNozqS3V0
O6e6OVuwFGGijSsj+myd4UXcNNzCGdjRMuBpl5b+PyJvL6ukDokXKbjzdjfq9+Fr
dhGkaG38YtyUPr+qDZ0rQIbLQDlhTH0017ue0s4wmX/rsbxeFeEh8rOPHW1bI4j7
GnYLX+qEwpmKnxr8yBM50SaK97II3PKI0YRz1glpw4PyZdDzxvpgIqnzVi71lN6J
BhyX79ZUYQxwWKovm/ZUWj2x+yDAAH7GycNilWXWZnhiv9pR3g46FOHYGUHq8s87
fiLGoW/0Bk7RFNuV6WlGhYKg9BoWAnTYgbJyXe3qU90aUbd+6041i+4aH35Y+/yS
02Mn0uOapTGT3ME3KughO9WryEM1lHMIvoS1ejdNI+K9SOhHtOhfCu9jurbx3YcV
mK6xZgu1ZG3bzlE61GzJOPz9MqSnUfYi6RwNQrAyCKOmOlQPCQINaazHVaDX1+kW
5YC/EKKWV0mmit5peAjHraJq5sN9oJ90u/rAa5Brc38Q36uJHDWGrJV5MKKtv68D
JWLdlbpPGOAvQg+04+Bp20yalAPy+kdfSG322iimZXCQCGT3jRNiFu/Vs1RXqlDU
/0QbsAu5op+CNDKoHvNbnEACojfb+nFn/CRMT0in+rySBntjV5hULzC3/Ae4zTE5
9xCaantco1V8Jx6u95AHxmYSvCTlC7wezuLB4S0QnCHsuWdA01bcnpExPjgGUhMf
iLY6WUH5y4TNBKUySYEcn3+cnGIyGpoSVLtIrjhXMA2nA6plc9XRBTQgfC2YvvHA
d+rURGu4tRm3jel5hV8gKo6JxCzOllxSnKxhNq2+DvxsB/G2tIWTmgJkSL3c2G9V
DjxBRy/9n5rYJklogCzbZiB6NESzTmo+tYbcEE1Gxlr19I+5lgywXICsOD8TmRVj
qpm/dO//fJtNJ4F/X+oGIZElRspqOjc3VLE2zTDyBqTm6SOdsEap5p5scbH5QcDv
TkiuALxsQkOYmx66U4krswhuLP2k/2gz0a0whY7FOb1i9Y9/lGPAuQfbdS4dDx9q
xgG4RM1XiN5vji5FhRoIGyfc7o2zioAywZRG3DXJyBnoLaIjY7TMaOYXA2krCHLv
nLv5jiF/B5SRO1oeHMEoacoEIRb3AB7PkhfNF9bB3KNMgGebuyGni3g9H3hw406e
tuLiyL5YERQywE6rFxPSpRfoXnlfCFiZeYl1fiAk283KqYOZprh51twt+Y9Vckdj
dalWMWdrjp1JMyqDA90TnhPxnYMsBplk4xlU9SNmfngnWUlz1JYVuJQHSBOTTqfl
KsbSQkG6PT9ReIac12zCZuQJ+3BJC0VrIFisrTlRGMtWGFPBUremFnieQZCPLoVi
zXygsZHz73INIV4QLUg9PDkldTC68YKqrD5zkPOUXprs6IYIXNL5C+qKzjLQXLQL
jJBB4sFj2xUta84zGMbrk1El+Ie3hAcIldGvNbwwflE3vCiiSPQL/w3t2S/ICZMX
G0a8xsGM6hdfa4ZYEvCzC6Zp7XblaPZhdqS/y4Y1JMbPA+cFiQJu39SwrPwEZo3y
cEKNOd1G4YhpotAjNf8rGJh5htCfzqOZVoFgW3zx02jeZNUQ/f98ndIqyhaEzvHs
vJ1wp3ubhWRG1kxfKrg2OOIouLumLv5u9vEnU8cn8tiv34PU02qBUOps+1WpMpsp
VGFkm+8WV5IIK8FHdDA5mYSZ4V0J4epi8FcIOlZBK/g49efS9HiRmaIHaPnpoGSC
0QnQa37U6UoBCjwMUS/Aneemo01vfCjUv9xFcUjprJ+NwdQHS8FRwci5AaKZaPAj
2PU7T/VJl4qHWNnk8P+6jyhlPcxOuNak435k3rKXkyAGSIkL5FDgIWmMU5wSi1fT
flfuHdAMjbHRfv46LfPU5eRbA1DYezvhv95r675HNXl+Guqv9RTkniunmnPxYmhn
S2wL/8GZCnxfjKqiG7utjfBY52LkFzCGkby4W7Zveokex7G/RwSIOgaY+ZGcL0TF
mBZ+8fJurJ6MUsZyfY06nKgXV8pfRXX+LmT2UUk8W4hRM4WjHu5ixu9qzWZnDGTq
3K1/QZWPvHqSFjC4sU/4xUG+xLuIaD/2FP5AslsjdKfvskCW6ir1C6ZsX57zLO9a
qhc1WzjJojKQALUcD0smgCHJZxHgXHBa/0ipRN35G5jYmSdCF61uUhua0I0Vml3J
8FredG0ba3x2mzUIoHGXmdJw/Uwpl+EoEtcDBWZGvo40eSu7bVlUd3iWUh33lCeh
vhq0tPU38Xk9Yo60s+FN1ZmOy7j7kOvQa4epk/THV9tzChw28InDZlMUI/qQzpYK
7Qh1tXOosxWHBShf7vU59v+vWZbZtSuMGHsEqlEKYFRDngd/TpAxMhvY6d8vLT7v
y/yFfQVW7FSAXn6JkAn+LiklwQzLKOE2Fgtb/vGY67CU9pCOswuP2ab7tpvH1D1q
EZHuHAnPNxcHU94FJ3gHP+PKuUxu7cw4tcScfI9EOIL/QXdkOM90EeZv03NHfjpi
1dVYGQwP7/f+gSGEAc05cBMB0sGg9v7q4ahi6Sc695d4dFNe4P2Pj37PiJj6r4Wf
yff0R7bXtaHLbt+SUpBpyPDGWkhOZSGLTqy+1s2XwY79I2YZX5E12cRhxsIaCs4g
eBNY/LShdKmg2u16aXhKlQy8LJc142blIJsG6ewFKNK7T4Usrdb0eFuiKiIKaAVw
E+q2rAKOy4nqNmlhtjMJZRR/dAcfVdXVUaIEYcFQJZXAX+k+f7o2Pyj1b6qsy2Ur
ca9QQYE288PxWysXeY9XmZjJtrFJqAsrakGuOnsbSduCmyAqNXMvdD8LscKJHvc2
dedqJwSdE32t1VfIG9ts/TY6M3ktoLiL1h/K4+ii9HyUA1N4vUcMwZ/mQcKvilfu
SBGlysBr2Rh2z4xINejmIU5rXLnkODW6ym+h89oLzTX2seDoI5LEK1CZdAL3Bnc0
QvExo74O1L1EQeX38LUtgTdhtNR7Vu2uE+ulitufr7NJb5ZTQTTxmRblVhDBFY63
DQjb6RwyqPrdX1CuaOIE6cVHEK1LPHKLZbcJwxzHjExeyU6wzTGiT3gLMhY0uBPw
J3lPNeRkouWQQ+18R6cAlBujovqbkUS5sVI3kzRh80YehsgbepcuUxEi8P4EHp7/
341fNl5o/vngrDoF3oiy94MTgGmlclQwl8UkPV74PFhynvT0qZ50yHqL/UJJ1OKl
gmZRwp09ZxpO4BsdZBmSdYJ0vCEmSMFdvA2nE/GKNSaLKlsKqbGEP3f70UHv8zE9
2127T7GdhePvBphwDhsE2GqcKoRWR9aMxcYYHrGVY3hixVXytNs23Er5sAgaA7B1
329yZtZCRTtHG2AR2O96K3S7GT13S84Kb/Epin5xmsZbUg7ZszxT3PH5Cotp6Bz8
ERg35UhouLLiuWDZ7eiPnyYIPfvuwuABo14iyCmX8B9PtcUlWzBkHCSP70S4Zoh8
3WOpVziL/oBOBLJBdtSR4veTC2Q49hvt39aFqjX62SryYacWEfOzPmxSCisPgVzm
cBVrI8W+pknZhYBYRoUZrmx3qo4pk/DDsJS8zs8MJA4qI4tVrLKa9YaRiNASm926
VKkPmeYylFPnrMB3anhyI6KIILXbMRrZGl/WGyyIZZh/uKxqYj3tZ9kWQqUN5fJt
E1gZh/E0S5IlR7+WaKdLbFMr/jjSw4cC8o9WFtZ/teaj1h6voNYtgsrw38Ezl/7f
fgkSNYaToZzVfAZrJF8WrmvBjQBjOyf1AtL5wkxXdPZyvhyqJ5I/+gsHYHTatqFB
pSyEdCdVYM3s7/8gmX5u/UVzb062ui9C+xXEDS1KVoxSDOidICX0yCie/Z4YE4TY
GLZoZtpIPGiW90UQGhBDqelF/n73STPQmrktDwvevlncw2FSwh2VkuXUY9Q7CE4z
e5mu21OJEu/c6UQl3RS2CvThJFxhebijx0zzUoeIZ3nRJxJCUho9i4CVvNyAKq27
5STaB9bugQQ4fX8E+KuANiXaxl3oxzrqkL70pLGyJIg51fY+ZfnLpPlOaGsTo+7A
Rnvayy4WSWohjpnTU1kD84wAO+13sYPwfi4mubG9EDE+QDwZIV15+33Pgg+QltLv
g2TkboAktxcIessUlcie9McUD6E1Wupy8fdsx0ZBCi3PmWVEfJdrm0DVRWEvw0+Z
w8DiKvtpM5sKFnIh92mzYrpye3xg9ebVOE7hxt47OeSKKKfwg6tBy7cg+9WhUDGc
seXvh3+pMlLsENnkUoaBQ7iZlitFOCHTUMIOO4IrEBz+bJqrrpFFeLBPjZtgKczY
Akr0nySOuQ7EPGLnyRtk0AHKmtyEqFql9u81LwaKAgLom91y0gkDlSIWkVCiBIjc
0pOM6LcNn90gCroGMAbBvA5ZkkHtQjrCEkcu4gPlCNywqvSrDMBdO0hp2xxUbGFD
XQOn1kfXihJuqiGrEvUQUot4/pxI/lrTNm6ditTpJXEuLCryJ+RY/ccfY0J7d9gx
/OTfRkpq/Pq9rY2fMLe1siFEWzM0ZtGfbqQcpBgZD82yDTFQQLQmcZLa9A8uatg4
qAsKK0tLJQrVqFOUvZdqHKcM7Lh1phLJCUNubduwbP8Bve/cw7W/V36zWO9qDbFR
/M817cki6Xll0PHyOlqWAtpwWMeZxj4+U693jty8J7607DGzJOEzml9gU6spH8J5
YgxQQdNRCQC3z69mZam+I1ttjcdD+YP1ZmHX31+FCtVnWnm0Ww0GHoBiMbpCzp2I
AoXw9tznP3xCx5FzuXwXm/0fAO83fIXZ44b9FB4TUk4MY/BEUyZx4sQk9X32ooyf
cxDZeJpPPuv8q/XjIyI8N9HcGujPc9Wlp2v6j+tKPyUquvXc+QLJh0pzcxRixDT6
1uTEFGOTucTDq10FV5MtjTCjX2U+AKAsN1ZVx51+HwcJn9ZSEOm1Oal9yXoDJ2Jp
RuchoF0T3Frclfy7oHQS4wi/ZcOdbgf/X93GgxtnaJwN2zePIsYrTi8w0cvzxriO
dIYKl6V98OiIQhKufbBe96+gOgngPzT4YEJ11rtuv+bDKHFfTIdE42gf1MwacNJK
ZTX616AOICzxNKtSPohsTqVKRCeTVcCiEKpGuleMAl3tx/P9fgb87JMzmt540sKB
g3YKWp32PeBzRRRXjVNZWQFWKly5R9ZiWZNpQWsmT4ooaqJVtyTLtDI3GlnGiaNR
wZwWU/rzHLK0brenBXbJpvZ7cLObcLMKC+9yPRiC3Es1bp0p5B1MUT4Wg3gtmnvh
RXQoeNdEbujPZBLl6hbrsKFVUBQHudkzbqUkj5begZ132rBqvJBvSCEFKhDLa8Hx
YVeO9kICdlLQk7RfOJP7m2vC6Le30hi4/NbtGjY8ihwqXJham3+YUnn1z37Y6BL8
25gK/tJsAi78rTL+TKDX/Km7jnSz8AQhrfANi9bvBcnBwGE+d3vfI9aqIX9oB0wK
cMY7hOP2ZLIjGH8ifiqo65XnZpdfDe5rkbF3g3/q8a5gzd3rYdtxfAQSgnC3tGF/
7A8+4aEcPiIIO8vwRyV0R3LheIFL7dn71HkJdJbuZ4/O7Za3FuSI5p57XOB1gd2m
RgFg2LzggziqQmW93AEq7TLV3UA759lq/SZu0bTCEYexqCpjR6oHmROqc5VzkkeS
sg4y1KdMHFK51E/M3QLfK1pFAvoAbRicaevwU1fggoqMVh2pud2GFvkr5hQNF58i
QuSjiCH2nT4bE70Xfq0OuQ3PCt9ilFCwGvOUGxtuTz07W2Fejkb0v/gWtkqir01J
0ImWMbgevr6b7nZj9Cu8Eq8bik3Zq8xVXq/i83IPyMk0fMuAzcWrjyetyDMjlzOB
62uaMAPO0x8AkT52z85R4IUO9cRvKlOAJoimDqOEViAwvVggaveqCQBFbbbaigSM
hJJrMOofU2pRDyB0XyUhJ3I+30Xbcp3UFkBrtFEo6wB5Qn75ZbtjaPpaJNRUYgs1
bBISEzsdmK7GMXYyccHvHLRYfWBeSVAyYXrqNfbTq4iWxxqRPmbiv/3wmgqLeh1f
lLX1nN1GjNGRSc+VRQQsxgs5a+M/u8JTA2//LfvHpas3B9bcK7CU+e1TUaxs/HAe
FlIQsWlR9oopjN8XGfbm2R8UN+QWwkgM8X2P8lsC/IdfrqLCWuf2tp1Dyc2PD+2g
pkW+KEqiMIDpfKlDoIO8DdMYsSgnfhFhM1RDuFjhw77k5UYUPVA2PSPFQF41Mn8d
hNgQbKY7iSM8P3bfJlNkV3MMJctj1Vstq1Q5BrwydBPMryY95r5KZeKFUW3P0cnc
9uw03M+Fej5rgH5p1L0ijxrUwUQKVgQxadn/EQ1EyVstG3LwspF58yEFp+k/iYn3
vnxXWOxNMF0isCyVTbSrtLe3cK0Vh/mKQwvfG2VIBK8rEAVs9p2o1bDtAuwHw0Pi
xnhCjtWpQfMI9DoBagOhk7L+zF3YHsSWTaDTtRos+SfT62GBNrJUQk69r4Yj4WX+
rpXLtvj2I9tL3YSZdT1cKn3aqob8cXRYgDmmIP08Gbkwzhbmqw+JZ0soaAkLWZnT
ZzCe34TIos2NEXTYxqK0hWLMQ3m1rvAoxWuxHPnoqZdahfTMRerycxZyKnNxkSc2
mCMJns69CBwvTrxs1MswFJIAdUAz0QaFCHjwYqqMsYdTdIIUjhKC7ntWfNYRv4of
aVYEMTiJd9gOffkf/V9/CqmcAJR4Ngd2MVGnxYtd0LUKIbfGq//Fe7OvBFFOzzTr
cy6hpe7czdo/BkvhhwYZ/MXVBm/2/crXE4bfiZy3dsP1GC2FSKGtRiaLtWONZiiv
52HLraV5J70PQyRO4sG9oU1kBtirqQN27SY8PriLVxxPuG7g8f7p7k54fW+UhpPg
/m0PoPw2sBUwZF8M04t7TC23ciaLFvulewYwUG0IgTS3sRyZ+JGsCO9prHeuPzn/
9iadIEXnWeNyUODCrBdRETyUpzUR3pn1i7dazmGQ8nWHbctOsRVsEch1p3yHmpzb
aoUzUbYa6jR+VdMOINwwm0Qb59kvvVb9ltovGo0D2cSi1hGGUS79zy0ZVMuJLuK0
Ne0UupV+wZyt3xphKY6YiQIYtV2K5IywFgztSdriCUlvg6QZG960+J6yFD1EKZxX
B2yWxAgqOT4mf+fe/fFpH/67PNxM3vo5qmhMzqog+oSKYRoP8C1DYN7IT/80Rm3T
fnE9TtcrORcIReapGZDwlulk8YMnYmsFfqhI4mBrqM7/jgRNJ9GWfJi4vkUlUNfC
eSKjlHwg6NN9coW3cugEhYBxvNh1GovERclozQ7zeGhsg3a3eTiWoWhBTKZSh5tQ
cwwOlPT/mEZOgJcSkZgZLRHiIh5LNQIkXHvmwDRtxlH4kTCbB8MA0A3kwTZ0J3CF
Y0BCOD12mwA9I9Y3A/GHQhFSGT6/T9ehNIOF5YdlpF4KEENWqAd/cbsbw22ns0cY
comklHWhLbnTVmMTE7JMCZDl3WgznnN944S/0C4/SfmVbqLIioF/HHdmwqrihzP/
4jkpQJuHPPIdHJryk+amupE4RJCb/0oHG+t1gHlhqMeYsglJWVqHDT3ntC8/7eXF
cCIidtXfZYLpPls+nrXcS+HNMSUsKxBno8r9/IylgM0QqCXM5F2KvANuJSudU20y
YAaf6PxFkRBc69Q966BEUrbHiH8Z/mvNPSp19j/rjJqbEDQiwJR3N+Ws2UnMY7Jg
DOsfiszH3ADwrE1u8hByrJsEC7MPYaYxT5gnhYbdLKrxfrFUUH6aYRnG/msWimJ1
6AZODfZrFBrQPFr+ffxelh3ksM3r4o5fRDHeZ/0BcEHEWzfMyMIE+Wo19GpUz2D/
WHhjaSvUiMd/IxPYl+vXCqN2BR7Pa6EI9ynKMRlGBwhUZFTALq8Pmt3DMOK4f1HC
mwotwU5UVdAkwXPo4l6J/u7NxS4cV6himMrNG87DBzh81uBkDvabwvSZ0BgvOSdi
2nr3c/cgox6Mb0uduOCZo+Aj2nV/3cxuw1IeRsewqcSCO8ilixcsf9BOmRFnSyYZ
mTPLqStKE1MgieQEv16jnBDzwC1BaJ0xgN6t8aJ1AQ1fZrBspDFC3LjIgnmcXJXd
a+uP8j9pCLLxdiAVUkKgROFHdzkcozsOiuLDKV/JHTLajvsuzoooQ+xYA4uraFwy
nQTyBR4Xh4dDde6YQ74Fp2Fk5ioLPn8V5JdrGFNDE2wgXynBoVabPnVQYcyphT7V
xEQWw0AkNUnBdPywDu60RjgvmbGATf35QAHV56Rzg7iHkmEPc6Hw/Oah5T4eQhyH
uU3rQ6mLweJC9cxv7w3c1obyLCQMkaJJLXs1lkgilIa9XZ0dpVayQnl3PITGJ+DL
TN9mjfNcKUPOTzT/vzMKkeR1K6yyx2sVwF8hz3LMionPSvxFdlpsxK33OxGQip+3
GKB9OUxcaYriXrks/17XleYHrtpgIajxqnlOZ5a9GnSCzl7SP7DlvDC0cUod8SKz
Oqho6JXo4mLZskkcv45mzbnBJv6bLPsiESOay/W1k8Yps9n09F3Lknti2dSQpvcd
Zh/uBB07RhzyezMKoCETGprKL4MS81SLWUGTqh0HJWfwhcoj3p0CdYyFgLAtbo1/
z13SmWedzYn3vSwyJfwfhAb4Iz1XUpQigEHzodl+nzs5YyjP/W4DXIvGNrH2GoXT
K3xUSilU06BoOorNyp45/4vpC4huX/NN4OsG1O4Cec4nbMAOdf6O9DChqrDCKrRM
ukyrr7aibyoF1enTQWm7Sra1vuJlX87Pb+q01VnPrX/gFujKehTgQQluOrnIEgyL
/UAPPWK+FKy9FrT3pp3Qz/fiiO6MXzQsplKxQ2ht5k+YrIajE7mb7bZH+S76o5Am
sqoi16Jf2bRk77fo77Ql1maKAnMrt5QK0ePIFRzaf5kzZBpP1SsbSfudwK2kcgUh
ptc6KOQCZHHKrDHHgDe/yU+/YeXd6bls53Pjied8vTo4M122CDz7qIA4w/DAcTAs
mZJk9Sk6UQTxKqdiHYB1G7HFb1dd+jMxBizQPUij1JE1jf8/zZtyUDnrjkQiOBf+
h2qjNYeTt0fUQ/C5jY46oPhkg/AXm5bD/PLXGGeuod8aPVpTrfx6R4Av5xwSZ50b
M+Qj5tGi8ICuEZ241FMYMtL1LHzdsa1kcAsdLA8H3DvlaTX2zd7bGGlG7eCi2NC6
YwolsVEdb8JdWY2/O4arqLZb3nOHQs4t6teOxhLzWn844JpW9ZcmQHnBwCWQNJW4
AvvbNBnQZIKAE9enPVzRrBtyEGGFwM1/fycBi6yAQW7kM/Gng22KuJiurpZjmB6z
edt/bwWGfQel9TYrMZLR/6DTKsA2DYj6YDKR8Y+RiQHnV549XbJELYo3KQ2lWRKb
KwgYUYkGPChKsN5ByFiZTm4zo0AgUHh5h4REPSoGhyVvhfHuo5iWq3ez9dGfEgit
8Nqbc8h5zN6kTXF2f8edPakU7jA/FJxuYZvL2BWmdHqsKUxTNEOA9D0Fagajlgnx
wtIVu4IjIb2MNra48ALziLqQ4GNv30jFROAeitPnDAXjJnS7/C3RE0qIPexOecPS
2xCEEp840JCBfeOVjohUZiW27HY2BpraOHfiBndFH+vv7j/sb08VJJcHh47fNqog
w6D/f1wGMZNGcGSC/b2lVnci4iICYlAsUQsGIehx0auMrD/GQAfintzLcEHLrAUI
qX5DNFTpdlQnsweQq/AWtQDdSS8QQISLxD0nxuZJdPcW5EcKXX3qa/E6mKIXMYYu
8Q2lQBbzsH0HDQfDsX8V3zbCgRZn7jC8imcYYLDr8uYI+HoGv3/damKufZQYBc/q
eKMgWZA3afAFSv4shRNSRmPeMO45r1oeXRLjHIUhC9TDEFkysQHCIbqI3nt8+Ysx
/A1JJqlNBnG18Dt//bsOwUp1HLhOxJaqyNefwMUrpjSyEoyf2j/ZXRvqdQHKtt6D
Xe824bQocaHHcKy4DhOZhlQKKR/PCggjwbwrn8q4JQa1LJKRsn9AzvY6Lif0DpAS
7nRdY7sLIVQ15/+VbAo5UaIHfR0ndzyPvQ42OAlvo6VJ+svbWCqMZC2sEkIbr6Hv
obUZ8Rzpn7R8ldfhreOBavl8+TPan9XtyVXiNBanLpISsyV8bVAG1n10wqyuY6Fv
O0RAp7GgAFfFZCRl1wyYNwvYmrVKHarf75RUEvaBR4lwMR3O70zR5SQM7TAyJ4cf
6wF0vQo+EobLs6J6+Z5OutNyIJOuJ4ce2wMGG/qd59QIA20rT9Vrg1GuzTaDrFlV
W9b0TJGLvFy7HZI4buiuPexRiJ6oKhLK0rJwFnsJALMZ4TSR+QU+CqN1X3Oo+Pff
Lj8q1RDzDMRURlPy415yAVXnLzSaCgSdgFylRRmYSD5lWB+mD6zpZdmeJdz8Babb
gt5B8FxOorR7kiOxH3rK8DIuYpdG0xOx4e+v4rK0BCaCJV4SliktdGOhXydwC3J9
JaUMb2ilLIXsaw7UoEuW57OqELlVvqEHi6sGhsmfCm5bX0zvcUIjOieZblboZHiw
hngD2713PmGptPncgLigXs71M7WkTPFGSzruUa0+YSoAaZsLTxZ1ZjlNyPrgBfTi
wxy2LAdwtbK87R/f3lt9H5weScCZmCWpCTtkKXxETOHADRpaRKueGnAMRjyky/nf
M0xUXBh4GqM8qRWQRRCR2ofzhNEBF7PyUMZVErW1nFuIvPv3xx3Oe64SzeUMSssn
iuibKfPqM37ttdY7fEdVn9JD863LfIWMLNVBqfNJ4XoRZl0R885pLcGp2Ji8C1xp
heWSuCx9Q5569N/CEOosiNEb3mLSlbFCSj++F1z9RznIi6kokr5j9sqB4+sT2wxN
BwAc/s+GQ97pX50ntnwLhyitEEkmMi/WyMQ0d01FI6ffpLwllCSO6vhcaV731670
CiMDXo0FjbBp6sXf7LjjHOX1qMYl7XF05TgVXIwCOzsWW/eBW6ug/GfasYuyonsH
BclZwR6AB8x26hoHBX+zDOxjAwuoXeolvrhrvQa6Ux6VeujCuWsfiymX/8ulw/Tw
sQxus/PdiavWgZUxAILsOTbrN4gtiffgrHNR3meYwTh+2C0uXEZqDYimyTAiCuqU
U0jGDx+SHWVRhBFdvaeW180brEvECtg8fXyNtjEyJF5aBE0XFc8GNJUegTXV2bvt
cHPzk60IpT7o39DnVeyXg3xVG+mcSRluPUwlV44AufGkIwIlTRY1twCaM6Xqdw7l
xdKeqaQX8zvabQPGGQ3B96mZsODeJpazgHzZqZCqVQiNSUACL0/FzKGnQ1ktpwOD
nhAwY++zKr61hy4/xllC0BBvyL0wnaogJZ6Z7DulvR+OpHRrVxxzmlUyYCVQR+rS
8wAYAEXc5XnLpV9NxH1e1PBZNHTfouLnpaVzmD79Qaa4JiGEzbK+tI9249Ypmdlx
H/196KpSn4GBee4diykAWF4KwCfAtEqHhBx2kRpeVItcBup0rQSDn6BMUxlZezJK
5ObmQJrBQ4TPI9Fcsf/t4CjiRP5+UZZRQ9CdXsZCVOCF+NdqcdUBBCizAA5O3GTq
dz1v0MKEbv8iRCf2bkvE26yp9pHALHcMGt0VcUz2hn5BXHRxKA8a+irucJVeGWSE
U5iEKHO8FvO43wD1SdecDxlJe/HXRINOCVA8n+ca8VzXbyJjJULLWKxKoVy3/KMm
GEBe3/h/3h26nBeDoaH0bGgaLM5es7PzXm7WjUtpwHRJLmRMP6Fme9x4UnB1IHMt
K0fkNel3hvObUm5TFIUwNmR7lRa78Qh8FQUEfx4C5p1hZ+4Iz4jBIDcIU5LAePHp
J5VkGMZOMNWzovOplhB21GUxThfCkvxLaNTdNqnCxoOWwRT7r4xxMKBI1DENX/P6
1ffEbjk5D+0xxo4i3I2Vpm/AJT7RDY0XKjzBZm1zOtjq4TjA/hmmgymI8WJW2DsS
GqmaPqWHqD32lS0f5j0uoOljB4kxw8crpV1PkpGj2LBYp7InbK6FcJWk1X906faj
5UeAzamvnCijC67J1W2pQk8Kcp+XcvV222BpjdL4cM3oeyXgUjMG49fwQ29/NUVC
iGagOUuTnxU0q3/P7IrMSjd3kf7Lu/Un0bMKANjb2lHs0VjD2eGpLwtore101fKy
x4uxng+2rjD4zA0WMiI+YS56OmbELFlAC3yrgOT3+7luo/jKbFzzipa2NhVJcYXf
xDmqWHSWaNPz/APbbJhA87+x5lVix6HZVwt4qp9/Eb+KJhIKG1QFnBdB0LXl/xZv
D6+P3w8K0WAatbVJJG4JD+ExJ6sOUhFrLJCrSYuEtO/ttN56VhrCranAYsQdjj7J
E9Aa7W/QCbt7Zv6XwvniCKnPrCsA7QBiRH/5IJS2FkHe0boToqSeNaeIyVV2GJXZ
IDzsBazPNsdb9BgpJeypgjMUSjbi7qGJ4AKZbEp/AQ0zdSad4h8pfsFpsVuDm23m
lWSnB7QZCRMrEDgYz1FPenPHVFAxWo186BmLOzLR6ncEQFelgLo82kAfF4Mfa/rL
YL6A5aQPzTCf5wldNys7HY3yY9aPbWBimTxCFznQCByNF7dp6nPE4anQr3SjjS2j
nsI2e1ERcJaHgLHEpp0TaAEPJmyP5VwUkIRcwyNvG9HqKWt+8PmBZvWWTizd5XD6
YnC0q7Y+MOd/7DLuOj6r1e71vozRJNGy1ZQ1WWlmnHA0YTxO77LTJ9Rav1JbbfTB
/QTJTG0hcx1d/L1rRMcj9R7F3C8bZeqTsjjCCLkOcmTwrPAoZ/xtNrs+Ky2DgKg3
A/zJFPvhrr8mMfzQM41ttH57HgBWKE4zQdBncW7MY93UcHTMddH+IywWg/IVm91T
+06JQZDtGIpI2t5XI7lKMvl+zWLHFvKEKdcRO1D7mA17P3Ycy2PAqh9haKWghclg
IbweJalw308V774dhRMMjuG5QMov2GGsbtRv0CgmGVLLEIPhkV5yxr88rkeve7Ex
241qd6LGRuZGSJNL1QSlfIQN+twDzMpOL80w6Q3le74k9onJEHU7CSF3k7ge8Hfv
6/HYUvwrC59duULfLKKjEQzP6WeS2WPflYUaZH4uS6Rih5Ap76eBceLKE+XWeoZL
ANTLeJpKAl1MpurVLSHWvzQlQZJHqGNTD2tFXOceAYO5MjuoD+/wT/u4DmXvStmO
HMKTsgAMiouHW1bc3SMxxGNCrC+tCwT3rXiQxTxahYUtr965f/a8JM0xugApevyA
64Mr9W+CQCg7HDrFVYXmyB/NR4jcJKdY4Z05cmzNPkUG7PKh+1jxq+z8ZOyy3gHQ
GHbxpQgRw9/Qr+VmjwriMKAaIWNyMQ8+5gxwNwbvX0l4LMzX9ONtFCRx0JB9T2lu
xhV/rb0Xr6nSwKy+GQ/IheVrHWf13kJZYakURQS0qWcDjwCf9FHvntcr2SE8mmnY
WQjD/TmZHOXp2Ga6eaVogn5HsvVPmgdbiNdigntFf60k5khr0I64Q7dJKy26CPdT
5PviEYStPMA1G3cCKIGgFP/hFBOc/tMraFav7+I0lmVa44xxecWjwai6nYC2IMtF
/XAOa0sXO69CPPiL4ljD6fF10V8jGDLi/TmUeCBLp8ORXmEG5tw9wX0fo+oaLGqD
yaKus5Gq0LEld0WX7xwwAMTOU/6sEiKLSeJ7dZdnGv74DFFCZ/pJaKZnYf4djr2O
xhLhmvBcIoRa45l9xxAPYNZJem5iJ1h8mE3mEy0W2qp+ALWAIQLa79FkOxqYJy3c
cAInauNOaDb3wQHb0bC+3T9ZOM3t+Inf0uuA5GJnihfmPBXQZGziOD/PEkSq3V/W
sJVBLzwxuRcqIvKzP/VGRjQRAf/XOvBKjZ8X6xKzM8lo+eQQBMhkSKK35/xFcZUE
vYI96P46/eQSuTVNonTJ6xfiJBNmptRZlVQYwcxn68gOhX5+c+ESDuO7ytFrfim9
8sELJPObEXK6eU1tR0tqKHtqXAsKg5po8uBXYnMFrFX7cDDaGcGFCUY1eYtkROBZ
1ZqXefEQFp0n1Bw03nQlYqSzCOfRSJGD/b3bE+QYJMy9TxkjbH9TJ0GeEeFhL1jQ
1gXuozRI5Hoyo5vCKXpk/kwFfn/aFWfaRTu0m9YWKJo7ZaivawNYELXIncqTBnnB
FClCRDfeQrBNp/kismv9K4juQjQGpKMxs5UHKgjmYvTp9kTr73mLQtpCUPMOKHrT
XgAWnxLWBlF5OhOXNq8gK3a3WZnrhJhxjO34QpRsP5j2rZ+bLWk7YzvhanM+xpI1
X5OnYldhf8x/aLYP9983vwLmLfWyLyX23mRIRZhuW2auqku8btLYIm9WY4EhbPo7
SYyb0c/BUWNd/u3tLGwwl1osid2uyltL1k78vEgK5Y11LoNjrITVBDMMEeMMsKo5
KH8rwZlKbrm5f4DbARFkyIvqOwJeWqzQk7Ti7h/lws7gvZoFy+LZQ8H/PHODnEr5
3AuazGxSPaGQPbwxkP5r8Xentp2iWPt4R8UI3BzOPA6c1P8ismIfxe+4wnHBSV+v
XZIWgusg9LImsiCxyEiz5f7SIAUX4QiQ8sRuvJi0mgycI2cIYJLgWDqf4hYdwnBr
N2t8bDO9lrqhiUCgckwd3hrBS/7bXpiJ16W6mDwOw3xLUW6neWpz3KPifNKNgvd6
qYtZB0JeYGg0sQOC7hfOuvwYLNIe1dWe58su+xnLvUyS55JjgqmN8SoEsFp2+vj0
dMQgeMwM7XjpjORDI9p4+9IO/fifGjyla3CnHtVT3OuMdOinvMuzp7HUTpCh33JK
UVA4M1yHL42OjmAqvIhWitiwthULdAhgJsOjcQzc8MdLR8e59gS9BQrSKYqiM431
8lP1z3sWW4qzBGHAiDs1wk/KK66qbl+W/OXRQuOsIfXBlpZ8HQ7l3FL55ZPDrC9Z
nx8Mb0Yn+oyZpyUSq9M2SH97sMdc1aVUE6of42X7L5nzKTam/xoiNZN3LBE10oyl
TRNFSgedOHCAT4x/2T76UaRIn6/SN/ZPpiIhrJq8JWG4hvmeaSijuApiBHU+2a1i
fVWbMEIs6V8w9xTxCwZ8sOZxPM09xXKbAposZ1CziYYSltoBG2utitib2v7fLUuD
Fihrr4MCmSNFDwuJpkm0qKWqbVxiI59RaPBcM/6lR+DN8hWE/4jeW59X8cgti4Su
/wGW6owl1fUst4x2MON/+4dG/Xz7UYjd4XcRg3ITvOrowpsedeaZYNFsOoHftj21
ol59V2gLfAPhGu211L4ofeIBgdhaboWDEZZVxEsZrvhAeNKiv1EiJknlb2oANJha
lOSTHpgPdANcADq/ohFxqpggUYrAPc5cG2l5vTrecLarNNLhUTOqdQJCOTePdFlG
VTwomxCAxMBgQYy/CBcpXc5Fd+r/O13QYQgIHsc1NTHfmirUHaBaA11FFubYciDK
0aZZXCKhqKZK65g73kjeezcrHD0rcadmOJNij2MNyEUuWc4DSEJWa400fBx/KKql
62ToRg9AnoLVQZyO37ewHit1Dtv9YZK9rKamXJIXnnqYbU+C8zw9dThNY/TVYjob
s/mjX1TiUS45gI0iFWn80oQPbs9nN/KDIGFJ9tQ0kFbybzSu2AbopIno/rhC33xM
diGLtE9J/G09SIPvqBzqmi82UlCFA+wR1uBVIkM7nvnTvntjvMcotC0OewZwnVGi
PkUu6AWWMY/f/EucSTBd4cidCjeBJThwmSdIGRMKTv6uzlDP2yI/7Yx+2lLOMoMc
Mlxqe1ryynwyI3F3BPSW+BnHiCHjtI0FtfNLxw1BuVhhY3GUnuihjKgS6DDQoPdZ
7w7Nc4q/swJFp8zQhL+jz63yWfo86hD2Smr+mVfa1pfCnXaaJE/De5txEUen/WRH
5nZ07+k5WG+jduQrfTUl+mFocip7r4jO+pVOaLv6cYFOuqlfGeZppJpGnWxANI0o
8cfsdZB1tkt/034fLLaeZPs3QoM4oLg9qHr89vc/tMN+dLy6t2hNzcc3uZzWVKZ1
m2iE84epephyS6kJpg7K8cf9stSg5wyA3Y/mZN26NcOXE0WseA9Py74a4TcctfeZ
ZDpbDN0DWPrjUnIS5jHHvQ4OeGQpYAWGaUxBHKbwAQBbA+phTYPTgeHZPXa1+QTD
9QsrSXKg/vKQGIy5YDeuWlwOj7IVCWfRGuw/eVLPTENIu5kLj7CS6aFlA0oKTqq/
y0XIB6SES82PD+fgZzouj67+axzwxuq6e6RMRHZiKDOea/izYLJgi/cM0xN4eMSB
P5in2e82cbd7EUWE7kU4i/J9LPc/vGZlrMQCmea1KJhjSEvXFPQeyoYHc2GEeyb1
BvdzH/dPbGulMfLM+af64TdDjJvmCbKu38NwHIjk0w+//UAKYGN3goqiwEf1gQdp
zSejE2/rC4ghRD1gegfEZAixJlzuDpy7/nzJn11NcEEcyJfMhvZEJA7xBVyPgryp
w9+O/Bn8BUwOq/b3A5j0O5O/e3I3NZT96o0Yd8NTlrkHyRrWJvpLE0MpxClfwesI
oSIJHGT4weQCBgHqavzKfafgXWE9DbTor+KutWkEQo1WK7p+P8X/FbRYA9XUdFPq
WySD500fM09/Plh5aH1Owk7aWU67EE3/fPLyyZG6SxVNmH/rg1Cv7y8nr2Y9rBbJ
cBejl9MY34x/DsR6g4CRixhnNJtRSbpFUhXO7eOhm2SBNGWoX2Ic3nbzJXwdBMOW
PrtNQQ8d9eeFBv5pnK4zssJp9twnMWUXIG9/PgEMhTAMoHiCh/x917HzCASALsHY
X1r9WBTXYFhxaP59wfkPkndGlB/Ca+IV764Hfa7bkUFWKVjoVgdkLJk7faSAF2H/
9XVoqSe47JrvNA01j2LOAutDtGZrpaLQgUDBZw3gic584ZgwXovOW1Ot9irU4zTT
ml7oV5mVNd7/vy2pAjwsHe8FxqgCeUXb2nFJsfGpGsX/sJhHw96MhKtEF4kDDJ9L
mEp95lj0irTvNYtibnaDS6EUALT3FMhzktv8JGcPHV70h/XaRk9pUsjdcfAoeokm
8vxNHgP+58qrKRAaHHhK+CxPfRFEHPb3dkL0bQdLltr7w1VMmQXJ6rluxO+kz9B9
BQYn4G46nMBwe5lt73IGssOfeHEoPjkSqKJa+12RJQDk9cdjq8fbqAejCrnJl27D
nPrCa8N63d1xshgMVdrGslCfU/981kS2wd3LqnrT48kprrZ387aO0M4onuO0rZTD
pqrU9n8TfLi+LU63NIOb7bhhjg2gqI491/vr2T99XT437/hhF0wcNqgJDjvF/OcO
rARDaKFLjGgjRoLFTB7kGS06tmlFyx0pzwGG+WioH6jOEWSY40Sd2nuSfOZnAlXW
AhWO5upr1zvHnrIfDl8cG27yalxzsvgNAmA7wmiuLtHrqeJXFHNPpZdDVUPEWSoL
KtlBI13xf9iK+gniHWqso0zRB0ABhAGJcXMrwgtCO/a+w/rt4KgkzbhbBg0XnOFu
kssJiEW+3tk4Q5w4PKtRe+mUm4V+IqdBAWSxsCdstYTBeNe4X9N/QGKyHEKzkENp
urogZeaSyyU1mmkUtbzhzitVA24ukQk405zq2XhAMStAEeekQod1A6ckcirX4M+6
UjYiycPnZqHalTVfsx0aow8ypN+zVzCTsUGSzRoId4tdNjcDSBH68z1zCGCv3ZdO
Op6F6iXkRrwRfC5NLua2GVlAs+rlgXx6QcfSX+9GwHybDVbOukmzwXJNwvxVxX5V
f73J1dnSsX/SIFehBdUIDIc+c74kdzHpbA/nxsOwRmZTtRf0jr01zcdRbKmcm9JD
FVpcMM4Cf4/QTZqQ4yPie+zfZqA0Fzqdm54JBSKvLQaTrrk2dd/WgDSyWn/xVWFj
lY4EaGb5MdfWyDNYeAXWV825dfqzSYyXn5mnMEnIorzcgq/lyyy9wyaxjjuvdYLw
UQpKrNPuilCf8/NWdAG1Xib0uNisNL/55aK7wYanO6a3ke1jj/ERca+IElU4dsM8
QOT1JXgi7yhDoDXz4XN0VvgCkQZ87FsOnblCNKOp2Yn/mb6EicEz71GEAoHrWdi5
XVRoWloHk16wKXevnbzNV3Ma/xzSv6qzKIGeGm54YrplLQeFsGIu0uOiQXVm7uUk
yhzAmcnkQtSrTMnX4Z9CjWynZEo6LHA0kF9U/FQtk87CfpX2l4bxRB4cwwLASIho
5sku7KGnqfa0XatpIUnYNq/ARckgU7IeXbQz/G5XDESUrOxJAGBfgCOCAB7uz09O
hLlL4XfCiLx/SmtC+NpuMCQ4t6YVB6fCIwvqHf5OPF9/PMeHHiruu3A1vFJEGbA7
Wa6VI4qseZu6irT7g8HSuK24kIJt0UNWAmMiGP9BHSHG4/FQwgiV5I9eIjkI8225
1PD3FCChX7FKnNg01W+dz3xAVssLgCTzg/GhK8vZwcLTh3c0a73wpeROtD942HCV
9OVFDiaJ4f6ELQznCCf0vZHUqCGaFj53u4o8TZJS4v6tHARa5E+6KJCjpkvnsCLL
gcdocU8aYasT3vjTTUgReoiza1gTIN5rXo8KtteBGwVJCMNoe/aR4+pfmCIQ2q85
JYyNUb40hKU/inuItf4eFr4UPUPhbCkSMJanNOQBMQVsiuha9YSXuf91kcC9DNAx
ButrMHh0gFtwb4yzcPaeBnU4A4dvw7KU3MDgIw+WuNazNSDWUGU+dUG3LIO27BfW
H8wwK9Qpq7q5vqbycMcCGFz2cGuoj4m7bDGUm7K5cPmGPGU6tDTnj0mvJtVuwAoz
XWW0hRoSGS8KNOagUoHWfzV1IiWy7BpvMAkgbbTBo3nCFx4NqCgqsFZ4fBkZr0tu
8QIuuxxilYG49rx6jfEOxcS3EbF11JM+c59UEcLx/7wPP4qpW+sU9urTrcrH7YBy
NvV3Z8jOAk0pUvCTHOlTxfkDl8znxp+E8WH7zuW3YyiRl+DkIB8rF3jWc8nIySdq
J1RWif4EWYTeTBWiTy8sulHKvV4BKBBLO8aI/1qkuALt+iMg4/ODancRjOdBQgLL
yup5mJenhw1qpsg6xfvevdCuh0sC5mQlnh1ubKjcEeHtsulofDL6PlkAQEm7i7eO
oSyl7mPV1ajqtQ/V7NPdO6It0edxekGVRPqqr0ZGXYjqUAGXxt3DVLxb8RhFDXry
gvUZD/5uL3xWGs74ZX7kg+WRLfzj+kbHcHroAi2jsogsFjl/gU5vSoyABpCIIPA4
ujqk+JEd1F9amYrBMEKu3kQ9cmLkLXGKb0oYfLwMyaAzkU+4xlkF7uHZL5WT6529
zH8G7wVWejaj77iBBEm0iZq2PpmsETGZKChmi3tNgcWDzrUu9vuphAU/9sDhqygF
IpT8rREGKgrFU+NosZXxqGZWjSe7za/VYl47nuZbbYSQxmjFYo8Em+05DIzKo0EO
56pbcUnS4lGdGpq62naHjOSOUwZmxjPphVO8cHyqIdaiGg1Vn7F+ScatA/vzUj6G
WwedtP5/51KgTzSkEfW1uuSbRs+I1AM4n4FcA63NG5GD0W0vapvUqNEqeN+WVgVd
eUrYbW0kyA9eFbTBO3EaIurF5lxwtXZ5nGbdzY1krNT82Cx1RuE6Tn9ZAamqoZGS
3ejDax92sSHOVn/CkQ41Wo22cmaxvsT4uTZloJoqXX198SGizyt+ppzwpmiZSObq
0p7rD4zH7Ocd7+zQZa1uXpxm2reONKqWPqr9Su5lXIe+g+ncbxm12S3F02cwkgQw
FoJ/bKmlIN0zV5X5q8Tjk/m/YfJdLkZKbzv0LscyDCznexyh533iy9aJFBNnx5pp
cj4Jr/vKYpiMXnGeAJiKOJ0btqMvYJlaDkvRKVB0SxdZccS3W7qb7AVHihPROhN4
9XTLyaCJLGGia06KkA8gPWJTDE3U+CREuPptMBHRXYU1j08coW0SFbTRhbr3ZvH6
3sv5CcLKtL9r5Lj88pZIeDt/Hu7Zi/zirs5Jaz8VSRfqNitODRI0Nqch9yH+TWd8
PDW3X97JgqTiE0oT4MWSLMzA8FGwT4kRH+MCyVNPa6bKt2z8aynIBZnHQKu8GdlX
mLh2p08bq09guGL1p4edE6B97CQl6qT/letCQDCyscn06NoJiPhG64RgR8iB+vN4
FLamShbj6/5GtL5S41Z1T7yLhfVeFuo4VZe3vNf1RMXbuu4WlbOk5wzittlv9gEb
sK2LKyv4pSSi15CkK0PRFQvRL3G6/K+qP5/HMYij48d5YLsZTEBhkPzgoDlVVd5J
sSUeBOTYOE3XV5DvsImU8LsV9A7lqNIwdMK3SB8ZPNuKYt2sKMNUVzEEP+GSs0je
g7wCBd70kKWBzBT9PpIIvzU473YqIX1saKZSuT8D8preOz9cOjhP2lHGOSZ+DWBb
6hlovhB24sYNjgcNiLP//xrRu6oE27Grqx5OV9rNQNEvkqQZlLSVgCBJQH484k/a
+VK4S2/dhsXP3ldw752yQo5ufo8dP82exyAXXbr059ECdZOV+15iiA4VQ7evYL6L
3Fm5/mEaMKPO8tMwT3E5ZwNaqilTdvT4sF0uQlCvC7k9ACuB9GCmSHREfjduOsMO
qzJXW6KU9i92Q9s4tjTTb9dUvSc0pPpb5Unu9jNQu55g+Jjg1hTSd1jaR7GKlrvd
eZv4vCJQ1TM+4/n4hvfWfHjsK0ERNQREE1ydjvBsXd3H9KFKVz9geSh2f+c5pd+v
6HQo3Zk2HyWy+ezqWnK809W+pS+v+SYXvNveWyMELZHIar1KvDT4BEBD+TvgI2F+
lWj54In85uoLeB+vWn/BmhcRoHG5np3/BLrmyFDelBlK6S+Amgmp26J/GFX8IzQV
luAw34YFx3adiZK4/FaNEqWOXZ/P09moJFlmfu/QoOdPhK1uGTZ+IEsr7zXyHQiz
5RDuKY6AndLnny9dl4gfwsvGCQXtjG+57RCpqPJs5SEG+Fl6SfyxojeoroplxTBd
DNoV4x140VMtsGdB9UnChF98TrfNaT262fbOdS6NdBWOF/og/+6myJpmrOBxchNr
v7dPojCFDgDLZeWjG14N5u4Ha/Vb9KhM/IA+A8VwlouMa1yN+YaUdswO1Ggllhap
8oVxM8b+esFfVpBEHaLYzocDfxA1SX0Wrb8jXsNaLgFqv1BY6URS/Qh5WwMxHaoG
mtL4oJwcKlQNP6n+SKPnIggo/RctZ5NvUlliShAgmhDXzWFbFOnf/PbrHHz3um1N
z8GoYuxG/OaqkRTl3pO3ErgE9FmCUs9/Xn64zW2UQu8/+J6WAxfBXy43yx35QFN0
SuOsytAo8UcAbQg9aXfhW+/wl3gBHTDeA9Aua7/6vlVJ9ejz7Hr+v+FrjWOJTt+V
wr5IsC93jFkQtMnylqhwb09jsCBwsRwK9rFMxkXZDi6K9PTLNnhGGUB2Bkg+sPNU
g+GbPqpe2r8cO6QM1Uu0yYVmVIsR7Kmsf3+EM1ylc9VoJzN0f9+CA3MZ0NZhROE3
ksr040M02e8ZoUHk4jqiFHpLESPV5gkeWh/JzfCHKMMoqYbdx+SbWvMjPSIMwUFr
nxm4Ruhd0Lv57wTvYKXddqkrRds3jUhlZcf1oCctV+LUGPJCV5T7Rs37ueCRl5MM
0hkCLk4FDzH9plbdSJtzEhCogcB+Kz5J7JZFh3DcmpsUF3q4xu0C4Iyi2v9z9vqr
2Jrsg1XryRXEHHfFNeUJOllunug/97z9uCDAnYrqgNb48TZslhUK4i/hOSsvlIU7
1HCnKrAP02j7AGq+Ba1CHy7LWYvPa+yySgMN7dT0/MjDG9m0NvbEEgxNd+wBzoDp
Zw+VpHy2etkdXD9PSKTBXY/cjEnJuPJhzRW2l6pO/8HVreUo6xQN7spPtQWdNukT
di4G6mBQ9G/B4evrLsvjsNIFDnin8VQZZ5kia0rayz1ylygWQiE5OktykmpghKPs
79oSKMZExeZyZFVKnEzeLDCCqgiiDXbS3H8nsO8gXMb8dfRQtQAVqO3MrT0iU1hO
icmb3UsZQjBB3LE8ki4BNu2cscAs6AfH6FmuXGf+GtR+0devPukM6qENZ/B8k2w9
Syzlwc0MJZw/f9XMPHI6MAlQx5GUr8fsoLMINnaSQUxO4Dhg+oZ75/T/VC8k4kHf
NyjmdIGnowTGn4IuMLngzxMS5BlK6eYB2taEHDaqTCc1p7EfPAMKut3xbFcROhYA
ZHdHOcVZxgKXdTo+9uI+Av67977MvtVTyIDFR89aLw9p7Y6KV2koipWRwJ5gfveX
xucDdEKObxjmU2G1vUFsXek560jiiPAK2ChdWmtUIktIOmbjuJz6iYFwW5uPyunV
zZZ4wjhDGdT3VtULWdl1vAd16zwUUlLy+ojRiWNqWnxKT4aRhy8qrR5Ybet/OVyc
afPHeZoyWiHt7mP2S+3fcSebkHeywBWatYgT8iWdZz0Mq491pNOOS2oz3ob2vtTA
//zVOS/htJYEqmKH3ic0DtX7kUXnhLkhF/JwW2vGuq3j3QhjBEBu20LwjiwerOUr
tkoLnhW/YDtzMMkywoSqoFsTmZmymJpYd66+Wd0iboPhmQu/Y5QXiNY2APSJ0sFw
CqQmmPEp/uy4qhEKGlv9Dp6hhqnQ/prBYlc3v7xXIawsyAyU1ePDasiH54TRiOey
assnpJga2w0uwX2y6e2AjY2P4f9iLE5yE6PqeDzoefFm6PQmWZBIMj+gyr4ozbc5
4TgPaVhYQQ/+2iJnKO3rUqK4KDB8wQ1lCoe68OLOfLsbmlUieID2Yhm6XjMEi5ju
MJfyrpE9uHRjMIKrpbWxcroC2vC0RVM+5TnWCFVRb1tiET0q0yig38RWTHdj9oGE
tRvG1DUleFvq7n4JJw10BZCxFqSwy5leD7cyVcWg+Hqrb31nWTKixW78C8cvHKJd
QJtZR/3M5PZ824O0jLbNJ5rC3sm4s5oRHPCj9TbWqqd19DWcqQ97jeKBsqc/t2D2
78kmwl+DSSLbXRbTxXPIa3eLXqWi46h3bSZXAPFeILfM76iBYN1Zg2UUXERtJ6G7
PG2v7imzfgOCcMRycU1vG6ao0whG/Bz33OyB4FYkOTlSxIZWyzBA7oq4q3R6oZt/
eP79lnqdjA3ur60RoP1m5Q1DPwuZVCqaSry5AXS/+PmhisfHzaRjG1ldG+ON+viQ
vQUosmKV0FTXMSNxgk4jGkIlbAXRVgTuq/EHt0t64zvjlzihRDUakBqEGJQDPhIz
Le/Zs8QbR3bHtvjRmg1xTKPgeYgDtNX0Eqq3nlnkZRa41tou8rJM4AhBHlLRuNLR
tDTwRsgrlM+7K5fLPtWDX/7u+dfTb9cFE3S785urzjakC9jeoiKprirwrq6vw/E1
Nap+65AGNcx/53rwFk1wQmmqTATF/lzrpBmfCd7z76sGTxfOQcI2jpkQHXcOQC2k
zCrF1iOSfEUMJtuQ3wB7WVHutTqOgNyVK1VKplmZxlQ3qOiaRZIBL/HgpNVLucij
98zSEXjm4Q0cUXIBmJvwb920pge1TiZoy/ijsb0dHGg4YhDvW7haapdzXFtljy8I
608EDoCjIksXl7iGbS/yOpJ02XuRDfA+U3hzvSP2Y8ub4LmQv8ZnqNu+3pyU24DN
ZFyFhseP+jxWAv3Hz/gy2DpaadnM0R+uY/lrl0cWGGIvxyJTT7nQ/xVd5tkEORjf
NBa1LSHb29Q83tCJLOZugt9lSLxpDbzGVF2M/yGX5gqvHoV3bK3FOkmF8C2NgWXI
i5wd7pTiEP2GrcA+PkVrMXTbPC9eAQSDp8xvDUjj0igi92J0hUeSP22eA1s3ZLIK
GWcOW3nBhUJe+xHB6PQCM2P1svw5lck9U6eVp9GExXqkq6vCB2OGUI43iyjbrThm
+itpYkEz2D0gelGbOIq04M46mTeAUlmeUBJl6ysGleqnUeqTTKqaXjZbNz+5J4MB
po3y9SmRtq/Cp8gPgmDQEVs1sDFFyR153fszEYYp1JOnOFFY/aiuAi7EZNPeta3I
xr3e9jVnsq2rcBEiwXe2enfR+r8yOwBTVmXHEMV4HT6lNjOJmpPBHis1k0dGsVGw
XXjQhzMLEs0CAu66VN8DMPLBd7QZyoh2ijZKljZ+w+VePrAFWFQUEqUlHlc8TIPt
xiBCaCaFitwbO71kbAFRp6mVfc/yzBnVM5wV5Vz/4pLAbDT/4PPOKcrywVZrn1pV
/GeuiRh/Jn3/dth1Ny+Ybl3EcMpCPCXyq41dfnUavnaHUZTZ8F/74ltq3++KNGrI
+VaD4T5cIxGBxMZz5rumRnjY4JFPo6radiJARoTiKh0CyY0pHFO5TxxniecjBXyo
WU7TbjxPGliUbcRtN2miQLJ2XTAz1/N9VAXB6d87O2On+6OAuHEQW1kt9CFPO+W8
BUPaEPw9t2JQd2gnje9B3ZRrmZUX4Sxd5WRcuELCr6DqRj33LF6kLEDhZi3mxX/j
EpN7C0fMBOG0F85IAX//6CinfVJAbPb1G3uHG4kq9wDkCIwpSFHwE6spxeN7bjGl
f+ccv72OICPWQtOxpJ+J3u1Gr94wVor7SEsWVVDhm0NHcz/eIxzwNPfcOwrjh8Q3
evjBUOSU/EjgdI3aTZ1gbhFpquGy3UQiSohVKhZTQAwY8EbCFtEPDQOLMoKdGWJM
hIbc9dz9mjKHG4f250p73JbqxrCWV7r8vPY0ARt/Hl/Vvb8v0tnpUkhhSiJRCqv4
qFSkBNM1XGFjMIXjZl6Bl3BOdTUMFNdxAb6G3asN2Vzke7zlOFVx/G0Ax2Ceglv3
hs7G4uUJIMki7XbNmDQyGi0unwjB8nRmSpgtt7l+zxjcn+ZYiY4HFI+Z7nHX6WJu
aWw+e+0T66OV5iql7IE72jRL2u7WPdqnW4+3Z+OVnUyj2TurIvqqsl5L3X9vkX1l
4JnMXuvArWc/8lzwg1YUH6rqnHfF/r+4YnorqN0Eib/X0fXiXowcLhVVsUjLTuWL
aV5aUusoBKvgu3mJRAgPkxnTYvHl76NZkM/BZGBXjx2V//rp55jHoAAzhl2T8Wem
HTyzncyQ3clVaC+Ool9IbsqLOePIRwXuAPkWf1ClzNoYLKXpgv0sn3gKVElQP2aK
YOdp5Up3i0DpEVenee3VQPYh5ayXCpU8b7YwZIDHmoLep+xIdGLC4NeG1zyYilTE
7RYCrERlpY37AxuNbwy+GUpPazpTjy+WZH6qUtZ02CSBUY1A/aysm7xO7IQMLdY+
ucdfB5iGhzHm1wMCzkVfHD6NQQkGTzLXOJdYIgeCupTVkH3H/mKlEDGen3Bq7aTo
cCHm/ASDlaZBzWL64DPl74LG69Dl9YInZvlefm39oIIuBOGHEhhquZW+nSk631Wa
RY5jiy0ZB9kUms2YTxG7RQdcdv6sTl6NstXKcqwr0hROMikJj/wyoQPuOTF1xL22
SX2Qqn8F3LkxkdNHKjqnqjp3o+5iwIbGBaVS9FkC0B2t6tmQvjtLDWaXSB79D1Kb
JdiZWr+WWd13NOqBwnucOTtrKH66xoQ+HuTl7azESii4TMHwReSR9gcQGhREB3Q3
`pragma protect end_protected
