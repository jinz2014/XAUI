// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BMnc9GMe+OA3GOP6XSgfHJ64HmdC7Om622pZgLBxBQ5Hs0rTcrM+FIJtrOIs7yLb
J3CnokbyF0jZeaMP1VNvHEpBJ7ShPmOekgVOQeEAUdQxhWKEfArpSvrxhKZrdbu4
9RQ0DoK0ebE8JYhUy/PLWzXOcxacHq2lfSipLsO4ryk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25568)
l+gznfwXaqsskFJ1HeVLWeCI6hAr6AZIVv0UYTV50IYpjmCMF0qpHn4vX3rTPuiN
96AwAz6zAtUBaGaewXSZeUkKcvy+2GaBnAv9IIGJVI/0fVrMZ1X6AtCOOJrE7RYY
WWCAcn9ka2qfxNbtV8ftGd/QtlcyGNhgL/maQsfnYNtBZMPm2ShLpq1DbXXPViE8
jLKAI4HOsRJZ0ynscvxWoZ+Wl9yH+1ApOFBg4RPlRMnxbtAPSmmxnfk1XCdDvUQu
qud49Y2XvX3+aqo0NpPIkC39JM8nw2YEik2IahEJ4oVU6+PPTQZ9nmXoSUAU4HdM
1VUawkJ0i+ziZns33R9wOhlWy+Otcb+hXquzW3VeKADlj3aB7bX16mvltaCA0PfV
JYd59T6rDuus6vSLbOlR3NwKFNelH1rq/OHNQzrne5ukE+ZiRa6Y8O/Mid4s/rMl
M5YJm448KyEzOr24OQWFerofVKm+P0xrRJsdyJUVcaeoVuzN/vApN+l0xxUPKrYO
3HPJAbQC6J+A3ID4NGuqIcPAReRTL5hu2h1VPf7bZk/a2P/qlpwLunMZEgCO2/l0
wA+RTA9hwa3NQZMbr83555jo5/hawF+zOCAvbrkJKsCdZxJiLFQ3nPoHOXm0uR8L
FI2nR/BEbONJDtENnKbjGypqsL3h7QfT+/br5ZCpb/zQrtQaW0GZHk+vpW5iC8MT
Rbp+k12UwHw5sZ60Z8JTMu6+UgTyGKnRtOhMBwROmYTkSyNAsKa5U8kb8aK3Wdzh
K7lMkg5VEooECDTFhMmrxr56sNEF2f6IgY/GR5BG4idAnT5ErA+SuhK8FjnNMd5P
dE6Eef+PKLHP98/zt1MoqgP0sa6Lpc9jlivtFPtWQBlt/+GhJyDRl8/QoNZIRo+o
1VtU8QKvVNBGnx9W0EbNrTexH66XKOSyw6b7EIlBGZt7qK6q87/ohSFzc4ml5YYg
hZ/VHw7ahLlE33PL/fDW4ohDvTZVfJ8MrM4LRk+Oz/ELO/72iHhY+6fzpipz/s62
qrqDSFXDKr4u17QYsKePxE6UKhwZuP8HNRlaEjFJdNETtrmTw0DB648NP/y25BQ/
ncP070U1YRXqpuZyso6rLG0MuZZRRloNPNb5s/7156n31VZc/G+kvk7ukRo8QtJm
nNssU+fxWV7nFCS7OdDp+jtp8AaQrTCgZQWX38ERVmxY6xuLB277qaGgrXd+YA0a
a7xNPNj0iBoHgOFbdDvH4qeYVxturPVpLiJrz/BfQg1yQk8OTUGR7gvw2D/HKHau
P3G+FQHFE0VQ279QBeENyI39M/nWcjC9CpqWPm+EkMXitAOwYDJDDteI1Om2Yl+b
4++zC5mBhlaNTI7tmis9FpjPA+vIu2pL5r+zT8rvK097rtfLaZIOvzHUgDf8K3NX
0LBE/hyuTX0AmP8LZIS1jUww3q1XqF10v/oxAJ13NYytuZ6xudHPUY49ANx+QPwO
NUjAlqtlLzDtTvBI8CPegRs8gAaFFo6+Pc74F+2xuMgtzD02vdVTIxts8fVesWim
ImFudjJjnaY57/Y+NeSxPpHpFKtE8ovFi6uVcjClHwR9MkSm98VL4g8MAIYjQz0t
Zr8l+dDNVIfOH60eteS8+dM5O0mCEgwFfe73QGi2/wu4tyNNLEmhZRtshCd48fDf
cugq/qtd2u7nU7cRg4/c+IX/dw9I9W59189XaHZUJuvHrpHZoqbtZ0meNFLfzAcE
NcKToGToheQGZzSFc6wdagtxtLFxYyNoQC8246BPaKn27OfzoWJP5H4/Lrbk4LAi
cPKS082i9xlcPDczFoz0E70RHCUS1f8u5uEKTdJ2dxRj0hLlgdub4H9Oa/JDe9Sh
Prxk+78oF++8/iyViIfzkNBTC+iZNxEN5QpsWTDNG1YbALzyhmWiBes1uRldzpgA
HmIjd2QbOjo2Q8PMM8gW9p52xdMD3S/Lk8EHCl80Jj5OwVGHmC0WgmEXecGf9ndz
FGNQDKIJKzC8TUZ6sFTzQmqTlQs3LLm9Qti3b0UbH/cbvK/smMsl327QTs2me39P
aBjwaxsGOF7X36MZW49t3rJpNVplyfq4C/u8uxd5A/kMA72Ajr4uDCC1LUQRh09X
J0IHPobqF2xG4cvke+GRKeu0TWIW45uBoGjMYCVIqquuJByTXar9Z4ZFQAstbFwc
YVnWC4Ai/5LlG9qVQR4dTudQz8ER9/8PHLcf6OTPvP4ddoUMQ4urrQdmZwwxXFFM
GFQgKE0kS8CVnNpZx9z/uf4/ui4hs2fTB4s2p3MX8shYkXpFh9WMAF3BfKZsyJtX
UFUkFSrsLppTN55yO/4CZjt9QXejDVeEhfVaaauBw3SFX3AHSIaXlRZgLloyHXO5
8nWsW7hv19onT+2/DxT7iJFvHJawHKYfb6tCc/Gvsjal8sDNWRK+oYR6uk0X2F6P
vm5gB8rNnXP85GblatUoira+IuDalMAxTLPqmxNjQQoqqf7crJu/FEjpUsVUEJKV
xsWNIpiLpRBrBHjwtljogxxiVtcsues8l9GS2vRKbjuuRfZlBR6AvZ8xBy3FuDOW
GbVwl7FJBhyozes5lsFl6batAyBfQpHhDddX+0JUAA1I3d3geLkNSvrKrzxd1wl4
fKMG74K7qN2TLNhA4r99++mh61TOTpCFYNLE5z3PEnryTUYb1yS1rmGmLYiXt0Zg
pSKHEPGJgUX419pGoocnGMS4CXYiMjN2DvPA6/H10CWWpb9OKBTtY+o8DnbWQIC/
zfGEv+L3nOslwXGvb3PQrVBXmLkTXK9K8FJ82whDaJKOBqbrmPBLRaamL8HsdgAW
4+jObhQcwjCxf8TIWbXIAulIh1BoQshbyiexB2MmhbfpqAzYNET9QZb6QWfG0n1G
iF8QHN3S+Q+hhq7PTPmvGXa6b2STQ7sNmf/n22Sv3Dl/zDk3x2iQ4QURcagY8g32
A2gEAnO7C+zqXi1fcKpb97rYljc+5+O8210ui26v1qH5fPzhg5/02iRlrw5HMHne
ooD4kqb1FHNjCnKICxi+WlUaVaU2gLluepv5wio7uOYYLeBrBBDRTU1x7i79+UaA
7x7W7LRkNkzB6eFtBddQECAVwKl78yV9d/cCCGXeHL7z5GiPTqHKLfSyRS8bxxJ7
o5QpeqU01oZ1bKtPVSZ9n3fFup57nMw9s5hwUJROp7MuJ1F1BUNe2xwPYhnoJXi1
Af+ht3jCKEIA3UborGk+4ejVvNHt3bZKZT4NWkjeUkyd2jiyesDlQVyWv8ZqDTfw
yD0MQPYSprRrYKN61tuV1GiVemFNQhgphHLEYpH07XjTUHttEmPOC8kSh4D21OBU
Jc1O4IujkOUJqnzTSi3W5qEDfNezRF2foCN2jHorlAkenisFXzBfzd2aNO2onaBX
t48MWqcChWbLXbUwbpekVEN9pFUcUeBvDqwuRVsasgl7DBNU7Tpqm7xP8hRBu7Kq
FBS+TviBWwt2+bWdS7PoYB+Z1/jKNxlq8IFmpet0fBshA0pPmezdoyOo5U8kUTqY
mk+aL/xK64lgXWP5g0jXDkYvVxLGjBEfLRhiinky+uDWe0e4kvR4BqkWtGiN4JSF
t+2hYHDxqHyv/oaut6zDyzeVWz/nwIAxJ2zehp7Mq4h6nSbtppSJ6DrnN16IMJt7
XIs2lCgGGi6/S3rdTGNYKOF1vrxT1A26E5I1JIubL0YASNSwT0ChNqtmpDSZcLMk
u6+U+3o4ixjTLO/w9dO17NTFCFU7sVc0TfOe59h3UDud+xFBX+6rMN3hBPkNWRoN
EMRYNhHZHV9npX3eA2mu/WXtQAlqAXjka8iLOILsfY0Z3JkkLfXYWFlHOV8olMV4
D93gC6DvgKtpMHkXe7ZjhPQgCZDh68dU4lPZcrQ7PJdUVwkkU+z27B8tKJ8QDZKT
bcljZ7GDo7VNu5CgxEnx4riQsSgaawN94ssLuHyWp9H8HGEIOqm0LBusquDWNHLg
Z0EGMb8oVyTqP4bJRE+y9QK7BnGIRM6oVziDpO2f1tbtREeD9kw5JVBC8upZ25Cr
qduUPB2s91OPlG+ZdIcO7LvcwoMwurZwfphHG+TjBqwkugeHjPHDC3LkR/0BQ22k
rna1bfRgl0Pwz2b0CQsQiwzcrbmqMhOYC0vKCuVHieSQZP3ZEmqhJyR/ERV/Jp5X
0EeloTcucwPIBfpP575MNUXHcdg8kMUedZ7hM1IM56bAr1C78NiC6HE0aijgOc2W
Y0/uF+cXAIs9NepCyaYyVDunJllAGdcjgeuLB4QUKQkHr0vLRFL4rbRSgXQafpNg
Ra9rG4Iqh4KV87mLyFDV93gCSdQI5DnvyoqGhRMC60MB4LIXA3l1sMmT2rsrr84C
6nfxSZ/AaMX8lF0mgou3Ia5tRMAnKutPfx/AF5cLsy0lyUxysD501qa81pydlw8L
M280Jn+ZKIbqzPKGJQ6h3vuyMYUuiezccX77jxVo7r9fWAE6LFXA2BdCTyrk7GXV
kLobKIgg1RAQc5dhUS6a8RATD/L4hlE+Ws87OaF7JAtGRQmEVcE/PSyt6gDHR1tW
vUJIouOt79fqZuq5rCejOryTf/acSmOViGOQp5OFJyox9V95A7h8Tm/3VOIrGKeI
HbG2dvMB9KxgO3QYs55SwhPBHQl1+w70bcPNs7jNTqOxFo1+UHjWuo2gFTacy+9H
qviRpmOxQMZSSqfZH0wNRPf5a0IiehY5wqqUlK6yr9ecM7jtDwmu5vrtfXSNPhuO
iT1DFMimA9UA5kXLsWHzBLrw7c1UNetei+kklkuAzKJoF6nQz1e3jrqHr4wdEPzC
vhxgbJjtqD2lj7nFdHoT4LV21PuIXBpAVXhr/Eqtx/Efkxfs0fLv3CxbsAoQT+l1
9h2psi+3IN9xYdS9c3/I3aOMmKB8S9rmPQk5JIO5SRLAvmh/kDB3bqoi3E+ss59h
yzFc4EU+Reo26A+9rHc5FQyMYgQjaenjwx7+NYl90FhRxLuMLyfD6rUOf/cqXzOQ
+HGaihs8wSScmdSMK//i5UqJ47jGf9YZt0kpMb9akFJfCbWlOegXX2TeomBDT4QM
X/aJgGnIMdK9bNCcF+Km3aycqZUnBFAxawZeTzRn7XwAyWOt/xaKfvUR/DO1Vwm8
GIWPCQnKD8FHlSev4+2ieahKwFc9U1XeZOAhd9FBGUMIEPU1bhDotf+kNvVcTOBI
uZBen+VHHqsjFdnSvbQP0dbzIe/iPZObV/x+gqwcymA9fYbjYISbZ4ufPOJzc1R6
uNuNv9LI+QD93sKCiGHPom1v5gViA3XriG4S3paBfvXNLOlWXc+VI7PQXt4ptbnj
Jx1HQkd9kJs5qnaXcNe/8nFywZt2WGjjix0KQM0me8H+/xc48ELR+3C3kNX3fUEK
sBiGY1afkdmNXbCk8D4j5jcvt385gcH1BtZhN4xj8lwD45fLHfIwK6+fhn0TT/o8
vG82ldtGdqGDogVe1yVLUlAfz4tLo5Urp4ilfnvQKI4RkkZcftd1c5HbGix/NP+f
stLEwEhwZrvIXAkkOlQ4ijEoylSYC23pMyoWb5EJtYy9W7W8N9aACTwuJftRRo+2
Kbcen1nPcXnjHpIO8nulooiNQLlieLtXnNz2KpKegzrs/ijCJAP7yHMCsywgV4q/
3lee5EgUCoek5IgI7pwunSq+sBG91049vKU3lla1bF0uTcGiokfvZoTzjId2fPp3
Hw/xRwhi9sukzd9NP2Yxf3XtzzG62VmYXvnq7eYXdNoryv0Af/Mc/qPYxkPQ7D2c
Tob57Z9ifjQRPue5qCwXvzqVXRrPd36YO3aRBKfnEvOGx2B6WEow+P/+pCiJBRJE
zYjoD9O9aTkfkJ7btlTh/jcXmcuNzik4dozC5K+Bxvq92a0tklPLq2lJg2OlIxd6
Rbb2NRYnvoMWUlgBU4/I1OGnV4GXaFYPK1Ul9BaAslW+JuraHNhiCBBQZxVNlKnU
hsczxc9WX5pbHClRe/5o9IELpNpRb1NryfvQLgk3aov9E9d8k7+mDNzoVgor55Ku
HT7wxnJPLgLkzKXeMisQYNUnVRsOOcuPtNnES8rVyFlRsfEUXraeiNjIkeb7HGJx
kTSDHaXR3VgRVLgOk7zg1U3/DYNdX6fVCEvbSFkpHqYFgF+qok0ouXz8C0/hovzc
n48mNwNmKdyZh3ilAstViEQhhlJnfGXtB/XTdNNnhVxb+Vy5s7bLH0w+SM+byCgW
iU6hPFZ3c/TVOBu7oFhyyhhfotyB2bEhwaH6KS0eHlO20FlunixH/BaibWCuezaL
k2tqpgEq/kNUZ530P42S60McHxw0ldVU9XB/VLgJ32Wb4kKzQ8o6BVv5+5Vvv0vr
qZy1lDPCndPc7KoCQdAgSlWkISJRx5vMAb1ew4MZ6O9s7FzcwfPcvRyRX0BxpFfK
WLgFRJj+V3FkzwZWHaZZxC/wusI4TkWlS7vN3x0TBuR7WMw+lsYspFv7zxT0rxNB
RLThoO1gxRGlhFJFsQddU9u7eXo+RW7b+UiVlZzQlwmiMbfprZDE2qBtjrEYnH3h
pb+RG7L3NpyeyvkDZvYQkVLzTC63g/lQRqnzm8jwJ1exjmPBD5Mtpj1XV+Mbm9tY
fjBojk0QYHPCGBYV4A5fHiP3cRU6UnwWI4MeFDeCwrYY3uX72CCXlwhBTQZpIoyR
BjtRhmFvFoJBxJo7StUvD7j5kCH1I419XAVB9QUIuaM5hZ2xBvZQsJRn3dLTPlVq
nO1/QUQRkTp6TAVsE4Oh/qayrvpBPcwHXFShgt8bIHCvTE9QXvA7+poFWmljiOfw
Rf42opnZFEPnmW6dC/Zx+FzcjNBw2VM6Ks/6hA4w0Q5QTJpAPzrHLwL0TyjQT8xk
7WcuGU8VfJLni2/FSiLJJCX4N7Hd9GP4aYNUKk1GQZP3kc/+XrcOdSA39jKi77Ry
Ql/AlftwRZ2e2I3S2VqSkq6fKfllRAFKZlgppnGXest1cXjsmkv0aL20x4P6IbVQ
FwrO0pDuChFU2qrlLEUlx0QDyhvb88CfeW7ltxaHuGzn4nj7ln7/XHYy3mYOjyIW
pVoKzoSqN5RBWEnQT8PCiT5JtMQ+lIeflhsLFlVpySrxf+Ql6F2HYJrmt0l5ioyc
UMOihYukmohnH/xKPmLQHV2UkorCI/hxNCJO6C51Mo8k/tSYNG4CX7Vw8nzUkcyw
Cw7PcJtfX8c3rwvl/zK+kv0sYJA3zXYT5OvXjG0SZILzYSkOsa/RXvYX0EU4FrQS
HOe0jEE0DAO2A1ojk2QMgt7yzX8+KSZo25HHNIOzGkkt6Bd3x7oDvq0AFeW200Mm
VzniMoNPrfengWXz3AkPwAerviT1jbd4zuXyrR4xjuB7KpzRSdMt94KbLA0m5hzd
NmGlx7vYAQYKAVATQu/hIdI1zhZ80TeA6hwRwwRwK9eSXejtfVFbLbNCrZQBmsfg
xB4KQGd7McQFR0Mud7PyG1BWt3lph8GLvVHIApjhIXuxmw/x1jrj9uKKpXnJLsIa
Qwm0N7aQtoIPcqV/tlQTKc/zsbNZ9XS66Kp/kn54ina5Haub9K3Arkj1qkoGohR9
cSryADCmDuQjMGUzdB64jyYh9fpK8xWKGz9HrdzapRXdYpc6Y/H2tEQ4voaLG3pn
RnyeYNWcibYidKxeXpEEbCWHkt9eCQLOL8F9SGj40A85ecCsD1i+Q0s2GRnd4VgO
hh0UyCAQjY58zkQ7EC/cSYw8kGnVS2YniS626wAon7ZusObwIgeHCz3gQIKQEuY5
BrmIFkgOdTSseteulum+NSCVFRcrCJDMho2Xru0OUFeylN62sewP3MYhEqujR/Qu
A9XUFB023dEeS5yOKUtaQF+Cp/yX7jFR3q918mU8qXz5ZcriwfmGR/Ms/Hb46hhP
1cNna6EMZFY01XUpAUu0AOexuPkTtKWYxW0EO8dqbc4NH6RwCIjdroYSt+p3GElQ
qTTkSe5w6rdgocuJ7kGDf5jy/Eti3gEzaeb38cf1Azn9lu8g6imhvNu/nrK7HOEU
e85Rcl9FXPwRbrwPA4aL6cOQUqTiEB4pufinVMe3EeJxr2nNMOgQJxI9MpGCatdU
ZoCLf620xq1wJxrhJwAmxsVC0vG+5IDsz4+y6XQqQ93KmezMGE4ltWWRr51ZSSEU
OpLYH8EuB2ByGQZ9uqBcqltKjT9lkftfJqyQNPTowDFoARoLOrHsAOBK2bORpfPK
nGzU260g2CfbjpeVhIhbvxYgwo1TWCiNzbdyXGtKCi7xE3YGTL4bPX3EKIkiuJ5O
SxJ00Yw7FkvPGQxGwCqBx/fPQ7g3kdoRLckMJ81DN06RB+M6Z/ViozpIGBQEugqc
SEHtdXEkMVfBs/Q4HDFbYu1tanVCZk66J6dmNLwXJJvuR3XCixTJZkZvF8lA9IRR
XSH/8AOKdQu1ipN65eKTw04sirOeC0pf+JxwqQW8CyvMbNpByU14qUNmUTCTyQuP
vln+mUeRFE6UZMhKWp3f6AlccTrBTfYyJIwU5VI5bRjzwESApflwvvjUpPfUqLpZ
7MnSG4LlSv50ZNtM37ovB/iGAFXpjqHUPjWB/vSbcKnrmE30bELyes13yKlg2Icu
uIYIUXJe8mqXet+2uffROJQwfHMhoF81II2KUrNgeWOmRd6z4QNc36Wx9FRYotNf
R5WV8svtL1smPbftFioVF0jJLknOHXFT+RBusMK1ZZdLefePbI/KQHd2Yg3GElq8
UY9ZZPTZFzvZDI1plDftwJUz8//3sCYglu0meIIQVyYILDFfQC/KZ9eT6sfb92Yh
wJB61J8MqHIWGVVKntiXcmA7zxwFBuOpyZaf/H77ZkVDz+hh5jQjYRUz3dcY6ycD
fyWYFkTfv/PcPumQZ7zhOLzvxzDtvex4qtdPsCVgxZhIriDna7ANH4RfVPbZBKJ0
KoiQnzKRPYiC/Ivy3l92xNTzwljkbHimucDwPjl5uGymaQqTAr7CRB6RPOzi0lCl
ZMfcmyfV89K+07YA1Z/dBoI76jY5MAFSTr3oGsNIOSfVHynZrhkorSgh0jw+KjQv
7U5gg4QU6FU/UuEyUJk8WNgjq1b0LCfh7cbyk1HPMoVkcIPgL6ftTieZlf0v2uZZ
oGHtBUgqK5Gj3LvFXskTx5wLrff2AOIM6s70bBhgjOZCnuaa6eg480T9MJgxpJ2g
CODIEgWa0WH1f8noYF6Gs+28uKjIDmmTnD4aRgrr+NUYHv6hVykIvI/yGin5yLEX
z3CuHE3GV9WK5T8ih1lngoiFn761jZmgzA7uLFovShLgIbhh3v+TKrW9g+EPlvwS
4oC/AK++RnvRv/l25POyKue3BtHV9kOStdDeLRWzOyIOuYUhSfVeGynOCXIncuFw
eUdncpJrg4s+qn6/z5lFUcHv8HrI6yMxJxTn7Ghx7WP5MV+sONMRp6x2q2jxrwkc
/I3N48Pdzocr/6y4D5aZVKZv02PTwvtYdWYyotuTwDxraHtWzrAjTMfdHJ0xHzM9
YLQdGdQ6W8ul/JgcXldhhA46uxvE7gbpXpL/+Qvs7brJyVBakINCRn5ec9NuZOAS
lT28eR38/Sx6vBNysbNJi7xkacnChgC/v//CUoBH2dCputOANGxPVkb/M5WRVTTT
/qpMxwQAJXPsIpMPx8Q0ZoN3L6mcl3hRzgrN5nT0ZBCs+8IyleWz4ZfC2G4jkfVC
/dxN+pesBoQOtnaF+5zXs1OkUDyM3/B3Lqu19Qxov+jLlJ7+xlAfOp8xEMnrYtKp
DjaG6iqAdxyXs3M79TQ3U9FQYDXoAalsYu8RdcN8ScqJWYOpHylUTqsFmLC4eHGq
5jjNuocVVwC0CNUgN2Oc7I+fx4XMAd/2mE9y0HvzQBvafdQ7XX2YG3ucDTJ3PgU9
tGv7fnZdZjcSNQCWSH5XQEIterVqtW0BcTxeKV+qfeWXygU9n42FOh1YxOqNtyo1
O0pHKtMJ08OxOMywjriAEl4zdwzB5UUOGS7eG4Yxup4P8cvAxXEdmN3/zoeXSP0/
+7b//Xf/HkoQI2501u8b2uWCkUtP6Jbe5FE4PA0GYd3AqpuvtRYDBzr4lSeTWv98
pGXp/id/VSpYjSYkEozRNHVKctsDsxRvcPBaNkaQY2EWePZRqyuy5uR6NHU9Z3ff
u4HgWkB5l674UBEgSn5SPPC5eKD5ZFNW0EA2VEphj2h/QxthoYJC1Sv1PX6zHA09
vsVpjnjnfPpesM1pWygMvEwddDTe1cb94FgrHtKp9MKq9CwEBFcPEqWMSPnDwFC5
FB9Xq862JvZQB61lBv/S1k3X7E83Gfw1NkEgEW9RtFSIBvEAoH9z36YpjWX2fWnC
TYWR44zhOk2xN60+YvtQ5RaermmN1gzxbVoPOZfUmc7Y07qxYMEVrwLOoBGRq7mV
3W1X/tJ7TmPSiqsr427nGEa/2qBI8et9PQc7X7nsbtyk3NeyZHUbMqti6TWa7odu
xO0BeS6yK9iX/a9GwV/K/YRlfw4Z7FmMLV9pNhHG1JMZboipx1xn5WjL7/2FhBXA
KiaTgieMmVtZluD5rvJhLu5VqwW48qNvBkXL4uq/ZITP9MkJTDQfhbzF7Nz5eRwR
jnI2Td0yC8VlVV+fx2VFZyyMJvECh8d3T+A0F1oroewhVgJ2xod4+ItNpo2JHj63
LiVEpEWrlcMZYXHM1YOIb1yqRgV2aTAUz63he+CTa2DFu1KR9de72GnheWApHedL
9cIAN1l73fomCvSA2jpwnD9NeLN7/BSz1y58kFTUWsdkpFO730FyquDPBopf4JHR
0txUbVFANeGzMZJRy/8UsbgRrI5BczzlEoJLbJqtVBLw9mB0+l2z6gVb0plLEVwc
u+NBLeIKLmm2oFxV0NC6tfo1PeuaR+BRviHA7UWe1p1x+F6w3wwD2oERZB/7rlFi
wH/257TCKOUxOcjz1To9v5UBNbwFEs7ttlkU3JA/Zv3E+TL+Us/msIib4FdW7XzS
7MrVs1Yl3ED5fRIklYhRIqdtORaoEBtUZKv7L1idWN0o/QFsgIaZ2OrFq+YB+3tx
N1+6qrnMDaJGpqKF9a7ERrWFvQq/rijr+5DD7NcW75M35nlpNwDnD9OK0qvYU9Z3
o+37hGJGticablm53tJX6W2facGLh1/TmvjxzrDxoodnkbY3YhtaTaXmEFPKuiYd
rBJwDijhmBciOtYV/VIBxBqqasqwgHOPoKYb/rmYUpZnWmF+a+VoYFkm28xSS4Qz
2ZsKFC31PhRWfnY+50yeaJlvEAYwSJTQZ/THpw1iVvSyW7ptuCbb07rhPmKyK6My
utt+/fEaMtFb9MNbnCGnvNI4vZ4/cD10Xi4MlywUDyQ01Zg+2zW5c1tZqoerEq4u
GUV8rtUDXhqcYkic26R7WeGsZB3uT8Ypba6PL+kOlVrwELKBASG0OTgW4/qNHWIj
SqmJw1O+JAhmijjC4Y2saRMllndmVwFCMAlHiynC2mjgd0Vjyhf49MXh2lzBeGXw
fFNeqFbNvmuKbDZMa1Ifwvf/BMSZBv2cLeU2a/FF3RmfmB9a5cfbkzF57nQGkqMO
JmT2oaZ+smfFDHUMXBrtVs51lqFCMVNlQ49SkDbttCKXH2uN5W9lY0f/MBTGOBTH
V8ECF3gFkO83FC01lrkWZikOkwG/tApGY4bjZv7ZG69Fjac0DbImdiXRI0JmICoH
QZe5+/ocETkOLFHBT5P4Qsa7vc1I3PUnc+yt3cdTgiA2o1uHLB6G79uS9OP2WAlH
RyamOhPpOWE6MB5K6dl6jY3FzwQZR0iOtluprZvLfKrr9hdajzh6QgnMT7/GsHT+
ESBl59SuLghcwhoS3HqRY6dTPj7kdq7ZERBG1zgm5VCLMncqHsaOYQY1M+iILgUf
Dv7Al/t2wGj/kP4ljudaq7xwW0/zR6Jr9UbSVNB581sq4KKU27MaCT6fDdI6EX89
tvTxb33XVVe30pbmC+Wujnr02IJvTHdhN/aZnFnMGUwaMKUVHBz7hNnDQ90a4Pr0
21kF+942Fl1lG6hTBbzNW+67ytsf+iP5qQsR1RvliMlqjXc7AVhtNZWoaxlAfpOF
qVuF+AOtJHG+7BO2UaLuMhpuwd6wDEBqRgaqjgVcQBj+4m21fVWNBTLBFkHelGfs
bwddBYIkGD4SX7FrLF5AwdNFV1jXtj4DFuMDL+VRSidF+nihAg5lkp/OkzO9cE6t
jL4/B53tsbRcAK4CqZkjGNwhTu21yS01tME7y/uoPBjlCD1EjgrMIUt6ZzXjbduC
cp6Uy753uA6dTHSwZbM5Lx0th3iHrrTxUuwP88nQQXjcv43Otwc+4ILhH6NgUhrO
b7ZDSjXuf2ys7TOEbNHUEFeW0bWS4EEwqOSzsDsH63y9NBmWiqXRFtYsFj/+IxSw
wLOOkQfZrjI53hI1XWiy7Uoas3CzOvMUu14zakaFn1HIhXXyZB8lXSUEDOUivDnW
Qz1Iwldmoo3r4Ccx9gK00J8A7D9FK1SGZUw9fEGYcy9nhAHwaF7KzmhBTJ3t/bab
P5CbVQUPnF/Ahd5Lu0cCzbtvDHozb28zt10zMNIIeGqDueJPlnlXrDCxX2/LIjzZ
yODXdQonTCnJiW/Rx8iA50pj4opMVISYTZBv00jJRHHYAbPL/x8C7mQgPYmeibDu
GHna5jnv/tIzdbSiD7dxzABbZiMjK1u2aSJCqtMPyD1IjAmNbjht6ER9GsuIf5gL
7yRpH7AbUkP5MPEMfphuiNb9fwFm1OI4LXGcLX8kqCRwu1QXH20KSAPmTPtEGTqa
4oWpg1sS2ERhden4fzOwfKPFRlevHVCYxwF2cVT2+CLr7IKKAZT9I76lvj3nsCOj
IgKRfiBaIk9yAyTxdd01T/UhkezrBVyMHyXll0J9Kv+KXlzV4iczLpT5c1vw5+0W
7yHhQfTEssYdAu4cPY7rPtYa7HacRSk6ZWa+EDzC336JzguYinfPOS43IwuzH/Sc
VI/NWCb20wPPYcDNDwixw1qxscF2xM6xLPtqMm9Q2m8ODxsiRlQcebwiaiKGXXKw
2W7FUvKDJLMquw2Iwe/B6OM/A0gJphc74yx14U+xzJehGdcneHfLri/5Zleq6SCp
Ku5dhMk1pZbYLBWjBPfRAgW9hrkUCjbKCkNM6FjfoNtS7xKFv3nibGA5g/s7dNtk
XlPDLTKjQ0SjY6VteT751rZeY2O4l2IsfEE7CxANdxg4l0Ya+1kCn17kbr2M3vxJ
DZxqjGImliJtK/ktd44o+gwVy3G8Hcyt1QdOe96rKRSG+1KneNqwd3bdJKtN8h2E
zyj9sjoc7f1Gg19JL0vlFFjprvtzpnOowenoEwwChdyDKzOJOkWsWbXKvdr0pWNV
xqEUMPqM0eF3/JaDiseL145W8SzGOA62xYoAGjnC0O2oUNK2JXeYqqCTCQH2afao
nYLQ3A0EHiFxL4li6LBajRyZGCAorDaz6/KeVhfJwHySP84yx+LNnMdcsE1rnoIr
ioJ0KDbjM73pygpamz+fNI51NoPvczv5HXK6cwu1MS15HJtIFrEcmZayve9RCcTE
x/yYHru2BrGqQhyPVnCW9QU7t1dS/NwHEwI+RSEoIMgy4JKszNTs2sGR9CDPJgkx
P+GuOG7+mr8dnYt9s6svvZtBkK+JrZ5Oi9SPnVH+3XX3erg5yAr4LS546HOTTSCL
EL2KL74fm7orkcLoQHqanyEtJbylsiq0awkinZ10zQ2j4OSG83TbxtTzqWDx7IpN
EtyIvaHUjOszVoZraOtjYwJ84JI1+9Cfu0LVxRVkvOr3S8RhUC2XQRwjm59DKPHn
Bq4n8nehHES8oZR/1NstSwKmglQUEhPHZjjp0UpSHh+Ekvkc8tM+pPW9la5cyZJM
r3+PmCxDViunfTdEgBVhKC42sGRbB4WYrSIdwMWy9yP58HOvQhgFz73HsZaiVorB
mobjsppPe9zuVuB9duD+PWfo61m53w6YXvaIeuUNWLHCr6qdnvlpx3w5zLygDVV1
YR5eq61EALRaaumCq8wY9LpERROjbjqesKZiVR4Y4ZFUxLScWTL5Cb7YZKbC8w7l
JvK8xoKnq8x4XIACqPIuwsOStaT7HpOCHXaIlGopIvQFlPDH6fFQDcEwVUUywiU5
dZLRU+V8aqCqBSH64Vm6Pw3vaDJbCsU6zPcDvKs4lUMqhAyk7bqJVsxAQqQhlOJW
lKl22hg5HRsa7RrJP8auW2zmUSuu6+nNXVDK0+oBpfsldjtl5cyl1sHG3LDtNfGf
lyBWJc0D3o+bOY9TTRbAgyTl0kYyCqwldizDajAoct2447wyO8rhgiJBvzrfs77I
nm6gqA5omfgHtNyQi0bTOmD60wQPW07cAO6jUkRjbmxgSCMg6jht/QYRCvQ5bzJL
0OdF8hd7ovzu/6Z78E5kf1AvSjfZbXZ9KOqZyVJDuVvy6NoTKSG1y8GjDHCTrvHB
Apq4OiTIw3TfFS326f6SH9+p4Ku2sG0xwR7X/99JTK/Iy/Hk0jeoZVsW4WO77K3s
GRIc8VwMafevh+3zIyLc5nS1HF5/vKuKL22i2CGm5Yl4hKoyZ/oN81ZhbA4plvcQ
+x6D/rzfHvOLJmeEJprdtR/MzR0+85hkmsqBkdql/5Us09bGEPn/AVyx5s0ggba7
StQAhEMemqm8yQ0sIi1tEQGHpc/qHyjNlbm3EgJHgrQtuZyG0sdr96E+6AtkE2GE
dMomzbWc4IyabqvcET+SwdjOEj4nvgCgcxWiYEfixJWYnpjEg3489GnDhuv2qnXK
fJs3+glDR8kPdQ61hvuSz1wyqRA94f4fLBJsS8AKwyIxLem/l2IPqv+sV7GhLRJS
Riukimd0zv8qADU+oNwao+FhqSx7M0UyVqSDVxfd5Yy34GnfS/a3oq69PvWdCxyX
ELavnPoOvlsKwmsqvNt2GnbGlvzmHPKQugcflqyzzY3cjPpUFYve6SBNP+qXaBxB
dKQQpENc2aJ+lR1xjQyObsk2Q828TLwvStkxi9Bxis9DzXgn7dcB1I1hzbu1FwcL
nTxChpz+FPjmywHtKSABPOpbaJwryz4wQyiYZiS6GHqqvOWCdkBnv7OEYIb0CVrW
oQE+arBW0kv08JPJg8Wn+ZfnyzlxqoUg2HX3LOz00IfPfmnKqlR1O9/p/svlNsw5
vAbBUK+vMHtS0TPSEN6kb/tXrZaykBjbZk3IBfhHydiJKI2Xb8HTQsqCE3buFgoM
LvUVUa6Mjyc4UdyCNjzSvmbaTXwD4VBcUmMGaxFmbKvoblbQGS1Crkg/l8EM2quX
GpA2cCX8n0koZejSxfbN6ZN5oWQd6hgbyysU+5TPYiSimdFLK/riTm88aoRJPglP
Fvtoic9JkiRH4Wn2XJ0w6kt/pXzHC0SnyKGkX1u+cCDncJ0aw8ShVs4z307CbEz3
XHKKvoRtyUR43TPRqXHvD6mtpngSeP6nKwiTt1BAgVgfsulIeQK38BL5OEVTZ7pq
sgJjs5rEGc6Ao4cqXHqj0VaMx/W/Slx5PQZQy+Pp+JpRfxRMtLC4iQeQf61kxnZf
+0u7F6TqOYcYiFbXyDJ/K/KEkJMVkqFWaNsFn6MeTcECDwCHzAcz797Nd3SE0nMj
cRRT68TTdmhn51D++cUnQErzSVCs+6KARYnS/Eyz0Kr/0z8XAaulWwUMo404V4br
mzxN1qA242MapRODG0WXxsJzOI081ifyU9+NfIfB7IEOXNZ+4bke06/Gkd2+XOaD
mNckYqGAMpbDJqSDSWVxqYKRsb3omYsUB82Jq0iCOp7HHXkZ8vnyjOtZt/r06Liy
UQsNZ1RW1QE/UdOBwV7424IQs2AqJ9kwAHk3bbCgyTt5lHEfBYaTdISeB4Rn4c+e
COgHDqzgjAy/BO9cElbwMu+gvxYPyUgW8hioZMCljmG0bPnaV4x0hwPllYtDucJ9
TMef3F0ykIwel1r2oNlNU7Iz9HwbH9vz/lKSy9ZrX69WktkME/hV/pALh0YgK2G/
ST8Yus41bPS6cWEiqPZFXOxzmzGRlKs2VLalNe4vlgY3J4Qm/uF8PbY36k38Vbel
hg+50dzQU73JVnnx8doKdnyjyV+a7ul3MK/CSOi6UhZ15MoV7PYNsz6RerM6CoYS
+JtJs23mCdOmheCdp344A9NomwCZfmB5zyB0xLmIdf7StYHPsCMTVZQucdiLOaFd
qgHV8QFTgVmoPLsEw41eIS8rbwarHztUSj2L1bYVJxeaFA+x7xbc+N7eGg1ISPCa
4GLmJJ7opqhfsvVHctbrFTiP5f2kSrDMxwiLpug5c97Ag95INTH9bAixbswNFTEy
g2NTx9+WCtxso+brattSc0CfORk388WA3oCVjGS4ctWAaqYYoIx0YqpUazkIq8PH
+WxQp7t8zB9PLAcLf7xT04OVrOI2Ljq0JcvuLHIsJi2U1XU/RPW06pDd0cNpyEgT
sf0NiTTWwHGFuVBZQQ1sNQkbIZC50D/Fh/zPcNZ+f26Tm2611wwwLsbjH06yu0zf
UMX/B0HbGTSqls7wegF9LZ7g/+OsoJE2nlvcuvk6am7WRWw99/48xXyiu/heudel
1GmX3MnplpWRUAJ+3qsAcL7zG9FaoV74Ei5zHsXWjCZeOV43UEyPz7pY+NFZZ0hB
cxCuJk5ocbUqt7CucsAYJlx9PpIM3e3VvV4zdMI7EDsvibXZ8hB6M9qTUruJYP5a
E2khMg/vr1E030Lb8oHoI1zGIxWLkLLAquBmsDuXnR8XV8QoRpbZm5s9oeuIZdkw
lHZXKmPtQuoNh1WefnCpw/h0T0FXBZ/YRqeApgYuXgt9KeYS1GtE2S2vJOw7luDY
akg7SCq5I9gM0r66RmFmLt9o1UWNKCmD7jEvVZ0rH5nVwp+scznN03JyUxk8r1gK
G8z6Px7qRNq2YKiEI4fLNbUEEk5EO7LyThNQELEPAYQxho1Y1uts17mLjbxB07w4
dOp92UHCDDHv4hnWnzctaBqzbhsTk1GX65paSLy+8SCZNvDGUccFtUAT6CRqkeID
hc+3ZeHA8OXfQItsrjwu06xSgjX5E6UF/jsn2g6NY5kditCQkwJ2fwpTTFKl5MZ+
qGGDH/aJrwTzMXHxU7UT8tvupPjdJSss1riwoSw0mzO4o3EtH7d/QXqd9/pFWFq+
EsXzh5JjTGkEC7XFxhohW4A9P3jLIEvbqAqxD1NMGprFljWMyFcqmzEayxFhooEp
fGqTXuHjxWfMnP4F9h4coJJ1Es8EY/tC+VQBRlRqYwF90pTZXnj8fKgfgSM+N4o9
z2RlaM2kfTt1S+318EWhQgQrgs8O8mkqYwRpRePGKdv2y8/IXNaNk1ZLEHIteowu
L9FhSKY7dKgIc9BOzPS1fu4EPazEqYX1NvEmyONLbS4KXMIFhH5+rIGVfEPfhSVd
m+orVQN/MStqUKKPQZqu3GCF2KC4uELsmXj/GU6F7nVd5JhvgYIfIzJJyWektp2y
+BUFj+GDVhZFiBCC3l63+CSmOiF0JhFxFnZmIbtwpXvT5eqC1Q34GRVLQP7v8mBb
pwNrCXwmVAtO+3/ppew40dOBwDpLjKoZZp/Ujf145DTVB9QLMqcWdvNzPzUs6FSH
BiRMycAjAbWc0jOyD+fIXlzz938V5OYq6bIolqq+PWrcIzi4fwypXjBFKzPp4b4n
zw/rhPOX5oMVY3GAFSdQQWlmSGohFsPhIw3tdHxpKn77WDdZHxhWCyPZOFDGh3n0
VZC4s3BJeB7tEdiFpvTwvVbHJ1yEohAp8tryZTPsEGL+BMQIY16d9jy/5T/RX5PQ
G9ttLvXOncqPKZr+aNnJUTQT/bPc974rxalnHU27l7Ds3rFym5RPDVRl3AWzWJ8e
KFFhpFtEsp2Qe56NZSNoIvW3YdEaKOgPluK1meeHTvfownKMmh2ub5TRYMdOBq1g
0qwQpoxgegQPhXNjwTLgoirqBjMZFYxv0D8pEkIvHqhiNSgYrgTaDK4/7iEsdiOY
9Iw505cuRUbexR7qBUqvLZcFOLcRFcNSpLlsyxHU20zLrzuErp8LXc6WN12z8rJE
2rDjC+hUsMLIVRWRFzkXizalV9eGj+AK3COvjPKtVGRvpL6tnPTB7UwwXvSYXtml
C5CZypJI8Z4fBhRAv115OPXQv5QoKmQmn7gq0mZ+GTlwzRsxuw940nl4t1lk4liB
mxSWbEYLRuaddBXhJZXyJXu/mAJkQ81Q8Kh/mpucUJKaL+D8HacrJJ0xGS7GFjfQ
bmoG7LZKLAAYnB0W0V+JIL5msNr4gz7D/HV/O6IAez7qDrvIHU39nt8+gj1Jdzif
m+aMwmFsJHC2AkvRYT/ztf92daNlbBKk2leXYHZv+zxbHs4hRX6PYazkp+KPA1IE
e3w6geGxWz2K9YMetUZHjFeQ2UQDDAoisuYXuSzX9b0ZPu3hN+Nb4bAel8ds5RaA
ruwUqdC4E1nczEf6GlBt05e9vPxYzT1UcoGRAhHOh+137Oyt2B015rbJB+OltOpL
JtJsPITxzEhJYNO5qOkrRl7n/XsMT4XqQ0UUHj2Z+L9L9z0eG4y6tECEWoJ6p9vk
9LwfxwObtHejIpgTxzTZVTg4FhUneoLUPzhxBuRwjO48Rkm0+e3RXXvV+04eeb/2
vQE+zFwpUMya8XzRgj4kRW3VatbJxtOsNxjDeg6oXGkGT+Ks0JnpZdkSOnovp6Qv
5MLmGkx/kFlZ1zcIynY0sU4JK8WksE8cbNOpKMbHncB6hj01FxWLCNleuR04m5Sl
DlzkP+76qXzWafirSShw5tOAcLfCM5kpTXb/cokWqZh1Q8l9bR+WBpDbRonNdgfc
LqqWn0evBcQ6DEvU+YhsEzxdraRpnoYcBLzEE6LRttLjaffnPDvrJzRqgrPAv1E5
pbzWiCNyOJ5qtrquRZ7Bc5o2YX0y+T1XL+X2O1LcbrutOz5+AKARWNBXGVztUK3T
m+Q+14+8dbpgZzLng0Xeh1WksLcOs9gMCSYauugfWKDos0iSIOEhYSsICMKT3f5d
UAiH7z99otEEz3Ib2XQ8l6w40zGcrq4P3DKSlvvD2WLeyPwaNiM+bnjZI+CzwkWh
I1sJC5iFN+uynrI8fUXylJCuchrZUFhzfgQA7tuMJSA+YF9xQqQukT+Vq6uXBThw
am0nDSyy5Mx976PmySQVMfUVP69O1NgcilhmkY+zJOY4Uf9BrVTe8OJqKCFrlGuw
OtCTzTtnXpOmB7y3HZeC9TGtLKtFpTDlIhVcT4TWCRza9ik5I8nTOTFUVA7K6D/6
s1WqQOx/4Cv2jL+NlSwQkg+uwbaI6K/8OezyeZqcf0l/CXPQd3YsctDVcjvvqHCl
nXOu7T+J/q+7uiw1GCCIRZ4NTU/iWOkP0aJOtzSDBof96ciWSxHJvcLNXqlAPjbA
sf5S7EiqVZiTT4Tqqo8AenlNAbxCWO3aRjzyPeKXrUXQKPjY79lMUtwDwJb/v4rI
LOqD43p8+u/JQiN4ESmmCihDnBhLHLTLOE4tUGlo2rLIztVpnGnhJXxBFgDbqUm9
oQccQqSYrRUdah9LNHU6Ljb/KsmtNQTBK5SmSVFhhpA/d46I/IzzEQ5BMIvW+GhY
6NLURETM/AH5agwI0CfcHYUhIARA7dAGOrVpicyMnVpiIcOdy1PT825M3NeMfX1D
DyOjPreDRvfZp4RUDVPKrmyGcohCLU+YDQGwQ1iCE/MW0XJSfb/bJ0Gn7a7tNuY7
No+UlhOOyuC1lGbiOJdzUc5BeGKQPKbd8tZpW/0vH+MyNUXt+wOUeqKSp9ouMpl2
njBfEHbici/5wrKvd8wLUQkcNLRdZYx72rdDoFv3luHuImJnTan6ERbXtmPrQwRi
Z1I0G1pjfvOWF0wE1iH+WYgGJBpxxUfYyErfbbOgx7H4XKylhz5qibB98eHBSa9r
nDpg4dMyKUqYAITODQbC43I898u2oGPhk1Z/9lxjUdpHToIF3ONFAKS/bdsc3nYh
LIunHbW0tVrticcTRYQrq2OlvX+u3Zv4ERxNtcofIHbyy8hMoOzz86tL11KmMC3V
rH+qHPd0FQXK4j6Vgf++w3YZMif93AkPqtwLwpxN29l8DfjOxtIvSZfR8KUuGlJd
DdBB6+afuFadT1zWy9ddSuoZJ7asiEZY4hGeB884FUsi4mZ6E9y3J0gbpwwqitUV
b9XWqV9PrXDyeIN4zv2sS4K596mTdnlpmOiffh4d5AGJrdbEsj8xEQc7CGbvYOIY
amUEhDuSH5euLnrWDG1/bjn2MhOR+weZuBqPN/crH1I3IH+pPsMDG38t3pNUMWom
r11+iMASwpPom8GAooYajO0QjoU/LDmtEZyxaDv5zUWJ64clXCuca94L5iPXtvgf
e0k0Xc6F892OWyHs3XaBWCIdd7l8otGLUI3pNTeNoZP7XsT9YwrJrV32hVV3/fxA
jFCbi9yME34OAZaXjqaMeoEzDyCw7wGMIGthrDpgMRQ2wb5J1u4asAp53m1vRTtl
WpqddlMlfSyw+C8qqa5QoMJ8lUeBQNtvkWV4+VIPtzPBs5seua6kP8dtfXuEurpi
W+qLKe/ck8nH7yYtvB06euD8wT3ALJ3CJ7HhluxaNcVbvkQEuoEbq+3pbQKWnvfb
IAt/i8VPp9Lq9hE0vVz5wrZxrZsZuJCC/3NnGUpdjQOV89u0yosqysIY7+ABr8DF
/Xr1Yp5w5XzCQbfhhWhYyL5xnBemAuLkZZYnkGW6EDG4NYHRoqtFD1N/4h0tYN8w
0+4Ynd0dciy1cHAgHTmgYZYgtTCDrgU6Mgf9DVcnCLZkXnKvtPILHPF4WfBHZeCW
Y8djpKjCvMq4lPUW2tdw3hI/LzvD/H4EdevYdoOWB7fJqqvm5/nquArwHkqn/LMN
M/UkMyHa4nncdPkz2G7ab3doYPocwkJ7jstKFN80OmuVRv6Qgemj7qgfiQjl5+G8
v/+kApdxVmN7CpVbGVmsB443Is3xY/9YuJku2Fjp+nmg10rd9ZkGGn1gs55GCxI/
BdMg2yf152o+ToteOFLzIz3f+K49MuvL5th4Ty6ijqclPUvNFW2I4aeTqhK8gTh0
g3kZZhRLmBRu2vv2D0kHopsha1lSPH/NpJ3mMidxCdI8JaFa4UoXXh4930RgdOe7
qW1wi7/zXjtvjv2/wwDFrCRzSau00+seBBdnL5Ikfv3XjqUVe4F66+cvc7kwnI1x
n8gKcv6R7IcgQqkLlQgXAIWN4liyJxrRVYLWvsuj5zTAsspQ64sw1msqMSefHuW5
b9VnlQQHALJYqh44JV6g949M0ZC/I+J7JVfoqvmBaewIZ5Z2sQvrbZ6J63yaNoAV
kIk1lIOsIQFYcjgii7gxd7TPfXtXgY4Mgn66hmqnTIKp4SOVNy62rBErovwaQcO6
hoCATV3DqJfpQv9WjIbFjBPcKV6YYmJHuWc8fu2nnUmFDh9mPi5/znUAFu7Aks5i
8u3dlFI2sL7BgZyaP2P0t0YOBEWyaXMBPt4jbxEZZYgB8YrYr9B9viqA9MTL8T4q
6S13i8y1woz/UHa7hErYhkGGwEHqZdS0p+IZdRiVNZdAF8es3OfoR6PuoxMhhdDu
ihYYWz315c+55lQ/6iHKOIG4R0XHIbdf/bEirN6qEU7MQxoWja90xPVO2qIP+VeJ
gBFWCyqPDb4IpEfPTOI/X1TTvi8xf/fFKLJqFqkkEam6SPMwB2WYb67Kg8eVOjZG
03IJdK/smadWN7GLO3n5rhvdas5s3DEsc9QCHDPBQQ/rnLaT3X//Uw8q75114tSN
cuHp7dlUYLQK6HJE8X/3IQtj41Cl9xhGOCo5CMetN/hZ0gkHxP3xmHsQjZ6ds43+
Zj9Hcp2TYAB28xfnx2Wwxg1bNdzzI5JI8rL+hTloyKxv1ErgK/uqxIEhYIZsx70x
M0Z4iQlWA5zJ+Ibzi5Ygph8+C0gDZZF67z7uy0Apb91qnVQxx4RqaVvf/0ZzgEcT
uSb85/DOGqAtttY+DNseuuw2HpVgaL5frX8G0/HG0ehlngJZMprWQp9GRBhNPiVI
LtE/Uf0hWw6oQblqjQrCUUXYyBbpESxnndqTztmbRXhKPwXRNAx+Ikogi45GG662
2j4+h/Tas+GBpLWkCkgQmB+jmJHf8zLH47uqIJsOr8lxSLP+GY5fB7obBGze+KUd
Ky8bUtod3WkUpkN3u+JEBSJkYQ+j8Vxryi4tI3BJ1JQELGY8fAzhnzcBH1c4OjZq
eki7ngP9CjuqGqCla+ln1kzUUE4hsVngohKWPs6i048daMhspdr6BYBFBjSBJYsQ
oFV/anZEYrZv4qqiqlPRWmjZyflrnJH/0Eu7pHve/x+Ttf8auDdPDjF7jKKlXW1M
2yi8Oot3Bt2sXGhlgivOJe6jhnMdS2owPCx4Aj3DYWE4yykg7yW3qXSujFMGZp7l
PUxa1TICHxK6dFsan0+aDfxqYS4OR1iXp4xBcSMdE6SnNJ9tjkVuPbgUskUa/QPa
vxh2ebple32ctzHnGkM5dKX6gIS0cJ5in4px8I8FhsfLsTZ4nkpYUNnX21T10Mji
zedGZ133FWcrs9FxUp6/Ep+F4gvA8jQXtnczoyOAZAf+c8TNp/wjAZQA0guhx+Rv
/rUd92ifFcaK9CELhpme0mgAuv4uYz5m7sR1MAgyaVVLlZ7yVEXihoePmd51Ha54
u1dVz8TVXXiaiidyORpp7GmbGqJAtOzfAp7XfOZfWnJqGZvvSOHxdLr9FMCz0/iA
Cu6gTMg4YRr7eRv6rSFu4wTpoVjGGq9jGBErv8qnm2H1E1o7q35hYTmgVaNTCQQB
WMRzvuJvUKbPWeeawuCDD437USSS5rXlfpWlio23XB2uFYUAR9tneqzrmB8F94tT
bziaZ9YdeJeWjFRzTwjzpmW1HRBvDqZkUIt+A+JpWp4pLNbfCJO4xq0pW5RMgGnO
IE1rtsQdYVZzci3G0SO4GBpMrJHWsx03gPotL2AtNYsjmQ1LIwpS9fAoqCDbupW9
Y9PKyx7CisSZCS+prj4eLY4k5KlsPzddOZ05TSa8W2cMTC+KHN4dqonwT8hTX4rp
j/aSHGczeoEZMOXA0cDn/cPoTYCTNsNTfTeeZNPXrhFjWaDGzpJomHyVM3Uo/ArR
g1URjiSnUKE22c4L63XSdUTv6ezWWnlamXnPZqaO3n6ns8zeT2iySnNi1T3HuYBP
Ts/idw+cY086k1MdFqU7mPL6MUHL+jSY0wlxaB8vwVp586h6MeoSfrOrogUlCt2Z
Oo5YAIjsKwz0Vit/aBJ4LO+o+m2aw0MVEhOo+Tq5+dH1TGe7E2TvGoaPo+PTHiH7
Fm/LLf1+6q3Dd+b6fOP9bV+0ZQWXIRmoh0SfPLKlDNa8PqhcjsTPvXQ57f2g8G2x
mXTtFEmS6x+PRWp1yah1JxWnNTWLHjdRImLr4K5A1vdqtr9meF5yq4jCfXzFhDa2
KQIezrfdKnEs4BVNTYCTYB1LnNrTOnBp5xpLPhC50+XEwmX+/US+YsNCSjhPX9FK
8Y2Wc3bZGwqUbOdHqFR5uwlq/k6UWgtwiydxXLRRcA6py2fEeeb5DeCiw2oFBMsu
lh+xMwkMsvkWve9c4JFx0rvsIQWDiJytHujeL3BO9tnGD5N9vm206qIh6EIAgSCq
mLrK+CvcdqR4cQO8MI4ndPMQtYMN5ug2RKhc2euGKTCS7+8Kt9O+gFtruS9TSdDo
Kr7Ur2iFZPt1Qx/HF4bwR8e9CuUEfvU4/7MS3+tj2XwsHzj+sT9AiyUezkUj+bxQ
gzUUZhtkUt4wejpRAn2CfjNOZJbcIz6jJ14y83MRQX+NFLgf/yJAapqzsOPRMcwe
riFU5wYeVOIOTta6aHCaa0zjsxlTeH12bB3cS4CwBTHIom/op5GUFmakP5w08+Kp
v0H49fFqy0DJE81PpvvvazLAiLKkRM7qMdPAhXm8rhPa5tMpa2OtO0vXqVmtGIzk
ZimHQdnCkKXoxT1B6yqORWILERo0rQ7Fyq3AkBLFgOBRLm3xlq8siFd5MX0mk7I0
ZZRBoTtmTlyq9b/sPSbjKeBNn4YB+FIBtG3OQei1bpYPXdi8rUIlI9saxLxZ/9zC
Qs9h6xQkbhSx/njjm1T4ca6CjWRu0PEjZ+jRLc86NWvQxJ8PTD7no6sHqJ2PcEO5
x0a7aF00u8jyYovVBcCggwi+Ls+fxWC5vhpKzwXIqUq23fGtsjnvbSYYGy9Np6dn
JM0zIrPcICV+O2eK5eugewIwXLoWu8OgbKJmAswqLj/LthXKNoR66R8zt3suPh9z
Vd8BzTCnKwnlx0w7WfKW3s/T1ePMsulGXRnFh2QGhoWOsf2fdPQ+hdmQ9vEmwYGu
GlUFzoeJig3gVGe8rT9+DzwRdTRsiGeO99nnfyXieNYWhuBWB1G/7Tc3qk7NoEfB
WVON2M6JFVv/8WlrwPkvjzm7xbSR17vFtgAR1PFxLiR6TJDf8+vcQRz46R9JK8dX
n6rjIX/LBDSZ1y6ZU0pv5jZWM2qIz7j7c7DO9RrwIGWszFm8O9j2yx4nssjYOHES
5RKPhh+eE0+9dwdMUDxvdV5SqgOqIc56NrbH936ny2c/RTAmuLEj6tR14D9tOex5
QFEbFff78tJtHuNvxy3zuKO0sZkLaQ1FUFmHxlrXsR/tGzu+f3132RHoldKyn3Vb
K5uC5ni3LyJa006lP5Cr0iMKRN4/Z3sgu+baLaHMwPM0ayI0WMau3tq1e4DYM/jL
7Ink/b29el0veOrbx+c/8gAD5MYecCJOdEXS/+sIr0r1Nbtflpe7yNZSHyN1aCLL
WcYJ5jKeiTSLBdJGY/SlYPdm4wj9ycbbigsFJJZs9toModlboJfN9NxoTjkiqUUP
Vm9YNM8cP/y0lcV5GQ4JHbMUfkjbtj2tBGyqeYgrgWk+UrkKhVaCbx9F7P9RS6+5
MhqKpDTbfnTR8PnXNT/Y7WgsuCYKJi+y0QGPIKcVgw9V21VqhsUi9eyjmN/Ox2jo
CvErRSUNJtR3sjeVfuIuc1Hw0PoOpi+OhddSSG2iXTbyXCUbEkjzT9JYQOso0+37
mkVO+VqGXVmvSLK53Oui/C6zaNsIMMZj2oPRtY4tAmuCME5MDfvdsE4biKW9PVAM
ssjcbDoe5SJhT6xleOgoTw8gTNAbmgKPNKZodBoOAyODvtLf+ucs+aVr/84dkNKL
1BXyHgE9cLLv4WKtS8r3KKcL5e8ZXVJdN/UueM72pQ8wpIKFpFqAJvKVMenwaAuN
LQ0haBjEwpFPf5YqztmCUS4qc+dtLzpBsQJfFCNQHwl5Lm2B2wU6ol7xNhNfHw6c
fKU8x27bIoW1rg954KULksWjoRSEjFoM+ut25J/GlaWv07ipIxOdMOVND06d+apM
CuV4SHvhapr0LZKVaUvHF+XkWfz0xUfuLrkYXubbY8Sh/iwJbXMlt6Sh0yjrnDu9
NOd+quCm7REcvfTnWOpCa7PBtXjbvDjBorQUH09DTFsHpdStLt3jL++MwrsiwPMk
gtmOkfR1NhH1p7wS1CaAtoiMYgAdWh2iklXIC1YrqGXfI/a1JNLLIa/ibBz89NB3
pdp6+iGeTyX5L+96zcBQcFITetaDZKXNDCutUWObzxcglMcqNkavQMblF7Reqeyl
eSa7JvQDgkfvqPXNXa13fRvsedBAQ/q4XB6pMHF/ONfC1d5HlWXCX6ekt5rc5sjb
H1GLjcYIoTGAilSTaEs41MevCpfm+aAM525QJ7w2jVNsDIKZOON4RUbUX//plNma
Xib7OKI0XBEUvnDz9Avhf7nDMoDeO4J6dtuiNw1N88Ybk5D3QoIz0OEv4K5myL7D
IiEjibJ7YhBpAvp9OSkfjZp+lcPuQZdYSm70YEz8jLOlsP8ICL9vBJbyTJKuVcVw
Zv0gsfJpfX3tlLL/x28QvUc55PENygvhCDzVOmoh1827k4/v8jtOGvor9fXOsM+E
SN5OqxbWV19GdKoEHRHEgcLDe4djn3zIjKRsvcbzwDvfZm/cV0HoifRmj8v5pe7z
KOkTE4uYFgtEYc4ugDcMhKtv/oDNXwwU2WWiiI1V8Hz653ZeiTAV9ppoMM5IiJSY
jhfol3+zcx1A8YzHhgEVQVOoiubEK1CUwYPlMX+IUTjC6RdOYNpNi+yYTX0uKoc9
II3Bs7TuS0pVqw9o3m71qCjGK51NJucfey9O0BZv1ZsA4p+f0OCwT5IgcJ7n+sVJ
0uJwWzDAM5bPRLq/z0G7Mb46eKNVHm0EvPPHKbfXVQOpEbK0jOhH5+Dgo3NhNsyB
gTJHifJeBbOOdCiE7V2+pQf42UfsqDAAi6MefNxmck1HDeYr257suHxAf6sqfNOZ
eNcy3/L189VpKhYhP6WsvJ7ZT4c9gWPapH6Lq2TICuiw32LNR8yBcfFBh8qaQ7B8
7ayse/Zb39bm/DxZMox5HnE1g5w00SNEG65x/Aarru6oZbskM8Wkyd/5o/lfLIh4
rBjGIXAMr5kTfiAHTm10J51ph+ccuJ6nYmhGxkHK5zn979QI5XvA437ClHSjojcd
pZz72AizMBCpFSMrO/gNc6yftR/akA9pc2CRego8s2jXtmfvcyv3ufGgjlGLt38L
8uZJVNoTu8f/CkB37FlN88km9oA90g7L63EpmqSOMMZ4gZUszlvDeomTQRziof0a
KSv3d4SwkA/yaNMJfMpYJVcvMrNXEUK/ZBKw5fMIV3cHQ9L6YDu3yVtA8qH+7bLd
/zdwkMTPR9okTurmZ81364By4yfNB957otMtPKkMBoimMfTTvdSR9Dc535nuYcZ2
IX8xofXEKO8k+EcOvNqDGcgQ8e++nn/hNDGsF6mbscMC1V93L6p3cUeGx0PfZ68L
s8XJmnyehWl+famj7QqCCByNavaOHXjXqF/gLFLc1OinyNfkRzkxOrRHRE1IppSI
ds9idH/COL4aPl7cjKiPpyLBO7/S61KFwPujOoJQ2SnIqODvgNw5qRDlwo/nAEq3
n+7qC/V+fuSJ7WEfAxNMR1OgCRRN9RZwzKM19tRzdsI/RRtpBEgmfjPzUW++0n5l
9s7W2KpfNCmr04AWISzhjTIJ6jpIAZAKtXP2tCLSOgdQBSZPKJ0EnF2IXGPUcceF
dI/g1qa3AkB+VPEzSc2OAYocgvDw1mXpOqJQ8PSOCksDrE8yWcCCycdUeTBrIcmS
6W+v+oAZdNL9Z6yUjwT3Mr7N1hhmy6NBF5RvBG4sO7YR/RnBAKisOanCFSJaOieG
58PjaY/4UP/K5GdY3QNocn1bXIq4pnO4tDLmoKiW1oypEauFQ/65ZdB8Elf3rbO8
6sVGKP8oTYfHg7pmq7gA8T3z6zPVD+D7gMMJ0bmMRt1TDYbVzPELgNVtZgpPkTSD
m6Bj0iiqn7n5UCY5BZMtWQJ+yPuu7P+l2uFrIXf/vjjASmD78lnQiStfTthRj60m
uIKEeb8R2SIMR+prdT/11cZgAjzO6nlhWdjmh3B58HTVasCRHb0Br5PLDsFE9UAe
+Usnr3McGIWgoNZQi/t+FuApMU/v3c6QjQQ0ArMcfCgGEiOTGi1/cgd+bO57CGZR
5Y2IHsIQVAdTpxPawRV6zekeHJKcDVQq5DZZL4zCkMpfO/niY+bQ/XI0yidGQ1HF
g3dI4pg6hN8uxjpsYfNo++41CJAEiH0p8g70JWJyBAnZHgjJHmRRvLds4groZb4l
VDuzi9/t2rbsnjWAh+RXCfpEW9HGpbN9XkbBfheNTvDGxg43arnLCpGvACzkguC6
RN2chrS7Alk62Azfd3fI8iM4HtRj9qfFtW5fVU1KsZRWX8/2hmGtUIaOxkfj5S/g
4/rVjdhtw3tg7RjFypoue3JPsWZdxZi/LyNCMIt+Pz1MN6rfE11sxXARKDeBY5de
gHrWlSfixBhHne5dwz/RPVrwBx6ianUAemrgcWkS3qxenriFkNtv3eNC8ZRAYasV
duoEYg60eBq5ZSt8bcYuI0Yssexn5qeZrDANR3Tkuu1ghstIQtJ+or8nQPW4oFoO
5ypeHsqqmqC0SjemGVZ+yO4zbUmCjlj921xTu4v0pG9j5D80uVpIhiy0xd0CC6rh
4ehP0E9kADoaPv4walX0rCyCUFb2rFndhFd+wg3Jg08hwtzt6W6oqkRXHZUvVXrK
VELU1RnVOI4wmhwtjYLKlGfI/JOgIY1JjjRAYn+SH16XbNI+eaRmQDAzFAqBMhG9
WCB9Z1o0QXlzaCdPs7YIOV5Z+LLv8LZwoGgRrhpp5Afr4bqAab22Oyf3peLWmhOC
ZGvLwE5br4y/6mJFZsA7mkGFMgk4MjAcf7mrzLcDrKjDJrkSjHgIy8ysDyAh/Gmy
E4dCUSbqRzwiW+Sh7+xzN6LqWlzEsKi4hAGRIGw2iXJ1fLQqfuRzrG2S6hYYvZ1n
t59lMSXw5SgMWWnp6bQKWVEyuXobQvGWxfdzEZMbds+N77pBWKybPS7+3zfTnHMC
4NQUu/osbINJEXOCROQufjgP9yXxEQ9/sJPkelOEdnM6omLSuQWFEtHSlK0MOujc
ewfw35+bLTyfOtlOM4bipsVfmHsFjpJHj02x5FTAcfrlPs7r/SGS13hbBa0VIH/D
+NJpkcCEmaJbVeFkUzHy2tYiVtvKkjn9yKAF9FFqqQqGyT3rWJbVPxZotE7OxMFZ
+5zHsXV3QiyxlKyrvn0WlRolyMlLA44GL54KizC4KDKaFeEdCzM47PVDogkXwCs0
/zueRlTa01DTZrM7HRH9QgSjk4UOqtwjsnqApEfo77lZUlnPXQwb5W8KV0zer9kv
Smt9QtGDyvURp5aHGF8PNmLIxghouTpjWtgWRFTsdaQ8Qb2H5dRSiz+WY2Z8FBie
R4G/j/uAEGQ7JPsqNYwlrxKKM0sn+xy6EEj7G1Vkx0WpXh/laOK+MJ87b3jtFkVf
opo7LazU1cOaIHbEn1lRuOg2ssU2y7bMxWmZYWoDozXfSbhFU4gLOn1aCy+0k5vP
UmHvs1KgsRTiVXFlh6ihhl5wqC/YrCFNEIsn4RzH8pN5DuRu7SdsBIqF7MXN8yUc
KXMb+HmVFkNx7Brk2NLvajSHP83VM206V9M3x+ZgVbM6IK0WOoad4Fqt9UUfj9Px
DcomrOX9EESrLj20ht4N/1BRmge/HlFK4qhQ0O74zbB5CXXM6k5XmB9O65ayfeKQ
Ll1anYQgYRt9Nkq9CKq29WROsDkd50tcXC/VmxoyBTXFyS9MB6V1LnbAY+PJTzBc
5lKWFzl/ZYCT3mcxHDwaKiiP3vZuvCyaLusvsQLlQpjyFjl80dNzTbZA26zA7agl
tf+ESUp5aqd8MJT7mhES0W5zABNG9MW6n3z2BWFCO9lugytUbyS40loSbCS31czT
V+xUhxJDcZk192+Y8JUh+3lT2wXvDkK4U8g1YrwTOv9jBoW3UHJcuBiSt7vuwAiz
M/4pFbFs5xzc2LLrTLe43hEJvEmkIZEvqBFdbwvHMUCoXE2hDoRQ8gLRp9uebjDD
VVmqmW1xz6dBf7Rhn18+QSLspJT1WcAr3hZ6HIc9NVpqlAkJSGQ4D/Xs/NmXCweg
07PVX6glNQUKu2DDruyd4oqGO36B7sRJTdMswBmjueS58kgMBtg+5rSAP6hi3X2x
27IeOjzNg9Xk5u6y41DcL4fgo+dDHxU6gN/dIi9NteaELVrY673U8Ove4RUD0jtj
Hnf14BkneziPY9LBQOx4c5Ie/iMfHuGZOZ+S/jRMTWLPxeHUMeM/RAwMg8JGx0bA
iJzZmCTTUIqigKe4Cc1WucH06iyrl0Uo6PLUY/m57FU24JLbMHVTx0k8GgP/aGzB
l3WQko8BhlF5mR2MVbHU/+2b7UYuGul0cx6IleB+1aX3nyIa89xvUVqbaVJ3LobI
KNgsxucD2M5YDelWIwFvt1teHEQKUD2FTNPPihwEMFUYRvn8A2mJLbMw7Tg1fdKa
W3HJuLNWuOmoHLUAg67ZtS3vqTwZUVhQofMnt2SoJNpzlpvWaJCFRIZq8PEbH5Hr
Q64UeL0QLzb2cWKLxTrAr2GXK+J0tZOKlc6jeaKtuO4fCROwX+8pU8hT9gA8b5gH
BGz8kD+jEj7OmkxmNSDR+AYJV30MajU0p4cKnS1sPxyG8+O8oFcjDmCSd7KjyC2D
/wc1lGMvZvu8Vd+EYD91IDk3OcyARDNOmABCAv0qxrw/zR1vLCxnO1vM7T6liJ9M
h2BHENJ3LrSM9WtwcnPacK6vwwrC+QR7gjh0CV27IDzPZqgFE4zh203jn/5GNxKG
yF5aO0vkIoTWgTBngctN+ARnesqSMDMY1G4iuLe8R/FG6eVmPy/WfW19/wKdHC+z
uVuGh1v4mN//y8GscQjoQeKCVh/x0q1dVEF4qdJcJMKx9OdZBoeWVQtW7nkL3kAT
4Swkhkt1njIep3qEjlZTqCe+uOkHrPrTj/ROwgECykAMUXLnE/LiIWDbuNfHzHKB
HO2BFTxQ7niYj6zxagm7tzLnX4Hm6dCDCStKxgV8SD7FIUhOT2HV7PCac/W2eSHi
9J2OZyfg8HyZOVppubdwHTLgCJuEZzmSY7aVgOfzLA8z4GN56QptcHonxfMMekHX
1sy6WcXGbnsY5uAtYh3dHsFdUwaQCZaJ532qVx8OXevgrJLWQCrpyUUL+N+PvjNB
OnFqi65A7tILlGgDyOmrfsFkx3xNljt+REHPoHkOFjthmBpBhsaEBmIE+l1iJJXk
2WG+uBDW+SGH903/DbkWkbuty7mmUe1tZs78TNOFea3YeJqGTE0oQ7yiRxbW+EZ2
3+OfCT5cU7QDgNKxC5xSA9/qY5lPRz3v5yIZj18/uEuXRkshBsq4+l24SCLQQMNs
srSpyxTRAESXZ1lG9yPP3Uq/wH7x/4tNX3jZktR2myTOPHZjnqO7aT/z8ldyNyTK
6w3to2PVcAl2EkqL8hoAd/IMjZNM5jA87ai7ip6ZIoTLEnAGgjAZ74kzAdDv9xfk
iBcHijh3bezuHnSzUW11R9DTQneSXNPkT11wdbFQoECMpbewh6Uy7x33y9VGQxjZ
jU//Qyjzf/ugANpy5yIGP5vjof3sayaRQ6D6GcLrmqixxEcL7ZNvM+QWvb/DTMf9
HfX9n58VEoX4yWkSxjbNJEy4orbfCYD+joH114uj6TZmYmMQmJrKFr3D11uDKCmM
cuq8tK+pQZPkQexgCgk6qjL4zWK94jmptHmkDLdL0RcVUsivEc1Nvr5ZrN3bN6s9
wqBtrQA0VQPfU9L1MEux8Axfk02BnPou+UlLbFY8aBOKT6S+LvK3bKhcnlZwxoxl
gJRo7JuSM6IBPVRlLn27ZXG014rgnAg5qxdIDmzCGO7kTesWtFEjg/vMoucx0MsY
KXJyImzFuql7WFdyMx2oluZrkLi7lSXtjisIPiAbveMeZ4m1Fn+yxklmtvVf1Hpp
TXdsUHS3fWjXJwlbrlgJbED1KLtXoCK1xIrAw2M7FP5e5g3M3i8wgr8+wzV4y0YW
oXYzzRSWoVpLhOl04CiYul/jelAcaxspYkGzh7/HFcD1XX5LyL5qu8HO2bbq8a9z
83rlQhyOInwTfDHA6fPpkLOQiqnG2xc64CXbmCOmDyGJW2YcbiapRiPZ8CSRjNY0
BzPx3phDSJUlsJIPa1DDlSkVtLsDqsNybbNZh7OlTLi3ev/BHFKPC31EQxyOTDMq
qEnRHs2PUl6VogLuj23jggsPqxrkc4VXnzJaVJWeyMg/9Z5sWgYmOvHGOqtSQ7XX
4R/oa/KYSCH1JleL0md1JwMcugGw2qVjOv1tioXpORFXV2HGh8oeHULrM8zskLQG
fol/koebs0lzLT/ylTQgClOgWfKzJcD89Tm20ZpI2R9vkXLYyywGcPr1LASZkkem
FdEFYWlj3J1D6BgUpi2mwS/CeuN8mOU+lqzwfndOzwSq0LQGybXf/0dRU2rGmiYm
+2wmlt9bmsaQRl/cn9ARM9PgeBnNScSLXT+VvrDr+rTGUs4Voi1r/N/MALOTAiZp
780waYDYRNgQg5GiSoz9JlCrYob998XjLuC8eEqD1pyNI+Bbn4oFIUXL6w5EiBjN
K4gxLST+fxc+tFVmunJsW6JxR0jTJPCbSc38Su1nP+ZUGh6iWzuo4ZnGKDioIpB+
KcBNPmL8aX8Q5DfqtP5Tdj1QZJiu2sfk6/HgOQBjfuvccQrTe7keXM/ssDimEfOM
yr/xfzuPeFlLyzBMFN+9FaqpfFxCOJCEzHuIwpythC9z7Ulweke7Orq3BM415Ahf
kpzjQ986TPs0TQYIaktajgq7t9EyIcynNdxvgytLEH49L5TNcWwknbAPSFr5yUwM
KL6/85mY80qsVA4UdnDtLB6pWkxfzQmNzwfchVAB54Q9a42OV8zzdbtzFU+Pci+t
/a2JmZhaXb8/gTvRwDwa+r84mV68Og2ke+NAZkb6LLDOUVUxFH7caznnY5QjM84S
2dmlHNxJr2rYlmhBZudfQKxaHrUR6FuxVnz5YV2OkOJ+eXhhH4Pm8TAJSZWhUdOR
0H1YPTup76cSDrx0gBTkT+pzKaJOmQByib7o/rC7e3daqd8RxtS1aQn2gG0bTxwz
RmXYnjQujzGqfO+3F+99xL6Vj8kN1iKLT9JuKlWX4xDq6pPaDFnvkJaf+0FGKNxe
qOWTHK+S82rokIjrkTLGwRKqi8Luen7p+da36wb75+E8e2tHzaHA2MObl4wLD4M1
8a9FXOnoGmDZeeLKiPo7AZXLGoQrNOiGAM4M0Rz+IC+qndmI+3I8AChzkSGcUUB1
xwuulC5R66+X11/ImLy2JfXlrc1K3uPj5X8o88dFIDRRznUFL4YJHcn+X9qjvXQC
y1dTz7oyCN7fO9a+lNi0ElEmNrSzwwCzhGwlkoj8rlzv9qHEXxkWMHq/YPV1ijue
TmybHD35LiefUTr5+EiUi4TfXd0bAk9Nh+8FsSt4+XjysVYHoUuQLK2gX2YVQJL+
M4OvWrF68/wEMIjtN8Tr9N2O4nFoieQ6j53l2p4Ud0SqBn5ZvMw4++22bFaly60T
fHUG2JXFkA9xRrWEc8vINh49BwOo9776mGc+J3G71TiMlVjvAtjxtWiI97WTMegX
rKE5hxPWdGPCVWK6ONm4jb7MpzhdglQkl75u9KhzI+i6nCCVIjcu2vCF4VIerG0t
P99s1OKBpa8xyhBPLINHX8VgA0CGYHZCRogxKwNRFE1jEGbOxw3SeZvJXPEBvQxU
XZxOBxXSESameh584XRnWot5o3WDGZ3daLiy+02qTangszQINdx3Q6efqNmUvf4s
mqDDleSvFmOIXjKnmmo2z0PqurBb2xQh9aZuLHflzf2P2WUeMkBcmyITv85MdLzc
MbpOK7duF6Yewty3ZJC6gkYSQQnb/293KGnLJJEA+kg1rPLh+86Rs67+/mZpP16h
5+b456F10+gDD5V08OHuM3nicb5YTYdviOZ/ZQw4D97vCQHv8J/uDI3+KzpiSX77
El13oJefjoiFDu80eieaW3eaIBUb0FQHHSRvE1zVqn5vmN01A0ePDuHTTXSKdkNL
ll2zNGK6ka3kD/fFr2XSy5KuNIqKpO4fky9nOZ3fgQoFPJl6PXSIbIzBUBEjwNC/
VlH4uNKfuOzRzfcvIXFNntohjkZ8u1JkOFetEENOcLOpZ7icaJUFFH2FLLUXRUcO
0Id0XQgf2+E2QH9d0yzcd2WBvVVIzSmhYAcfI8nytvT3jGFSBY26Mcji7aTV4vz7
GbmuTs7m/VB8SgIyibznl+C+xraSrWq5KIVBc05lMRJt79q/w5BS3woU4uN//Zus
Dp0uCKpF+R1m12hyOqKG1ZvO0Vvd6PN6Hxni7yYJLhZ+ZE32bfqIOh6i7yJCCmAE
RutxwtAm0fl+B5AK2U1xBjRMH0yWmHAWh+XopVK2INWnORSF060WWghe8gpRc7nY
cXABoyKcYU5SQbJtcDt5JwmvS8reMgkjtccHoYAsq4YVsEjebi8owFZ4qWuKPeuu
ukSPIllMaib6/w+Fv/yTaFrTKi0EFZlu7HDGA30PPofXYiwn7gC7eRkIO7jzCAie
i7co/NYH9DpgmDh6AGaPll6o8X+K1Ss3AVDhMf7ZEcfEJaRYIoTeRHnarnLsFFW2
/1CSXr7CeyeQNCWM/IVGV8CECpn0j7G/kT10UF8c5lsvl2gHjxc7XW2588nfNFVV
5lhGYrMgPOe2lMb5IlB5P6ChbITFR/wsW0e9AL6IeUk=
`pragma protect end_protected
