// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ajmw7c65xH9cmt+9r17zw9LG/gKAtQI9mA5H1P3drROi6f21kGOwGsv3uZyEGvsc
MeP8uTWf2F4T4IU7CaMImuU+PqSG1Vn9NJPFy98OpIBfxue0UimFp9/Y3qKOv3ns
XW0m7RZretwd+dOK0KFyabFeD55ZJPIDbPhqJgdwegY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8432)
TRbp21qGo7g3nAH8u9n2v7+9/hOUMI+oqTiiTjE98StMsnq9NKvlh2vzylwEQdH2
1ESh5Qmew3CyR06QZxlW159sAjuTKo0QwNpsyDe6JRIlLEu4DKc0VZiwW/q+bTUn
O4JvjTdLMzV7Qm+c+X8GE9XLpaP/Zbd19+j7onIPhHVcl4a9bu8O7Y7cGW2JKJRU
8uGeOg43/5q5Ckne82axG5OIICJQlMGhJu/rlUtGxv5eexQIUTx8JCs0Vok9/1Uz
JVQqnKCcBO0Nf4av8fuHeFoaUKqODZvus+l/oe15amWXoJ8wV9q7NG1m2d8yIR4F
iGY9x3jpOEjQ1fqfSMZKvKk0d0u2VeHmvaxLt3KQkZKALLYIrXyWbrvJcmejyoCc
NHtnccq7T2PQk+VSIlX4MCyLNegdHqXEaZcN0Rt9B2zfBBjAYj/uNp58laL+52Xw
DVBN3MLn5A2C4wCNcajIxBmPt00B1HLE5bQPrfTxfweioy1xzT9Z+9HqkpeNPYEB
ybzxx8/urqTRc2a2Zj2rH50Txs0Z0702bI+F0Ol+V4rQfvnQs7ENz/erLutZ4K5e
HQS8qn7W+e2m9jrT3MKIFyQQprUkgM1A5CYTXAPzxLtuGcH4hchGnqeUevXfgN+c
ZDkPW1tcisuEFsUgSB1IMH2BD7RlMcpTZiGLkBmjOeil1qKLIrSQCIQyODbueO77
0ikA2uPv5/S5gCSKUBgSz85X5bMOkoe6KNzNn4mS9A9pEcA//peAAD2hneU8Slmc
BKaVFNbfpZU5be3B2/XOEmy+Mxc/vnzbyzddeUHb9huMTj8qJ+p2UkmdmK2wCcGS
rbxQqxgfewq/h2QBJs2oGqUp/xmqliQdgi4Kij4Sxy0xKSXQlXgJXudBtuZ0kmSK
LfuLqo+SyHjzOzRcnq+vsFS786jk+k6N0EU9ORSffISPphHIs1ad7qA4q2dwjo+N
4qCnu9kyrLJXKrkHVBK3Iqwiyo+njnIGw+/nolhtHbv0a92wECnYmS45fgLPSmdd
oy05yCtgsmCQZGn8kA0pfexbVhMl1NiS9MywNvQHqG5vizWlKdWwv5F4e1lk56vd
7jWTQ5L+q9fSC/+h9rSjZhGyoXo3ROctAt6n9jLG16stGn4sgxiRq/1kuPmzzfJl
nqZotqNuCD+uXZflwKsCZxmvZ5hzkrUXEY3cEmbu+UekafAYjLGPFwsGt9rv71ye
bUYw1r2f7iqOfgRQdnAoyG8WqQZpaclQDyTY+Cuf6REXmWd9T4cWbarlhbvt5MJB
xwipScjHquEqFks/FS0LTkLBzkNxAIn0f8X2wdBFL7/rZUXZV1epvzqEBz3P8lah
5k5VBJ0MDspCOZkG6hpsn8U8N9+Ktx2WWJSyx1z6RZArWkKPcVWVcZI+z4+DyZZb
c/ndjc0KtPaQTCqGZpcvTvbbyWBpgVWLjqoWBsApLKLKWFERMLjwo1oVOygsingJ
tKEEjAstd2Hai4AJSw4yLr10IrsaPaaQ7i7FPBnIqd0A3hJHHVnu0X4ZeUgNb0eR
xnMXnw3nBf+5z0Pj1FvddezYjxJiSjuzQ2mRjRtZQR6AtxfXEFn0o4lvAbkukKlC
oycMsmL9JHAKtz+zkwaXpifx1ucidYISIRPL2GKZtO0chliBy6HKU9ZIkmCBJyHZ
fteEo4y0T5uw/2B668pjE/u8FUIp3tQG+lMV0Eaw/zdwk+OJ5NXHKB0/Gfe0bKRM
Mqs+F1JvRwYgfdYMV1aCmTBN/ZJr6N+gS7EdmVjdHnhOBId4rC5AzAM8FKMVfBGT
SNJ+0m3BTgnnc/a6h/SjM+BXvZKr/fHkWmXdlP2wOZoizKyf3uHF1GA2ZAgJAH1q
3Ij7UxBrf8namapVeCXtVXi45Y+LCz2MdNHbIeS8U3Xdj6ZdBSNSz+xQmPpHyEe9
JeGVCWV71zZERGSAGiKQRjyddKKf6Fpk/w2knIvurNsiv5iJ/ZKmPGgm7t2CHmAV
wjHMcV0rwSpWg65q914ZtCPQmLaPTYIjdK22HFEiYGTiNi/j6KzI3C0dlZ/rzXVd
I8ZF9wr/sMBvpsHa0LUtCsCIXjiT1LrlUjSkiXAg1PZMHDmes01ChKBvieNi6LqM
c92Pw+8fBp5Uc2uXQ5FLYSprpRdw9IQQZ8h6UxiuE6F35xRBFMH5iXlfiI3T85+5
vFMRHx3InxVVx7gl/xEoiC6H+K+TYRID+sGWMyqjogSTyyyLk+MTPUixh9MSCtew
MfAY5O+bxblA+42M6HPD6XOoVP2FjHI5pp4jJ29hiUStn7ndXJBYZir4k2swM0/W
HRbhdHLas8jpQ4xEqyTwcOvAk8VAqMn0uqL76QmydIYgbQf3pdvVT8kx4kcHz648
BIP51pqQ6U+vI6GAGT+a5z/a5N/s+VnYR0In44Aa5CUV7bgNdMV6YkBcA+QNsXJZ
44Y0Gzj7xY+51Y2pVh6nfwI3d3NNt/5mLp0n3wh/Rhckd64Kj5/u+14SZ8GNDdP+
zPqj2R4h0GREtA/7RFV0RVbgcbnZbnHAh66nlfr3kU8lLrunPPYpfmXbwWbeds13
uIFM3iKog51jaJBfcBRwZunlOOjPx8PDB2ximlmLuTdNxAWdXaqACXdjglMYGbgS
oKPUfM3Zxx4DO678JDd2sdndpvBr4wn0ZUOO7ZbNQAKfpBdiyStq+QwqDSRCr3Ul
9ZjAjyB6o+ZN2BlKi0JT+L5mXHHw+aytMvnLQpv+V1WWKmskBAnRlJIrFqnsvksx
BBcfFe9uctzwemsT2bHPkvDpNZlGxZu+8UC1BmjX7HJvGkHnvhBDSNVGGNsM6LSe
uTZwJNSE1h+MAapAq1uk+GaegQG8Gv7SaPiuUB54bvlfD2PAh10yPYFMXx3BQdT4
LH/FycmZLB7t9Ma9n3Tmsfh3GsUF/E1sx0/a7bA/IxKvGBiIbhxj4S66USC3dxBr
lyJRaUJNueALjejKoqrLLoyaJkMmSuRD1JKH8GRgRhBJ2qzIpEuDqx5aTsxbWYYF
lplejRuWy2/ZrbRS364rM0pKSoJdBS2FiEtFvin0BudWfQIg3AgmaaY0evD851eu
zoZlat0YD2avk3mPb/DHDMyGfERFGZoLIdZNbylGDPfqoy7UimwmY0lh4eoPX67h
NyKRd+rb9Gk75ur2DctvwCZ82Khxw5FrqTNcF5HHAqyzazTozHmFyQNYsZKQUfFX
BRRDm4md71FH/xNsJwQFKiJnup5fdRoSbFc2/l5bktwx4RXeSeJhbk6XJUgC8L+K
BJ/3HKGJPhusOzoLsd1Vi3dq03jsMuIjom9cKA8E53VaNC2x+WmGgG04SjqY04rY
3S//HcrLNDdcN7MQixO4kSFw9uubXvmZa3rjU86HUNTsRDwsmAa2NliYONNK6zzX
/5FiU70qk0TjU0lSv9Rsn6QtninAI2ZPDSynvdey3w0YM6Es0hxDuNiBKQgzEWkz
6O1E8f5ARdaMNJzKaSOK5ynaOjBpOVZtLiwkIOaqi6lqA+osFgH1Co6Jstr7wWya
cY37jvMSG+ZgnbdsDnbscJLYYkNIYENX7zk+zorKQkoJeJygP3GD7qrxQJFwrLOO
R6e3zC1A72GGHMX9XdUpdFZ9e1S2NeZUNfT2Cf92vOwmKmROuOByvz9E1m66Ak94
GNP0Vj3MupRMFO/kcEUVl9giy5HlnanUx6hxOiihnoB37i6T5IDWGJP9/udKJdLV
iFai/IX97SgHKv/Te2poXJACrjB99z9tBwxhmQBo3L/3G4qtCGXSmxHL8wcOMn2y
Q0U0VHlk87RtmqdBS76UEgla8LGIuS0sxNjByQDZ/JnWDuhzf7DV3yYt3P+zBVis
y3CplVG1R1UEzGSp7u60Ogy+0vAtVIR9bqc86tD37gIPz8fhT2Pr3i+ZD+0jMrjb
Kjxl3Tm/RO+LbdBxYqRnNsouU6g+1rZSCU17A7OeRLhzUmm/rv2jfN+65Lskpdhs
Ay6sX0gWiYr5flASYZJgsd0CE7La9tSW27N6qhaQOk5BY+oAsOjGUksAuInuelut
ANu5TFjUp8M3c80W/y2muBWj8uNS0RnbSRl4eR710KrgPjxvpPEHW8u3/m6QxJYp
1XcN1zCps0hZe47vEyEbXEQZjWYFprnMTCsvqE/Cq+UhClyA+fZojeszKwAkGqWx
ZOhZ4aXg6+zAhMtGXsXRc9mRp2uyng24ZC7kn8esisGJMGjVRQjcbySUcrwtJucy
AOkYMCKAeDP/zJ0aR+t9up+M9M9z7E1I+F4JkB+jmFERUq3XglWiWlDrx7yKzaiH
SQC/9NhZFwTGNHzv3CpVp1hfXeD90gWXV2QqS0taYaROQksEhfd2DUNCwmcdcf+D
+SbdYyn591iCC/dEU9W+qwdGQsInSHzD331gM+ovgUCDPQEfbCuz5BX5oRIcfpHS
OA0EZ7qPNXR8wNry9JEnpx/3bGoSKz//qFTwHYQm2aprAEXBvfDShKDZc76MbBZH
x8CRCGJdVyXg43bPKRdKRnf38YI5MB1vhKoBbgf4dz4MUkF6r8oSkNhbOama+L/b
bu+v0WRfhxMr+qEjJCTfQumW+fdMhJe5fAgkAoJcjbly5rwC6FU6Gvlin8gJ6ciC
INab1Fk3bB2de5oykfTsrU1eV/fy/EOBwJ3oM4cH/cSFGI3D0qLnDVh93USxQFY6
49GCdj76hMnFd1HMo5Pd+x84SV271DWnKdKbBO1Vao+UuCJg2ySx8GvWjgxFf2l0
aT56Q/9a4F1uryDqTMSLCyn1AcXrueQqcFhuqbO/ADYHfhy5vyDFHQAmozOedUXL
VYXTt+kdt9Rzd6Zp0M2H9bGyTRUBpCE1lSAKyJeerW958fMr8ZEYEVn6JbXNuj7M
kGaGYt1IcnO4AhXiqem9yrN8a1zcIl1m9gRgUBijlkmR4IoRZTs/q9mIX08yA85L
ZWdtOs2UqGGGE5Ye60dgeak9fhxDP+i2Wwg4Y1aU2rGqMDpo/zToW4ET27Toj7BZ
C+k79qX7ryybK3VJ1bJQoPthqsJ+i4ayXshlQgKN4Z7RvpuMUXoKhezwJaXfykAU
c7zjrQHhud3/BfKzWnthinUPnrADH2Y4s+tETP5eTKdjqh6Pk1b8a5RU4cTj7JEE
KbZbSaoV1hruQ52m1qQJUdgVbhlWo+yl7ZC2m2/SLFMwB6VM11Sx2R8lM9D1Ipsj
btyfSBr3PxqnZM7fO77JyPSbgs6gcJoT9BDACGRpnCZ18g47nag1rSgCrzZNZf93
SiXnMuxKA1/BeKRva1uNe3bBqr8ZpVM7L2dADLbANLlHKhfc1jBJrrB68cm7CZSE
sXlfyqCfEETvt/tTTHB5ILHVqTn4qIklczC5lXdv2CyjbL3AE+Vpr8qBY7PEunV3
QFbnKBc+hZ1lEI2sbaqq+V/1gV0wdxkTfin4DspyrcedMjD60nNpC1+3W1V0dft3
IUaotV2eZoctU7F83zuNePEWiL4qqu8QQwJKHSn3dSFuHcToMbnqylBjW6b4oNqI
+NxUaBDUvxXHCvWrDFl6Lw8rezJ/qdYX2HQKOIo5q5uzhsmWUUTqax3QA9/ZPj0x
zloKArsGMqhfCSezmrg/Q3xEQ0Zcqked21fwZZ78vl93B6e/PBTzH3IEG5H4tiT1
X1fyZfoi3wvZzQpMBhJsbj/CWcwYhbA3z5FrPNRBNijYUEUfLkBIrh5q+80O23LH
R6AKzHAgJ5LbJq/kPqIEVvJBdIGJW907OfNYVA8DPy1MZd9uPYXfZus6aIMUryuS
Pj3TLpQjihCcOD/CFamX4Ejc3Hjg4kyswqVOuJaMBuP/4pevE09roglY0zJxNNGb
d0KqfK3prKrZJPwQWmMSUP9l3VYFrkJWvqJSVHp3ZKIi7DaTAiiWcnJwXVYOWYp8
aFIH9EHwOsx/aqpVGLc/xlZYQvW5BnmRYr5XyIswZUupBFPQohxwbpeo4J/TH/Pc
VTWVXt0rlLtkxnQvpVw5bwzFwTZ+ty6HkQNmzBriD9rr6cXvG1P9YQj9dvnwiheE
zruVuico4R8EiwgWQ7Y3g0MylqdDaxgVuDCVigsOXKoCABD4JZHV8syVNFobvW8e
zY8qBg/3uAumrwac/O6SdxLyaZRma1x1SFlq0sUYBhpSqd4JSODhXNy+STcWZm6x
1FbDPqqDAKMP70Av5TZKZbCnnvHfQ+ScDOTW0oNiJ5BxeVHNzO09dlgQKcsm0uZC
Htq4/Z7qClAii5lQC2sJwFCXSfrRmgNIVemUjNZg9gdhF1gVoUODqfRK3CVDP002
/b1aiYvRHpE8eyWcy+JrP9S7aUEzRg3jHOBpw6Yq4r7I7Q7V92Y+hHS6VPQdX+30
7jCmLKbGs9qDG0xD59lM/qJt99fn1N8RyDFtOi0ZFA5X/PkwJ5f1OFipZktYCkSt
GaGjnvJfe9r6NSBlxdDvwP7HelJolQWKHKtbEfSnz+31aWxSVMcQXARv1Mp0KHGY
BgB8FWdfVUncalsl12vpGP+gByd7cCR/k5f2JbVeKPHpLI5a/mONLmm6pcIMi8c3
ZuGAdwb88yROrlsoybtWR06HFgodqCkTgYZEP+kpkWLVZxl3ZBXs7Tc4AxxZT+qA
hpcIPmuRVz8sXYvPYk2Bdr9nIPeyqKe/VxM1dR+1XtH9lPF9wKfqhSqHJHYZziqu
fZlVsYOH2H/C5JJl5onUx/1hhyAs8Gaxj2DbzXlTvXUGdZqa2qs2TLwLTjRz+CwV
aXQ24hiuWooFTTuKYnrELYz5/CLxTq1QVXD6VTAk8k1i1AAt7HfWZ7repbyGHbCH
+Qc47R86OkknLIQ0rVWonNByTbdjnBzNXMnCpv0LFm9tN3i4EtoxR0vnACY6Kgjn
xgCntif7BiYYTYzmdkdzi65Z2W7S1rNufwvUesiQTDmqQPqAa/HW8FTVpgy7QY0/
F3XlBWQnPXbMEAiB47IA/JAzXX/VRA5doh99hj8gd/ZV180PvStaTvKAKLyEVl+M
qMLN/oS3DflqYZoZLE3mkZkoVszufuSF8mk9FhOynw0xpeNIa3mKX9Y1Jwe+74sU
+bp/RDPje+x0sHeGs6vEFnhmYCRmLkzJkGZ4ppO4/xZ1Q5ZLbtwgOlWeHHw+0Pjc
Os72QXz0tlTRApRogRkGWykbyvCQheigEHO92k59ydJRP1TOvlqIgZWldvwmOuy/
EB1A9BeIEVFoLWmwAcp+wPirTsedilcLQJOCwOrteVmcBXxgzUPAWadz7L+b4ogp
KuJSzMam5f4cYGGxLlprLEfrT0RW6YUEW4tTrHV0NMMnHd5+GDpTifpP/x7h8BE/
MHlRwqSkr84PavMuj5TKZFPXINSBXU3PLDalJtlDJosfyjguQXvVLSk8DydvUMnK
89rox4Ibj3A0dNnHCmDPCgrvpbshI9y/DQ3G7nnZpzuOGDyTn5uylNctukEgG0rJ
p5vPnMcS9qTal/QjPeaHBIZpS/iN0djTP6UcdZojcKDtbc9PCOQr95PK4n3BTJNd
AmMqrvdOBgnrMKT1lqenmpXDovkwquhJU9GV1vKdNelnqs5YxqGb3onIirCx00mt
8qwK2frt3bRZMNlT3MObjngbUykN7JJwYC5+fVt2wmfXl6m9PT0nA5U0dSxpKPWY
lpeIYvJ4MTf5n0oqY67ykYNXr0xqZ7s5EYgYTc3b3xkrppQzFa9tsxKdqeEiprOR
s61m/KEnVsqrSZRWUMw1Uyb9TMqhxEP+T8GNNgPbfuCJzaYfZE831gZ2CM5rSGjx
HgtCuEhQ/2UsCANFxwruQn3MR1+2YgkNAUoDX3NBEolmDYj/hXskBPVUyclQ7XUI
ZoRCZzjf/kqwZ69UeIbk2h7md1PkhnfvdgvIdNW2RFTflJlW207i/YNGjLgtPYAW
DizDL8Rnr9toGn3k1z3EtyCz31MW1xp3xOoydy/wbsRpNnwI4IfgyWsXf4dC166r
AkA3maxxUzb0FpaA0pDDEfa35kdNiXqdbHHbZIq3SPs2FKmvkjLv5ovZg8Qoh2Gz
K2pihzI6FfU/dIXrOQ9E2bW+4L6HdA1MmIhINvh31P1tDLjoovkzss4YTd55ULFz
vBgsIgrYNicGC8ZY4f0SAVzbgAuA7i9gv8c12y3SVuiyGVJNPSH4bNzkTVYANt3D
AascyyPNHZRfO3olKbP6sn4FUWhaYdrqHNaiBrPcNxbcBKHPGTNPiPloisiXZMam
O2+r3j3KDsPTbTBaSA6SKJ74xjiEV/1Ti0Xeit2AJc1cAHSic9JnAgHi5AQOrwrg
PHRoKtQNAWSp/m8wTtvG6OdEtItoQ8V2EKbsmGiFD5Nd3fiKvfxwBV0T5M/chLE+
TRg5+8A4KZFS9qXA5yJyFO4tvehV1DNfX+OfHW/AimLH2x5Q53rg4fbeFd7zgtMI
zQXJOJ9tZGXi82Dqbcv9pReYy38bokQZHUf1VA0kJ935yOtXWmL2aDwuuhoYpOQ9
InB82CJeK+OHd7Hsswc+dGZfv5KPxe4FkFp9XH5sjQPWPoIRJe8D7bWJb8kBvJmG
FF54JnwEtUFMdaYYIWDjbSD4RSa1FGRWiAuRvR1tn8zBrDpjtoXLl9La1cx9TS2J
k4hMZV/mVdgt0THw8GAD0FOEPP3f2l8vGIwTSmBfX0XrXNfgowM5R5IzEgICJbG5
pXx3sFwGMCgA4BrkH0hoOgs9clC3gXZULUPVmvFzAGOFjK1TjMVpcNpaKHroRkDK
pNStvTHp/4aJMaFl0p9KlPMLMZmIFynUuby56+jTSgsB9fOD+Rf8q3L0Chq/5wxW
cSOINqjMWW6ywsI2FWyh0eBasr2Bt2LU0xcLpHCONDA9tIfKkqVNRyu+nCAMr80K
ez3z1Booz6jcNqIVR/wMteFHCtj0vNT6vFuijpKwwpHXvTD3As+a3vXN+oWA3629
L9O/Q8k/geKz0Dc2s60C+BQvmbLI+mkJZCDqdodYX/6pKXxK1wUH0+SsFUMW342q
DhI7vxY6r+uLUzr2aukVKsteMhK3R3av2OBYUfyZ/v1Y3ZkpWRZo/4fn7SmWJlgp
TeQzlb2JurkzKTP7pA2pJRiLUoRhMy5qS8ug1K2faoIi5phZhFaSVOVDtmv0UVqt
PG2tEDdYHj8nLJO6o0bta+UVmwam7jrntTZ1BCWhPCeVK8DxsRVUJJ0Q1daPB0jE
vxl8foE5Lk+5+cuYLnaxGpwhsXwrMGpxy/i5PRcnM3fqd61HfYdeWX9aXJ7PHbiC
D6GXtBjR8rFoj5qYo2FT/NagS3Y0ZwjlNr27EkBSUgalxI99UJ3obGNh6tGCgvUU
toOVK2ZFDXzA/Zw0T1sE+pH2C8DPZBcveieKM9YkN7cgN82CUvQbubn8PC79+a0s
6WZFQ67hUhDPsN6BTqKbrhX/16xByHYYTRJWADZjDcfj4z2ynERd1z+CkvN8P70p
M0bKcWulm7XixiVQfvLpJkGQCFwgojfxieED7vHzBD+I0ujTtJpMEIAsniTkLK2O
Y58ZrWbNY0fflnuy6DhVsSe/QCIewBEMSRfw52JxaMW03HdGKLWzPKiH3ijR5rCK
Nq9DZKBwSS/FZQIhyYRbKoOFZoScmXl71l7y9M54kEiO5KtpJTOEPhLxbhEC+xBA
O75+gxzEgbwnibMQ77SnHKWSjY/LRFyYsDEhZHu5C15gNUYOnDFZxNNEFYB/VNeP
31ccVFsQTbq753HVG5TGqpsGfxGeTIJLWhP8jUM0GyF5gC48g2bcZokWLk/XWwPk
HxVnpE6yhhwaGMDtoVy996r54ao592Cm/GTFN7MBoAONL3EluDhfGsjR0UFrp1ZZ
GIKXmz1cMR+nz6ihXojwLVou3slXjudhB+UuOg6sQ+nCUHoXnRZR/0Prf2tqxTmW
VxS4TiKMQJMBbZL0uRGdkflnujlJnx75r7KHqkR2IOu2SuNZudDiQQ6R32Am49Qt
wtcqnL/O41asJvhQjSbiiGFjYZqJ+xqQy7wdoJPqxMF/sfDcZ443uw1k1Xf29uUJ
/YFy5T4fOrn4Zc52yculTisYd4W9UKK1mrsphDWvQEi/Cei8kd4D85MFn1oqbn/e
HzJcMxMPFgYOAvC5DE6BJYzCLyN2mRJXAW1xq/4MzfDgZ8b0cHsUWTJx2HK4pEe9
HzWZCC1bQyPgmQqBHS2vWANDZVxh8vVxXRmYYSX3MxWvU4FA2GpQjMmuSLwgeds2
FAY7fGtPSLu3eDSlMhMplhDgjsW3PAG6JDn7Ly73lZStuxa9lUoWN7wr12EAkXWH
JJQ0ZbgBdI89sDnw3J8RHljOnGdIQ4uFCVeW0/mgPftZ5IaY7up+JPIg+IxpkjBC
e5wT2NlYh9gKyhVknsUA5CPv/GChJT8Pi+3oH5oAARGgiuwzzVPT/IElBRbm8WD7
sPK7uCYmT7xVcFed8+DOG5vSqxJ56qJ/dGcC+CJOCqDMCGJiZdgCFCogtvcbZICq
5jaqbrxmWPmBswN2Wpbo8Z91Z+51RaoF1gjogPpUBQWnU4FsjtyuUZyGY/b+rx17
C3rzsLMrbCBR+KTKKixQOxSIZ3mMwcgfzCIE1dGNCQpjEf56BpskuSAEd744OyuE
2fAhFLZEkdOwo/Q9jYB84FaPbe247gu1/0khMANF9bZPFeiQGIC0dlOt7CxdFDT5
1Rkiox4bV8ljQzeBRj0a1gSGyVGOb3aNctae0gQOnMGRxE5D8CmoY7wZ04F/DqYH
79m+7gNh3oZ/97aYJYlobxOpQ2Wr3kKZnCbX5Xxul996/fDRRuKbPkNYtsCQAw0j
FM/4XlVsvVp7fxHRGISLtk0gl11osZIfyZcHIA3hhIs4FKBb3Qmn5/lSQBa6LX2i
CqfVq2tFtQ38GNFEzIB0sCVqecg5BoPl54O8O/WlcC+1DMqxolnQMwXB4FhQy3IW
6OJmAljYFNrzMCcWnxAsiOM/07i4FEZXsCA7NSmWHbJ7ecsIRs6uPWFZjp7g40P2
RRdH0Dv9FTIRGdU9HHyLsac9UY5g0iP7ZjgC8vm4a5ehMOxPF01x8a8TxsiBdyLP
a0fjy1El5Y0VnPji4uyyxozw//X2CJftKZXTMGqUVvze6OMhC37kvmH4aqOxM/o7
kVgIvDkaqKqXnvZbxNqWdgVDkiPSHPRP0xOvwPFNB7zZvx7Z+JcfnUyhiwhT5dbL
GmGVmE0ELaTU8zyafa4klHeQCDxvNM6HUQoHmQlM5DRQ72zqvKyfhM8PoLQTAxQY
0G4gRLY2nWwJ9sAcN32Nm1Qhk3pdmqI3jql++miDKKE=
`pragma protect end_protected
