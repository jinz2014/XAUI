// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bRmZiwNt2uF6nFdIgbuEEYAE2rCWBITZlmRS5eP+JLY6gqNBco0fEGKWdJ3lf06f
NTUmHf6TsF+TS7kNKqt3xWosAYt12ddszsY87/fvfm3gGgICWgXI1LMobMGxlbop
zqgegpf9jbHuM93hgt1NSZXtl3qUIlkeTN4IaHziGdk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13232)
rGVPuMGhWqD7KVaJdP8yfsPd0CJqN6PqS/FUKCsC4qliAI3o6xj5IuzCs11fC2Fg
0fe3RjJtzbn6smAZaUKBXSj8+XFRYGsLZj8qUeFCVwQO/gWDPLsWayeI03igvAgj
1RSUEOKRsd2qSV/PoMWQi/LpsZDfTCEsznVrtxPJztxailBhadG5KOorvpWBCxa7
QnCwjVruxMDbpiv3mBtEt067vcmwRNLveuIk1XHxzA0827e+EQR9hXD2nTJ+DnmX
2q/0sNwTfci6QqYFNetFrBmvWOtCOkx0YOTHc8b8+zawDASKEQA9eHN25+qhuD++
MoiRptK023WKd7+SyeBOW3XS1xUjrfJwEaJW8tVAXFFlZgt5/07UzcLqp/jxwmIo
JWQkkDP4jq6ey9dHdjxR5qwTuUQEEgeqZ/B7lMYkvj+Bl0fD9p+uSn5PTIemYKS4
V0uzHJj7l7Gxz9o+EuwQhDwE68IsYgnTwY3w5f+kZvRkUhXWpGxJXP82I6JUy9mZ
Uq6M6uEgQ42SBHCpkEx4epV1XgJ1Y5Bp0twKVhOYfacU1FgnephXe3QAySF6tjYt
9+i2efhEJPMC9gaUSfjtYQ3zvk78L4+Kr7faIZESeG58LK96El+gtftCim26oe2l
cesDUwMJeUYszoN8EvFn1BmANE/p3kBkL4jNiI3z8NrlSih+d4x95CEqQtCJimiK
jk7KggLnex0RewuBqqoRxzorw1/cD+f3o/duDP5uBKgT9bp5d0ANi+fuCD/TUD5j
MxgN0IhwpsF/yNnJkvzv4otsQh1A9RWGMp3GVWdVj+ZEiPdlfEQpr3Jfs2FM5vj7
Yd16FL0onVCgfLnfsbzCHCcKAg28CzrKP83bo4CwEMpZS/diMxw6VxGMGRvv/z5s
r4QIfgfhrdA3d4My2iNgXUfyzUfXp3c5ZJGcFfnfCGGpKGAb60JMwwRQjfEgwT7T
8AamUZW9E8K435NaOccnUMSfYA2gDFl3d/8jw8N6Fh/H5kAoFOQsAb+SR0aM18AA
4kMqFbVlUgnCrogJUFpaHO092L2BStK/OtUAj5xRT7w66xwSsSul9pTLDgpaYqug
DLq/m3RAc4bdXS+q6ic00wUWoPskORopL4cISMZslKZhEPT9s2LzCuG8cQXFH7o/
M90aBaAF2GKpZHZvzPnWqHQPLigjLMD+JvKOjygaq2a9eKV3DrsE7JTgonrOQGo1
kSEj54/4W7/o61t0bJnkHFIpImDAKG4P6AtjV152CMxJrdl/Jr3NFE8ASxpC4G63
uivfNFt5ve7QUFI9Jxkq4S+TD6ZNJ5enWVvgjJmGYWl80iQp4dgnB3NwXknG1tPb
6fo3V9GXHqGygPkAk3b/s/vcq++qSBpKYhnHapCXlaHje/tGKs0yaZmmwPZQZ8zG
zHmrxZFTw4L/NIMYNngI7iZMNO+fJiWlowsUIOJJFPeUhsqDxXNnZZH4s0A7ff8u
z+ziZ3N3r3KdW1AaySMyBQZdh43S0XmmuVeCfnnvl7nN4nUfk2AJm3sz9MN9TXBD
DgHvCHc25VkN9XV/p3mtYmWvwxfEg+lXjQ8opISHxDRGw9UH73VbRuUIinr/QcOL
7JSwLzfcI0cjm5BFCFacFl7InaA1zoDhy3YNYggAi1CG3J4VhPfquZTBlkcQPn9M
q7MdT4csIiyC5PV3N7ly+Pg2zQcKYFXOTiQP3lC58x2mN183JSr4nE5CgYh2kaLI
zdiaI+jibapHWZePC0+C0MK1CcO0YZc8YlVtjIeC+zAvNwSaR1zIQ29g0TDrQFHG
vT0JyOMZro84MHCQ51fDTgHm0uelE+F5CT/W+LdZFsMNBlB/ZSa4NK8xpHheHEK6
vs7CAtWiHyzlEHA2ms2SIUvswP/1GK3DWEZo66nXerwrpoBTZn3eEhTILGU0hqoE
rw3BzSvhHtYjCFo/ZbFPdFy3VBRsLAElQHB5ndDtxmir0R/HIow9htjQHzEKwSzE
kGH+NHFnJQEa34I3uvjQsYaxhblmPBb5w7tC5B0Pvv+9EJvUkFA2C0JFqjoouhS7
a2yF2iZNAynI5qC9FNk8r9EL7FHGMgJkwsl34QgggBl8N77xzoCew7CrSB6GMQj9
cerUgUkes23+MznMIR6bC4vU+GyTVDyh/DkVOhkcMRKf/Q9DVMN6EPduxsf2Accj
dZJA5UtusqwZRugjHAqBl/x4ki96BtGYf9PcjRbIscLaYjuldYuYJVkrFoUEb9ZH
HffzlmxWlrqqjblGSP31K413LZovOemwonnJTO5LL4lY/kCfXbrEozWdVxOQGc1T
V0ZHIEDMZLCWSITJMETJFpRYubAwKnY6UdJb5Pcc20mOYwJzwDujh90FN+Awqy89
+mpRRgeYqIhruVFLSG/9Rl+5wA1r8VReHpCX3+7qLGjDDZxS6aeKqVKARmwx6t6t
S3tX3M+PAkqEJ3k2vni4BjAP9ja/P3pAUiWb0H5+Rf0YRUy22g9T24lpr16TYGAo
MKTXkXWkhmOSGFZWkOFCBjB5o8xJVcT8Pe5mQDvIBXqDaoKi8meBYt01aLVJN1PJ
zwSrHQslYt0S3h42UtVPbzP4ne+ESMN/zbAClkPtgrH6jUsv0FXHAjO0SuAkQiXn
fk+1z/q3V1Y0NIjFa/eYwZnRp/lfQodCY6YTurBdLBZ+w8C5Iw2p2mxuBUa3U20Q
i4BcHRtepZ0HpxnbGGbOu7tm0Fu6JB5CCHl9+bzqtaJF7oVOuIwZn/vk0SlfpI6U
/RWH4YUHrk42gFiSEU9dDQ0ui2cIK14WYRVwUUcdnMsWj7yvnx4C+ldMasG6W6FG
WJyIitHc2oFZa/7LnxZTFyYJpcVetAkThelKGXsLjbn8bV//2qrvkG7oT5BPlr75
bP1Dp05ns5nBwLwGytE16gP93jOyo9KL27LScpFxUp9WjiKIgFlGGKmCWGmdFncJ
SyDwoQpjM+GcDXJ8A0zE97m6vNeFFgmJWKdUsegeTmtlDDGgdeklDXni+vfhRpBs
WOmGmLercyIusAbS9jrNbSzQ7opwY3PNb/iSttKuha+7E9GhVfGbrU6UnK6RPiY5
B1bkNgdeWl0Q1q5c2TFXW/pAfuz83LV73mJnrOZip61xXdkBoryKrqDCnhzZNidP
SuOuu4TpHVWDLpf6H33Fnqi5Sv8E2uJ58F/6NSb6uBWN30kyO5GVMgZCRutjon4n
fiD5cjE8/Kb9oFRq92Aw2DlIR7FvxQpeiHsPJ1GV0RcwVg98Qt2F9dtvAcngHLt1
rYguvvjxTqP7ukvnvuriKSuqNccH49gMuSfC/YQ+zVTDnfoPlv/Tons5AZEn5YIC
5hfd0l+RIv4R4hTrTKeR/KMJA4FwY5ASyQEkPLTERh4BWrIPTvby9I27WgnxcNv2
+p8N+VQiMvHtYWhpiHVgxkVRwyjZFFkUmXmT3zc8sQHn5/8WWlFqMH0w+r/3bpS3
bhenT4mprRQuPpK83hs0pUZzBBSAuEGNhRBRRb7NxjjT6mox1nvh5Qcc23HsaGRS
GRTiCSLlZK32mI08OplSX7BP7NpEioq0mydznW4MWgtEsl/cvkyO9xbxTmFZNLoG
CZJVGl945y924qRQxWFrEwwBpP48NoqL3aZ/R2XS/O9+Ijz3hqyUSu0ACVNAUtzo
3mWiAtDtJZ16d2X6BjMnZJyHWfT5qzxAuPKlywTRxIh4EYasA7HJ3b9mKSXV6NVK
wBGHUfr5d1PPjOA0lWoBRrC3Ivs0evrOESgthOQfMfuEjrOJVS3AplSpJWV8rYlO
L/l155gNMi06fy+QS79+awRUpIozDtGzy2fCzSmMdZOJSrwCEfau2ihjsJZ7vNfd
A12xjHflOSTmKysB9FDCx2bFtzrusBfeOXrhxvII68UBRVJUSo3GteQgcgxPTCE1
NFYOTS5mrNQ1y/z7cof6zIvFAkAI86AEQIl3+j7POQE7EEgVrGkWdQhPJT1S/9Rj
Er5+S1S4xnXUe/f4k2cOFSyy9hJF40O/VtZqAAfpKEfuwCDP0Mp6K4W5jpoXJKHA
OU1dtnXhTia9/ZCyVNw7+5XdLZNjqGJZG60YAM9f7TazyOrX3zfUIsSo6XXrP7Op
3KgZvOhVQoBRyj5cNPqA60I6pEXue4cXtr0mDxNf60tGeQUn9JN/EZr+I99o1Gcu
drHIm3TL02UTasEn3KwHFOlmOc3sGWrnmmCX5uzqAi8Ynnp7BHjIxJsI/P2YLqUo
XlG/xHwFk44atxg8b/jMppSQ3CYvce214jYFLQSiE0IPpVwJEc7hsHTuKcUTw7B2
q8jvshShQ8fkQ5iWeo5kZnzEoRO1JtZasEQQGNnv3zPVr06pKMYZyF18jpmY67lI
KaGxJ9isF6nrgao9YVqgWCWULDDuMyi+HZCAF8GEpkWVZe7YrBPCdiTFAbUYruFz
pSfuqMOs9HQdaY/087NR+0DZyAOxPgscRyTyUL+bNsSilDTuEey+h9vhM2+ic9oR
UZFf995Gt4nCGubEtDEaz1aGelXM3xI+hGNtuK7vb4/m8WyLhOpoeXSXRBbQx8ps
zOwN4P/sBj7J07Vz1nnWswlZzOjlXhYJMmzuqBpB/lSb4TDjOAe1iYymM33374Z5
JEpxd1vEBJIB8ffEr+Wo+ebcCuL5uXmu2s3C4ka2D9b60L0+em5vhZgxJVQMS4Rc
wWWdbRAdBAu0Eep+JqFeD0UX+hjvVug/ZJnieZJpn3fthmehqOvAZ628Y1jdFfXc
wM6V4SBUN/o8ws5YAF3Li+xvzJVCab6wOZKZ1fOfockzxZBwptYAvFPKlPhOhlpu
DVUJ1cq+lovbBk49sd50NhfTWVjYQEx8pcbw2A3CQXvy1OtNvm4HKnnz9ZSRupOZ
U4vUOSZzlihFQzrcEVr7k1Fc5V1moRvhGhaUXgNaOWIYFQzep3qInn9039XFq0bU
oS4cTb+YL+we5FUiSI4b5i5/leoOxiV4PRcgHy+SWhuhImdYuQyiQXIFPPQuilhY
yYWCgx36Jr3CDCGJ2xxmfvEtd20kMA5YFdNJ9gMbfSTiNt+8ryofLlG9+zWejwLL
4PeuO5K8mlT7b29qIIScfJfDAEuAuX9QCOyAVAQIB+0Vovf634V4WRGTmrjYXh6Z
7w2vrbqNS/QmNkww+PRmQfBh83JdYc8ZorALv08c17zooSvf/IBE3iCXNgJXZAxX
ZdKe22BzKccoYRJnjj2uWWeIuA1CTrPfcFRaEZPHQW8ircswhFlgqwWVygDwpniO
p9jBpvOmh5sKKmh140aam356LiERFdTU/tZDuswXyG7A4VZMzqPONr1iJI6mq44P
v373OOvn3hoUmiF094ddQO7W+e1uY7RzEMNdC2fZ/cdk6i2sTm2cxjd2GyXAyhgJ
+2C2hsp0eVb0oqvFqdJ8AZo8Nyzpn2gsR6JjynAAiShDJtbzdR21hEzgSg/enrWr
VseJ5To3dhXuakWKEA0ZRE88ydJ8FhAfwBAgaG9mtJ+Kxmt0TfLhzI91EK4eoQCo
xddxFwJ4CzkZkEfDTEn41RiJ93q4jHASmtHidA1SYEDmkP5TzWfTwimIWgcpkb+H
DYorFG6ZVNu2Jp1G0xUEPv8rw8uWt3G4Kg5M7UvjDc1mVvYhFCZs12qLm9dh6fCR
k8RBGi7/LjkL4pCGvik6equAFyX6uwMvae9ouEdTLaXxZfpvenXKiMc4qynM9Jyl
9tpL9CokRb1T8Zomcqv9X8nXNr9viTJuecN8hLvKKKkFJ5tgscJC5iRKbY0L4FQI
y8u7kzaoEoVV3y03ve0CyPOjKGmKYFueNgyk7J4/wezTmN82PpV8avIAafy7rWVF
qqr/JhdrC8yKi1aK8z4qCUuEuBv5ryDlAi6ML8bDYUzEWNcRqVkDxh3GYMA2TyHU
5y5f2e4yL1lo/sM4jySD2gfSwdcKt7pI4hZADgx43EhivKD1EABEdoKIY5XVaavW
QgQ+QsUDwxuycKAICxuEyjbp7RwI7YWWDIKfesIrfI6ZFyOXycxx5rk72lQMcwtN
2SvuAakZTd0d4SddOECJ7qIAGdTB6dT5oGoqFiltJNDVjzezTohgWqwAt0y5JAkV
n5XcCvE7BMpCrRuilBg92fpc2bUgU8dKMEpoB/uZrB7+R1RUncxmV9xcOp+GhtH5
YEmgiuOUezOXsVln/wgtSirTZwY6NoSLrA6zpcJ7qX8fskB8nRq9XA47i7n3P8sp
aCMnVzFwbmGIwRIeJaJp3ddYZtovyZM0HmGIKrxm9G+KREKTtPqCBUirkwDvjaW6
t0Yh3N6pX6Rfwjl5koE37XVbRHNcyJ4ZFA/+GvBB9XUFwUcbSLTdR3FvLtSPOVka
QDpr7n4Jsm8nVpGgr7LLeoSXjcx+VEIhw0asm9Yn0lp57R+h93IOdagUcj+IUDq2
+twTyRdDo0BzTjdnhQUrmIvBecbwDnRViRA/jyD55DWWLSmGtkRKOWTSqrVciLyg
y/HFp16ESreN1zeMbCmftMR/SkAfvaAo05NdClpFm5aogRRVwsNRUyAnvfkundDK
QK/pZkEFyQGISN01Vu/s5JYuxixgUSOG7vTgItJSxydP6rqrW195aQNq8O4/o1v9
85HQuNBtsQoxktTUJdTcYJEpkQylr0y+GWzBK5C4WsxoFFHXhv3/aRy5FQ7VENIn
QpfSsvKUdxbAwcutrK+nM3vtirJlS5IUPlJxN/l7o2puloC4YDpiucT4FfPZ5hFK
TRuPLdpWIQnTNw+kmu1DrZUTFTlF/NYFZ7umVho44Gf0ujGVNwY2uS+9a1pkna9U
mRboe1FiwNsR0vTDAdASYZ1Glebs+RincLALBWbjK3+Fg55QQv0DfIIn6Z0e+MTv
Ay2XWf72YQhf8W9qYR/IqLez6vgux+YQsDBKEZSft8ljG7+LOB7vSrPwFN4wSVpw
4Ph2Lm8HW5BNGNzcXQ+1Q0REMumtFh0u2pdwt/u0A7xio5ttVXHK81Vm9/y53Ob+
k0yknTmuEBeO814Tqk6IuHmlICdsdK7aAI7ktgCNKOOSHDYBgmBZjueCKDMrkrh/
/PMdNnd8nUNGBNSWADwRZqBQY6XeiVBW55T3MMDa54kP7RkFV85rn7Y3VFiC435R
Wgvc0Lr6AbPMZmnNzocRqzX5JGXngkM8RXHRtHTX1akuQBf3q7e19iOmAf7CxIia
FWiqTuMbUVjDuIQ0EgKv5ON6UwrWHEPrHBuYrkxho95O8cr15+ktNzxBBqLDWOyT
nPDzION7klYw4ZZmntE2ZeIBPxjgOlcKkpi+R+3y4zVR83MwfaIpP6rQhTM7R2/T
kAKOi+9AU8/AOpTw8FXKHthGn0LZFAYirDrkiXoB7QHecfmM+ka0QNPrY+bc1PEm
vRfC6m45bXWcBjz/owhjOMIBxFWHjhrnG2uTHhJdmPgXVURWpxd94ErpzQSUOBRd
p2AcIrP2wSZUFdKQfaFQXYUytidyjoSYGL7/2KlDVPzMAdUqXHmWh5X5nSZfIW9I
GXfBSBtLZtI4csGib5CMgN+rMwZZ32ReEs2ty2D7CnZyJVPI2QPlXP/RCY1kU5dw
nKqtydZqLfUS5Zccjv2E6EiBmwdIhle3wq0hxmySwSVe2XZl4IfCd7ejHdS5ZSNX
vZjxfzvr9iheikunwd6sJRLlOfmRD74RQbYuAHYUFDpW0wyeX5wwhrCSD98b2Qbr
p4MF2cI6DtPZ9KB3BYrD1XUNhjKc8wnGXLbJcxDqV2E2PAeIb6dYXIZuB1NCgPnw
3WUAHwOLJXxdiOTZcPFG8p7i8UuY7iO9FuHRm41ITtQR2DxZuCf808oYAXjsF2em
8VE0HotnU9ZwJ4DruLyzY9Zcgh1yx3TlMGlv01Cc+vaQbwLWaTTMrW8J0rYSnhS9
8jFSO3bueAeN/0RPQceRUkORaNbXpblbeqDfF1mEFN9FpUGbuxheZb4z/4uu2J1s
lXbyN5ihSZl+VQPRrHFz3Q95UrCdo+gfGzwx4A6C0RroV49YTzgxHsDIoKUmjeAf
B9dF+rqUA1F/1QK826rwYv9ncH+c4kgsnpSSxwlrfxI7SNgWcV5We5Mfgi/0a4RM
KmVMpDiYKVwDjrs3xlOuTTXM3poC49u9Wk8Fmyni3X2ZE/RXrPjqoCQfGpWjcYok
ayL1bvH/rb7fTIJ5xsLhKodnBBE5SYeXkedlQ2lmJzkDCYZY9p/V81PmW9QECq/G
ujrvjrVHwxaztqh/0E6W+q6KL6QyPludCdDn/8H1LEP5JtGeI4NUPn2FQeSEuzXb
YO9I+QGxDUNDHqEA3sfdaizRN4wYiGde66nBzXtcFnRa/sFhmoDEk5KgiMiJJhn2
nQzhxeWVdOjWmgIF8Zt7c2cBsnTqcvoLPKCcobtF//L0ako+TVyDAE3TWlI7lGPS
d+eSgKpwht1LD9rwVFjomjB3C4FiRQcKFCZ+FSYs9CTY9e70iuoL1fR9NSEBvusb
1ZmGx3+LI3BAkDEFHPYDTVqh/WgpKJcjgaql7ou7BRmfiizQqI4oN28X+Bg2Nc/A
AjmFOVNv4PxJW27T7I/oELMQgo9uj7yObS6zpc11oqZNsy9lYv7wdQve7Qwv5fwb
3Ii6LX4aeuPws4XM8NaayyS6xIV+/EkuIoT7qZXdLtc04xwkklWm0MOZw4k87N7u
0N6S2q+OBh8kTpIDrOe6BFkGNfIviR57JIH2Blx2r6Z4AKXAv4dn9NRmCVYHPEkw
QeVqsuKgDsmiqjt1G3+DcYtX83ccl4ojLeBwpxgS8JeoRf49g5SMVISA+s7OkFUt
lx0rL0CpVLanEwpwEcvr+1L/7xaCoWrNzHmlyQ9BbUBgnzQmbazFsbxaDbnWr92K
ICSRD11yIC069wPpLFZD7r8z5ZXE9v+CWa25qr12sXYIisHPP7+wvTYaQKSl0a8w
dADWgx02EHO1Sxtz2sRXwWpewshV4YPpSLJVe9EGN0UWFZZ5XNfpa2/L9tpL+TC6
WB/aKm8GyILpr3qSgvaFbY2eJTsbq3/QKF5Hz4XWF/5h4R5nmj7oU+AsoY4gXbg7
N9M7RpdD3J0ODZL+8i7AAJjY0v5mT/ky3U3pP34Lj7InevcsVcN0T/0Hdpq+57aX
gfBXuBEZnmcyGElsaL8y1lN8MCqJ3Re0e0zjpqo+m0j1F7Iw40b5Dxs8qFsx5JxW
xPLMpjtal2i3fJa8A3ervvGgHdp8NcM/5eFsH+uPj2eBf71Td02BOf0DJUOxGJRr
ClScL467+sKLqjMljmwiRvxvLlPbs8vQzWJiHeat6u3DcBjWsfj/qjyujJ/xygz+
XtsQQI7bKNyt77Q3KZvFQgBN6kA87txpbbpFtf5sPvC890hRjM2apg1lp3tWOqUt
5a325pLwxgVboD69o5wSggJey+bSoFzc3dsa0gBywhPf4Y8sKRULGt/uDDUMhITE
j5caY5ZGnzgBpGavU4n466bEM7++izMriQG6euM5UXkQTvvACYXBuurMGd9Woa9h
PPBk3rAvMN2rfwDCiYV9lS5FaTKs6ZIo/JAdr69kuBW0vJtK/+rl5iO7cRhqVH90
v5YSGQQRThOzBxTJ8svfBrMuHIqC7X6pP2vwU8v2I6R7X3/0pscSIokQQ19XTkIz
Kz/BZpybeWFag0vQ9VSX9pM2kn1wqN7sUzdZFc0yzFLs52pgEba431wqWxKIqGHP
azI2eyB6h93mjD552EvNwWdAJUGW9Mg8Z8YpJiZRwos4Zcb8DOCG4yzQ8RxYtC+O
JcdbYBIzp12Jm5MIxgx4w7988NMz+Jyxn3NeoqShkwUqBgNUSQxJvfGrl6cMqNBi
+xuu+MymTlt1UylrNGiRq+knGO4P3U+UsPEAhqmvKaaSaxqAk36rc6mAQQwjZy/t
ICt5vbNOBZFVv07EUvo+0PArH+XHZY2xiDJHXF+2lhw+DUshtJR5MZHK+zJjMGRR
1Og8nVJsR+R0SfmFKcB57FbwrHuqqrxrybaS9+Eua93rY4L9NGKyyNZYzG0kAYXu
9n9dBWqpqektldmjuY0ohQnSfaLPhDFwLkfQ6wU5XhGIX4sTv1EVdijIklOQltr7
eogaIpbylJrz59Sg8GevQionZEgm0SbecMV/mm/ZgkejX3gCJWmmx3aZ7JCoTJL+
nfRvieZeFQCcCT4o0p4gYGh709PXt6PfGF2KQZHXHspqG8kSCWKoYezMCYQFyMsq
XdK0UywvErE0Pyhb3i/eoFG34J4MOni4Bhm9iVj/Yjl5zEwrEmdojsoGBpwNEj1q
eb8ABpFOAp0wZV65+nNPKPfpCaKT/C2J88jEsXuOqU+NHwMddIHvieeQ52RPdgL7
MyYXVsYmrQbpNtv9lQ9MLtchAyJlFZVse5ZvMfWg2IbIha33SzlRyEevY60fLLnO
98HVsD4KIUvcnBmqW9vn947Od76Mei/8CWUnPYwQINHCCjkn+l/ybpu8/cc16IKl
wLeYu5JfsrXgGIkRpc53/HFBboYdyZf4GjqgiVKnAH0w3CDURiVuGgYoIUnmf/9p
8Gzsc08qw2+bSoG8tVJIvlL+7BALmcRgzFqXjqyz4JkV12QJa9ehvDj3/yB0CagE
ghuThADXIw13KkifBCUMZJHxxQBb+ylPFyWUOPr8JlpV6BBwvCH7dpQiIGggTx+x
F8Akbp9c6/x38E++lwXHJEnjU65kVZ+9cU55O02a2/UIGTQ9a8WKb2NyxT9oYV9A
newRBtCWl+NJfQknjg3GIyb2/hhczVKmdF5xudz8uFkZBRpSLOQAcDd+h1l8dPMM
vq1kwyPuzSnZFP2xeFKIeyJhWzyEEUxgbK+P5/HIHRZGeplsC9HKSg5+tPF80/my
K7CHELCSzoozy6faz+Vw6lSOdU5AQz2rINx0WFU3mPtbbQ+YwOvMnj9lOttmIaPE
1IvhuKCdJ8H9zNmqSMAxhi31wsJUTCSffGplFy3Lzj838ofA+cT8JBANswkZdZaE
6yzkoosMvxoCZnqNxC/6ycDyJYXLGxoLU+rqBxs+s/B4HqOXS5gZi97eL6ODaTQH
5iAYmNc18VcIscvdEgV+oY7Sg4jgRfOLxMiedvGfNGLz/gLNsYencnCylGTpZ034
nHVih78981C/Mn1EhzpEqcw0s8xFOI5dkdYJP0Dh4EqlUd3zatuNyeqqJSPplIDX
t7IGvqomotrc5VEdhK5Oh6Cqpk/v4SibrPVkd05qiZVBVo2I2phemaBJhect+yxs
hNGCyqDgFzByGfSVBWKs1JUAIkz/pg0iBiG+aYwjyyHltGzALMt6q1pBZKKSmfa7
MGKKCBVBt1Clohgne2Y45zUqB+N5J0/s1dmEGAzjF+zzMj+kjpL6yCOY2nL6kx67
6/FoGIMNMA3lLv0JsL6dnJ7p1XluOdvjkQXKhP0O96Ett5aVRNnvWPFKhbASg9F0
cuBn5kjfA0kc+VIEc6OCEOWsh+pWm9enA8t6qkO7JnHAFOOvDTZqntgTLtPSOgDa
VK5cq13h9ewXlbdiim9aaZYLzKlcF+z9pNO9jbHG6Ql7DOZUyZiPMwfjqrohtWMp
b8yS9q7INkNXcnL5Ej++Nw8oMgsavA+IT6VXJnqE84h0lSzHYfYl2gBVNAuVgYo0
6l6jxeCbRT6ZDTWuNv7xpm9XHfY0lBFPoNCKsYtUGsG9joalsz7halH/EcyOeabF
sm54T+QwA3FLCBxcQCydhFXY4gNo0UjCjOGJLnHzmSXSLZINPQYM5S1JtILuu4dv
PzU6Hu6cROXxauFpXGskPhYfYbH7r9h/J1C1iyLM+/AP+l6kdN+g6H74TSLJosPv
s6nbfyxPVcQ3juDHtC1SP08wJLf7ktmBR2XPzkniGlzLbu7eGFYEnUW4nBK9oDeW
4BVZnwRIXyBYdgWQTpHB9NNOtU3pub/YLmml3BWU0AajjUPoJ7RkgPLc3Jvw90JH
30hiSoP9TUQbdgOzCnOb8AmB4P9JyWFBYAGBtcKPwQgFSF9LLsyJ8kQ1/XbBpz54
SLnP+5dshRuuSu0eEI/gXyhFeCBmyoLrNbLkr7hNYpEeTFNrOprODLjaBOwbEDjQ
JmyFqgq8o3YQHPQECm0lB8YMVGK6xzOPNKBkvqy/hn7R97GAbgpIZP2KtrYHMAiY
pZEfmXuCmFnEzgW3l1CRJzqpTqIVfMDxxDKVO5QAWOsEfOiCSCFEYU+Tv5FSKr2Z
QzDfErdX8razAWdlJ/FUQ0lTxNUEBtSAUE4Zfy72a8lXFXNFJu+q+O2Qa34qSmLe
VadLWizxpqJqOKtttuHkY7TkGpKMaSqErLkcYILyDalS466orjS5BcnYVsuCUfwK
vsMXsVEuhjW3lpQB31UzJrxkDLAgteM01OVOzlIkZN/arRFe0fsJUFGvcPMDlqKn
QW4PTeYgOpZG8TZhg/Hi+1gwl+wxauI+Wr1pFo65AScVmEef+eQIAPwufqLgM3WH
6cMArkWQwvC/gZf+aUWvzohyKUV44rVLyfzXlWaMU11AyO2M/PxfVGKJbNzbHE13
yqOrfRTdXxiGnQDTwkYo6sz3jpKzwl3W5xrgl3Ou5aQ6jbYISPNJ7Rwbu92Fsitv
tYX10mPB0po1QhxGPc3Gkj6aW+X5KhwHWMdW20C63EsM2mbxCKqQNyyPY8uoloua
AMh9jif9q5cS3MHsrNw+QVM97RYbH37QdsxVq+s/q+eE8M8IJsbxve0yLy+Im2C5
R2e4BDB0c9DSjOCBDa2RH44SrXJws+5ny79BrvGes8JlnFaMEHCQ67xU+r1L6XZm
in9JYzkHEupiZieZ8y+dAnwMMVdLhV8VKmbZQWSovPY9xBWwDUZx/wRKbjHUrZ33
YI23vbhITIi+6OGhHrRPl8BhjQRDUMp0Jywe/8PsZSvAAbRCIGQraeKqVfFMPSme
lzlE8v1KvXhr95FhKdrpf9BwQ4cjUB2o6ZxbBLqXnnkr0G2BwULzp1inK3qLgD83
aP2H0D0QeL9WJVr1UCC1y9aZyyge+yNHc8WQEw4GrHMyJ7qgXrbJQAV14SwKv8Y5
z5vufGvyA357wzK3aDFEDzGjjUp4SFfBTASimGvEE+hNwUsgjYBQj9XQyet4j47i
pkNd278L1b7Z+0LjTEVfiTEo2C2Lv36drVPNvidls0EOi/jny0tu71IC6mLoKwqL
LIN5aPwqt77fjxaD4rIXqyzegc5lsC56PT5LWv9lVPYJTl3wBvMK/VNjAmujyNcx
luLtcOVrEZlIXk0IZHov49FpfPCiuNTdoR7n1rA+De0u3IKAjLCCC7ruzOHSNjPm
Ekr9enXwjXKJq4uWR+UnzRcf7Ki2BJiY6/1So9KnsiWtKBoQZz5rl67UyOvgbc3I
GGTHiQvq64z4Fosge/PsylcRCN1pVMSySCJ8TcwPnI+f6MKmvKhynpoSNFvMiUhH
ftbrozb9CFNgcw0RG8AH2eQmOYbFhXcYgD9zU34H3Q5WDNJg7L/Ok+OSg7p4Gqrd
n7BaZUGpaxqORXN2gZKYuKqswCCtlpy0Qn9rjsSF8dzC9QVpE0AR5PmegVCiiM5Z
ToRkPVjd0Jrm6L4XAthnUUNW5Jk3Cn7tYH133Ije5YUUB97wM0Qw56+5Npzxo8fc
cGwrMK77Jc92B483AE97JfoZzyUyRyoMra9HBT4YfcFAOraEsG9a2f4S4fjVTBcB
31zrtsO/O88OZum1/X8p5bpcLxGYRAukFlbuytWMLnlVCj3UDJ+VYnvU1zgxti4D
CHyACGqu2VGowH0oFQvIEJRLoTYQgpNR7BJhdi/RUF7F2249PcxM0xzkSaHNUalr
nnnG3V5/ksb4Gi17qVf6skveLHIlf89KCYNQnuXbF2dslXIXALN8pQoy/x3Q5Ljw
8E+E39p4RW7x+nV5P9aDrwzzDOAT3KAxXflX6A56Jt/PcA3axHOR177jrzHDVdGI
3ocx16/nvR1dA+Sf5QP8hAERnHiDz3dd99MfGCtbxb4vzVbubChcB3D0ohSMYl/a
skkw+tH3PQ2FdHQdhIYWIH6vY6dlAZYFL2d1rlVVo+7AuSZzCwuhd/1IXREyyjIA
iSE39YfXloPyZEfS304uV3MfdYfYebkSeUY5iR5fowSen2Rj96Hqfz4m6d1sVgeS
fC4ZoVtzidAaG3BZ2FhmT9QZ1Kco/ILv62kzehDDQfPGrQ51+4MZUruRFaz9b0t/
se/Xdkp5c5L2YCHu7eYF/pmNyghuTM8F422NfdidxMjP7In3oerejYJa6BXmXVHv
t98H2IDzb816uUyEtXlSSzRbgnuW2fR3ioPAHeWUDe3J6+o2LJx3xSE6C9+cGq+1
T6UWYZx0IWo3TM/iaqody+x0nu8ewCVTr6o95MMlNrQbbW1WDonUK3Gy+7TF6rOA
6t+SnZnjVslLzJZVEihGA9fvw4VZJNgFhXrfKBaYRrHELSUo5Yf7l90yFE8q/ki6
pIBrfsL7gpJtT9ubwNRYyHxaiqCorFLH+C4bQqhkStbjXycCGzjkPecOwjgN6ItY
8m1w3GUnqAXEr3azRHUBV3s4q6qmP60QXrXlzJ4KwZlAzd6D5oVaqiRjfr5e1OTL
u+k1vH//oVLh/Va2fFU2OsDN1GbFt6mADFKkeCXEfr5oaFwCI3rBswuyzfDIDzcw
qO0WZcV/fYvMKNlRxewjHbeHSWNkEKdCiIWHzwnsHtyjwkl78IeIcwzoJv2I0smD
dfx6TLFrRbikm2M6In7/L+MwoR0qpKD8Zi6MIuIJg92tbSS49BC269p+pwcqkl6h
vyoPdV7Az0SZYGIZ463bUV3CtuG2dUvUjlev7NEG/5myQLd34fuCA4gvUqPAFaOs
kCsb7yXRlbcdINE+VkSTA0dNM92tJzp7bKE2ksO2ZS44bUgzjoMGNG/bDDCSAODh
jf1VECppO6RVaoYYQbm+0ZTfnoVhOCHNU6bA1/OQ7jUlKzPrP2xI6ThgYHKvmSOA
nt99UosRGXsz6vCoKJDhLQoNaK9dW3Et6o8liB/4AQAYmHFc0Yj6wrfm0tQ8ZXxC
wDFYIlpJNwEJWc5luFZHK0z/HGSoX+Y/Yhzzf72go0+9eKtKv460nclq9AVJqXLe
N2Ly4bF4CojWBKk57SaAmAD6/EhQJKHq7RasmgA/n/43ryDOoEfyKN5KyZanAnXb
dpLR+rjNY9cWz773xiii9B6qyti47P0YwICS22ja9JcuQoX/ijQkjNHNAlK5Ew+6
ZpPPerP9D6Mg0ZQ/gMEJgDus9v/o34gHbn+j63XNffvl5Sj/dP/t1fsHHaS2qLv+
Qn3wOsH2RcxIZG+eOicuu+FuDKJTvnumPgmyzQxlwZuvRZnfIaahaV1WMtfZLGBa
FajtYSFDooPAPynW9wpJ3afkg+EypAt6wo+1kPGRp21YEfsLsqam85NBuXXFsB6s
RsBA9wu+gMf66ex+mJ8TijD2V0JrCP5xx4VqCrHsB1CCbr2AqyRFEmH14HZGapx+
zAnvHmVXUxa0EfBAJgH7olnHsGrJDe8iX3GWYGwSaJ5gfdQsCAhXcON9LL3Ia706
u/KuyjMQMB6u5sfuRTXTyWi0qwS182lFphMQ7lRi7yYMIh2QuvKzXjNAToDzAcwh
2onhWy/e/03EZoOY7UZ3vqSsqiBBrb/zPnujxPmucxWeCHgRiYNkbzhnHJSKF768
7O9UCggbgXIXmtqZXsyKr31/NQ9ttkRB2+UlI961LNusaAp06UKVo5fzij4WrMC4
EssiqO6bOz9Ip6Wvzkri8qzeDJTzL6jMyhQ0Iz3LxkqPwd2FjLXg1UP5a0dddwXm
4oR7XpGwbnGCtUiLcPpnMTrTKvguNOW07Wi2+Fb2DQIFR8dTHWNgkC7ykWmFIguQ
KszVgdFjtonwrIo9GyeMsk2TRE8VMFAlTraPQxH/8leNDlfL8cjac+nIT3JSO7E3
QelMe84X7hh/PHGAoh4fj9gIcgfnIDtNsJYqyHC2Jv4TOqtugC7R2YCsBs7t0rg7
F+fqtQMde/53AvSMJ7Z0rdij54GmLb2uEJbMjku52KR49CM82VhEI99V14A5MRsL
k0wXfsVK//zV/SNjPj21l4OyMHP1ltFt0tVkHlxuY9wIp1o7gZgJkZkISWNmqZ0I
Wo+iBybR7iqeazq8FFPhhC7Etqae8AcVxLE27/QifYh7AUCZmYDLsMurTXzgZK6a
xTH0OreOb5HNFvT7ecE3L9puR9rvaxYJ9z3peZZRoWvxPC0rNzritgw/vvrypM33
JCJsMkjnOgBGo/UUmDUrdER6+vN5XanPCYokYvJhJU3qjSznCe4vf7yiV29P8XnN
+f2qY4agatK/EEXfL51gXo9rh2pfApxdOqCwBqJMKIljd8DJVGtuRGaaysJjZA14
iaxlMR03OzR2ZXYHA/ujrclvtP9/AmKWE0NZb7IVox6UuPVpuNPZ2hK+Qqh5uF80
YbzZEd3k45ZOLTq4RBT/qg7HF/i+YnzQDWUMb1fmoZ4lCu+3wzfJm2ECsPZg/SL7
Gko243xzG28beus3SYSBNPt17kPnWWCeT84kmRGqO3I8c/Z37UrvawevkhrPWZcx
w5svooXC9bb5EhJmdQ7DQyirQmvV+RITG0h/Xk20L8g2MU1H+tsxYzeUk6jlyBrh
coQY+PXmbFJ2iYAateRx64DsGl/sKYFI3Zwc1hmeI+Ds0moF4zgmguSm/8R4b66k
CjXmjt3JtrqeUZo9/DX7o8SbVuD4OSOVe+0isHF3vqdogwjxjlTjSoX7qkp1zWAV
Z804OLTzP6DkkH1YRIB1mq3DDUKftrqlrhYp1GT9fF0KopjwUGhWQtl5rdF0BQSp
0Qb5BZjCEcEiHBVz5HLk498Ox9w4sp0e3V/oz2MWeZMW15OYVIyd8T6lndrW0ZMk
Ocv5O4mPp7o3kOh9G21HWono/VteociCTrusge3gZm2Z5x4pMr3Ds4MSaWcUVeWO
Hy2h8ozeyQxFA8Vz/K+Qkwe2fXyPX0lNpW7dSRvTSUEllKTtg1lH0J3IDOvq5Sj8
jFaHbCkgityvpcScbgS23/bNCBPg3QAkGVf6bVIZYj9omYG+RCjV5L8HGWNGfcot
2TRqyE4u23TZ9FZToRnBqMhZsy1sVxS811VgL0ZbRigpR5fdxSnJiL0MftCotmmm
YfhKLzquxJKGN/m1cvHjhyenAUZpCFnISfrC2LpCgzedr94bHum5URKle7ost8do
kF9CBwML38jURTZ1xYiQjH+OzTS6YZz30qBTckYRKf4cSyYXDQAJwQerK2ijBKnH
9FzQGzm5zLcqOyL6UB8TeDP3BSHKxCijJ0pFWJraLvCFeEDNHuhJHd27xG/8tFDz
IOEcpxd1HJ/2e1QugA+0jjJCkeG3rksS6LaWgOtSpcSmeaijXEIlsxR22kq6f1LA
h6f15k6tFET6MZXqIoJrG1cwYlxgdmzANcNlRMyOIyB4e+JHWvofT0NrcP+6dKxW
Spg41etfvH8Bigi8vRLmezATcATT8gluf+zbODeQFiZAoAN0LMumx2TGpmZ8owUS
3jytApf9K1U3MNwIDGzwiDH2+kVEFzQqTGUJXmSyuspNYVpfETi9AJ9UQJ7DDK2v
MfQhg+1PsmN4wwwFIr9bqQLz7LPdj/4qBwWKODizCxFdBdxQQpWf9vSInraK1ndh
I4l2gFCxGEDYrlbwzxjyaekMSyXtS0Tsjz5BoWspyC8=
`pragma protect end_protected
