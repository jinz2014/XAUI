// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kTzd6Fx+u2toD/BFghn9yD2HKKepTvlF5K+GBGRhLm+N4K/dpVigoYllPUgI45Vy
llfqkP6UvrWUL6E9tX284D6LzTdzDemQrzFQspu7xgHB9z522Y+nGqbxPPuX87qF
a36MuG2YjaHpnXqixhhhLCrI9DVj5JHQ/9hd7yE3cAQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
F/f2PrqOwwz8dXUfhbHcgGpBZ+f8wuV/uoz7Ov39CpPKdEVfC+1lZbASsmSoJZQt
kiCsjy4Dxr/5LOi+GKM/50KzyM2i3V+wz+dISxnuYhqaSanRk1pS5mnrZZxRUeoy
UDaNbXUSOFhFQH990i0vAfsQa3Ya/QK6UJPugtODI++ke3G/dkDHrwE+tXnby//T
txprXYn4GwXnwEcqqbuhiBZGpGXt4j6VVCudv3tWlXjdMH4wUXTae3T0VNNpH01f
1fkJCPligLK5WTMahAyUwHQ61Ox+PSxoit6pN6B7guMW6g03cGAovZim6ZnuxJfp
M0KX7TsagKs8g10yeZ5DBCgt5E/l+Oh3BNUMLI/3jYSXNyc2lRHk0S0AHbG1iQgo
qnv48WFTfWaixT7JbxK0n7iBVrLe4LrwDsG3LusfbUXp9RedCyNHWlkgRTHMcz/z
aCP/3vdQdRbjtV/UcjcooOSfoO8zp7SYEb8U1lUCuYWz7cuVT5w0YEvdJlROGqKM
CLSkKrsDGqRAEoQEZ3Odmi8q61jqsBr9StdGlUIfHhjPKNpq8sszGMwTfDQtYfph
H7MMxbkygpBtfy1Wpcqt3R0ylSvGO00L20WzFMdK7X8ieENVyjqRFJzxcky+1bmR
wbuxcdHznH24X03XZivh4Xa/WEcyrIUxjbBpfX5U7qjymVG/+zMRT8NsbdY+VK0n
23hiehTK/ho5ZlLPa3RdJ7BB+ikJUyndJM5ZEe5vcaDqOALrYfwqdhosdVzbUsFa
rP84u2wk1TcGr9qdY7OtlkfUG8T3R/FMI51Fi15Agux2y87ORjqhnyuza6vVcv1q
pyOyf87FkgKeTmAt1JVPrPYWQhDLIqR2G2OMG9jrfA0BdidHaxNvwrfR5DEcHiMK
CDboDcKsH3gD/7SXWl37AwOvZUWfCGf4An3TzIk0uUABMDVceybULO9aqIh7cDDE
bue5UkPmeE9jlOJSTRp3NvTkrqdF4mHFOAFUYfQxTrLphzswxpu0PG6eorik6d4U
x0m10BZTVQ7iyNAewu6G2N+1RHjujSkCLHkhpXxbxc7eFCfdl140pSfooMy6lkQP
txG1dYRceAshTPHV6GNxbq5LE7Ko8fHGJTZddwuIvzGuad/TKFyBu9SBlhowBahc
eRrdfV70fCaqtZGe/arAO3B/lXO9OYprfb1/mdAqvuNEPP8V+ePJle+xqL0NbCm2
sebIdhnoP0MhOb6DfgeDSUycJGYLaf6gAtS5se3uQkRE8QIgJI4Q9cEtrvPPUgDO
7BXQws6R9pDaVXaWcOZcaKzoCu5otkXKJowV3sHu9ZquhoNu22W53v85dmgbatLw
A/KfODb2mXVu/NF6TuEx/dw9K7Ucl884llGdcFNI7eySoxhPCopyDESeknqmmSft
Ka66qFtUmkswA3J78r/kvXcUE+fX7tqNH/LQqiYpD0fyn4TwIXgQ0pAe78M9V0/E
zwwMHYb4l2BMHCv+YRNbBzZjWTRnRE/HPQZo3cPB24Ey1Tl/nzotcVD2ZAkyitRI
BF8FWPY7ZEsycsKQzCGyYVJHCYTqr1w42f4EirYo6PFXoZu9s0Glm7ESMnoE5BWe
6ujlTl3SqOLug7/n1+Q4KAlstjJ6w1xxItaMCOM+IVxx+6WJzRA3J8tkwMPykAlw
AqvpIx32L2r5BzE6FVWyMLSnH/m374qAOJxIEvS9EhH0i8XSyKIswqaOjbenW4vV
eKV1qD9yqwYYaFG9xwu8f/Bosh4aXGtYeMQ93+7nSesCTqBxuA05Gmv16XsE81Ez
1PJ3sq56bCVn8GF00/iEUdS9dRxySc26GadOb6foLqKNemiS6Fjf38ak+IqU0quF
6vfBNNKOVsCxImFJ4qLc0eo/GxLpDuxmZcYD4ELXg5jcNV4/bzYl8cCqEZ1ePGK6
8lfMYSYKXLNx7SBMB5+zfI+cNSnmgsOhOalJvWgoFW7sBGBxmbyHBFp53IrQSuP1
BcVJqGZqOsoR6WVzIhD+9S1otUFXByziB3r4vV8owqRPdTvJ0xsNKIHjozgAgSzo
FsPIuhludm0rf5CQYz8hmakm9EYG9fj04IDG2Tg51wg7+Wblg3lqgUoMa2pEUML7
SiHj+HEeqNCHClYdUQ7rnimOhnrWExRCovaGzxU2yAJOOqJCNxca6gvQ1pBxCEM/
MmCHF0alHGIYXRwsHIVmCTsRkKUQpOOaNVu3nFk1yeIGN8CJGyA/OS6DHRd3tW46
OOUjrVx6/w3em1dQsWK3wYDX5t2R0dtVWtgrh0sFuprCWZOPCpHWOozvtkkxkAih
acygVIO4OArfGSN4tX1AKQHH3CLKd/4yxkuN5fEPmMVRlGXRCaJCUp+u6PI200+W
TLc97m7DOEyWfWEEWUtGEzB++VgHWsfCN+zKX/D6z91WCudH+MK00iBZyKMarnt+
OIT0YUSdSNU1nku8tAosUmEoSBso/wKRfru/eRZ3W25JH5Iu9xat1YgR9LlRgzkf
1W+rj8+ZkJUR9QF/Ma+wncLa7MuS8i7XgPJRDDoHmT0w3S9E6sZiECoNy5mkD0pA
WuaYDNzriXx4tjStpbkjYY5YQ5Iu61ZpVxhZXMgDvL3wzu7G+kSR+aq/gs0bzvxL
f5Hl6e9MuUUDFDiTJ0C1o8ayILqODNA8lNpwaTmWs6djKz3E6GsyRq5ucN20y9UQ
tMDd8EjPV+vVSkGU2awlJxyxNgMblvaSMgbO6X4n0Zh5N7739IypCaXgWi3chxZB
1Hxy+s4RPrlf8Up+spgM1HR0glTaEtgLsc6GY1yodx9Av6arZslsu6mZvnaNaIDm
Rf/6MWiIRd9sD2PvZCVYPL2rITcjVfDE9ee55k0PXfxr941h0H3YyABlwSpgJ1cf
PQxd56uJ/h4J8zkCECCeZpc+NpzgfMvZRp6Na8xyMhXYPJ5qrVbBWqrABa/l0cvX
2ZWxTGA1I3tDltwY5Z9a7Uhu+aXw20AZpE2oypHXzw1yj2mBNZQEa59nSuJ9s/hx
BTGxSW0p6c+Ld0ZNAy6BSrckb9NjqraB9L1wkBIIwk/YOULwx6fgGkytWpD0Md7e
PMif2kfPrWHLpgSzetyWCLnkJIz/oCql6lVDI8nhtZGbZpewpknYJjoRsDLaKw/4
8RCydY7C0oNxiR8lN149agKNkjxqsBpYbTUpincq9ogS1TyP+D2JT9j6TskMD9tc
K0mapqfifk3wzLFKwAORH5N7Apg6dMqwytLdDnfoWQJR+MWc3LW5ssU1dWtKVmmJ
G9z45wEn/lxP4hlMKyKut+3mZSZsZZh1KQ8I2c4LvTI4Iq8D5AoegyC5+ns4QIWs
iyBF7+SYlIAEopz2CPCk5B+R8VZFpRj6JLN934IexfKjNnxqnfUE+GNMXVwfWjpb
lDqmLZ0SRkBBkG6qXlZRnifJfS8hz5oLG6QDVP2CzAoE+i+8LzMUJ8NXQQuFgBfP
0qndrmgmgzVuTcTiHpAGMpjRvXKveZ/ouzHLp5Nadh1m7OrArFQYFTSlxr1vmyQn
ELNarJf5PKNnGmMmcTqAhnDs1g3RUrF54r0hOMFXAH2nbt0KYBnhAOeWjRQJi1Js
07RNh2c1Hmt1YQzpeRIZthzui057DmGICL5LLwPTXB2jWeEwBUDHjccqdVDvX/ug
mT4W8C8n6j7URMD/SEa/cNs9hDiYCQZD/GUhMMx8qHrW8lLyuEkakWtqoP5k6Nv9
dZ6vRqY75MiVTDnVJ1ZX8XSRN7cqGGmZLQK8Ja1idYas4HwCCh/4Vq7euU7054kZ
RQiKwFaY729lyk+piVNQkxujYBJE784EV2HlaJ7JSKUXfgZlen4J8ubradq5b+7h
5jyTKROKNbtUOcrZkjffzLZhu2e3UeBPX1BEyM06Fk2N7Ynxahnjua500wW8KO20
RE3C3rXS81Q6Nd4CCQ/CxytduNpoJ7tBN0ckEKvkr9K1jeEvSLvl65GK71bSY2M4
xGx3l1+9R0dmeobl2vn4H+v/ubb9lb0jL//heDpyKLHCPegsJ2h/hxg0b/hwgkGu
N54HWdtG8Ngf8MIAH5MMydxGRgsmMTLlJbFv3KMIrIt/cXNwpe6tkHBiMe82OFak
d6h/6P/vP0Ub3+jlU/9RXCaO7AczA3YESDQjNQBxodKpXHeaGuSA7EY5m3vvxuvD
lH+52ZJ3pqU0ozO7cNC179e0YdgSjbEDEVgvvWyMRgyJKH0BFSJdZgxwsiQxH4jR
Nl4PT7MKxdDVZzUTzg+zRW7vBNUKtIMkZDYjCPdn/G+Cpa+k+zbnIUf15FTXWNPy
9GSSmItmb2zGf4gvNU0FxLPmhyX3hxy8/3G4JoUVuQbbpmG/+9O0r4eLgxQlnEB9
LNl1IWmYgKxgPMCL2E3SJdYKXhrrTEy3LNvvTgzPUJ0NE4evRn/LYTjhP9PrNwYD
2keRDHb3TYwr6CaCDQ4t4X9RNpnDJuXTFk5Zkk8C3Y49brOMRg3IaT6o8JsLuZFG
9/tg0k/JddiYmqQhN60s2fYwOiRfDtPtSTZNntmGOp4gtNsEY4lcSdqwS54HGl5J
wDKeijDEd/7JCMePBoFqfPUxq1BkWVQajwrZHPg2Aoig0zst3PTauHPy80X8PEWm
EIAcGlxU+yCMknWlN+3aZH0xKEwk2eAuM+UHPkHP7iFizmz+nn7XwloB8QJgWvBP
jzBGo0Ccf4ObNqH7Ym1/m5CzhS4J9Ptlu0dVqZ1e8AtxhGqKmh47tud+qTPsiPSv
iIE6dT4rqwH0Lk2cZ9buJKmg/UEVYi4K1noZhkNjzzyEP/FmX3SahygtDczZ50lC
py6q1kQkbZePX+U7aPyfG6iaZoo1KknzyUZY90b0HXJ4M+hQkn/jhiiJIt3/fnm/
7P3uCXHTjlHkisZvZsS0KrbL7h4HZTcqGiotswjcdocssrgh0Brbf/YHYxbGIIDE
nGV0sTkCBaaKpUlUIpgTDPRufq6/2Zzljha/KP/UUAqR0AmDRxCZak05hgVrWysz
+FpnLUEo4PZKNrvgGPdE44anOWGEWweCBc+J+R+GhRyc5tq5xFJjhSBiY6OK8mhs
eiF8CZXKMuZ0O+OelA7/hXIVOVD8nIsF56dGkX6iCrdzMjxjVq97m9xIPt6tFUKc
AOljYE4GmWBUOvDQeG+Sa3LmUhn1/vTs3AEsfO8nl94HVTj3mlrOwGuPWtH7E5t3
r6ZrwAXj4xVpPVviFk35uEW9yFdkbGEjwdc+SdwjT/VQ3fImSmkSFY7/BdVd1Iaf
kp615Gqz5ntp8fprO6QUsPCPcosQfvo3pBRXYw5THK9V0vNI4zsHUEnmFpF7UMku
/bhOFl6dzhw3NJXz+hazvdsQGX+pSMX8RY7/NQCUzvvzqkYBwq7VZ1UswT3GI0cY
eITVsCYjWPZ/6lIC7lmUssRhkVozQEd4CJ+9GKyN4ULaj+o45jTn4Pdye0dD2s60
rtG2HA2kaQZm/Z/uZWp5xfs+FuXzxF8JigYxy9r01jaDrsAC6JfARqqXMTyBOrIK
C7+s1m8DnmZIPiMF0vzgxI2AtJr+EyJUaA2zxL8oyD47OEULnfbDShYcm2HraCHv
/UGDPe6CS3la25tesOEcwzYJmMcOp5z7FboPn7wg/Y4+ndLxf5CXQbreEJY/xDLJ
syvdgt5yuFXsBhj7LU0paXSlDBi6pqloclp0V3ip+zZDs6kokT3lJebNA9OpCUy5
bjI6bm9h439SMk6x+kwEVN2TojYuPj7xvkOjTAC6yz6iKArB0t9Vb58ePcQ3Qayj
0fxdpVs1YxCDVmokWIzl1yu0ZCxsS7spcxhia33TFzdV6L+JZwAHqYG/GVAtmn3b
lXuJ/5rEPNymuA3w68ayIdK7Tcv6AwhyFzdy1VFdWYpt6mYt039IoDijCMGP2rWO
p4XmS6rCNxCXhMC/KAXtTZxBqov7r6iY+Iuhne40JecH+AN27434DoMiE7nAn3q9
TYyVCdZ8HANSw29YwfKC6axc4A6dExBqbNIbwAlmJBmg76qns6FL83IzuUKRQwOr
X2DooUC2xwJawwwgRh0ILMcgs5cAtQlk/HTk2prA4l/Sk6ZSwmP2yMdOhF792Nex
Y9T8/OIiDVC0hgGJP8qm+CMqC87KoDcpEVZPRbfFxInTTmGlMZi3KbK3X8m9i3Ex
o5ukT6JmAnoBv+PPg8uUKRwPKoQqt6Nb3JzTQxEIT+l55zK4X8Kw4Kh/EI8fEdHK
UqJDPO1GYeCaqRin7ltf83HqUSkQs/CikihQ+KZUm8H/YWtbNBAutbHPE1Aqk369
Ean2PKE9Mksi59rr0KVCgVBrySNlJo/wm1ICj6lfsAniHxLfRgBksbcnFxTv+Uet
yvwPW/5eLnd/NvkHDPYupCO/vKIcZ0ejTFDbH2Nw5lOfsr4fIOCE6Spz3Dj6+e4m
iQGt6VVS5ETV9IQ2i5b0uYsW1Hmc0g7TdQqM7rpCOUz9MOpTGv0/yGH6287E76I+
7FfiFDN4nuiGW4cW5m9IRAuI7GmEE0nDHpbEsxfBAkLw33xq/EqD3Tz7fcY214Y6
Vr6gSihBQvjA0vLiDyXxFZOoEnVQq8f9ucsO/xjZLW5/OnMuUYtnuXKJu+jUNSU9
MJyzrKBqvJSD7ksDXr8lN8futUZ0yuf+bqgK31/cAERY7xXKxObIzshK4xf/RaXZ
LQIN7N/KhMfzzJRG2ccRJ753Zwy65u0cdLr4jIRz62gI+P0DfwYIcvEeZstFeZ9k
VC+1Y4VAWiMOpxr344mOdsf6JKxTE30WWdA5Yzv4oI/kZZM7wCeBc8px8U4JjVC5
4YUw2kf9H999wBCrWiT/lfMCcEUhqZV6S4fLOFUET/KPH1XmQxodCge8HguQv+jP
P4YmJrXhGa6vS+GkX+nHldyBb5s2q+APp6ljMQUX6bYzomjvxXAJFiCuh1mW/M4N
ft/lAdEfxz8mJBaGymMggmwmogorHqis0YVqScJdqyqyZgcrs/NXzYxK6ygTKk9U
XArwRh2o7dkhyESTFQ7kuBnSV8t6Zl+9ubJoiPKQ+gNwuGbJVKC+mO8rp3SjsKfE
dLFJtQSL1gZC0PM6He5k9p4NSDq6sv+nvUHtHm2ANsZmDSJQtjFV6R9fx2f0yj7a
H/BNSiWE45BPEbB73BPOJxd1lQy7UDOScdpNO7ZtILL00AoL3kEuK+800MLTJ4kf
s4XsLkqR2WAbV6KZWJy0jxe8Fi7J2musHdj4WLTz8vfuNZJT990iv2nBgEE1tf4A
WKiAPatXiJSGTDXay+S96DRLwFKvMdBpd/vFYZX3mG6lW4HBYii4gniLZM7+9aMN
pFds6kJlHXGMpcMbSYjzSokZ+of639lS8x40e45mHjsFq87jyly2fqwva7FiIYCe
UGHd5gzhZZm/GNjiB1s3+uNcW1QCE42mFAtW5PFyp1e8jKzMa7xj7856G4tj+J1Y
cUYmlqOwo4Y9+TyLFz5pyJ8x3f289Vg6g6jS1crcsURP8mRDCxxbVo2k6xGIHOdk
oocWkYRkb49pJeRMDoxEDg==
`pragma protect end_protected
