// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gfeL74a+9FPKE53crhxOHukV8pprQSugdM05e7cttrAxQEgEzbUwM7V1KcoF1mYc
T2xKgzCnB1CtZ9rJ2F71Qq/1eW3WZAXb/zcY7axNXRwB2UhXlL690YpGSW008hln
AA71o6dwJiQ3e+ihCpADRnqmBe8NyGMfFy7VAm9Vf+Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 42576)
evJ2FOg5HfY77g4ksl9tdTMXiH167j29DfGCyRzSUYeGM4oqtpf83z1u4pkbjbmm
NmsFwm7sSII0HPc3cFJd0nuVYCXqC3D/LYWS8sxnDFx5BOVsx84NW6tfIR/gU/Qz
u+hGTk3tlEzHCfJVqqsDWDe6hgzvMWSCBdENUBII6oyI2hFtJV8fq9+61jNNyu2n
3yN1SKYaBdRU333ejk3xCsvkPpLsehdbfDo6auU/57BWs3SjkUQ/6Og359iVmN1N
0UYWf1ZqNMqEfe96hP0BZaeluhoFO4GonJWl6lrBMDKNMiirVIrPTUbEonZU9CsC
32pzncMduQmPA4tfzh9OczdEOrvMXIecN3KqEWil+btJmlC7y0xTA6qLuq6nWHWc
zQKdVFpk7cPdVIEoI1fcNQA4Ffo/a9BF98p0uFZEHddivEFL84eZ3dBfxkNDK9gB
VQN14Bk3AZ+7SNtV0DTG/OTh4G+5pP6pouhq1/BHnkiNgzxvpDR5HmEg/3O0pS//
1alrzaXKqX73EeSb+SM1yHVRR7zCJyW9A4XO+QAt60CzALWsZBjrWQzFLRpJaqks
hlGvz8+XtdadmZYg51AIAMOqyleEBH6Kfa6XPoMUW9lKvExp4mWkvXDk6mcCqflc
XxExz/3sVCSAPtffLg6AlAeM3S1ZtrQq20EioP3BULlPcEJ8M4YMXpd0TrC16Mij
EOxqeipmFQMLZalLu2KVJkqcAng0Sm+08yy55TeANdtDsbRsUzYb0lBr9GdOC72B
XwKrzf1e5RogjL+ExwHruKMubFiU9CY8xav8J5ya7vidSyvb6nmolA8EV5jgmbn2
Lkr9Z1YJy4fMWAZYxwo6lDthRZgqWBjp8+13ptJ3j0Ro4wW4vdTujYue1G+5O2K5
OOcBfkWbCUHWMeAOI+TujU5t49k3zXR743HZW3BBcmb8XCgeA25jS8FmiQnalNHv
I1S2KBV9K6a4zSw+tfD7gTNy8KDs2vN7YimjYFqD0XNLaVm8VcaoG1052VMWiuNw
uTxWo22AKxdwYQhu8J4dSgKXLC7fgmkQbnLraWBIMWysgiG4JSUqvVPxinbPVQDN
7ec57/9jAWK24vPEZlQh/zJp8738uFY5gD9gp7tGJmqasvrFytIB8+n52PEdbfLd
gbxjD5bOguadA9IMsS1WC1AdrRfl2b7UjSPXXAto1nle9eT5E6hGRKiKWFz1dlz1
hrLDhZKUKlG9soqaZEGlxa7MVNS3XWgrnScdCF48JIIyjDiqU17m9a8CtiQSSUMU
sIMuVFAllDaMsuH1KmZLJvHUSsXPuk8h0SvJbQHIA88b4mBxZmuwjt/XAXsn4jZb
yFPI+gF05Ir6OCGsB2VQ72Y6vcoxGnzuIHwR/BGm+2vG/1O13YEkNtBpxKj9JAH1
nktxwO61zujSJcyr+pPi2lT4kBzWbZha4YeotGZnnMt557GDWU8Vm7yUtN8PcRcd
f7JTrbzqcLCx8x5wR/eFgtDix2L4jwPgsvF2RAUeoCkuFQGJ/oVoV4TWlTUrDht9
7bDhxxhf68YmrxCKpZ2XHIIVjnXgJAOGopF83Js41tQNET0QPbpePDmWcqs4gjeI
nf6EBjwSrt9a/OpQ1qhSMOGG3kRH+Tq7bRS8FS0d3iVH7hENbf0LeddFSC+ZYfFn
96/oDjh+LDTTepqI3cjkuk8/uyEFEMHi1Hy0dlQflMX1bIiMtll//4sp+nnp7ZuC
TvwtfW63aZiYFJeHP2uA/Q4UeDelB2c34bYJDYyHyOd6xiUGxFRCfYul1yiUdAL6
iw3rE2lyW7jR5L0bVWS6bfIJZFCps3+eEhOJmAG8GO/uGJS/1lKQj0kqHuTqLCYO
aNu/6V9f8ZKCUbPS2fs6HpOZ4CiCP/opXejyNbilKL60YesudxCBoMAiXsWNRU3b
LOMuk3fL7eRWCL9Gsaw2qRAk0oBWiFbgbQpq5ng3AEEI6YZyuecFhXrPoLCkvQ/j
Zrl33DlDp1sDVUHJFsGuZGKb+UCOWQ6O4CihnZmMDgVKRDgsRaeXUP45VgaeRe72
7psGMnqlVvdy46rPrYqna6DeBoVhNXK20NCm/3V77n7udbqsUpFijucXNAAQzS6I
k6e2KridsQLaMsDlKXFzmXNDwLIqd/Q7ntrx4Wikhg/qRHPLzV1fP1688hqUuksf
ZpeBH43AqBRwuhdUQPLPkarHRNEpq8txINn5Wlvb3uPqvQ0FYFRKycPqNSj7OVQ5
ACn1bcS67WXKqN3kHZrxtsN3nUJ2ndyGQwkq+Q8C+DZO4P/vVHrOclzPliJJFJgu
mHwYRxpgi6XhFmQkXlVwiHW4P9OXdAyC8gSB+BM1L6yVmmC+8VMpksUYUJaRn9Vr
SE/czQxjaYG6v2VM5QHgnCWSdwETvGyvmdPEmDutUqE48GZF20ajB8W1MioWZ+Iy
Xt7Gc5yf7c3iMilVO3HV5IQB72HTMPQeknMjufSmzzcbY0j8smc1KyFW6yZPSm27
wwNDvPs9M8bENHBO4I6O0xm2/6XhwPzez/U9pwHmsKOSg8KUpkbmIJfzG1ZyOUyL
urEVgur9cvX0YpwxCd2gaquu7o/jbh6PfjhBw+dFI6FYh7vERj/SYC+jSXXD4tgW
Jlqx8C0RnA5fqavVVlUqQjFN6MxAziHBjHcO6IFIbrj5TdO66RwtSwX9ubJ+yyy5
O//z10OlePbR+KimVPRkGgTF9P2sfypSWAvNEjvvPV4mpt/9WijAcgmC+DMsOu4o
eEaxmzkPmuHgZJZ68tjoT0liP9auW5fslcfSOFmvUg5XdvEDLuREYGrWjec2w8RN
s5rvwV2Z6nMb9g8PfFX4AaG7Mu020tpAjcAhpwWA7h3MeWZN2Mgds6YVgXPrVdpK
riL55blVdttQTTugT+GLNGBXDAwK1DM49xlrC/SylWH+beqIIqDOkMQ0qE6v+nUv
KL9d8NyoXbYDEOS8o0hORGVCDqZux7sE9Dy5/a2j6PBUiyxOOIojjumXXu7L0eCs
qsaNKhVGEily3rgPMaTfy/XRXAOEDX3oYYBglCKXXrXaOLbKyO5KL1/Sv90Yirwg
mv8kiKzTdGpkXfbn/KvwbGsL3JGgls06lzn/qi1EtVitWUhoam8mMAfQ8MUlGYqz
yFXo3EDFwW/ACTuqOD5cNsrcuwNmmstCzKRhcTo5ecij41qgY0BZ0R+lN64QKiYy
ozB78nVkcxsIuD9l3LXnbJ2nefnipXWu+t2PxdjpJDslBbIuUiPwOaZo1tygm1I1
u1yfbwXk2l06KzI8AbOON1rXL56msE+tO8WLzpA1FeFsJ5BQX18YBLeXKR+QfPbb
nc89xo1qx0nwnffgndNvTPG9n474QOsbi8SwWlCfUmN+LddNLc45aHPpBrUJys9n
6ynikxeDfsS+WTXYuHPhIthLpfmbos9ykFGPFtQspghWsHcbrB3uPi88brf7+kgg
SNLMIKdCGyfWTpariDHrESsbF5Q42MsHFcpUTCDv8i2nH8rIxx54fipEI+mMn+do
mHzG8KFaRdru2ZlUI0s7MaRrah9UgCozThc3tvss/uahzMluJ/Eh9ZrCIQUiqkyt
JRSoRMVMUo3HFPCC2c1yzcaxoNyyCTdTr7c1uqNt7//bOGjYpmhlnfPBNHJxK6+H
r94HK7oq83MGLUy6oqs6j4GYFZ170X9QBXh0dxiPAb073yD9ZxnZyI0onZh/ZA26
n1j3lHqVJuDcbAk99PDIJZUXjCz3iE7DzinqHij8DX3yoLfyPoXisshYBnKO48Lc
FuXygXXVkNvPoS6MvPNa2LMU8gOBlBbP46j6x4DN4OGiOnI8oEt2TcYY9urRsUeY
izh3kCDlysk0H03rLMh/A1nun6nuOyY1jC1G8tP0k+H/4hF8m4uE1+xI3PIbYyuu
UEBJme05BjJ2Ej/DdaE5srJB5GcLdjsVT9EZmlTX/tau4KPraL/ZnudFv0R6mr4R
p8B4ClIlNy0jW+ONCAvjr6dbzKWqlQBYOGZuHGbp8HV1t3/LG+Hej7ej8WR8J7kK
XTNzjgJaNoEdPMnfeyLRcKCuA4PfuFWJbJ73SiJ2LNP0VzJtSo8mrngP/3jGKOTK
6obFrzjnCQk7ZGxwK1iWEqxKuWIsMJsMMd/Xtm3crYE9hqgw32LqkYMl4yOiu+0u
OM3v/n6X0y4AHjT2yfL1TKdbu+f35Lz1afHyLOSlyLdZBtiITex+dnQiVlRJ7/JQ
umXnd3964Po0oR0o0gBqfW+BosatBCGWDbyrdwuBPp93gmIkJqkbHub16bzeDDoT
0swzdjKI3jEKdyzistVLSGmkLdiGHQpY2bq7PKy4Sr136dPiUi6JBthudNLKpBtJ
YDxlpPbez6jAkYBPPoAJujAc7pnf/LiWu+htXHBqoMpIqKdvX0ZOZyco7QId2qMg
VovamU9GeLZlftsvNE96TG1LIaYlO1OTo1tFlbOJpM/oI5EksnrdC9gx7iSSbJYR
aWqL0/GN3mdFKP6xyGNk9YwO/2TqYbwCP8z/LFW0w/eLR8MwlGqZnK2zEbCuvzN9
yEal8IsEpv4tlmGxJjYrcFLfnkbRxO+D/I8s4BcHBAjI01zCG/3g6Z/ZYnYi8W0c
GYWbGyZmEK+Go9s/8MpQG1MCtgcjwlwa2XqByTK8jaLd6I5xPzu1FmImnYWcrwNW
4fyeCf+bGYjyyNb6+3ZBDob/O8antXlATQLUnnxAUQw2N+FSk2jywqs45Cvvol9j
A400UsklodzuzXypWmpKBcZdjDFVGev3w+je8hcT3rfrt9xNPgUNcNcJmpWNyOHp
NrtPYB4qeWu7b5Xi8gRenRE5Ahf4pKWi3gKHuAvXVGWCxRCYuOGk9gua5WD0V5F3
HKR8X4sRC5GhDhnulcWV454Bo5/BBDybxdbIkJlpj/DsP0XVtB0HTe2X/J6Mumgc
IhYp60wsNECPFWOB/FvnsNjXRApcvN8DyHkI166K10ICboDboqaaNd/vBbTb6RGN
3ijB32kM7HjYr7lxW1R5Pm/UMfCqnmv6xCnp3U3MvB+qGyx0LpZRwxAsISjuU2dg
co5n8PkKh3veGVVHINrWLVmIglDt6cfJgWaGNja9yc3IPYBK+3xqVz6H3WeFPrjy
9PFpU1x6vvVXtR85UzEnMTFlkijqFHVVvUvEEmSg7eNvzyj6q+bQoJsbH5Nxzx6l
07hP1DtzAjAIZbPc8ZYXBBxKDg7gbFwCK+L1nqS37rhQqRAF6VwVTGFWnrOnQivs
jJb1GO/Yx/BcQUgoYxpf6oa1ZxI0TsHW5kHPNXSRZPjrWJgxCgdCb9B6nk7qm+wT
tUGtl9OYTlXCfMlfUpHfY3zrjBKRNLcWZhPt12yu2/vFyBCoE2iyax0MM8tD+hfV
m/F3PB7oJCz76vMAZXBDr8ePlWetYguOrQ5E5UMAuQtfF1yWa5NLShai+8wd+oHT
CLCT0IYGCsHrMyXjbaqae4XvwQOmHwY4woPft0lmxY5UtU5JMFRBBS7fdes9FO0P
eBgN90DUOP0XL/6NuclECmt0hul11pp5VeeHI7BGvuKqC43yUbaZe6ClM3I1lK7z
d7fl6KnzvniWZzHtkhkgVUy6SiR6voW2ClOGGnLezNtcGdjO09/56RgOOFkGWglo
hPFhgDiShWkdzyn7OGkwqtr/jtGl0bt9N5s2VnvsenlUKJk4F+cUZcGPCXZ/LbTP
u8/myxMlXQII0+SVAilm2/zQ2K/g6gScZIyMFlx+XPz2nD1RgieedThwoDQ1/Vp0
fDwD3xrhO92+iDN8w9u4GVP8gcJxpO/2A9Ra7WBX1MlSmKiOGXNGkYKow2bsaHnZ
1yLgxpG4CB4wD2QKzGYISuB7c20hVLluNI1J4mSgE74q4dUGTV5St7YYxH3Xqv0n
brE3xrvzIImo23+XGUft5AuIlGJTqYJd+gWr7KPZBTjTsXaJJ3TB8F8awJHW+Laa
cSv6XFkOldmz1vw/WALVe1UIYbv/yFa1ughjPUPQEvYlJzFRAgbGh3LBhc1f5qWo
gSD0gq64wpvzU9Cvi02B5/L3eFh1wBY5JXuvbULOJoLwcOtc4dh1Pudd33Xu7Ams
GiilUOuf+9VTDUxjL+kbuvv+0kJaEf/v+p1wYPhKfbaO5byl/9ehS6qEZdxo/oer
21XRci5RWwWwcyPPYyNDWptTcx/V9uCAPfi9z5FN67CL3dFkMe0l7mKxgZUNEj4V
H23IFTcwcCkGZmeI45S0l/6c++L2H2JIMx0rhogbo31qpsaQxB6WM9zxTYjhI7H3
deaYB560QYE27AqMfTILNV9I4AzeXn5BJBGV1cHv8Y9uN034l9n/lLBoAEAzQf9Q
7EaLEHY2Paj1vZJrXJgt1IPYYbJHX2vN7DYBNeuf4ioegVFjxMjryTZH4wDZhm6u
x0sd0JFx2E/bH49jGWukgwwaIqdAyFTJK3gFUx7IvKSUPiITUwXs61IrGOwhLOFX
4oRwlsKR1WBgNsd2ylzwaqBei2DS3Yg2u56evZl0aumRcPNEUJssPPOzpWPXui/m
eiwjgXdn+C5Ts0OKytSJongeyCTC+93tqLxfSaJoWPSPPaJDPUOrmK/d0W/h6deD
kyYStdp3JRS5BTdq6OMGvcKXyszmhklv1f/NlVtB9dpCwkPrIjIm2pMxzVmGp8AP
IyMqrmZHTcWya6bAe+TdE6i553TKvD4XQ5Q7QVIlugxml0MdLKZYbqgp5ZWh3IWo
4u6JEp3itmFakMfjFuNGNv8ovSL+JLWkvDYa9XOHOr55GxQ7uWDQ28KwSqoMrJ0Y
YWwxoqaWd7E2nNQI5XkPco406R6SiVi1chLV1bxTE/MRK7qJHa6VAcSg7jdXGu15
RrZYhDVAW11iiWOHDoUcn4zrAEOOsifVs5MzWDpN2ZpY/xEcUKCBeZZL1mlDlOkx
drLIvEtLHXyHGCkJDVf1p90/T7Fy0gBMhcw8MsRRkVMjKZhaujmbzROp26uEb6Z8
ufPWfjWZQN2AsPPxaqeMGQqRsAdQ8rzI70rWTjHd3nW8htDjV8/RRNO7AhkQ814Z
BnUqDKEYhYCzuFdg4uWsHk6vVK8+o2s+2S8o6Px63phVcakcJxlb3y3Jl0dVecPg
W4S9/7yJIueXV0lRXk4Ig9/nmenVNFK3wACalP7+hiRL6vvKYR/fc3Q23Yze/svT
cNI4DnGKuoJtM3tKY4d/Suk9yA932Z1VUgvRW2DOAHJxwtUDbe2DUOiitdypbWiC
LCCEw4ST16LCD2zTWfeUGaooSLwGAazeiU1j3Mc+SsXXpSEGY3jGZyKtzidD+W77
QzZRHCMigdg9vywxQ98ighCpcpOx0ePiRwJRUlh79D+Hro9hZjHWUqZ8TASvrEij
n7RQcJPq3/Xr1EvoVOGnaujgp67miUBFiUBayKeOMFONIaC56SJVqiCzM4i8oNcO
0lQfpHGdt60/6BgV/EEtbOaQ9C/KrNJWWM87TBw+s8pyenMU+xLYeBsUSTKyvshc
g7HVv8rpjUbwbJXAg/j7QheLL1382S5Q4Z49pt2Ud5PfanHvAqZjHVt0Y+ZYBng4
UsVGhJphzetuj1u2tKcIntQu50kiPykvSTzMRj3bbBxTVBB1ms9cuUESiiq2F0XG
wEihR5zHpgsiARAmvsIAQbXGhc4ru/N/UDv7MrjUasYRe22tzFB7r8+ay3ZY1pHe
p8vR5WmXtwSYjw9+y/kl2yrKPJOmrY32haPZI2MUpZcCo8c0mNWjCOV4KE7S6tGd
oQQcKCAu/3jT2sJztziqCkcWEp0hvw8nUU0UdFw7ebfPlUYqaYipa0GQF7FrByR9
MEBQz3xCl1hQxNEAGQoQbMJhczhD9Dfk1y+j/SCwPPwJyNyDcaGbFmZWr8Bj6F+M
3xItb6TBE9gF7YFEwsqPGGr9ZBTHMD0KW4HJl+dgS5JWs0SD3jOi2zD6NeOy0xsw
6pGFJXFwB1/FgzCuQQlS1Rk0fkx+REPvNGwZpKfFtO8UQEMTaVFq2BLH73z5+0IL
loCd9PojlHsD3MPOz1AKJ44bxuupOORjYgAbO3wjzZIZiW/RnIUb/RyGIZkVtmkz
g9dlstcvTE/EVTcew0JNsmq0rxh299luBFf4xX1CcG1w/IcxL+zuOC/2/ZgQXYZk
TjTQzMcCZbKPZdLETiV22oi6UxPF5vzEbX/Jh31ucggrjUgGTNPyhlh4wsujH1KG
Ii1kftrCoKL7LW5XS8CrdOlkTKnHSjTV5J7tevddqwQzNqEeI+ROb/UNxtREoOaG
4QTEAOObuf1fNsb4Jdt4ED7HtadzTC6dboGnRVS8ppbafx7O7QpjiLfVrmloVymG
u/ZwPw6Y1lkyferqPht7rB1usqVyGRUcgW092eCS58+0zWHFvzTnT+7c+0qmQgUF
UoF1aOEKyH6O9+iP41TIU8QhETOHGHBp7F8CJ1Lzj3Q3nfFI93wbfTTu/g9CXGD/
Hm06MfrFc/8MYxjI9Y4x+PlcBjAOETxUhQMLdFNLQzE0EpMZMRu9HuTEN4Mj4GBf
0dAZfgBi650J9m/heY1LaB09CFLATxFZ81+h2D1j6ojd2oaRXuLsjofxAxhWYtgY
IRu8TpiYtMpTz/qD5vRX39WyeJc5bmLKU0mKN7ygt41GMxXmLSToSUhLYvTuSERl
gwipUsRJ1iOm8kAJIfS6iJ9Ue1DqZrtLagkbjkEHlk1KLKNDBkDxhj/0zXwE14h9
ngZUsgZSs/z+jrCoiIMAcS66h1paXUe8nW6c0D5vjKoO6KbPyOY1sv46k3f7gCQ0
SCk60WUb+phbDbJeperwLu7j3Fj4qf7Hq3Cmul80ovq2P5rG3px1tPZDPDILuh0i
XyQfv7e4qU3xPWMZrK4DXHPnsFZA885IqvQf43N0fNDHywFhfeANZ3xBhnDLAHBv
xGKSsIv9JZJihKvJ83h4DRGOWkWoYGpwrjreQl7RjGU9+4PMrgInwrWD6CRPphep
Y7olPWJELFro0A3ei7sFt5kCFJ+ShRIc+zalhZmxFUaoJj7Kiktw4uuavHj+7HIY
8aENyQucc1WevSh5Zc4s1wLn5Dt5ggnsw2gtHOmO2T2HmjqVh/6rITTEKUzqbIMg
TAiCYhb32OwBPBFSsfZIqFVeHrAQ/2Wj9DkZ8lixeuyfwTy4qxijBD1MIuUkIBlZ
BYif/TSDPEEJ4WAy/HYMqgcYHi7DkAIezYquRE0g/h5WuFwz4wXEUWWj6Z7IdByI
E08mbY8OnCuEsja42keQcVy0L2afj18xLTxRaqmEQOTYgPOG9ZeUMFBzFDDLwOA1
LJHSLHABX9K56sRziXqTe6bdFFabSJdx6sfXqlznB+uccIxQIQLHW2Aluhw7azkP
McK3LweTdT5p/LxSvIgzWtlSvBYdx4kV9SOklNOo6iXTKVB9prrrRpM/6yvrAe2Z
kcFKZzkzK6qkku6S6XXHqqJUaMbx0Ei80HqILcv1M4QdWBhyArAGvKQOLq8/Cb5z
PEABbtegccox8c2hbkyJvrsvQdNC/Rt8uka68UM0d5wqQTAJkypXsJurEu8gJvrI
JlH2s45fiVHJXQuM5gClJ3DmQ/r107eeE6qRyJjhieVZa+zPdvU7sQJE9YjAV2Gd
WprtWhTbaMfMrrBI85RvW7ahdd4QSSadf4ZcTM9Z0QRPPfPtNYmmjQk/busK35G7
ds6QcWiJDCQH7LXg48YBfvvFPdpji6ww5Onbo/G3EeMyAMyxsczCiE9YtFgieL9N
xdlklo/3Jxd6pqf2xtiL85zfZOAJuGLv1xcasXXBn7IuQwfKSgbXILkI1sD8QrPj
PKnugEUNp/Hw6YPMdEqvl7xmQta+w3RNlFXJNptZq2VkHso2oquaonBrlpkV1WRL
yppgdJ5qznkdYsLxqFrVTk6vrFJH3epdyVKVy+O/nywK/+TlCKxiFSEXf1vXeL2S
816ZIkPSCc8kxQsHQrHxbikj4zMx2j+8dyRESWN8snL4odjpjiO8ZFDuXxORRXHX
QxBQHNe7krx+pFqkl3kipEXEASBfy3XDmcVBQ8kTymOxeh5/FgvPN1M7MtADdZP+
Cq1PRihItEizqIVTcv94LKGA31j/8DRWiBrGBTl1y1lCF2+cK/m8MGFNtOO4ob3V
fXVJAzE7tsc9zriNpg9mZPzUg7NpVkpD8Y0y9qubwzJIyJMRIZHMHdY/VUhcCysE
sSInnMB/puJVJQKRBHW9GsLK3diaAuNpnLMzKBaDxTRCkRrPS2940XUh2dOZbvuS
jS6p7xY8vae4o3YlYMQS4sO1Asly05cjYO0bz2bxMI6jgqhSpbHQRc2ANheAAa5z
OLwt4NjGfKQqI/LuS4RU2gUozVBnicmWghcY3U6YNGqS18OTNleXBq11sC0bRy2n
iEt/whkxd7qIkXuI/c+ACu9Q21Z6tr8F4GQMcg3mjtKpajMXKm5zi7V1LZtX3ka6
cB/yN3EzWwU+hv50yMlW6zKjJ8dh9jHrQe8oqsUI0+TAQJmbVhLcq9URzqRF9Fw7
U0xjbMHnQ+HU+hSttwLZtbY2lznmKi/bkJEPgy7epXwGdSjtiolNYlKO4XzNUUq2
ajkxeGm/3rno/3C/41PXwrG+GBoVsrcH25d2dPqTOyMzWc7FA2TNI0JQ7mdAliil
CVZ0/9Lo4KtT1tYLfbqIRPjYLBhsPDtxj4e4ZtXNueCpNvL3oWdtTQ92hSxmoPKk
X4ssOT7Fo7UBqLBDwv80l4z/97za6vDNTeU2edPdZFBopINKRvnpWQ1bdbiuTzP7
QDXZX86kV6l2zrYRkLgRG5zwrNM2fCcWUOnUE/1k/Pef8YKn/fdd8/c6M2htROQj
kGBPMyXTEychBjeSOkBcJQHh8j4HCiruzt1ffUN6Eiv/shc/DbZydNeNguvU6EVD
thEmONQsu4iMnc3y/h3/unfgiULp5MVLaZqtd1FNYWmot/f61Ji8FKK1djr8THzF
rGYuiM6c+gZTaa+97BKle7v9Fi2bF6+zR2rvRYkfhbAVyX4jm1ncuRTgTM5AwZVr
FLVvr6WSthaSpVcouDemLNIDY204t5qkUSqFT9EVdApRog69e7+gEgj3a1sqQdVH
HtivOt5UESTm97v1eOYHopU/swHi88h3z1YYG1anTUHffNAV/REl80TEduGS4p6c
XlWSOY0/y1JSGsShOf70ukXuxonKCNhNjN4wuozh9G3UYpBKsV5F+Zn1BwZ+hzr0
xcHbyxMJsXXKdHUJpdo8Kj/VdbNePdZlZmrzckG5DfTlkeW82GivXeipk6hA7jqm
uJkcQnh+1DEA1lHlq0W8b9wi7SqyFXWB9MMNLpitHsrIYcwJxD5XcEbjIRaUlzY/
TKchdsgIzdFBCLTE/g4qvLOhkfOXqVDCTvDuXEE/tSXA9GQ3bKhG+gArJryAZ+jc
psrky22xUzQ1zXCbRIenC5Pobf6aTimlL7shSsSQ/1VMpgXVaWwD+1ZyOn7QFBXr
pyjldu9vWEh2WbAFshZvTFisMpCj8xYN2yvn3avLHlt7v5YmHNiSRN9x9n9MZPgc
qQi7GE7f7Z67kSBrznGkq1pwva6si8r6Dh7KWIASlQzK7yMH4mhpxwKqWsxLCA62
eBSP8DYxvYdrRr3zWDxaDSpN7SqJy23X5nsVJeUT2qAs3EkYDlu18IGx5bQXspXV
JFh3l/I5RdXsffETRT1qhTjOM+3/aszDwx/lNzeZw0GMYpEzWb7fKwRSyXpMSYYz
ypAQT0HPwSPAfesLhH6ajFLM4Ca/jHbtX07T2nzepCE+hf7rYBXD4eXuw/ZvOXWq
ay6LCNZBvpMMvJNATysJ7qUmUl1Ezo+ucbxGc4uKOH0hjhSDtoCTSNEfm4LPBUSn
atAK/Ogc3A3odp0ridzza+K8b+Y19Csy22Q5S/049/nMj6ogOVkVMjaEBqB05TZv
BzEQHlONwUFARyYcIz1hZROJgem3bDBkJhhozJDBCHtEZjlaotujl1F5DBiAomMo
JSDPBJJeo/3thpSFjBpg+gQuvXKIXX6vWkxXLK0twD73T9RTRqtFPJ9k0+MYjpYj
2MKYF4HjkIFy3qsRjX/uENKvwoG79WVCivEH2VDax51A/A59sK9PtBZcU0pin/GP
57ceySHznqj9+IHCmKHqmN5xHOx96tuUDUHj4+9OQcevxwgQGKUsw2BNt+a/3x5x
kCPiVbybVlerUBeD4FriCI2XFqu9DMFE0wkaZZXvhmtrR8IsdV3XVjUucdwwIDXY
7OydrfOo7LTr9ygfkgKWuf43tnEQ2gTEawUD6Xrv9XBbKNY72dV4tvKctjfTjeM/
GOYdm2QRwOuAHoWvXwMPidw9U3gzzFQB0HBEZVLgcxsqSEUjnygaHM3brSdHnHgk
CXZIcdv5z0yBmt1hI1AnwKExuOWilMV0u0Ess39nv0U68e3q/oCRe9xo7DvrDiW2
9OHfJ+iwEzP0k18dWKjwKWjl088Sl7ecU55oHdj9MOXF0BfSGzdkKN5XVvCeMf5/
jd6nrgAaB7Rvyv3eKO9YcBDaxDwANhzQS2vnEXMRTpSk6EyIYUY8SwtRTmLjwYL0
MPlTSDAG2fl82knJJLOmEUhX5Er46i0eNA47OatnSZIYjeRFBMTE8ccyz0Hu0TSl
o3TLBPe5e8qlmBThWeBeMtWhd9AYfGNHxKGgAGRK/Ql9K6bUJXSP/1mMu7A+73b+
/upf22UlpCSzbctHcix+4xpSImREj3EYXPAAxWCi43170kuIvk/xNQnMTXC79upL
bHXjeIWED+9rfoJ7bjZNfxYr9IH6aY/K3J9DCYljOWFECAzlOvpbuaSfHX1bShrh
4gvv068uU+Wn41uuPJrFj81MHKoZsdzWVqVF4lJJkUSwD4qX14+ktDCprQvoeM30
aye6HHaIe5S4viinDT4VAMGsD0TWazBtBX4/apRoO0UVLRA1tLHOTVxecLEZXL/n
AUW5lRZ17p1SpHFGxjor4EM/WthX2L4d0Gy9mt1QWMUTCoCZGzHJNEzWhaO+MSbH
Cmpq1SoYYBOvzPnuZExzDSZTlW9BZdEKLxbVyfzsCHdgvslGc65zQ4D8aR5GUB4w
Ub7rZVeyxYFVlUalppZPJDM/BK+X+AJIZ68xxBCYHjXwKuoeqdO96jCkIkyMTw5Y
lN0Zk+o8QeXvKGcDzk+V1ndl54naE6W8efixGAVb97aNjHS7iZDjW40NC6CHHvk4
ZR8FlAcDQOeR9IFTf79aorLDrA4w2c0SVy8DKmFGK51+tp2SrZfw5wAVr5Lj24BO
/17b3BCya7+iYYoETltT9fQmtoG5QSHWHKXowmT58KPDTmf88z/xo/WWXPjDMZk4
MkzYaLs8rj8qiVpLWW7sXFHeKN3nYi4iZKKU75orApWjLleUReKVW2s7KF13S5zW
wEu5+fYfu53Y6/9EsG1chHTVeXBlCVW9Q3vCl20P71uiP6TRHCMoMls25xIPKLsI
BQs+EfN23pnyOcew10Twmxar5rYlIf6oueoYAbSCHGWAFN8hab5awkHx/2NsvHBh
ocCqlS4FpyCvu3B77QjaicSMEQDcsm4aoM9mlWuJln+mwFS7M/nda7iKqW1hyPzb
SaAcOynqhpppqw4OlQWyyTysO5ITwcj1j06MRlumMmUTL+hn4fmbXH+2Tr7ojJn0
TryN7Kj1DIRvH3Bt/8Z8rmi/Gv0hM9/iKQBGVlTxMvxvqcDTjtlLnBiO3x8FGXej
cYlP6A6tIHox2Wb2jlnD2/IxVnQ+dJiW7a2AR2mGWTbxqXttwIyphLRFRdoxFp5Z
ZhnrlKAtTxpRZKEdIDxJi2SlBBicRit2amHRXzgJHub5RUBAIA/7eY+t/rLWmdCL
XuEsryZZgnFx2XZFWa+rX/AohWnWSo80v1uO81uqTHAB+2x4GOZvYj6ZCis8ecQJ
6GKLsRRMpDqerJCoWL42Rdk8XM/1LBvKlX3BWcxGEMlTvKIcVfp4wPE7cJqORpQD
mgoeHR9NS5u88sRUMRKm582mlrFAYtzcqQ9nfz47VbaYXd3fOHUHpzpbcAYup4dV
y2y8Y+25iMdQDKd7qD1U4k+e9wB4Zfddf3FTYrPGQ4/+04+g14FbJkGfXkvLFgwB
JgtocN1oOetZzJnwTf3WOWlZEpsj2CilYibb+4Fgv0MFPHmAVqi5WbJT5dbzMaU8
fFbaEQ7MP6rqY3PyHBCTBtp41G1XKGhm4AsHxMhV7HlzDwlZvphaXlJ013B3MXdd
bG9YvSRvPaAdJp/MTrKeWZR1Ko97fY2KG0WR5ze9J3Lf8zCmfWi2rw/Cjfj2LNsS
YxMhcF6do/5ce1HQOFFAHWEEuX4OzJeox+wvzuj4MqSwvHUuG1j7SdegjqhqzOD+
Hog0i9N27df2bq1lMjnvClW7Nu7a2zyu561RbeyQ+Ywq6IjOCe4nNchVLvFbJAYi
MrMM5DxdwDQ5puOifA8dkDvBYNqHJzmLFFPHzQPz227FYWmekLY0gXnzuM4GDgTt
/7AQubB30UBw/cZu7mOVtzNdtBheqmtvA8u3ZkAaFosHjKImfnZJFo4W7gFTnI1j
ETyNFcZsOgZUGOfNogvNbNJRUPJx/GP2iyvccvOQhmkQTqagWv3/B3IxGxDzMXt9
jdgvSM6iyaet2E3YzLYSgcGJ7JIsj+LgwXA7gUblsbzTpQszqKmGk5/9okt4vv7A
maPlpHVQ5MhFilFRPGwo2PSY13uhxH+cKgmmyhtjJlosPbSGuveCNAHYpMObvG4b
xVfcezf3NuaXes7JAYXG+AkMPmkhlaybH7euu/MzMINLGHIl4j/RqwpMpcdUlN88
NMyNPkU29DuwBGhX64Tymia6lqmQ3sx4bB4BgbsrRyaSyHEqnxv68nIqoUgYltis
JeNXinUQJS/+md22dcQZhOFkK+3f0TuvzTJgo6VRn5MiAYoLYpqqMzM+3n1QY7zo
VxVD1hFjKIUX/fuL6ai4DN+ABCEaFSe4d58TJwhTfNJRFmJ+f/8cj6xVpvF8Fxdy
IqcVCQ/xzsLlwbX1HntYwPtVq4Tx7DZqMFBaTI5DLlSZnlUzN3SAUcI1vfQUfytk
+d56CYqlUFNssstKfKZen2hnan4GH5dXPM6s+R0+KyasNmypSS8vPA+/g9VKmhG2
1iao/HU8sObl3bWHAlPbjPvO7o4U8Rbgm3NnYJU8sw+7a4JJNWn+DSdMrn2dyDtO
O+Alw+hRhoIP4vFLBFHpZfebpSBcqwSa1rzMUOS5RVXEnDGNJgIwaNhR4EUwC54r
W3sGhn4GEgSOmhy3c1zuzcOXmJOfD1aSeGGu7cbku5G8JiALYq+Aud0l2kj1shZ1
pzRSvR3IeWFRhrZXnxLfKaRhmM9/zRh8n1U0kMb+uUBLL7UpN+uWv3VKAtebQpP5
BHfzUnPG9tQeFS+D2e2JrXqLT2JvzhXsjy4BzBRRX7qO5Y37GqJDO9FKfFxRgcSL
mU60osBLMW7YGeItLT0Ged8ZgBPZGgB8g2Zmol5noBxLD/bmm69cjYhyEDiial8j
tvql4cP9g9eOSYDmGDPTUfuu4eFqW0tHd/YRxENYOsJJJVHZ2VsU5x5H9P64w2sx
TcyaX4NJ9g0Qp9fTOEWbJ6VEhzzQNT23RpI+xBvX9cgcwA4kO1tLOzylBIk5JIGo
D+4jbEuMNeO//D9CU1nNfLMYtnhyugRmxW6tf/WDIkaIJh3StiVw7QQt8gwpndgU
DyiU/zeZ8g1x3EsWrEG2ayjnjtIVkRLRJ6oh4fD2Jqtj0fhD93pfKD4SVwoAQLat
ffhPLWyjfiah4Zv6w2f79CpWsbRnzh6DnSrnKUws8zCos5U8n6xkRr+bgtgUPnKg
bRAdQJtGh9W6uSHBTVpULYRAqlCpDDVEor04uvB0TjYmzFXE3fBFXPUdHeEd6WOW
ZQQnWU8m18DALTMAYXRvcDVRVW8S0MJFrkr7JJ8XUgdlHKL8qftL+pEkwZInASMK
ACZ+wezBm9QdPmkdZbkgR7ATuLxBUCCbr3h1iy2Of8w6mmAvU+tjs1sW4c0WAaMm
scG4V/CrRLzatGnv52fvnJvIYu8YYQ/nEZstoN25T3eMIr6JXD8J2r8Hn7cm51J7
lqOqvPkdFL7EjNLnpIVboJtkl95pKuGVrgnbdmz1AQR0wc8lN9A5VyaofuVsHpbQ
yWROLsD950Z1hZ1Hrcv8YvDJawIAenXbynWQ+32ThztaZT2xU9dRaao5HzPy/rK6
vvn/4F10gjD4zcigrBHFkKEFOgW2iRFTVFVcWt3Nym7awafXhHiQpRB5wAZGPtLT
ItgbDp/qIMN8Uu4/YIHYrkWA8aeqEZdKhausk6Pe4Ja6aMsDZl0iWV5vVL+dHmIm
mSGm//2q+tBitRCloQPGCHtoydPOe6Wy4mE1YeGtTUJwtLtTtDZqEAgt+QS/H4wW
gCwC9NUswU0bAufEtn3owlmPc6aq/AbSFdPXU5uGPceDM9RxOj3gkyg9FkMWgPRW
9kXT/OQ0Pk9fo4VfGlWdq9evVhX+UCVvvJm3hcuacsYDoOPex7nbL8E9LIEUYXXI
HSyKfJlPs7xtLfDSDY+MbFLjFdUQvLAqqD//B7WMXTqty3yKSqqv/BFP9V9aG/Sh
ETeEo4w2WLOliCzb17sHohBQ3opMveadmqiCkDkQc4UYtQIHGuSJJMXVSbogONpX
d2XsZLWrUgN96YNfsUz/k7HaJD0fmSmt+nuuWPFy+SKkDkPZXw6PAxSf9bVLg7kQ
sjUglP0WZ7X0j2QDYjaIXoLwrparH0u73CBTos/i3dPryTW0HXt6fgYI+HBHLl/5
eY2Ja6IdI0OiUw96VVdXpxuH63fUFksQGQ/y0QJhhZ9G1xorCAFZYrcF9VVc/H6u
fg0UbmHckn9fIWYQQA4UXwmKQ88A/2k9+9gvHgc4BiVpSdiWjg39WyVpGeHFG1lK
BBJ6m4LG2C4L63h4VESVwRudbCLQSoLafWkSsMgdXwyqgWRZK26jM+qNndKxxaAc
gL0O4vgEQB7gG3hMyQ+vCHM/WglnlFv96zIA12bAari6hUmdKJgrlDAbdBhWAFMY
ta6+2oVby8r6CwkMhUd5GeGpcd7k/mbkjwMAquywHb9WSUGdzjlW8OL32dffw3Fw
d6XcQk42hmgz0P26Mn0HIrc1uEL/q+eXxOdGnUo/HcrZuJ6wfuF2JYVf0kGnOnHQ
XnRJbVguvSEUTeAXV93s7JSNsrzSoyl2AJN8YAL2R5cLp2FqsNHDbx5I6SC/Ar7M
A4dLJe/X9u/Mg0snSOCOTNGZot/yWTV1G5+GSS/9K3gSSC4IKTGaQq97L6VQ/iI8
HIeWeMk6l1L+IcfvGWwJpio0jVIYaZdqZi1MJkrJK4jsssh3+WewFkolL4zNMy3c
WvMD3F1hgmqN1tKkLRlyZ3AMbMO4T9YAdEObbmq11ScRMEq6w1oNiuWV+fSpql13
N1Mi1OxZTYcjKv33p7bVxkrmGqXuELV2YQsFbRswlPs8gH4z5EFr1Q2NkLEUtp+r
fySxjkalFtO+vFKOK48myEh2OpbeyMapdztdTt7pagI96jzpxRvzfwCd2HdBWQQS
SHESVRaQyLYBeSn38Eb5VkO0FaySC9SbN4vGCLKuhHsn0c+qGh034btBkV3wyOHf
LKWzVqqV48TKf5AiRsfBAoQGPY7csClpyyMGdUd6zdXo+e8dOt595gD87sMgQ0ac
D5iKaISvRAsQzQOHFqOXBvC+uxf0tlqZKEMEZ8GSLFaZ4MIauhVAQ7EGeFd9Xg5T
wl2PW1aC1phymwE/7e2NrnuNpm3orLp6AHb9xNWQvWIG3lnrt3zrd6xr+sGuzzSs
PsjSidOEePCV0wkN6lVT0BB+x7U9BLUxmnzhhFZXduh9M91IeLRqNsMysdKZ07kw
u1/d97G96c9qkufizvRTm/L6PqrJRcBNTrAzh+MJOufZ5p3NZqwjBCsHK0MiQIiQ
bSyKSAO8fCvHUprm8ohodrpy9a7DxtmbXoOlQD0MDVNjPYhO2OfdhRFaC/gmxXUD
3dHdcn7dLPVa/yKCdphxQQ9QFnXgSVI7cigib2h2Wq9qfcxz1IJWcELfRQGsqt1p
MYccu/l2kz13k/AY4/iBod9uBEecxTEygNtRaP2td/oHv/iLv2hNNLVMTi0YrjL/
gVCkhFYKcFnCnznS65WEw6MN7MWHV9e/xlnQ3fX7PlcRDC/LgwS9u2mSRI7Iq2bQ
fpaUPe+UANX1ELmjdlId7oUwDseHk5Hrv1CsLsAszXjszhEZ9N/htm3owCZ7k4jJ
Qf8+ZUtwKJAH2q1N+CsydajDdB0kEpctuGIoKXo3DdE8XQtq2Jei9Y+DVaTmsdYx
lPGTYcH0TMQ3qBFXsQwiao2WR/PDgxmZsSKsngoi90jArr52AUtCWwsBC2nRCcNh
7gaa8NLpcpMvNazNSQgfVHnvmbwWdFLplU4A5lJH4Ncul5QAkRErRttNsQTh8J4o
1WdJqVxyK0FXZVF4gUxArTWqqoGmxBm6hZnAT3+c7sB79rFYGRc7670rGNsIiCwT
DHiFn4q5+DS70MEt64pU97+Ys0+b1tF7Gc/MbQc6jq/elPB7vFQAxKZBex+x8UKD
1ypJ/Rc+mRVwPFT3DcNM+YyX+CwMKp7wYIvyXoDSXLIV7FdyYMRyhZb+XmZlkNao
6dtulXiOU0jBKF5MRbGWVfmwqpykBPRxWK/orkTC5xIFaFvqGcCLXVw6KbmA3LNq
X8yhCFKIO0LjRqf9Qxw4Rem3nC4mZ7cqmO8VputPJNkPSHoprRC0d+Kw/qcr4sKn
6mfYxeQQYyx8OCp3zj0ouNcc4gYE/us9zlp5yAcCBrKnDiCqx2kde6T99PkxTJ4R
aC8eWEEp4R82hIMRSeS1nTgCLk+5f5mPXj6srfJmRoZbac7bF2ZGN8lLjTFHywQG
hp9krIuO/YJzajwzXt/ZfLu80fzBcMzuBXaoHcu55y/pNKLtx/U8LmRU1EijiLK2
3TRhmqFOzYfN+SXzAOtdDMWW4PjE/dLDUZfmKyZQQtL3aVz30WfHp9r3u4SnINU8
FMScr6WWbjq8wWo7/mPAdVXQfiSZSF1y08OX7UXorylj9ChUDU/IjDOjIE8V96Oi
hDP6M6Xi4pMsAI9Wc57CyZyTy6MwLmiT7Ln/JlKNe4b8OQ3l+jZh1/w3ZWLhvSPQ
50jQ7F5t4TlXV1d+6Xfy7fHYc6hs1BKJpzgluNEdAuqbzrFVFBIQyYIEnQsc/6Fv
ydLzptXSQKIGuNGF2tNJPFdjoduC1MPb6jCkvHUYSmDGC/Mc7wjN5xsWdWQJg43n
kFnuOPDhmPDpyt33ZzgLFwX9w89S6qAm0djBRkJgXatJP9JRF0WBa4x8/POBC9Ku
eW/kTpWQjYHVmR6ov81mzZ4kneKqcXUDaYBE+6eNG4vCjVAkI/vGv1v6OJWVID5O
BoG0hoZwm0CrAmxWYSeOutWjsrf/5nPyJZVcTS+QkhoRIKpf7yWbs/F7HOYVw3A2
B447sNzVHYIQYi9TIzQ8aqIq4Sh2nZ2X7bqSeGRsc72Nl+ZVvPR+WsN9fzrzlCZx
uWLGjAtEHbMj2hwfP/fEHEhthKr3phGSr4KTll3JaeDlPMyutEcskKE2kpvqnRMT
qL2aBQPbzZ2I6STGBpNSI0yZ8p9xLeGB06iEchsftX09N5IJtw7QbD9Z46vS8FWx
Xj7l/Q17ukJL0zz7kHYvXHQLxyoOqn1qvnOOvJGD9RmaU2YIkITapepfeInU11Mx
Qnunu6Owp5DUjiT+eKwEdo8ASg8H+nDLkNT3Nqwiqo5Zb//hzNBldpzxXkKYXTx/
NAhY8E7OoDh0nF2RO8siKUYHZF+ueolSQPeSQQkMcrHrioSUht8RH2v0mk/LMPTJ
gpHs46UEf6a897Sui2Ez0Lr+Us2J3CqgEdDiBqrtDN8SvlMqyXy0iSRHMOHBsoNl
8QRzcvjRXx1BztUf+mbRRYBRZKqDdU80M8N+1WTWlTmY5XfXihqDqdM4sWe41xsl
2HvAFfoGy2MOkB5IyyCrqs8YuVeX5P7/gBnlwGofJ6jJxfBggHyWFRvMukAgpM+r
7VCjKXRZ1McY/Fo/TTVASvScd+7x1xQ3XtLHwSjgLn/aZnExsSjTmxNBE27wZV6o
nFSSwhBXDYUaef3PShB2iQcDEaLQTQgw3s5YH/ZkgPqHuPDPOJgn9jd5HCQc92Gr
5/l5vTXt0k7RWLzKXTo+YqEr/ReARwZXJwVcfXuCmA1YU2YskwTD1os7TsuXdzzO
+DGIPMDOL4Ye+abikKOyuusXmzThr4EcX2yeII7qRzTHcQ9+4iWcSFeishYKy6Uv
FY91mSqw5J4JFaVH02TI58mOGbWmpkrMWG0GC5SyffOAksG45y2/wNqW245jRS2W
4AgeTblUXx3QExsqbG8FWKe6Y5kZIRtQETjV7AIwx/YBCBdI+Cdd/xsnsEOxUs64
3DYQlZ6/m0qZYeG0ysK51gN5BGjV3svkkzrZiL4ReL/0fZzrHRSeG2uS4l/b9FU7
+Re12QLMQMBJI23Piqpru5aNTCLnx8oyDiMiCqsOvknDIGH5ganDRcYe1OqsIeSl
Pg5J+pA8Iy2gCucLZm6xrHsGl0sCn+fcgUXNNBnt94a0oHpzCaEu2YthQVQ8syA3
7zlTBnNtYPhAQ1mhz8X7LNt7farw+/muHNB+brMDIvM7/MzzyxKcbcV2xDxEBzSv
r63VCrBFYLTiAJFoTn4C5ZwFXlgNBk+9hcPK1mXoJ9Jvp/ktpF3y5LnwF+sVYyCI
mIHeJyPw2iwagbCANFfImemmd8AnB0n+FEIeyyfxC6irCIeZnQSlA7n86ZZQ/QZP
OQnZ+0cfPrZwBGF+EnAIeunzzj1QsrjFQRxnkN4dAM1mLjFswwdz1kZqtWJGobuh
d9X9DZwcBwXr1aWOmfLRAGAxwlaM3Bf+cxtv9hHopt40bdtky8mm9azuLkne5EMZ
pg725ieS/9FaW1noCk4O5vwZ/GrCIklCotBTWqmuQTtwkv29DwHmdFvSJmaINQm5
VYQfZdT8Xv2f79UIRIEEJTD11uQjOJr9z7vwQWn3mhbXSvYGgHZNhi67+8vTd5Q9
KODfAc557oWbDyEdVngnmpYmiP8LbmATpPkaIqdBzWHeldZ5J7DB+rOSoASxaNvJ
PAJUZd000OgT/P9WgyMeBnIzNCv1A6kMjNhPO5QN41Dcm4/LTxqF0K7B2VCXs5sK
f1cNSdJiLKV4XVT+D5FQ0i7RtcxUISuE/fNPPdN9oy4lLUe2n9njDmXRdzya1BLv
jg7jINNFEgu8nMjJexONc6+WTX64duUyyJrF/ZCO4fbV/vwpdg5XAkMmCeGFmwRi
Pp1ICYewM8jnSUHV6PsXrYzQ4gY2ciRbzwTnjawjCJNBzQ+2yducxtAqYpdKEebc
TGnkb+Y1KHy9B4FwmLqS++fioQWQkkr6gpYSU9sqDiD7z6J6LMsMmkNFKvS1EIx1
KXE5LT77OAo+qunCHMNJ8SOkIippn1QjV4gOW6eKfqRkcp3KOndkasn6BoBDePa2
g9eOcWcYFX2pCVwXVwtpNfauywPzCmUYxCFrGcGipyvwalCUT4d40pQAm1nYpwif
45MpV3FsZD3CUXZLdfmMiX7DlPHpR+A6qNows+AV7psyT32ykALlnUJxK2kS5de0
d4aSX2DdtXB260741pfIvvE6L2rKX81AVi618oJ6RXGOvY9lt59OuAnMoT2iWFe3
Amy81OtS91FKhT5MY46DatAIKg+B/cv6x2aDyVcOpjIz6lOf5s/C9t6J86W3L7IX
bnMff/xKTofqikUZMLx27zvLKNDrqjgtd7yhQLs/RkzSCbieX7iUiK+Zj9STN/52
qTZqo9ZrtF9oQkVoRAqvC7ayl0c46cmdQO6rHepRPLNjcz7C5GwcJMxf0FCELHqf
GgaSEiIn28C+F/nc5gJu+q6DuRln8RhlJZBx4T+3ZqkbgDu7MZVNv2IrCihgUY6B
M6eD2zTYpFSGXHs4VCDHtzKAMxZYU1mRQz5R3QX9p4KyLtUpxPouOADK0szEwXK4
FHbEJe1sxC03QHiZugHN2uiOo+FDuKZueTzF2W7/9SMdFkPerKvgdxds1gUf1k3r
oI7utyy+ChyqdHYf7QSwuBk+CIQqT6sCizzbIXOVswVZMpvYsnPhX+TskK81rMct
cy/Jp12Uead/r1ZEwT4nBG43ypjuJ6I+N38AaJNqKtnpXsIpIZrEXxFSZOj9uWqv
m8dBMuGmuuvqmW0vFW9aklx/BFnK95n4XdzvyiQarU3AbIStxu75vlk2ULilFWNF
u0GRTRKqBNArV89vkGSrRrhn0ab780RXhp/x6t2EZN8O7vfZvCdDzrrlWL2TEBne
x4UKXG5TP3U1K8fzHjTrDQ860CQ17dGoh3ogV9rGwykRjVpaXSLGVZFjtzb1utxe
2t+mmhFGWf0NYNdgrF+PB5iiq8LVmXBst2KkWeNJAB4fi8yc+IEp5aaa8wdu+uRf
/ORcXOjKanEpVsxczuOZKbZ3f/770yYdCTPADOY0EqeghWXCtpcB1DdF1RVHJU2m
cgYA0eT4SrMMZnTbIX/ZS/33TOeZLdbLcJ2WyUQ3Y2i11FAhUzOdd/M+R4f42VUI
uiuFDaIV7LO+VCiTohIuIbZPmrXwAiVELko2JsqycfTzhsspJkhF8jBw2JGDVlVn
IENcA2Nq8SbjoKitwYyHTIob73VwsBts1qqDZ1VoPsiDFt3L3pvf0LxnKMeIQnzA
+7GBOqcqJ5OeDLpNLuJusHwhkNZkh902M6DOMnCSkqKk/gGjPRTfWnXPIjIJbuim
l2himtgeuYDZISA7kWpUQcq9kWDAy+rXBtD36UMoviiYBMO/r11Imn0EDFCY5LLq
i5zPODEWJpCPbUnxGaoWHA+INB5SY7CtQ8ryXuJas92V6olcjvth6aWv+4Na30FY
RK2Egv/9/WuFqQlkHcmFw8lLLJeWYPYv1RzwsDSWBT2sNqxvG6GGB8Ggl//3rDCn
HM/yptGTUpjmyaYsdYSluPYwPr5EoeSLEe+P0mJSB7k7OZpOlj83wbNedCDgC5bw
3ljiNvOns0eWpWTS1Lb22mEFsZiLZ4I7sj3zfO1CziZGB00t48eks1VZaE0ufeXy
gyp4a+2j/rHs2F0Nxn0riUILndGodwAw0mFAH1ay8kREaPFlVVEwcFu6I/QwNIYq
J6atOZcuMpKvU0jspmSAbE3Aae53Q2go3J8+r32wyJijh0X44fxBZdFqtWwZdn1U
hy4YXTQcf3KuORvrA5QkyJa0WpMMQponUl+d7GWPgxsgPt91HiTkG8QCf1B+h8Gx
dnV6g0Bqfv3K/oTW8jrcK7k7qOHxKhZIM10gHbfWC2noZ+qgtBeLI6vZIwnXPsdz
ZZXjHhV9ViqMbCx8VKWD6MXV5JojN+C97/eMlTwi0w/K/lsygLsAXcfAa/NaDVqs
69qT615T/ywCAzB4hQHgdrZd7bkAOZ30CURnpA+jtv6rxHNyY8dGBvtSPQfhnNNb
l1TvWh3gKghJDJkuwT3GZ3/Pnx6deomC0tJCEVKh/URXtqaLKTYEyYast1Cw6abe
VRbqjmneprga2Ipt8eYN/EXvwJYMDePYbRTwRTpgKWoq2eiJ3DjZdx7Ig6+W5K/0
YtToxTzqbne2xlxl1JdTjvtlDexYyR/KbuV2TCY4r5i2wdz6gOK9Q5KiyRYSJZY6
RB9db8cZRPeqxE+aRcarNKx5iahoS7XywQ7CA5AoF5K9/R5MpEOQZkg3kYxsFvJk
LD28hg8FFh4LJtLJyvAMtRRIfsAgmd4XVIxJPCsTeZryp65uTe8r3aXnxGaD8JZb
HPLo4E5lO29bhXNBEBMdRa5+SAfnkDe0v6pCvPymz27nwy0MVTXeQ5+UleotZPOl
V1oxYMsvKmQvkREsFKJQzqOYMlcQnfCpSF2hDXJS3asP8J9GSH3+XJN+HHxyVpbq
7ZPUvSfimrbkSo5TGIm/Xna33aWA+k/ks30DZY7cPt8FRTXkdz8cc5IYIGEflWuV
ofAhYljMG78xhpExJquySEZHQQLG2Hc2SE0Wn0hUW4/8MQvvYBDHdaFnyekybpyA
3fqqOgFoLRDvwfep2eVczs+7x2XeKVd9v/Gz8YIgt9EV2a5CTOGKCSuY98P8VJcg
Tke45An7EzAvyHE0W4falhczgpsUDuMVek3SG2jgTqB/mlwOFyVjBp8lrP1zxyGO
Q4FaAbyKBswZ2Qeb2NbjMt5igLXcVCbpLjVo5bqTApeP5xRuQYv1Odned46AToDT
K+VcXpe6wL+kKx/l1BLN0crDnRO4R9S3pjXVABI+R3n3SpEje77f5OdxVBHD4IPO
CMGZ+7av4lZyGrFmodjdyea5l84ekS4zmzcMVZ8E14WOszfqF2rZfXaoADxLs/u/
mdustJ/zJ2suSS8XrifKP4l9Kfvj6jgImrAx5REaYdA6YA2biHUP8bjJA/NNbvNA
PNpcOt34/J2iKvDPKYCtj5Wm1jFWSppYBaTjFF21Gb6dNWxE0prUsWc8G4vG9KDL
ZXEqPXXgxuZ+xFkAsBhD1QJoKvcsX4DpBCr5/qLQvnbGV9ueDScBcbQ4B1fpPCxi
iDKp3ZYY7Z76z+xhtjKpxjW/9XyMq9OMWbldnOADxmnI3BHgPVM6TMgoh+gILB5b
VSvD2kniApEWqDmSZ4qt0tmLLU+WTb9K5u28kcP3iSfSshiMcn6MmYhvbEd52t52
PlH3TNV6GdLF97HBB+bfYCy0+5wfutLuGb/MbLGZhfLmAx29lV0CsRtK3+pKOEOz
7fqNLbyC9s4bybtBucOdLlm1cCLn0AXUvd3HarvzzSRjTljtph7hHWboILjXQSEo
u0ZTL09DdBoL1GsB/9WmENIHLOi80aP4U36ckbYPa/FJ3vxycahBMHtX/hiIhgWY
R1pNy6i2hMSm1fDK0vpqwgKdWD5ciVG+/qp5MLn1DVzxkcRmPtTo3P60Hcj/n01S
gaTFb2wHdZaEu9LLxSvhG5d6wDasOx7ikwcweAynpbAk3/Y2Pfkl4k5omPj/FfLh
Zq9Cq/EJcFr6NI1f1RJe5j1nFQu2/KJ6CDRI2CCWhrbCrTs/HJOtXcOq09ARhkAN
oGLhYeDCVW03ZS68uRThox+OX2qk6u2ZHAnK0O4U7upQKwEKhw1WiN6i2RvfMwAT
OY68PP5J52YI7kkcB6xC9Rghad2EWkvTyloO/lCf6JHM3K2i3/fRZWdmh/Rx00nC
ljhNBPTdGZPiNmbC4BnYRlYU8klWP8rt1PqrH9C2/50c7yqk05rYxK7hnRu2PykY
NBXBtKUV9tGfAbQdz07j71yiLO7bvdHlBZOo5Lq7viWPVtAfWClUjS8d0YQGETU0
oVxVXLm5/DcH17D4JgYazkw0kFE4QwcXCyt3/ybbT6igfYHU/WpZS/PR4OkfRxk3
xLm+dqo+y9b+qh+6Yy08CVKUe6sV7TlzjnWEb2okLesYnUpsaXXrGFpO24yuc09q
sQFqf4dp/VQBj8rVero6gqTcMOhCzqmRFUxw12QYHZkXAfAhxjfwbXP0NRyBF6Tv
ZwdpNwr0PfGJEW6ikwqhJgzzZGKaOEp3A2gYKC1Q+2XDQOmex9LPP3Qx/DYJtiRF
573EugycfgdXyhzfVoiDBcNnHoOpm43nBOrtjS44+bucvJBXnyV+WxtnYx740tlV
VhUPCzXgLpL3bpnlPsCOdZ/W5HbR/bSKdgrSyUefjZya0w0nl5LehuQ+tNQjb55d
pu+CuUoAl+fPQz4eVO2zsw74KConBh/O3vWtDwQxeEDc4ZVRAPYIGNMG+PVu8oop
BhzquEvmrUrqczYpTHOjcvnVPFOZmUqUDV1Cb0EpZPbu4aO9Hpmmgq+Lo3+cjyzE
DDHRWWk4PVvvrJT+FCUpxUX0JKacgXpi5Jk7/ebLzAloOGjMemJRrLRFY8BMCLaS
CTu/IRl0YOAmAbksyF6c3SRaWMkZkIoqgM+gi9DI89mStaM12WLcx6m2ALBXxqI0
SDY7pdr91Lyy29c0K2idswlsj/06IhPtglt8MfqzR2ms2VWur3YnQtzv/YzsjpBu
RYriZaunUhOi+O315Jmy9jxsPCrR4TF0+B/dPk8TZBVf3UWokTjBCJ05YhAn2E6e
arYCvWjctMsorcTyt0I4V/6FNFxYC2nxxlGGMTpEV5OJhqi6tWwaRNjCk7LyemXR
5iLy16DJGgkeDhvBpQWz61+vJjBSBd3jn0ewvyJaicTSdEdXEAbNH4vH9Fi1Qmdz
hTlBo4gWZ4suSHi6uovnGTnpr0yygbA0nz2g2NwLv7z68uma4miO5yoMTforghKo
6vNKrGO3O1VBDD7WQl1sNX8z3/RvobCNPW/j8/Bq6l01ynRvGVYYM523gQUr1ztD
pbrAssDtd3dVknFedEexEEgK9siTMwc9H0EtPgi+oTr3H9Eb6uNfB68W2cs3HvkT
aFR1k8uWHcGAjBXq3E1GAFDdnCIAtWzdVmEQiLMu2AFm5+KSjQMCsstiAsdPTs4q
l9SkNiEpfgjzD0g6zewW8Se0jxabBQ47Zp94o3wnUZgjA3qEwhJ21OcI5qzWU/Df
IgEJGvcelK7DmHtQPRVtpI5yO7bAoiuxvtRcxOritDI2WAaYs6E9y8JkZqTI2HZq
xuUwFdGa0Rh6NZATLApTcNXZDewNIYeavKXlvbNGO0msmE1crkCe4GTvfeGvZ17O
+FgDxo7pEUGcwwVlSvf5vf9VNfwG+GTusHfoMUPoJoWtJLn0v2Cl8sVZceApJ7zL
14tIN8tUOQ7Mjp2ROjBWPYWIYlLOpgnzPFwIZ2Y6hW9jZ0IiXFvwIg5xDZo+n0sV
3y9kfe8gSC/wy3QCiM+0k/BYxa2WIFiNTgnGesBSLR+3PhvvyRq60whzsqAIPO3C
+kdC1NtAFySlygblmT2epIyJvnhLdSJi86h8yK47jPoA/xelkLyZRJa4jJz5BmT4
brxEHiimiODPbqaCblefRL4EDqNqGU+TKexn37jUT4a2HmWbBJ9deypElXg1X5lz
AcfGIVElj6M+/nhozniwPNovg77uuc1KFgcCTAohlBH9lroNI64n2AFkuijxvshh
HqrURnra2SUsra4l/YEr/e9i3iw2ugPI2wTNeJk56GX0axsV1m03sEso5ghWvmla
hfOnvUcUG4q+bw+cRHdsv0UXJMl8rhRd4vYOVIKxupjIwAKuPNeuUCu+VBO/3Bfe
oNL/uM43cRmdSZ/8kfgo7eivG5E8NExxGXJ78pZA2mnl+jRD8VeC8lLnGDWKXjlY
qjErvY311jfEZBgZbZlgQYmgst3Q6mJOoGhfqFBN+0PoxM/bzjVNrfip+ICUEo+O
84cnyDgYrhDLOs1pXAgNmklAtuKvgk1R5ync28vQGqb6goayDAMhFoRS4Lnfu+A8
95/h+qFutA8uYF2kOnW5N3nflIaznD70OeGFK212Dm8R69zuopzHrvWvDTGMU9sp
ZoznWSSrbbWdFpUsL2MkN7JYKT1FeVZUQrYTaRRMzARCMlJ2LHJ5bP9qTY7D7R6C
w25hRU47y0diYZ8xcEqo/A+FUctCpLYXQqcI1x3yARD8KG5aqctd7WMpJjIH1V2m
4cMJOVi/+txur2JHzgej+uXsxQ5Z1wWHzbWawb2+FL8n0VWagNGMvVWQwt0SxU6e
f0Z07v5lrNvgKPCsXCd2sAwPwjQBI0WZ/J4dDLg30wPY5HiiPmTAsHYxzKHYmj2e
K6rg9yK0acHJGs4Dg1nPW8M0hBWh2ZwGmDkk8u4KMkXSe/UqtsNyYwQfhHOKqi43
ap1WdKqRi6SzKODOQ48Nz5OPqcr9zGKpuhcfvwXvscYaYKJ/oBrCWoTRBpiFpyZ7
dgkFNa1Lf6IBJcxSDMHc1WbjdYWr13lwyUN+bpRGVpv4hsTGEiAakxL1lyaB2Tnj
4nwrd97Hs7pcC4vcuBtDRIfz5aCcjd0qHw1IQvbHEbukZu2ar7hIu4gKDotMqMoH
O3uPgbc67/KR0nGoy7Dzlob1fknXeX3q4B61CMz5UYdp7SbqL7ba1HRNClcJmJSF
sukN3lLw8Pm+HPhH4lFeZD+4uyiFu/XuBtrbq82+BBeretlzImqwVr83+5vyck+b
mYOKadj5UxtxT9SZ9GlLPaTMew+HN3r5S/8XMO5ww1E3m3hg7nvC+6BCvKj8yMTC
qKkaOFLe0Jzvf1a4vEKYdsTl9dLVQ6v+aMwLSqNKn6jPDzTsM1Doak3N/a1cMjFo
aJK1vCSkjjnBLbCgMC/i9pQ222gJ9xgOKyPEHHZ41wmJ3JvkifeSuSxIUYbF5gfy
a3fgqRBpbrdr39fCHd9vJgD3xHZv8fVzJBPyrB1DJF9+6w2un17UtBUN0waSxBBG
NNqC0vfAbVZk7HUTRhnCJgwxYqPJUSf6aiLqbF9kICYmtkjhQWjaJ45p+8VKjEkE
nNwH++UWZTxO65mJ2HVAjcf64ZV2OFVG/a8jL8xdR5CBPdKRtRheJ2IncYk1sjS1
YidbpvPoaqQW7eipLMMgYfJsPq7wMxidxbbaB7WqUGiaP1XlmjaKLrYSPLdIgGud
tVxbZHe4LI6rSkCHIpE7b6N8Zp9qnEXROmfMg27+xsgwNgow2+gqEjlZXECVCK3B
JeFBJlytdSlaVE8KWkaiMO5e4A+eQDVGTbnXqYuN03bt7w68flYLwRSfgY3FJkui
K4cx2O+/t/yIngaINzWJxQoD2zhDUl7x/7u3MuJQQ4PHMmNFdQU2zCjqnPLTLDJU
kpzpEYhko+sGzuZL7H+8gptsptjU15XT7Q0i+gIxfjU53wLW5huplGKWfXto3scN
C5zF391D9YffiVEi7NDSiNpu587uSn8shy96qKal7+/OoFdM4EQ7Ny/K2G4AQaza
eaBPfSzVLEYGp+8Fn2uMf9lP7SoHopXm/3VYTvgvDgUQl4kA6KEkQ+RzC8nZBVgp
0BEG4oZjdmk3OLqnzGx1xnTBmQKhynCBeg9XOTbaWag8NbLwj+drmQmxxuzTlCk/
0BIJaRZ9fnHQtBogcgljpH1BnIstfYSSqckja69t5ibSn47fdCqYF6xyWVw0VPgV
djbqgyHUkOE039P1IJ9B03CTop3PPl8v61DoiY2vwqIUwSO+/hxDBEbDN1S1GSM/
aIMl6yKRKwZQuMrAbxM2aceY2pTRNsoGyk3XdS1oDLmA2GggoQ4YhqLkVSyS/TnS
B3W00uR/4pzZXIBT16jczXbHjyiSJsQuGc7Eh5nGuBONaSbn9OotZRK/bI/q2pTg
NE/FQQLT0n4bx57gxyL/bD8+9bzmwAxylSzNDw1pvDtOSJpxghgH21lXyc66Glbl
9HKRbl6/U7jryF274hulCcbRnxGWjy1XVBWMkCNxJFm+sBpDmjOShF0ZMuXC30xA
gaJf77m4ksUiUfM21YbCAlRptYwWa9RGu3aHmCYTJEOF26UTsHiY/g/RTD4GyS6k
s+MBzYldyZ5jt9c44dmlsyI5+VeVGscJ1UsqWsy3wek0/59VHdnTiSbyXhchAyxs
bpaHsUH83XLPNlSYRAstXGfoONF0SKsC1QVjqr2iLhBs+RhBfKkAXqcC1UbK+oTP
SMZAt4VD7PdKbY2Ku77BDtWca64xsLSPviQu1PbsNW3vnQMpWej3ri44aJKmDUJ5
JCIwRwM+2faUX/kfUp0O4scTp3M8L6v6Rl536s1jkCwyTXPYKR6+0TY6Xl3NXrXa
GVuFKrLUmtSxixQfPxAmtGa8lVjW1tiJnAlhfN/iqEqO288IBaPbtK/zycx69NIO
Dsqm5s8otbQSjqIRGAfA8WgzsDlUK7zk8+GamJLjmDzFAs6lchVYI/Xrw8Jez7YC
YnlZRmrBEtHMM+RMlnC9eyRNnBMPLLeZnpavE0T6rPGkWnJ7bf2n0HIqA0YRxbIn
QAdfvtLeSpGvVZpVhrrLSqA1R5rprBGgpq4lgvN0Qkyx/zkJGe7ImYIsNA0QiBl4
VrFcChrnWPqoKhlvhzVCSsse8I/KPN1IkUKarqkRnId5Lu3t122UumdWVII9H4uc
au2iZrnF+c6nZpJuszQsm8F1MBkUi+N+1RD8mto9XBecxqs57CXzdm5+BMyuU72S
QvdRb9obIzKquoCzMd0rnlG3NHa+46Ca8jTFcQQ9B763IFW0WcWkmJI0WLxUzzov
TRQRDSLmtrGai716EQZKGvtS5aPIbmxD/ihQor6daERqpQ2S210DHjS0FCL1CZmA
Q5Ia8Xz2iE2PWWkidweL8uXeEC83MrB6e0iZQ7P1YM9gZtL/6r1o5ik88q1NXSIL
8hOSak1I5OitWJy6bV9M4RvAlavwd1OazQdij0lB7K0JoC5fDpHn8yyKLAb1ksMQ
VxVP0LwAAS6j8ijzMZGf9oVlBV5qU1fv5JCyvDhbUE+OQiE0dDJ1GpGxhW6WrdT2
LzDCov0N+Ymxyr7qq0eSRlzBC21uurrOHaxrGfUj6s9I0YFAg6a7B27x2h+hilj3
GGboQw9AFyfqf4SPI24NS/pRO/G4dFMSEp8IoegKJQmbNHEVoUHZjnESXejZoOZj
hQ6IaP170xFcL7hcy2rS39rJg3kVKxyASNK6IYE2hbkgbcBui7I3lJqztszF3EsU
mjBy5iBt0SbRPABF6ABVkIn9IoBhCfYCvIqQhkw/n+srlBOOMoUV0lbjY4ACYOeG
Kmz/agXnnmXFzwuSYBFhOG+QPNT/sfgDTHIQhO1yi9qDSjer/4cZSbLt8N6ywu9H
xtS7mEPlskRVpbtiVV5ANyt/IFY9pAEtBAMk/CT4zBfJf5wD6M69FNW4S/dfUDJG
U9a1+ux1cbtI/HlxO5GFdElLGuIJuw+zLslaTakQ4ETdUMjw8dHMFlydYrVGGwZg
Ijs10Mg/C2j+XmOeZrpcrRn4ZSxkPBg52DbBloLKO3SK4x7cTXNaLhae0Bg+azB5
5rZWwBoGqmXjzI0er3vTk36OZVQRCs5GsdK1+bgk34wYcEx8GTXjkrP3meCXo9LM
v/6MrBk/83j0eroZiD1KndB0w6TyIsWK2xqC5/o2lBRL1eggwIJdMEXJwrOcE3T5
Kl/1z8txWaVUXwHenPwA+sQoY6fQJAZ8buBDVygd6K7zDNOEh8YjQ8Ly1LyFdlKZ
YqO0zGXQyOO5+oDHwIj+qWZE+TOiRkB6DQGzJa6kBm7I/3hUXDuYOzXIMqJ/COBw
1174nd91NBWtA/KQZNfEPU43rsGaQRfclROtSZHUlzlc8lPK6Fz1PcLtCT0J4z/h
dVU9HLkkDNvP+q3/XHgQtrR5fgq6bEyZd7VyGMJadtr0lt1vqJxcUbZvjIWuYHOG
FFyIDKgAKhK6xxYhsssMYPWtzv/H36ZHWoTXdJXEbm8MUD+fy9e2mBEgqMD//D6W
XE+//14RN4P4slp2++a+rscdRWhMPZEaWOeZ0r0phni9eJeFc5YB2QXcrKvWM6jp
lfvWXDrkPt/KN5PvZGPOE5Tzeez/7o+egLBc0q2F6VL0vzXTqQr/LWAdBmnkCve3
N5tP6e1gcRPJeSzxtaA7SlhdlPmY730IWar8pCVFX08QOIPv4iwuWzQPBsm5n2r3
cKPZL6FP9s9wzIe8teu32x9ZQd0EvCWCWdEwkS5ZAXckqT8/o9YyiHAeIP9W7KsB
6eWQteLD5OzlcP85jVH68fLEYnym4Xzztb/EnIcWLi4WAXokziSTn6uktHRmMRHF
j8Sp8s9J1krnilIMvbIFHaw4jnGLHKPPSZ5f1DVt6Dd6DYH7Qy05JqYypPPvEqjx
mUaRRZRvltUGeZo3eFx9jcFDOHbInQ2WUPi8H9GttCSImCIa4X9NTCOBUEpak0ZK
r7whB5J3udOs6DViqfMVDfWjhSOhYQQlA+b1lDteOYw3rfw3Cvr3YaRaA1iJJsSf
+wVjDg21l20DZBz3TrlreKlt5FDjbV5V6PWjvmVOFLMqF6r0NJEDlYlm1pJS54SX
+d1eVYWLi2s3PR+LznY1s032xs5ZGNcLxa2mkwwb3QqaGI19iO/ReErmCwsU2JUc
RQNPN7Vzkqk1WORRiD4XZaegji+rUnI36gllBGWvKUU4wHhR07a7USFeFQFEPCWV
LU0YoIHScDh+9c2LNWcDbi4Xr7zdipwPDlV9ZiV1b7OwW7MFIxc5nCNrAnsFrz05
muO2UrPZsys5ahbQCJ8BLgzHQ9vRCXnzV/sjo4/CzXr3DhZ0iSlaHpKesWEJlTnF
kUxVyxFRqapap33CkObr44JYWUCMTcQWzGlfam5Heq74V21knCwvd0jvnA5fXT9S
MXj8Qs9Q81bbmf82l06EFCUnylAnth0raES+MyPbbWFdxe5cLDVAYSxFAzScZ3/4
NZXm7FvCwA+ptUAh167nY52Awpw/ao2alvDjJQroqUCI17pLbrraW7MrhfL1ujvm
621+1xEaSEqepbweTEF/kvuxyozqw984whz70Ej2ZkyNAcoSryb7O7SB7I3BrRKd
C7H8ZM+o3Q+8eh3JfnQoHyPfCzcorpv2J8SuHNBImpxCqNH4d5MC2zA29oitw9iJ
QDePwreZ94hX4n7E758XT5Q1an7yCsUtchOQFfBQ6D56k2EUyA9Kj/l2nQYX66/3
8V2gtdoBE81zYHle52jiMAYinEsL0SBTB939/niVbYZJ1QRUdE8w3x2X7e2alPYU
k/wFDDKvM6gubpLtxdyIyavVOIuEQ7Z6eiBSir7kocJgDXE37ChGRL2wQWPlxtDH
+2FV9oF0SCw1kRB6ZaS5QNCJDu1fI4DYutTGbs37SLjzLF+Mt2HFv8vwJ53LRI4p
hHEXOE1T8FPpv1x+9CjFYZf+Z35fLIejQfAK7L/Yf9tjY+nYP6hXXugIz75gxcaz
gQB5K5BwJ4NS8VFQm8tCoKCjE8FoEC1YP8OVHKYchqGizCvhmgcz+p+iobFvj1HQ
LPA6rIKMolBTcovTGYwHO/vMBGJsUPEX/U74tscOj/M9kJrLS+6Z+5IJauqSSb7r
ac4mL0oDnG9v04BdkSBfI2l0QLiPOGxsjrStNu0RP0gG11iO9autL2IHCgogBiF2
BYp4PHadUDPIQqWTWVDhIQwMTzSM2zF3qj4lUL225oRH4gDXi9lNT04ISew1vA8Z
KO9pMF0oRbBMIO5nPQDMmk87WEXnADY4ZP7LFqDRVDMKr9Vug14f7JmsA37Hh1Yn
T6FCV2zrTJlR946T9hERkkE/BsNWbRoX2L2OhBpAzwZCMbOtIZ94iBhh3Jq44E3C
IR8SqHrEGjGb3xQp8GInvTXWsqY5rgCY3klL274dI9fhnwoD0rT+bkMsWquG3rEK
9LjBD4t4d6Vvn5T9WyDB+iBkS39uvxLJqjOcx3dmkhp/ZiEKP1cNxBGnsuqJ32jW
YDBrrrXvf6G0o1NV1X37Qeq/aiO2aU1Bqk0ixUYsIcakTWz7GT5P40BULty/QOEo
sWjA8XJTsOL1zA4VrySBjAL/qdr4cENfz7l9xLxOvl8RF43X9o/wZhukbxm2inRn
UTwmmUZ6kmnBpZEl+W+Krv+s1RFsSX5zUSvd39nVL5p/VImQMoP3swUjse8MRSEI
4TcQ9aL3zXu+DoiyLc25F0kvtk9XQ0+kb8qdJICjS79Qb/dr1HPzQ2Izf8s5qc9b
3+Ia2WmNoKWZYqyIrqckaS68QVZq12pkMK3c2JwFjqVEeBJu6LFWGpL8vbjn2SZj
++unaP+ppscvMiRDvn9BpvhN50KLgz1tAKO9QOtgbsjuEg+/E0KiyuuCz42cE3jQ
WGTcWIMdGuxoVxmq0ZvZzUoEZUMJMmz5ueKlipC57TIi3vIppAQxjcmqC4/7BIiD
UdJdueHz8I24CvY4HXCqdQt7UyXiBB3PuYhV5QZm2f4JMisAyK2W3LIFeIeOy8Qc
Lq87xctT2BqbRFpotZul7PjNDqIKqdArXjfH0n9fCuW24oBRa33Jx86iY7SeyRFz
bd9g+2kpHddolInE3M96MsOwDBPmEinJJwCyL97fGkiaWdlRq6aysWX7S/DZ92ff
JK4/gG2I3/ZnaTZNBUUWkvAnmOaw/OQafVJDg8YHn7USklPT5pc2wga2jZoswC+K
KDr2H/dBB7MyXloAGVyENcEBLPWaIUSRPkVCyxbUMsWTeP931zCRDu6vvhxciA0Q
MTmXTP77Z19zI3XRjS22iStaK8FYhK28LF0N1RsT6Oa4GnNoT+CQAtB8Q47H4xHG
s8NTSyRwLoJff3w9ey7Lif9fNfkLqGbP0qLWBxmgCZ+P/7qXxwnnuEuB6//ESwfc
aDeGiM1hoQJCovbCBNHWVm7AzASy/3qa55gjV/CHeR361JNWwKv+8ew7vqBbUGGV
K0nc4bArmydgc8yshoNhOmgk16Ea9w3qzWP0sotzVkGfVFxMDOc4Oy52lG3Ik7PS
y52YCrWkWuiVyxNV34F1ojyYLVzAagFMg7mlBYVJxHpqgTndzMwGwMlFHZNhPFfo
38TRbn5W9g0IprsN3GQhEk9lz1uRLmiI8zaOcKNX/Bo093xwoX5mSOyjvnlieWVp
xNI0gqHtMaV39op56UrLTB2oYpilryQb4zmPpo+zBZkNbyh9ejlWYgSt1jpxTsTT
ne/+SxleswQJ8umh5vLa4Na6a34iRRwuw3b+7uF1RZHTM01tFlb6F7wcePQnG4If
UP3JECudp+A5dUsZWjV9l1e56yDYAeyxUulg2+CQeioAlfP8+lBMnVcZ24QpUgf2
nSxGfHNTATHs9k0zj12Y3l5ec2AyCp5hc0ruF4mSJ3VeewqyRVYbJMXedV95J24F
Lx4DaZzWy2lra70IHhoGQRMQ4Fe5jfjmJMXtfzurS+S8kHXSFiGRNRoC5huobpp4
/IPkCSKP6N9AED3DdJLj64Hk3QEU683efc8uHCD/PTyPqYdHrd5XBuAu39EeCMxp
He+coolkVAeXW/dikp2ENbWcFqMqntEag1+qStKPT8IIks2hm461nqA3Db4Cmm1j
A9aD7t7/Adr8bj/g1wBOKVgbWBslw7Skc1G929ZuYH5RfzMFZvTY+36OmCTMx2VB
uTCmNByTbnu5Ih08SR55yxtg09sIMpwqr2k0szh3EvazC/f5IQ/kzCk6EOG7b1Hp
a2yzlMaMPx1UpiJgfnuTUSPVhrI+8P1BCE+lT6veAsZJmZ/stxrJHg1kh3SVKdWa
cSalKsDzjXoWwRVHW1AKMS+GkfNMCHuQOpznQ5kNThHmaru43MxLheRKRGeP8j40
NOAif+ZjEV4TKkwud8cJs647TVzltuA60DKEXiBkYXXz1ubGTvDVElIMgheNBDPL
2oSymsmWiVX4hDewAhPabU+G1ESOMtdgzwoXeGYgaUMPGfmydRJvRZhVZkwIQMsq
ToPtvyOKw7QsvWBWilMiW8zklF/ilW87k8u0ckOOJ2CGR8z5tcZccMO0pjNERS60
eCtG1DJiPDrB0GpTsKxcXJxyvs5GdEocXYHZKa6O3ExU/na5FrZRDgpQMwl5uYn8
A2xsxlU2gyxgj7gEAgHUoHYcBaePxt8tVLf4KMvOt54Rl6m45STCbpB3Ixls2y2q
7zvUPSmX2RLBv/58wXBYgRmVsV9wwM2HmxV+s2JozV2LdYBgWrj3S57eNV7BjQFt
Cru5XQ+fwlBnI/0xe81qW7zAvK5yElKRjeOdD2ugdedhxWrXsWEAWbc6FBz8VTre
jtH9qh9CN2mrK/xnKhYpQd/X9sKko16zKdKDzHhRBSl9LpHjLjgYqRSbwq3JZoPw
2LMPvmszObwP+4vCW1ETrlpmgXlWzws+/kiIaHU0y1GeCmT8cGmhZi25085yYr6d
vFNL1itmIxp2b2wVBYV+2sRlSySwiyBlgDdJku3y6BqCRh6jCBEAT29RLsawh6k9
vE8ie076tGs79QCXcREq/vmd4yy/IhV+QOmcXni6GCd/5GK3hAigOJbGnVcBKJgX
2VREIIWqdnWlR9dXzMv5kxn5G/y0G8+fWKz3Y4HIlyaQtT0yILAKqKmmThny6str
wXwOjp2Y03aUMJFZjJjnoFMDE7vKoFZVMwLmHgRouTbzTxuS3QeTi5yv6fdMkhFc
bkyjZXk0U2A0mNAlc1zbyTXhArHAYHcYpGp7ePiVnF7nGTs0bdAxTX5dXMvWSPmc
oieD8Y2LCndlAdtjT5w9kiiyCD/Db+7urJamuc93DnoGaVNbRe3Jc3u+EcNGTSII
L9lw8CIg4QfwBe59vXjrHwRSGDURcl5SkbXmJznvTzhTTYtnPRNrICcCIsC3CY3e
yzYGxgFTj+bPEAy7CdCQcQoQfmXJhJr/zASqywFmAolamw7Pj4eyYZ288eQ3RVDx
V08HmycuTA8v2cxh2ZPG7syrAQB9XMyYeeOh7YZXutbXPrr+zeZKdgJhV36Hfj7d
bG0tD3s+zAyTmmqV04OadcVj4Ma+xRS36Chg0YDlYOpatv0de5zsJa/6SN0TqsCc
YxuhHUjFu3qvzvyh2fEZutE0qEfVTbMd89UU7pXvDjxpHc3K4+MwsmyNIB/SnaMP
2592DWwJ/oMVf7wDSKmN57wwfJ8xnKxTKQCtWU+N8BimcnW1T0cX6nFQUXzC3DR/
YFngy2k7CcJCO3P0q0xWZIvVWhuoyhHFhgJyAEzdOJ4AcPMbEDynWFDgHj/tU+xj
aea9TSfhA1kFJI/D6BwMzd17dpzvW6igrOu82xRklIOe2NL3aOQebipRxhxwS2WF
1GeFwGgiPAg77x//kE9sLSD7I/YehJkg5itT3Nlz9lb0otgVGoxP7id7r0ywuWpr
AfIKA1LBCOmE4EBT+akOV6fgCvLWNrJraarb8l9W0EO52kZdIQ5x6ViIjlH4VbYr
gqewSa4QXglujf8Tj+7SKLQ7wLPKAixo2BFHUHC8CgpKrMzy2PuAX8mJbgVHmrWt
k4Y66DcTLpRPISMPrQ9cqEBehQp8YGHicStaxZ0w9sXgLp5cByjn4jgkGikqqhYg
eChEvyRLoCvJjh+dEOEl7gQWixvHRN5mhHJqjdV6rC05FGwl93xtovQqSWRAKOr9
O2JYG2fQZh1ReiXekSyB7DmGU6P4LrsZ0xUcFfOJIQT1vQCDBKBetE4MW8aR00ao
JKvzrK6/2oc6cHy0bA94ce+RMBWINu+Af3Jk58WsRbMD73v6PSbcX+2EIxWNL/dF
K8hNanXbt/MZfejHSIsRBwZ52lc0yFjvzF0zBdlnET8RV9BB/SnrU06x/mg42fI2
OsoTf0R3fjI16cRzfVd/WosvGjk3nxxn4o/ihsY9+dqcE4gBiQnwvPc4mGEc6lNj
aQtEwOLfr4Z+g9kp0BQVb2icUH+UL/ZI/GUco2E0+xag8ehZrQ999ZmU77scmhnT
cV0zkGxxYtK+lT+jNlwE9HKVUA82QaPMydmRgruTFaVMJMF1MXKPi0rKQg/YPSu8
qWXjPV78KxAnBVfet1Kzz5BGWkm3lUP1RbGqA3DbIC8yONtRHp5GCJLbYDOKcbSa
T8NWGoZlnvipRqvOh1ZMmeHb6pYSDDyXHMqsDxXPTNrShH0UffqZMBYLz/E4Fc96
tzBvMRxUuyKxaQ8xGhPIEQ8Cg72TSwnaly3RXUh/KIw8zu8GjSWY0CgOvR7GNjLY
FqoiiLwK0lPV60W8HmqFsaxyrGSCJpAsc9ueZzYzmET1JbFqsRxFSYPqTyIC8Zix
GVuKjk92Fxk7Otru/IQT4F0j63Llab028mJWpFWPBprq96SQHZIR2XmLZjHeolLi
cXwfhzz7qJcYQcXdKyJJ5pyXvIjoOigf78cStdFz5C49lxxxNNhnU7HC3lAH0FCE
eqdxvZWeyqLLDPtmqUdZgmmewDRqjd6Gary64GpPkzHYFqZCUcjKiigpY/lhQNTP
Ytr+Ir3x0D3onqh7b8KeMKLRtUBFNZh33Fqw1uP9C8jtHgMkeaMu8fwa0LUewcpK
idRXCvOnNnFb1TyWslSq8bDtEOQXzJJ85Gy17vYPc7XSRe4H12EtapQGEPo8fQ3I
g5+CC5TJZmt1QV+fYc+Ea+Pr9oFa7jLF9V3yZa9hQ8Zi/SBvExVEzIvgf3P6WiO6
Ysvle1MJT+QQyxYJqPvGPudQmzmW8Rnp3/q/qc0gMM7tlacV6raM9m3R3vjHLohQ
o/CKnTcYhcRuplp0qwkr7vPx7X5pcUdi8Az4+xFPxVLNn3QZhd4wcsLxaZIqVZX5
yydiLxgsdVh6wRdYyuNG4dip2XyDuZPm8GL75V30jyJP0RSJcydIRKIIuWQGPspN
fi/q+qkn3NMLiTrt2MEU+fAdNrS/TlCtBLv0SmIJMRRyyqonvYT/nwEiE8KV+ew9
RkkGA7MDHmdurVEYoTwYQ4bW8FCtI+enFLOOA/fX7flIMgkDCsC0s3Pyj7Jtn2DA
KE0UbaGSRL/5AIu7GuL51aoxTYQqB6BhOYOuYUJR/+LBpRYGzpXB58tJ7ZT3ac8S
xTGiCBxL7Ayw+reCm1LMxJlppm0ET9kSF/DCmrSgVqtaDFyA18ceRxNAxxtM7iIt
MWf6tjfg/3IKA9xwimV/OrRqEFQxLMyhPjmxKfIf0LpUYWnj7ShpdyGLK+HWnU6t
U8tgSMGBY0rh2QuW6OBGLcD3v5a6gNmXuOll+tdfzSOVSuyJiYXQqzIY4C+0abUf
S67yNVQvCZ8bkRhIPv/D0X4OkS6lTGdjddYBnR/8tky4nxfl8rG3pjFyuqas94LV
fNWZKljk07R3LtLB2Ym1Gbf70kheTTzDTyDZq3JwXvFUugw2kIQoZLi694CYkUJq
bvWqe7xqyqTbz89peSxFSTOgS88mc5hZTJptLyUJ1FUZQ+dcgI+KIj91GC0WrA1w
q4A5/SVSzTk6H9wNMdbl/yynCLDwk7ZYQT0PFJ2zDjSyDoGd8DYct4iwjLmTsY9l
sSKyHu9e+41FTzDmypjFKkfzMq/ZIVNZErh0ArVw+pDiUD7FGx9+i66UasvTc1Vx
Ke1x5x/JtWyCDWRHq8Y2NWr9t0+ofU38b0n9tOjNUHU2VpeyDrQiF4UBk8bCqkg2
oQkfMqHE+2fRD9bU1TK8j1o9KiN75WfPVHr04A4R+SVzP0NHpvDfvP9hfDLVPSIQ
BTQlysAqkK2SuriOKi2vskQ5AY3oYNe1kuyNN6GaK3oszNgZNWs2jpv2qFhVTdjd
WkDTzx61Kggtu9MY7JGfCY+Qrmr8R0GaN6XvHjTYHywJK6xVAGhwUrW+WLc/PLFO
HTDEZ5ULOoPHGxcHwx4QlOBCygOsGn+7x9gnSVwr34KIlXWVnopcMufw38ZwyYkH
nYpHBdlgWJ8LPI2NRMiXjl04GZYUoa7cBL8Mg6EazjvV4zoeRUlAfMgBbt7/brSq
Os/fhyWYnvP9yq4d9PkEv0H5CSlDZSc00xe+3+9IywnmzDIwRuXnY+6RzZUPydZS
6URSk3dv3tJEi6eMREtOLE5UsUeU8+mmbpnDP8R6m5FTvHVK4YnZqsmyB1K405ui
BlVONe3YyfZjk0gym3an7O2L2theOFrqWS+x0LEFg/HB37SVgVX8Pmu36gUaVUia
3JBU+WnusQ2eNvpRcUzoVZ1l09dFFwn9S8NxJrirci23tbT3mJdn55smTGner5K3
74eSfwrl3nOVbjoXNb7YPseRgPZR1BlXyVelb4lTbnm5YYsfQwHRmfrNtlCG7Bwt
/p1aeHicWp3JXt29he59T8qQ78tuUbfCUUA3RVNH9f2tUMshlZdPhGP99gpvFezX
W7D34jsMDoDApcBHCys0OBcl4yP9eSlppviJnlpZeiRPYRZ+himmu3DQnFhl4BtV
8vTOX1vCedB5MmwSgLmcT+8n8TC+xeQnz17FwjgbYngp1AOgAgU2y0g0TQ4ZlZez
Zpx8D1jfRW9eHYJz30XoIwRUlKxD/feXykDaesagk2sPb4ItJsPuQeUV6HY/HZnE
My4pCPf02nqK1Na6HkkD1BfZcBUFzoJzZy28Q8FT05UCsnwYU7OMMYaYMwEW6f3I
inY/pwrantJoEQjROf8r5JzbBzGLZFmY6XN4o4hEsMKw4gIQgVcIo+3YFSBrZA7R
5R+wm7TAUN/MV0no7ztupsHD1Xsd33TeEcDy7SqYb396LYgJA8m4o/5w12KzmpEf
fwkWENIz2RtdVB3/hTgBogRQ3Yb7TIIMoQAGg5Ufx6NWiu+aHqsEFKjOfVgNC9En
OnKtKDl20zyn0sfXM9e4YvNXcvMOKvr4ueEG1V1imzEgpi40Z+xQF4pjvr4I/e2L
2c5ko5xRIP1aaXsPBA0tFb5/OHY1JX+nZ+lK8Mf3MBiQs3Fzp9CvxOjwC6HL85c3
gJTE4CnRZv4CHKHHkC4Qar/H/3RZXSlJguwkGSYXFypWCe2qroee943k4iMotNub
KgvG+C9w6qiIQVQAwjFoEDdrK8O93ZKLeMIvkp9Nyi0T1QNhNjzMjmTjH6+RXe6p
lQRfauAdTlpMOcMiRS+D+Z6OmUlcLF+ZX71FOBGvoai9OaUdoLvcd5Gx/Wbn+wEi
zvBA7jkaaXyAFwTe51DoBDG8D5rac+fPlVDdmOCfN1f6EVN9ACMwPEWNgiUvgLVn
EVEpLMWBtLzVC5UQlNnNNgEmZVgcWEy+ZxBHeWmz0oaGbIN6aosKIC/Tz651ynlE
Ag6VT5EbLnaC6tc8jP5CfNMfd2eOjqca3ABEfQNNuWxxqJMINzFjD35BdTKqpxlX
60Gaybgxu+MiGRDIL+dJDkMCXGUgVgVdNXi/nMeiHsbLycmbRr6++r0LRZFKZAMd
4yPY+avuv106z5od7nAGen8zc0WS6LJwv7fANfMuZpfniGne+jM3srB+4+S/z48/
rmP4TPuTOAySWdt3QKqRCKcwzV/wCwqZ8Ap1gasv66CcJMKipGanMuPX0E9tSaEb
1M5desz64C2z24zn13TZMzcJSfZ1hZF5TW5jBCUFeHivM5Jo5M5Jngz6nHTtxPCW
8/Ie8TrrBp96J8qyg6lbpIfxuZwqBQSI4p2iWjXR5flLdr/7I3oF7i9xacD83o++
YTiGl/G5Ali8V0wv1CMOzy53RQSRe0VVqgrksU87jmOPXOk0M6BpMvHfrlRJuLpB
ME4KO+QMp78Lqrh9kKhTTVOTKnyGiCaoAkdIWhBn2ju81rHW8oMV+DHeeD1Dyf+m
BISswicjOOT6ojf5IcpqWIY375PA7siP1hTr3ju7hD3mExwldATjJcLJDTohz5IR
F525xpJHugkyUH4OJ4saDqha/AARS69XBe2xtAaBTdwB40F8C9q2VNlJMomyyHsk
6eO5WgWyBap0FEsXtZA1aT1mjk28qFkWSI+O+WJBnDCTe4QCM8GgRGwQGc+fzGYX
6kFRcAOAknQSgw8yJkbXhKX6c+ZAIiBtdkONo54ZVHxg+EWV/PV50cOXTZh4eRme
qpSSb722H+Dh8doGrxXYKMICuBw9f/cBw4X0q0kVep8CDLnkECQscOn1rvXZ9sC0
zaSwmlQMF8nJNcV7Ro82/H0fsmpK8niMasym/L0QbRvW23hzb3rAlXWiis4WTZse
9wl/cbjGPnOWzxXkarAqGGp7dBPD37g4eT8GMU36Nl5SbmUB1AI5T1Q22vjs819O
20mayD+Eqnm2JDJMbqnjEnkEBopcPTiwE6zr6PWf/yXRrguhP4LleE14c/gMbEPh
JqRCCV9AzifYbATPNUw6CvHb9l+YVRGvuFUJjgVPQOMBP3k72YxWk3QYdy2mVxci
Y7xQH9OG9LDi4X9xLiY92WVjLhv0UrS9mDoOSESlcFW5pzaN9cWdF0NNeCVKOin0
DWeDWd5MQ3H42zX45loUBB4QiUWHH3OC+Tz/HCRFqZgweqe0uE0l5smHktpEtJCo
fslL/6Pm7lF12Fcq0yXZNNBXfYcrFwTrAvz5Lq+iGv7cUXePFJwgFzk/mE7nMLju
rfmnmRPLm4PWHKrRzHZZ9Fyg1xtIvL4977RKJKQIFG21K/GWxSadjyOt13iAYWFF
NAx+pYPhTh+fwd6de1XgCrkVMlfMcBwWMU8/xYSgA2TjcF6X9AUWynFAIZvPLFmH
Iz1Uv5alMc6nkmYbl1B/X82tZU4eIGCsAJPzXt++XJUTxqwdNxNYQZBSs2VVNGH1
FCiWhakAm9TT5qXuthtfiQR8/E29UQartZs67nPHwRyfpzIuajduK6aTbD8SYmvL
8UYAHHek09d0nET9DTo0kYQVmP3bkUamcSbJGzoi+kD6JIQaXK+9Spbk8oBhWIUc
X81oUMZe7e7KidjLwqAz2l4Cx0+1TzftATgZkItW6XEaunCgmr8AvbSS0rw5pD9i
3yGbhEtMfcN0PW4BPtYaWvWl/9W+QnyFaaa/JZRrSeGzTrqhsumH9LaCB9wFj4b+
6C8zVw1heQqIyJ1b+aFgfv9YzVtuT6D+oOoyCcuSluWTNQtpL5RKlbeBAfdXPafv
O+3t+VZ8nnklivOcrgHO7HuQ5YvlU3LFwkeHaBl7HpLQsjmPUdKy/lCFYTtas6RT
1ACNyk18O2s8ic04GPO6hbC/QVsRQAmS1y7GbML2nEl60Cqhg3Zi/2iXf/I3uZqP
UT+MqZB0uqDeU0EmWLNjwczFOijUCUsF314RuUQfmnzVlp6jFpRrsU++6ySgAnzK
b/2pgNgb3ZmclcUJwlst8vSt3pTmyUaylMSw0Npi8CoNwiTJtOF6JSFBV70YkAti
MZgBtYjB9bE27wepxplmrW/18+3HzTYRpjpXaF2xlSfXwW7U/DYHt/HkHiAsVmyL
rLk1oIdsG3NmEefJnS/8LiPh3J+wMx4Ka9Aw3ixxtrHMDMG6ed6xnBN0R5/jYLvJ
4pxA7/1mX3CzZ1jDZNjwViBSV+OPFDTwnkEu7jhiPSXZin596oJAhpkaPAE814XQ
lMAD0mHnNghUSVY5II7xpZTv0Tw5NyXEUFqewvgSolRg98EQkUQlZ+Xo8qD81R/V
+F3PTeED/xsk+526LxQVokJmE6OsvDc/Pg5oNcMIgcid37YYZzuSvObr3tmORVln
OiMlTm9Eo1AxsPxcCjjjFU6DpC3OoYTWTFu4S+Tf0RTKuwkoZGAV3ZxgDuT5QMGA
+m5dcSDRc5/sBN3+rMt6uL7X+vemeSYg+8JTeh0zhyQgtX5oBmcw1P3d82WadZub
FslM3JOIMJhBAUb4Lq75gKjM1gjX1ZgHXF++ixb9C9TAGSPibhlQ6x+BN3z/S9Hi
yV5uXrhqPzBlhJexwx0xs/2QPiLJOwWMV6CGmv+ylu1yj1XA4VDI906EJr5AE5Vn
+2lEm/S5+35Oq3cF9EVlvlQt7wjCYYFz6IDY/gJN3jCzym2YIxkrkco0QRUHnI1k
/VTD3UqoFXlLWs6O5Zbafv4GUCzlIHMgKK5DfBMgWJeTWFuItLhQCLBdqo6qkd/4
spzwFodOhdR5ZLS22ZpPdBwXppexfSR4qZpN7FOwJ7oXkchiWCke4j7TtSWJRHw1
GPrLaSXXFSn/gWfu7gPJJegdPc+BiqxraS/N/rjD+DH3huMVeTcEkSyI6U0kRaz+
Y+o95AadTd6QDif2ISUZxRvxhfAJ7Yi2piuae1uVVchS5Ditgg1OubnJertlVHmu
6+Y3xIPeTKvXxzkZorgoSoFcbjfnQ39/OgNLsXlxXtEvOQhkJE7/7QSd3ot3PPtO
u16yjBwYKBXVfIntwTGPQ9ZB5yGIVzicpicJPP6I+mSW7ZSVHdO747EzormKaMWP
D+Al0I9mFpbYikkBhbD6tNuqpJlt21Ojpd/IeDAKoNFC759wzygMY/hTtVQi2mdP
NmiA+gvMnpZDANBZ3/tSeKoMTTTpL1a2gblalGymVqFslDpE9yLORQZhNtdL/cS5
0lCBXPMR84m+Opj8u1iEpr/npsqn3B/wektWAzKrXp/dGhYUcXt7g9vec9v0bQwf
n5UO97Hc2UtwFZ9aN8idHXmek1sYtf2WUPOd23E1o5c5LYMKek/KeczTYyVZr7Fu
i5UVPFIJ2m4yvigNJJmrSAB51rYY1qSV/Tl9u3KdUPZn9fU9n6oEfnj460ORzA+O
tGCMpBKl43z/lFqECZV24oIz3kb55b/2hovx8/1T2PMc9PlKLAxCT9DHOBhoyo5l
mpohGCCLQT6t0WZvXaGYnardaFcCbF7VNcnygLsabBm4IH/MTgIOZ79Y0TcTu2vA
L1BZjyFLGSHk+FZoVCxcgKUPLdwgYt8LJlzhIAvJJctebu+VmfYjzp2ziaoOZX+6
JBk1NV5NRI6eOoE+97QzaAvT99wK/IlarjlXElS1YyGKfIdRAb1qMxrlhMuuoO15
IGhwynKtKbDgE4QcLHPpKYrsDKfvEeyboYgiW33xzn05loERZDk95Yz/vuvZMxuU
zNtwQ0ISYJe/7dyampw6RW8+MhLM0/rqNmiSbwfo5UviajtuZjLQmFqh6PKcg1pT
bjbmx8dTJJIf9sxgc0ZvsxjvuDDKGzUuOxD042Glt+YkSSPDppqokFCh+X0JXJTu
zBe9H8KCCXv42wTo3GS32bpyQhvARXN21GFFC6UyrhO98NwUiCIcJUf4dffrAJcD
J5GkB9n27VIcDgjJDgyauuJuc0Ame0uxtNRW2XW1IS2+Du4a0/BQ9xNfyxJoeigQ
/ZvfE81BvFv+Dk7E3fku1mt5VGJdlVIwOtH43FhPdw/DjsDMgCQXxXuvD//xngQU
1IUiQJgVU3H4HgzqiBcIg/gHOv+F1wGZHf/nsCtGWzG57I9DnY9HZkPpC2BdKIkO
K1DVpKk8N32hJQO3/Tq+C4xQAfHUXdMosv9qHpFzf9UYEV4EzN9cq539fMHH0U7i
qERNsecnFRJJQA4TwYx98FRjSfv2B+21w1Qz29MeDsiGLaxnoutLkFtLKsVpeoXU
dDCii6+OzrgpOGpKlJwUStapZ/7CscuegGvWJ2xfb33hYkHwKIgujPSYP655bGDy
udmwE7sZgwldu1KnlyBR21Y5BnUL6VYy+5X+Fh0flLNH5d6F0IXm4xE/ByudCMfM
id24dWHIMvEtonDh8sYAnsgH3p/xjo2SXYYn+f5VibG/OjuXw7corww8Fa+Rbv1j
1eu/tVgqgQJRPi8+KUMOn3kA8ke9WOHhe0bFKaO7gFa2+mDqjGz569CfjAvXEbUz
2zAuPzxPhPEKW+xCT0TC0sw6ArM/MD3sXy/5Mhdi7aY3axltnSO2TKcLwmvyVGkl
P9Ul4MBRbuJX8Di24BItta/frSzTwwSSxRYiPVnxzpnww0mS8k5Zo4f/pkfJAXg2
J+bHACrMmOaOWU1U8RzGXs5tmkWEv7w0db3Xbbkzq5aZ9kr4kDcWQT6yJy8Ws3/o
tr4phL9gssufjV3uvJWbtMojB+zTpkB9AoAq0X9o5pNvS8s1UsC/nyz3XOKWz2nP
gL8dChZl8C8i6F24xkPSQSUew3LmDvhAU6BlfbjHNoes9FKP6hVXd3PKBnFc6fqX
GRHkwieMgMQICotNYXOzA+UnzqHtjI/8YDN2oyRjRjTd+wbR2u46XCCQFN7FppeE
SnFbDrS7GJMWUy0Ar+XJQW9m7SNdyNaow3rERkLyaL+vEmhqlJulXCOmhJYkp++v
hT4sChX+oCrvNMlw0y6aqEvi3zicr/bbw1BVAo9khd+5zezspxz4Tl47duHvbKF0
YNlnfh1emZpw4utbVbongCWDppU4hgRDIUDZ3Ip1S2ASZJIMITLMjUXhaYgFbJtz
4L3JDs8fIOfwnxRt1SGQ7n/P6teTkMUJmzn0Bz/C9W6KSkfhPJ4abfvZyhZqSrMs
/JINwozFcZUP1e59c7p+TABNRNpw6IN1DfCj3IeeSKrxulaH9yODB5Q4yvE9zN9e
KfRZ+2aAjoFTaPXANrbSNcfIXk7uOv2bASiyUrDgLtAtERgFQhZwUlqrxJmcOfo2
GkdyBpSpmjGMbYP01RbzFINkY0/tlXPiWZkIfeJBBMqLn2nWzuxqRnS44AhcYApU
K9pvs87iPnzoE0HnXanNf9NjFDendAIQpVwplq0fOTm7wt5+hqfEwU6PFQhSbkIt
UTpAY+1qrsUh2EPL3SUDyoHiqjM6VSrENPXyY+fiGF7CsJdr8SZvX3aKkf5XwogR
GBW5A/DI1uqW41Q+4GwwX4QlpG21aVqq7BROaNfV0Bd8CWSxosDJh82txNyV3JU8
qkemgo3xKkDx/TvFrLsreCTWZU8OlrU9y+D8xaAV2Ao9sJglJcNQikR6L1YwNTGC
WELPy5EAAnRwNRdMPDrLVn6ZqYGI2yIBduKniZZVjb/ie5B9y1tCohrH6nVv56no
DF9aNoO2oNjU9cfzexLV81T2uvk2Jn+VIhdrOct8w5eE3uW5/5hDrqowM8yZhUph
A6grMUDU6ZsgUIhv6AkseIbvm0k+alpae4O2uCeODo6NjSGktghdGTfS7qXFADPV
uNxFocWxWPEp0rNwYzKuZIyMqKn6hHEQVemUW3YAdBQi4CwkNR6cPe3dgpj3TFOD
QJLrkbrJ8RXfovnA4qIH7avUIOwvynNvKB+cg05gDt1ybPAviPy7K3KN5nFAoGNU
gX7o6AuqziH+OGvgJawFS1gSYGfpTkBDE3mnG2Gxn2cXWbwjoB3eMvk4MkYPUNBb
McEWXHVarcucvVWUUWoI0prd3WYxlOE0jJ2NAJXtkr7lFmcBweBhxuvFxILoVKeC
0483T4ygH4tdakP2F2oDc5eO1cW86Y2ky8CgmVPa1U85HKqboRY8PbRSyO1NFOW6
jK9sjXloah+dWXfVJwKTp/pLjLnlh4sWe/9AmRrqGHPmgQSYrBTODnXXO0vzlSeM
7FV6FBP794jDSSw7qeXXK5hdSjGjOX8jW/REGU8i2D/nVi6AK6f0rk/f5aNo0pJk
dN799CJ8PvmXcICsPe1StgN1W6sJUA0BI0g2+OdAa7Xxm2Po8rG5q+dcR31w79c0
P4O7/cf+pnIihILluMnCY6Q8hZyrJWBeMiKikcVOv/dJQBvIjXqHRgSEJZkRLigr
r0oj7c6cwq7wF4mhF8nO5+eTlUyDNZHlGqhcEkaEktI/i9/guzUtsC3gUtJhkp0C
vRa5nO4g1K4xr5aZyvXDixRtskOSOj9k/7JkmsqhqPPDjoMffnQRdJoTRk7heMii
vm2F78ZYK9G7/sqpClRZaOxovlExWoiDbolDyy5vguZiM5Uc7VTlQiVKl/WXAqK5
AiOBOZJ8A6SSeQ2yhrNQbgQq99W4qxbnARG4JEfBjRGvEASK+yCd0zMQFNVskhT5
F4aUFn7/GOQiRy2pQlhs+Ha6sJjuXQGBvm/d9U6euE1ViV2UuNqxIIFA26zeT7dP
/alpV8mSBZF/YdKP8EtEgRs2mVNZ/4n/dRbfpekFCqf/myfJ4YL+ZPP1Q6yxwEFy
W3VZYpqO+By8NOgL2RUuUR7/+Hq4h9VhwDqD+DHf6C7Uxtz0JTPaEeDq1EkAOzaV
klboCmtr4dlwo5xvwIGdN5LKDecnkAg1PuK6f23ZUm1ZeZCWqbwWRDY5HhrwMCf1
yfxVdxNrQJ81bTfHdos0QVTytQPQaSvb8FwMD0Jmmps6WxFYr1RbgLq7VeKSnzgi
Dp+TGsl5JTCkGrvaLS2uITfubM+EX9/dM8HskoG7H6ORfDT3PhukF8+fiBlIIYu8
QGYpcXvXpQsLC2BUrruu+HYWSBfEKZA3tnX/IbJYh0+w8brg/1lysnJ9AGvClR3k
WtjGXRTBIkPGfUrrzsfm6at4Nje7Z9wroKibIT5TpNfCCf2juQL68vbN737XmgLx
rgHr88uFGC6Tjglo4VH9kj9cnSWPutmpAwFB0ihTpb5sv1D7GqCdDQLZMwVPEdMn
aasxF8sE6V1DTT6MkXELrr5t3zc1aoC/DEMZOFxuyMuHdS4fLRlYbVvyVn3EHuFn
/DN1i3dssgiwkgprVtEAr27GBII7AzBrP4eKzhcolmYdRSIGa4/m9tx/jfDGyonL
gG4sikCcJ0TZ7smSeLufq6CsQCulTAfeGBDpwAhUw7wmJdKOfiye/wBLG79D31BR
EiMjvi5p7O142N7E5r6BwlahPNyc1HCH+7c7DTYy6er47TUokEcRbKRLLmdgjdVp
tWYvGo4WvJT86CJaUM5TuxBT9ZiKz2aEHK+wYic6CJ/m2YZRuADyGQG1drPk5TJt
aA5VTjuG3VfXe754c62nl8rvwOYUiX79lj9hBoivlktIzpH3iGuZM/0cufZ/Vu4+
v5k2MVyaQ4mrtqH+QuOJACm6x7L0tfGRClwHtwFB2qPM7anwOsYMLUtkufs7ErCL
q1FdrYr9wgABWJBm0es5jlR+zQhLCLXekvTQo43dwyokwqk3AAVB0yAANEgmePTH
LceNgpDJJ51GH6pR4pl/l2Um1sTOYRp96i9Kxx0z4dA1pGL88Ha5d8zf0lnyk2Xc
Gg2BxYoUAJX0Ui3II+fjhofR7Lo0dA3vk8if9BJ9ngI5K+JIaCWQgbk9Kj73SFLD
Cgi2JS4H/Txwh8SehzFyysC0/pEYm6dYzi+F9t9EYubA/oeWmoOK0cJ2ufnU2V0N
A1+CHVopJL+c6kwntAH1vbFaORQi6Zqae+lfCYG2k5MsxuiMaUwMpltIFEugiY7q
2wSTXWk7UYSayUSBIN+uuKHmjQcijbBlyozPsjugl+iKvG/6f4lr1HYvhOtKc/xE
0FODBsms2fJ3dofeXCBH3N5IQKS7fUCxDiIG90229FQEFjDsPQgz6IEVH3U03EtZ
7Ab9aIQMPamRO40E+ijKILRSZJz0xi4SZKrdlZcf6Cn39aBD8e4vQV1P80svvzez
jDZj1lQM/DR916fgfdg6WJuXDpLLE37+arZgrSioTdkiq4k/0Q7fra06V7P1QJjQ
IA0bi7kQYpZkVFws0PBhD7QHIAfw4TcEzlJQGXF3+x/42UhqTmv2h6Bkkvv5Z1uU
eocJZIUAZcicFxPyn5wcXSpByyhBExyMe/GZmj44yGHO4t06glvhXMMXWMkAG6Ro
ZgG149NRVBcFJ7lcDlauMTelcP1nEiir4TcnwoFk1pDITdsGvWQniuPYF1BKZB7z
UOAjzG3+alOydGo30qud9Kf0VB77nMr97c1H0vM1hvofQ0sgO87k8fetTPdBBefq
r6thNQ3rRiDOYBC19cJrmVuqbJJAPWjpkDEBCmCAGASwxMb10jhRDiegfPsu+acX
DJt8hWvovq65Mpe+OPxtfuLD8rs63vF1QAOJd5dvsd0yaNWuPE07KvZGMyQ5jjSP
TFZ6pcU1JX0JMqQv2s4TujBxADnlZN4xuQg0fTXU7X6euJpT5cc8p4y6511jibzS
++RTbZ1bIcuxlrLtnHCGXqcjflebgTfvQMWPQ4lJHVKkK/r3XGpla34OmI9c31gE
+TaD8CGBL8joexhuQP0hq0S8cglNTBI/geQDj0scuFwtD2Bfb5Bhnn74xZATwBeU
HLQJcnmq5gPOFoaJeZURoNYwS/lGuj/H3eFdpqWV3k1wenbkzIs/kPMMpi+zXvkA
gxf9GRwijhF9SGXf8CcI22O7ocDkyrgwiR5RzN6Mx8xILGk1lPtJNxPe7BKUgHZy
dRnd3T1bVDbB56xZLeB0OAwAFacQD3tm2ZRFfbx8C6iRs3kTYnkmNr4Fdl8atjtP
JOxxd3HmNfyhP+nq2QaLzDCA7fD5e8IMD8VASJDPetnKMv+XuPbbTqW/nUsq6NSO
bZmysIyQH4IKoyHh40PMKl/Ui3op6Brt+V7oRoYoQfaXuTWMouIwKpARFExlWGJR
/3eQPxVeHboepIdG/5HfI3XtLEcZfNmnmtpo2pAzy9vFx2uJq+oXoTjztwg910jm
F3EzP0yw1iSezeUdsE+iCRcQQBYFHjFK6sjUMtGPykshpoS4WqNcps5Q25F9BrdJ
eCE6QO33L89xcVrt+r24t60k898pvprXcouAsb9Jyy/eQMtrdtgpqaka2Q6x8Il6
3WKkuo53b9Im8eSVKs9g9soWxZ7J/F++kLczT1KjxbokeuukhhG1T/fQoLX6mAFn
3rgLUQBDTGXfZSH4NWPLJ1Y5kXO6qVQkLiLhnVFHueNhKMIr1K9MT4ya45dJOPJt
ywQb5UTKdz3D3YqfZ6AZTRa1EDw3nQESv2ELsPq6XRAuZj2Y8fBVvqYqAzeS3d/l
cnu8qfeEe7AMKR2LY4DLWHB2Fc9hbG5OckbiqyqOfqAxW6M9v3Pacwmug9nbyBF8
4hJS0TB3bpGjsfkPCjDmuYOTevu8D1jTw0n9rT+PycL7EiMIwbPXlS45hiYKSgI/
i8++6HmiAUtoElLze0EnFYgIq/Hpa34htFGoVxCVhxNirbQ62DXYK+djfOZ0WJ0x
qDXM/VobShv0Ol2X6RoZhxBh1B0sIPCL1miRB1pZtFQvBzUV094uvtcS4KJa81tO
IOo0ayuh+oS0KsbU+F3YPfWyGDjJE0he3+cmAwGfWDR0b+a+HwScye79y4ELFCCr
X6TK5imm5454dq3qAx/m60GkOfYAeERr0Fa2XHkcPbWuCJTn7BQKoJrrruli1Uub
8M9zyIEgWN4/qznJVn/huLpBvwK+b5D6S49keEwkBxHkP/SfbqbomeePEfvuXLHV
Xe3rWZ/Yf9b7WzTRmw6zqAobvv9McjXV/yZVG+DQqUp7jt1LQ0QUOYqNxZr52MqC
iIA+EsjsnaHq5gxGZabO6fAyhrEAvkrkMT/CZZ8G4bTcG3bDtKOS/tDc9kUtNixl
q/XMverZHVcF+ICwKHUoEJZbKB5jb3XeprRIv2x/vKa+KKtrRcMuktO89LpM4rRj
fg5QTnROuA3BVZ12ERtbUcOwkS9aGWNLYa6nQhih/b14fbpDNzVBoU9PtbLo6r09
J9TfMSAvsHpK6FQ3DEmDOl4TXbUWxceYEuol7wTDICsTFFTnFpKJ3in7biKYhgEK
DlN3ILmrEtoyjrCE7pTfMQc36ZMMNYYt7lth64rvWZhrtLcOvKT4NnsbyTe8JbOF
vEhlUCNki2eh+fPEeVEhfwnBK90T4dwtnucsYnqMJMoPhDHMWboKhaYfWjG+SPV1
0rvg7QMLibjS2851LG3UCAUiKfspuFx+5vYSv6UTbfK73hK3Yw5BN8kL906kbkzR
ycjnmQ0ULz6HLDOOf+2EGoOCJ7gDQ2raGFmB2kSrDx3liGy7Mm9ssEkFSvgburag
bA/LI8JdPr39i9S3L/E04NeT7kY5n1+eHGYEruJLSNVMNq2iDkew3jxYGyHCJ5vu
LXzyP4HTJU1yjFNvQ1mexQzCFWu4NR6DVa19gNQ22evrzXp3PD7DqamyqIkgxe2n
H2bP3wnsk0xoyeZIsyTKKWHPM2nj5JFOp6GMVvBUtu0Zs/dRcWW7RVBAFU2q7u2n
+oB344QB1oMRBrLUCdZ34Mzm2lnBlZTPAWeFQ6HhqTl3sls//pOQg5YoIht+Ya3k
bBKYOmakSzAcrUDDfAk3+xFxUQi3K5bUNE8fOeX9KJpJk2oCrUDUOEgG9p3mjDWi
9lSxkj0+suv4RGHkwSza+3XvfXdntMxFZCZKwaAucPnpPtYD4dFi25I91uQQZNGo
vkAjKKh15bp3h9TicXVXXhilVxGRQ6mwyMV2JQ7AHPJtO1k6Pg1FQDwNJpAqOADE
wNg8fuVMjM2WA9KFq5KFVBYmCK4hOKr3qshgrFtcQvj5em7KN48E6Rfzqn6bg5RK
ujcTS7icLhLPjdLr61IxMCvV8ON1dQ3/OSU3hLGvlMfnncb8tOo+Q9UevKjiMP0U
CvByp1/HzHku7/8remsDcV8/wW3zgtBXlLx2u8WE2zv0vB3WrTAlca+7Mg4lrusj
ttTDEL9VRdVu71Hv325Lzl7h8iDayVN7zEjfTjMoOn4kg+LmBIzvRJV6ji7LRG+j
Jf7kFv7OCEZtvGIfr0an1qQLh2h0Dfi1fK5PH4qskdBhL5E+KK5WixnY7lqxR4RX
sqtkk+rZWydVcrDgRAK8CQcPWvRMujBTmjjNtn+mpHDW4/r9Gji2sUzdh4MsmyTO
RqyLPPAk06Ui+Ywqt/SD5i8fjowUBtkjor1my4LBXCtKzIVaRGmygcs9f/CLpeCn
QGkk84QQTDdoIloPEZaOQpIjB5zEP2Y58BpGETOI/qKJFgnpQ9Gq+Ddb2uO6sFXn
+ZCo8DCvfsxSbGLwvP+ReqG0Cq9rnsd0DU13TCbAHgTFyrxGXSJ2SHJJtZem+Uuu
DA+v716eoZnFBDxz7vuKWNX+79GoMgySN3kE4q+ZZgimcSoN/CpJc3ZiD7BVrgQ6
1IsL1+8wCedGbfaZ2IRk+n0m4rFLNFIqW4sTtT0R1zdL3RL4B4QJnnaAIsT28dPL
ahZ1eVLUGfRWWaitwdMb2+XsON/x9/43E+N3xebtlq08Zhm9UjnmcIba9ZFvI1Pe
6EvOXgkFEJjau0PBG6mIyNaiRZ0pzDVLB3LPcsDRIKtjlZFqbqDZpugqUpEhdYxv
g9inGi5xm2F8yMlK+XJd9dNBq4wEtp08aKRsbMP3vdyOtYLYhNE85in55CCYkK0C
9GytGsXYr1b8c2Z/d16fyM/LffdHNDhskCWvViUwP8HFi34hPqak/irPa6v+8Anm
lOrWJLxAOUapeVaQjF1Zqcfl2ndn+BPsKbC0vP8buzxTdqW6r0ld7Umc/3sMxX8C
q5FG/oIPTRN4fwOWBTqu2q0KK5NdniD6Tfd6ehtKLWenEHQkxsC0W3lUmRsLEL3A
0L598oqkR2EYfcrF4xEqwZgWrlxt9ZnhpTSEwVvp5qhlGQsC1kPXJaEexJ1y9v1n
ttiRh91cw1CbO2auJtorfH1I/6oXJl2oVfHgVaIG8C1xgkyqe5U13YoE8FxwvY4c
WIEqQoEKn3TtOFRhVlFy020awWMtgWD3KZK+wDE/C0tvca+/QMsFMQvlZP3JL+LV
qIKfQut4dSTG7/hYCLn6/cKJ6DPc/yCn7nyITjbfEG88G5Cz7tPO1LlTOzP692wK
ONrbSxnHuZ8QA6XM824zvpkbsDkNvojOII/EZNEupOdgQO5lz1dpC1wAz7dtRBaw
W/oiZsEvzXWXvVPl76ZA3iUTRPqMWUQnXlZ4snc51lJC4u3YBRDlIOojFIEk6x7O
li2Zz4cN2EJxkMGtizyVih7CHb4Or83ek149aoCBgWg5vpr+JKoS4xSl/K7MK7Md
9ZiqoShbF2D+hfa/I1P0tS8awBK8/du4A4tq+Rgo7+8Tq1tz3gFTI52pyCQdRJtr
RwzvD8A5IIh8BFB76njgJLVy3G8B5DJuFzG8QxcXC+JyasEJlx5pHDh+o3psCXup
JIazANJqB3TOo0vnEC5quuhBhUd5Zk5+D0vdJrDKs89LkHEC/mJ1iatDVYcjBgzZ
ufR3XJ5DUAArNJLRh3kAvC1nq7SVe/MkwhSdAa+Ad31OhZXk9VmBSHCk+hjUE6jh
/AQ1Et+XhI/6yuui5sYkIIvM0wQ8Tb5V2LD1kFq4mIAdggDny/VIYQpsamFOs+pM
mA4ULqYDVB5q+H2hx0kGTwv4EKHl3iCeR3CXOF4uzbUOhFTaMCYJAjbhSAO0LoUs
H9ivj2DvL1QB/Y25VSUStQbad+LCcfQRozJBwHoi6ziufRHP/xfOa6Y2r4VHfqbW
zamaNyOAJx7fzDFF7aMlNnnwoFYKf6EMMMGxtzmGq88H60bhBrGjqO52uK9VBS0/
oMpzQ9Q2TMSYBJ7rndk4lD+rUjtn2RZiU048VtUhN8BxLHT+l5bd1zvtiZjnm5C5
RJrREqeucEp98iN3AWcan8YRiPKRqXC/MeNBmw1bSMBokZsgMmtIfX+5AtG7nZAF
LBARy7uc7147bax6RmvR4WO0FRdjpRGGPOFDdtONYUbjhr65zvdjJBK6KIML+zwK
35hs8GiyUWDV538cyBc1QXa7Y6UXIQw/xnCVjCKHUDQ+JkeFtf2Cu/280hKxpkqg
EmU8D+ihFWErWlGyAkN3DPBifSMYiIfWcKYkO9FwKYeK15sali9YZXhadGlqtM1V
Qhgarud1jleXXnDrjZIBQZ3JS1pPr//9n8ZwgsLe4Tburhywqbh6lvmAC9jJzPMQ
gbEh9QuHIIcHYbTc12bSBkqsPb+RfB/i4yFhSruWXsJ+NaPhwFyd5khRzDZ8GNq9
u4YehHhjDifBx/c9+ti+8tWfn2Csg1uC6iF3fPW9hCTpEHfnJvwukifOKpIttiPI
Y419SdBJesKezrowNrQMINQFOC8qyE6DmXfgMNC1sC6RQCaM0jw6qfdoKtb9X1LZ
z6Zg9tXUbUR8vY0+QE+pus93looe2/K0eTHOwWABuZ/9mpNWSJrYPg8pb14g+tpb
tK6gfu4AjhaOF2S8cCQ7OaLxNq9smys8KHsoHD3Jb3hTjNwE0Z3ZKQyCc/AzaMJR
sstVzjJa27Bkb25nyTWPd/rYhtEccxaZaH6ZhhIMrUduF/6wy8lhKIXSIrfrvphP
lPvIA6MmpJWXBsnt2qUzVRRTqG6V/g8eRRXoqbqi3kjDHtMmVTulSVstf8ZZlps2
90PD/ZSnvQeUl9wl4jHPczUsyO+uHQS2HkrPxcGtWU35bfgelg6ouniy4IR1RR01
pO3dJl2O6aQfz0U6j27GqvCeFbfa7ln/ERHiRm24a/viumffAd12OVmBPMDzZ7CV
9BDIrDHsOQcU9Kyj/HvHSQH80ZNRt9+PMHwHCKAsONgWSEG9IUTcS/zWv/n/2yTV
27U3tx1OEDogVm8t3XYxvXswKHZYLTd+O6rQy+NVtaTBEfsirS2AjgdUz8sGFp6C
CLCphrBX1Wm7aj4L3e5q50ooy9YEcniYy+SfnsN7iAA11oGQEHqed6yjaC0lGOb8
wgpCVQ/uy9yepAaKq8SPtF136fkHIhVj6ZOo9f4lXS8HsH3oOFtX1qAX4ue+BuAP
hPZtYHRe6ZiKuuJC8u15TvJ4lvbgSLakrw9aq1/aWk0EPfKp0O0V3MrXaNJnuPhN
Or1cSEnnXxyWtyvYkY83RKKcSCKJf8JfjqnGwBkliLCZsXY8b3e/7L9hxYLrG2LR
HE57zmuIegspiem3z0LMmutdY2wroTe9Wsbxidb2lKsRps7FYRMmye+keClcMex3
ZosQvCsfq1HwVEtegnVYzS/YDBuU3SkiPBu3+eAwsewmARENRlU1wATTBlLtSpTY
zrX6vLOKwre7hHKcSx60xL8S5hfTjZg2nsyS+LfK+Lt2tdYi2B1HBbr68lh8dmJW
wBx5slYun8JWoJXBefa6YJIGjSi7nr2oLflKbOgojm+B+1tzOJ1yDtxprJq7yXQp
w6rR8Cuu14i59XF7xoeFGWlJNKIHBYyXTJm/m3QTFBpJBabQp37p4tJFi97Gd3IJ
1AKOzopQ1vCiHmc0IjjSZk8+i1g3bqq44tSyCiBXZphDIjJNobKC91u26kMwvE0k
fMjNkhYEJgJxJHEyyt0t7JwkOKEHUaRMSxd1sdWybrwz9F903UZi5OvdVr3api5s
HgEDMe76aqYySOrza1XP6udhC55cO3jonNiOuON8BCLTSuFOa9bLGINjM6GErRUD
wtBnzge0Km4Sgto+qC+IUTjljDUrauJ0lHetXni0GN+0cMBy8tklhfurHDxvtmkL
hqTJhU9CkkQ2wTWTK2zMgVpfzRYe/vPEdJX7VO58oExqM3LV/taEfMzUXSOxJ1Zo
Cap/2ShLMJgF4xnUwhC7QF1/wsFKabmPzPYvR8fqmw2oZFX/cOvLYjWn62m06a2h
2UORtzqXFuwbQzjJiI53eZZg/V7VwkA6CtdzjOfaltL9faDkXcpDvT2iPakb21bg
v0CsxxyO77mWgFfcQO6NinkHUHJpSVu/j0RGMOUZPIqzp+MtpwymAD2bqU9gEaPs
K7hYFAPax8LicIklkCBeVmQdp7w3+k0g5tYtUjOJhPPUIQzxGI9IKi7OoqgL/yDt
qcgxGQNNAiqQTBIV11Mldac1O7dDlqFA/YE33UznAh94DRe6X6Wl9clPhyUBDIhP
S/uBGzhyGMpA1CicXjYlkgE8tBBkQ2UFB4GEd954belWCOBLc1vJcGVC2D2InwbG
s1O3IPSCw3vNr5r9UrxVyYRRbFA4yKmpRAxgoG6P04vzmK2Imt1yoyFQDHhM3Wwj
7M7q2VaTX+xWDL+MCE9SR8JUrHuo8qeWYXNmfkC5o8gU7QcL06uU6/Uys2zFgsSn
5GJ8enLcbt3v+yMGeeLBSBwYMM151dev1Q6+AdRtii9WBHUsDGUY6j5Plc9e0lKM
V75thbG2NiAKVZqetN4P7kcPfkWXrEQVYJ7zsPN0TFwT7X8rqnPBtMjVQFcBaWaX
3bUDcNGNPkxuvXX74jwSc6lWFlYMRpJgxcg2NQ5/Sf/E3xWgWMGKRSm/mJs+kk3d
c+dwlCnRxPoYoIQtktETa2Qv1yMNrhxPX+PvASetkOfJE7e74V0k8OdzPEwhzWD4
vP0jzjDJ64kPluzek5hFbeZ+4fHqPl64oNlmhqr3HEM0hsKAviPVyuwBr9BWx249
NeYMO19OQok0+/86wPm2FyNdeT+H1UXloHBmNZBXETiEggi2kKNkZvxq5nzHRBWm
/qq4FgSHViCcUC430va8SoH4nd1tyOLn3Q2+NRlNp+8I3/kteiMjvYtzXkx1LE+k
q498v6rjTag1xWV/EZESsl2qBfmhUc4rbxNGTi+Z6RK5OMmzrHXf2NfGPjOrqpdT
KL408RVPQnt2rYQwk+kQBLAUG+jJv7H25eZJqYA6YQu7/Np/0ILlG25zKuYADuvQ
ybECOhRKp4uiqqhMjjzwmC7untqN9h+vEvT0m69nUNazq5cqXfcLbc6E7+anVcj2
A6UqONvfhyUCAdo7ejxWJs2ZkKPtDqjprsxCvwdIoGMIuZj1lOUhdu07uRTscXc1
`pragma protect end_protected
