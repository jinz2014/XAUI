// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D4/yIp7dL3pCWhp4OzgIY3STklolPOiVtgDY48o9YnGTmL2+Q25tx+C6RqBU1rFw
oOjxZjVn8ohGklvwVkVo7hIFKwW1sQtbPAh/Tu6DnHuXHUzL6YUG/PcsgLKo2N+G
GuOAcnTZCKf1J7am8fuEX5z2ztnLQDvcuLoGi78bt84=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11376)
W1cx3adEoVOldi18CHuTdNObpHX1Y06mIaPrBcKByQoEe38LxfoHsw9tKxOpEUpF
xkSnwadBEfmLB5PRavF9etBikkPIYLe8OJo/AJKHk922L5+w6PlexD3MX/k774nC
HgTxr8uiA+1YWJsDHqZGoYHqBOnqQcu6+8PGC7qfZo50NFWUfHzKWUuDGFUdeY10
j1tCQbE1UbOdBweflhilvussGzjtbaes8Wx9VHNCBqpncxebzr7/jcuu+u8ITs4u
W4zDcS/XEUm5gMTP09irVX/HHcihy3my6KX7flneK62FYBtHWZBiWkZIv1KZ4Yid
twXVU/BI83qNj81pLogaQS8r2kzV4SqD50/Ul+QVwwxdvPpSCBiNY8V+pHFQkSDL
XE0jaFmWC8L0ZG7gkNeyN1Uc05gWsvDFIMvleaFMY/xxY7MWPnoNBgxEfWCqkeSp
qwWlff8bIr/5QePcFJLdUIoyiiyDxLA452R8hgIff6T91h3o0iA9kMejejSN81Gg
JX7dauCtxI2Fo5rpPRYjHdr6oY2k8vuDty1cLDCeiKDkgl3nazZ1Za6Ap5AHBxl+
vtflOgrUXFbmu8EfD3Tb5iANS7r2wFc3YiwzgI0Cr2qU8TRQaEtvEXIdplmLrIf8
8EB4+GlN5gTc7HvZd1EmoSMlDojilIMjv5Xv9tGIkmaZrLfJsZm/n91NIjQdxT6j
a4NbUDwzIWcKLEfwsGiWt8Xw85j2Wc8T4gHfdCzEKNr54BSM5dm+M1HyS935z8+s
z8xPCIu8Jr5EwSNiVSuBBJbVGiumlLx2SbdoiMLkfT70zsUid2jpPJwK7k0Sip9+
NB8Ros2MCbFI7H/9KQEELF0YQdNjqXE6siHs5UIGOGoK26TyQ1cL0+3FmMT77h5/
Q1C64+EodeuHpGQIAv2bmlaTsKc0Yet7WGOc3Wq01cZa94BHByWNrP0kUJfNDJZo
Qhw/2pFzCBYt6Lt6LCx+94pp0g4oOHZtfy3bccMsivROSG0Rsbfw1ruY6i//46oN
r5m0YT2Lc1Gtl+FP8yRGas/fhhs3B4DQ6eJGgxHpcj+LfVfOEXmVq2K+nWXzee5l
5Nxcadhev6MancZYM7MZRoQkZSAP+dIkx3FmCd88y3IY8/jBJxkcirOQV+9XWJOU
o7RRCg0zausW5a4waQ7a+qWthcHrzf1LhX1j2JEMREOaVYKBtESMg4mx9kQZriGS
wjXYJPvXZ3YhnMvhMXqtEEfOadNZfz/kH+GHzKecKmVFUolb07z+bL/Qjz9t4w4o
v2arzOlk9rfrd75wQFZ7LdP1f9NatonPuHJ09b//FSX/XXcoCdXcFp+fOCFiKWt0
F+WHA3BXyALN8WjJsu/VoaHTomSdKBARrIIV1r8I3BJDODEcSP6podlw64iNOc9A
0epE5X8dve/h8PIQTEf+sxX1tq6VZUeyxZTfbTyEi6wz6cUczW5KSLaBvdAsxwdK
uxv6GmhXrn850kupp/Gu+IL4RjQungxtV8DrlUIUpWPyRd2klikDAUsHB154XR95
UxwsocivGF30tBXaTnQsrWTeF4xZN1FM/3yVgpYTuFUvd3Frbd6a2dgOg/FkI9Mb
wqBB4bEbNVt5Sc4oBCP1noBC7+RVBxQYwiQ1VKzq4uk3+j0b+f3rGpsDuzlXKPoO
q2LQ/710zbJ7IlwX074Aq9s4ne9y5uqQ2Y42R4IJU9YacnxlZ1eYpVQQrCUq5xig
g2RAP4+cpDiuMD0ItTuf174cR9OnO8/kwem/nuxVgM4EgJvBorQmERyVKlQ3Dom/
FrIV4XHoTkmTR/pyRMTaqoBKV1o/xpLbR2jUTAkECL/MKnMvVb0eJvG1IK9j3IqK
ZaurO7DNSAD2kI9xY7h6dJzX77MACQ8pxNc6QSGmrV+ydbpYZkLVVevCMlWQFeZ2
zMPHWY1XklDQkKVe9xZwxr7yChtmWP+MruVWM9ZQI5mbae1GmhZ8mL6UmfLhbpdP
BJMSxJY74OTdylUF3D1V4uYDa3IsnU1hY2R9+mgZew+NDgMs4upvJFhZuNkmVXos
gWZ3mPZCVgupoU8WE8dCJ5v+70C3wh525WaQPuIQQil33c73fiN1Jzkc/PldVNi2
EjM/SLYFZF5iXMOlWvq7bBefr/BytdE4YegXGkXGbMDIANz0Q0ejj+iLJ1VMRnD/
cmI6GhE89/X7GgMaibsu/7DgrWYcYIx8T64SZ7q8Y3BymDeAaEUfyzu1bSCta/Zy
pf+DK5SQQCVZe/k3jkMqWSeWqvpELK/CBJA9S+mIkpaPhFzBFWDt7cec5bz4MpzS
Cq9UaIQzHszyNK13Jh6ezfuLSXe+5womPO4ruVpKyHjJmNt+g+YQ3w3jwBfz8HQe
u+aDYMgGW0+/lSPfxv2c1qCfpH9yYurunrHPjAqk7lEQDBIz/XWkMi6gRGiiPoR9
i2buffKuml/7oYVm+pqcgV4rLhLRRsYZ8phSse3pusxSrXgLkhMzDYlHTu8iMuJR
VVaRXqym9+QmsanR5sVa0UgFLRIfapAUmH+/TznGZVVQ8xLCs/d1IuqeAirCg4Og
iE31XrGU6MLDoGnyRA0eW72f7ZFdaCn5ho4eMLO+zqlRTaLlgktDi7dpWd4Bz2GK
9pMMgfPskwKRmXPeCRlhQtvh0lAr6jXNm/XomZ01sFHs7zpjpB6YchJmIGfVm3yL
KsfRu14hoQxN66tzTJpRzoEdik8HYvBpwgZ5f20t8RAgjKtR8j4pv8T3qZuer5C1
9jzyzymXZtLhAULiNUZu3wyBmPlWT82fD4g7ZVeta+dJleBctDB+Ep/dAM1984Ch
lgP8Jpdf+x7Csq0la7vDGoR+RXDr5rbMxlIcg99bojJZ+uGMq0b/ZxSAzhoQW44f
htTKkMZn3tiiaprFzsxfKeWM7k4ubwrWqxNChek+AGWpiNh4hTRLNYH+GGVdrfn7
XJWUA8zXOUJH1q7TFcd9tJPgLVBY+pzzf+uaKWM5HZB+MswPiH4vV1FQs1ERJEku
Zh/RqwdQx8ENJcg6I4jZ2dShaXbB2cmalXP2GxbdMOH6uFWCDsWFtNKicCBjnCNL
PPLot9zVtGVJ3F/t8wdBuhknjE9Yuog6GlVTrgKgI8a5sBrw7LK1KKo81wHiS9kv
vI6JkLBb2a3VxdaimnXTO/lIfUqUgnmsaVhwHYKFIOPC2Yefjt5Cz3gfvRbEEMM/
fpHY8Sxzj+8URIdM06k42rsXDAKGY+58SqFdK+kFZvuCxChk2sTye517QYq9kYmn
Ef7vDHfbLxj50HszIV7icr9kDWJA9pniOCBig4Hwd5samcJNza7b8FWAYUTKFHGW
M4O7r1oo9w62r/squT5e682GIJJ6okZLb+MqBZePiE1waA1xmAV9dshixzetC23T
zcAf0PlZK8cKWpDKEcUtQkOkK69dd2MoJwKC+DI/4nGdblV+GZxHQDOkgs7OH3sL
g63v+Jx1jiiAPcyi2/skNj+Cvp0Y3dTJSYG5CGaVi2RjCNMnJiz/lqd6xv8aUv2e
DLPCEniGkvFE+2XLGYUD+B0i01eslLO/XRdG3XeEZ6AVVwtbQ+d030QTXMXfvMUa
qZptI+CM99eXdTDoTrE0sTwZqgzu3iWEkg651oEIZ2gr6kjJH0ldyo1TZFzgqK83
Jm+Vr4nEcjTMCaOZCIJNTBllac4QL+ymscxqS3O5JAK/JEgGv1EBFLW5NG8tebye
EAMLgobC84lAQw7tNW0tE5CjgsOeem8o5JmUvEnBmZfeDsZN0KNLqpkZiVJ1FWzj
93Aqq5QgiuGdOb0mLDflRaoOo1z6BXPawHxxx9wkF2q5dggXxBlW2hHn8kHdXmrf
u+ZAsjiuQfr//eJLDREWCzNMYskuqvWHIot5KH8dnG/UrlChYe837e4sS5CckTVv
uzjHzATfHoLbGqGPCyRkZM2rb9L8AEBNrLhsP+gingV8pjtWFgz9OoFtk071noKC
M4prulZFTPhjt8YOxRzPsgVqwtmFUbr4ITgEE/9ogJ9+eHmQFPRwQddPSDmX/X5H
DfGfsbXWPgq6zvGoGqzkszpWMFGWLJc98a9DHEnL26JrLxQVllpfA72Vuub8RDAu
wlC1dSzd2QjmXdpzuwGlInTwreOE4UdKZsSavFV0Ou8BJgcGfvfRSh4CgyuXNGQZ
AKt9QrDnlekvZedpzM9zpe1qUsPzC+Fib3giLOEN6R0EI/blL0CR7J6r98FVevw0
6UWegt74Kw/EvgvDD+ToaoYlM9pqdCqqeIHwR2Qs+niiEX9gBKqVEdP3vLcIgmt2
4ZKrpXMJMXrjrapRkeNsXWt1Al39BTAZA/nDm+sczAlgl3jML2VzC1I40plrZcSl
pGHgr43n94VkbnQZD2Iu4IrW+V9ojFqYFEeKpHuKlEXFT/0T5+ImUk1j9xGhchY4
7fAe2puNX3yKaZvtMJYDYfn7sPSbL7WwsMrIPVCGAgSDD/fQB+5vGzZkDFgEo8nH
mW9K/xP2kimDTVTL+AOHppnszi1G21I9PLBwzrLEwFMS4ePjw5v/zXdyTxAAkHcT
8pRN2OYgLm25QZdXuhgZoyGhBWKRX/+NLyWA/Ct44GqOm+wItdw4N17dHIWCwNU8
eu0uyACrbn8aUYzwNibhkdf1FQUyIzzjcPEF9HmOr0JmqJ70UYmuIcIzxkPlGNnU
ANqX/YjONaYHA/7PZ+TzR7zjGZArnWgHF/N4vQXd1IPzBc8hxQYvdfK3i1LLkX1K
WAd/GLCAeUe4c6u08k3NvCF3UQ18Y2WdKAMjmZFDtmWSQ83Z9LuKQMadqmBhO/aO
X5KM4gdxBskcO3txserAvdodR5fNqr9/8kQP+NQ5sL/hvSJmbvXzw0XnG/ip0dDz
7a81y8o1clK/Y7MNINf9XozKZQIvmbYauP0mFDgOYKj4GF6TriW7ip97q92RpcTl
n91dzrZt582ju70NJdqxWGu+kiqy6llN4HVSZ1D+cml96LDsrBMJKpwPFHSOOqAV
zVO9FVQTorMV9yOnLO6+MPQ/UcreqvWX/3U3G3DDddXMWlk7W/8i8SqmCXOqvF3P
J2XzA0gfNTD4dY2OynCxkAIkbmUtai0OVf6R200HRNDikKmWENoDzObQdvI3ajNg
SUYoJq/S2aaNpEZZlSSrM5QnT9WvhQj/zEdayxczHoeu/yg4mPpUNF+lA+Zgl4QH
FIUmBmwOz9+FanfJZ1Qix8kWAkaQwPCYdqNJx7SjnhqrXEfwpvnWu8FS8FGBy65o
Jn5V3xyAYRrOldi0vPobkZIbS4K8cCRv5ti1T03TKl9KvVZySXY1moE/S5lWBChM
5FrpoPRC+SR1eOrmOPhMqJoR62L6lgvEbWwYxME7mjrAti/iugQqiYwcNNOwWMYC
kWhAUaRKBxFo/SVz7r98npaOsPNszyAsetMZhxtOPv/wU1TmlFv9HBhq7Ye8JIZu
HH0bfMxWh5CSD7S2SFPXl3utbV00pu8NU2FWTQsEOzLXEDgMccel/nW8K+K1AP5L
S2sWQR2pTH6/Db3aG1jrWkFmiYiXPVePOAS5ab3YbOaUecA0H343Yfb6qkeE+FeK
tSFwksyZ+Qbul22fvzkEqaKTnsq3b9Hlr8VV9OaxUIdboeZ5a/zmxEoiwSYqCRkg
YqJHzpyr1l7P5XefmfxJPpCW1xqVdcEdus6SELmOAMCmliwVxz4ySIiYQ3Ot6EWO
IB3ejxybsEj1iQ72Jz/n9bmuZqpTVVVKvUN3CE5rG9f8Pc08XGMm6z7a7YN2n9/b
szYIav0YN1CEc5TxbyuTO0TV32sVl0Imia95sXgvdiIIGiOWZg8xAdMTKELS90mO
j01UElUCEofmwWnF7cD+rQPbE6H4nw1FA9nFPTEw+EwktArjTU+1r6dITnEN3H75
JQEvu4t/ReTi7UZUqPh+D39fcV6zB7WDUpnv4RqbUHYpTpRBSOPS22JsDUCK7DKG
uaqDC5OhkaBIiTLKMs4CYlinC22PfopDyw0lTBtfx9WfcWLYLQVZrizHimnNzuCn
Ocff1bDLebHA0p/qkOl/B59RO5vVpok+PHR6DBoZPmm6BazrVFERDTaCOSOImrJU
VfH6dHjbXKI5nNgVIAvg3Rd761wWFq7ttLtKdE3FwqosAfDB0DZjQfdfsoYPk5fz
z0eEgRur2JQMpP5f2aVlzqIw+yn9c33uSFUxK8hxAiFwNxHlqlI3dQJvDCvOe03x
cg5AKI8klevS34aFf9WdmI9ZNilFrF0Pw3YdveJeYEpLszjbTHasP0uAC+Vwv2b3
TE7Md7poNBiaz87HaX+c0WpiPpRwJbW2SYyhMpOE6fctxTyvqyvxsHzSddLEniYj
W0NVs7gIswXoKkkKXJUVwbwVmEJa2jFvX9uUQFb8oDEHoM+H37BCbzJNc85cv3+H
Y94YR8b/rnVpz/14gzk1MF8ypSlVoCwJC/qa6OOwrcdsBAs79LDJBo7GrnvRaW2B
0PCR7GhEU+7P/vZpP9djqkaaW9f2lpyDjI30tndCHUy2E+4DennGO7xZmcFAWfZt
QPrQsN6pIgkoIunEk9srS1Sw+hD8unODyWJEGJVln2CD4KWaAO1B275KmkFjNcu9
xrwyvLRlYQ3yLPVthcxWcznv8WelF0/7NRfAq8N0joEYsBBJVk5vzHo5gco6wai+
zWhpfaXjRkFN2ne06rn8vdSZ9c+FmrazwHvQoZ2X3I5sy0bo7JiNTdmTMB0i3NeZ
Vux0WiqnNlMDlpiltajSfLYDLToD0R9RAr28jFE7wu5nqxyG5SBcKKaVY+eww631
HVsyFnFhXfQhVjQsNx8PeN22EuiXIfug6Gd3gbvSBw2VzUgPGk7kfgSFAsn8fgDo
5bOBo2uXYkVjQPKX1748ZTy94D/BeR8KRzPnJmtTGHlnff0jfzXgSZHicERZmbFI
hI8j06yf51vADPtnz2hKMLqJuqb7/G4hk+zE0j5zmI5fa9Ezb8DTv2uXP6cFVkgV
IZcW2QH4ghursoRDNZWpsUGJi7lnPScM7WmNn5dqQQgObx8feU0m9kXHCpShH35O
VOs7DEa2LxhO/EtTvoGd/BV9v4oODwFyGAbjbqPTc5Cx1p2qZMXaN3YasVXk7ZhF
nEUoWPe6wtpT7iYMDsxjcXKTZ3JmXdmxYeVO6yrZZZy8OeakoEHgOqUgiuHT4s1l
GKdt96WV1+yR/tq/EA0Y07zVse0ltcAUH56EyuNh4hLwoTm5H/4Vi9aWKKt/xRuS
Ytclo6Sz2ZCfUKcwiVGaHDL3+26pSjNRDtu+/4uLuMbzzu7DZYkqlapky+leTIi7
478fnfs6orfg4+Rq0dBz191keZsG8OGKeKXhHRNhKCPr7hFPTQ1Xc0Q3Gu2TDRCf
3uuRY3R7cU5aC828A5cZBCXWQeh46SaTqdhOFeztId5dQSeGMk2NLHisPHnLjsQ1
h3SVJy7vYbIAPvjwXRd38lTq8xi1G54AccmvKfD0BhZvHcT05iPNI7gDRgxZegge
foubo08IdzI2NNNlLC9Twzoq+sMWSOrMpGb3cHxURTr/ZvZpaXC2f2yLgWUDS+ln
J9q+KLIahYQ/N60uvvzMHbMZJNRH2zf6jw3Fx/Hu5I1Ixk9Ooso22SkL8l/+OKnZ
olkVWwx9978oQRYAfaRiM4SqPJcjtSR828+Y23M400wgZqUzjqRmGWPMeQlUfD11
5GktOWSPviXfn9GNTyPf+RvqYcS041KW7TCryzwYNu/KhnGR2HMz40i1yHFSEMd4
8c7QQoNeemWpMUOTPGuXENz5PcXdVQXLzgoAdFvZURafmPxYLEH+e+9jm74+Fosz
Jl+E/TZApjCjvpQBvsiKaYdZ5lCSgbof7oevHwn/e0FNsEwCzc3xyl63dNCU4v+G
Y0vMy58Mw1nLIalhX8iYPdD0s0WArip6CQTtnx+TsOWU5DQM1Awb/f9rjjwgeBDq
5KOFY9rRjxBs9GstY6eScRThpjpcXKQGVm0cPed1i8TE16vBjyWtDS3PlSkx9Cce
BSb4YM+6b8hgd8oG7gPGZsttqwZOEv8hY+lKKHYrylBG32vCpGxUo1bHgAqJFQw/
pWiEwFCFIo2WFoQbhXU2kvXjSNBYZ+IiEgQp9k12ZAx7aYp+oKQwS2Dd7S3dLKsj
vW90OK4yn2Y3TnHJnsXwH3fm2IiUP4cScyOxSqrldZnun34jzkkhkOO/Kh780ETK
Dus2L3J96ucQUm+xctzZTH1pfbnch5ICx/Dwf5Fxv8Wzm5AG40IwdyYdLr5RsK0T
Mf8zQSTR9ukLxhlJD+sZwJC8Bahnb0YFQNy+w7oSe0LwgedM+BXyPsLuT7WmTY2x
xFDyDqrpdKraepILJ4CmDGXNXZ6fnzPA7zmYIq8kDL/uM3nHGjQfGAeuhw9sA4NN
Wh+0rl+WNzU9jRbB6ObdTslX4UzGyTOee6TZ1YAlyD7LoOUMdvN1roYSUEXZ6ETL
xmVZ2rWD83oJ8gnf1ZreJHG5sE9p0IalenX60OVXgwumh4I3AlRhGSN8tTu3pORH
xupK1w3EBX5/2kdPyRmTY1IyTfAbnAVHmWKNR8OTMiHX1SFPTYNpIwoG3QpYOfcI
ocg9u4K4Lx4JRD0GC66KdovIzbwShR45h/xCzwJYSDNtXbCt2/Xu6WRJi03q/SuV
TsPDWQz4aBKEBjZ86TdEIkgIA0lzEq1E1J+ePx9Yz7RZURGw33/dxoO1nnylKkyV
nBtCe0rIl7de4r0v2rFSwIk0pfNCGJLsQgUKSalTNroveUcELB7x1hKrGIQ3W5sH
tzRH93zv/4G93ASRlSfaPN/gRc3VFLNBIckuKHwOKtCx+PCGY9yufUSaXi6fw+cc
4Dy7JdMWGoHh64uUqtHivawJdwaOGWOm/twXD6dHYQZ1mUG6ugSw6PFyggeB/qFy
th6rNY+FLfJY58KpLmXdTWblV2CytjrUTuHJddzjmELIrkz774DXm07YIYCenNKf
FXVO/JU0oFs1YVIEszXVMxSwOpiwJ1+OzSP7G4ZowzgNFvGWfBVgAWnFZ7xAAvBa
Pbkg4+QoN/0G4YYN09mc+DdQv/bOJETyg2BajbN55BDMYCDZrC9MkMvW9Hvtynrt
ob3P1K9dXDKrf2N/nD6P8GeXG7ykVAndyKpG7lHv2HyECYnzpMm0zWKy87WawDd+
NAtWthe7+nWf/2F3IdfMzqcEz2rPvN1MpmRWuA3kTOGp2lfIdi2HpO9t5y2YERF3
6od3WdqL8z4ejUXWrZMiFdRFWKuGKOqU1uHKQhhAyBEohklxuAxGl1WwpPxxLB4C
W694rCwYhtdBFcKAp78uEFPHMsN3FD5WB69Jm4wsZOubVuYp+04WFA8seeQabdQL
TGOBtwiXD/SPZRBZKOxeNKr1X1NpKAzGQKfAmDR4pVrYS684wH/Iqd7kCG1Q3Aic
ORZYxwDrvRCvxWXs5K/+PNpAHoNcmlHM+Sz/jfeM8Pz0/nBLZcll9L6A1F7ClMlw
KDGpIK9f8ANnd/XtS7AyOtBJBTu862V+Xm9CtM/qN69dH7nbZX9jKegZrYvDU8zZ
MHB7CsEzRaiot9ZHsZm8iVP5gREmAahaUHWPCjMbXCPMItPxxGDteR5Q2sF7/95B
Hkedx6lRMUfsKiqDhfsC+SLG9dfyXoGwyBsI1xh4gJeFUHL34VNtV2dFbMOVUEor
KbmrWzILbGXiVs50I1/XySY5SWNl2NT0k03yLpkS3xnlnPihIj2UVStOpU+4i8Dd
VHnyRIajCd3Youa8ICONFOxRl3Jmkz4wxnD3lJF6qu9rX98JTdgG0lV6ShQ9nNz3
zAvJjkxv3i7Vm8gfedaUraDTYuEtdFoxpprP9+Hznodr88RKWUiuC0p4QL6qFVGW
XXeuqBfQqm+m0CRp4otlZ8ZLUR84QFj/AoVhK1SA8ojWoY7Cix72RLLj8Zakt09v
lxoGF39v6g1AsuY5GNo45bf+/+DFxsTfC0/cea2TDYHSFRYkWSlhQssdsdWn7jWw
c0mKTyitKVT6yrzkotZe/A1QnkT5kSWJa2Jb1+kRehHBJaVKmKp1aFZShSab+Kgs
YJ+Hpx7YbJBBUjrTgEVDzflLn2mzzrFnAKHQCj0Ol4qqYsO8ne94xaydnlc3betB
mM8rxXINyITmptSVIO97amhtd3Fp4oRaCJK5kcf3DmJth244E4Ax+/+ilzIjWnjh
pGyGhavf4oowV0DFRCG2VNTn6Ot3f88RBeuQnxWE8kqM+F9dYRldKvR/v51ja4Py
6igOblfywcmwK7towNpnqzCouw1QQScM1kzRbLHEGrGkeJg+ufPTU12rxCs4LaWC
2S32c+HSPSsbjzR/xo5+OSJsuwCTDPCe/Tg3kV0S4WJYwvLhAJvkfpozje3CCI/i
AXvBmojH9YT3rbD3HhJrHuAnOl90bYU5QFXl7qKsyai75u+SJCKd0nhO0qGfKakd
gpCxdSU2M+jacfMCd29/Croxre+YqtlFtb2VQy+fyRFT0TvIYZt4TNzmdByP6omP
8uo2jZNDaT3/HhfLmzq/rjzuG0CQZynt0zINfIne8SsaDhsEaOtd5yiVDYiK6ht2
zx1HsDaN9L+ZJ2m/Ezuc00C/qprIIHdY6tsrVYa/VSXTVMNHSmxZypbBZyazLWDo
WSiXQpzdlqfwSFwGX1a0bvemQGJWBVAJ5nOzOB1oOG/rEADFDb4tUN/WpreBcFye
pNYd0RPPPfBKzb6GzXRXXvgQPp5qmp5XAM6urnEHr68l45uK5ktjsg2inV/+hB2k
ikfIWKYvQ6Bx+JOho0am9u/Y4DwLU+n9lDH+a+VohhiiPxNGNvd/j4xHm2l1QK+t
V0N0/hNzngbJ1iWchpLRQ/Iz5MHloDZ4F4nzA07dUh0WaNpZjFwAPz9qZEiVB8lj
nY9pMb3PPVnrbU+fxztApxcZQhXBBl8f3eeqVXKddbkQlx5BZPRldGnWPOBOxwRv
oFygg1Fj+hgZIDcm38/bVzTdrpm8v2zuRj/JhCKXu4+RDTSEHF94GUNX4WP2wnP8
0aVBDQZg3HwqR6JKUv1Dw3HUfXfynBt98Mz2FSzpSFAa0yXpGXeVWohW0WclFk/t
E8/aUsi7xEqqOeDxKvxGFBa+L4jSlPJdD8kyWgo48CDWGh69CF2ANU75o9GbHsZp
88tJ2z5gldkLwqXLvJWnIYfXCpROsVNlHvxl8vFL9TtWOUcn1XXfoJQeYc6lnozf
plsw1CVkxT1GdBNx5BKzAWQ9YGRfzeOYIdqub5vkF+pVrVs+RRBjyavULmmlAcBx
9Po9wYNMHIHJ44Cmt33NRcBqbly4W12ObSBw36N6KizqmaMKAmORGlnaAWZ/qmFv
LHQF23NqgNbyEnXzP1sBHrWGKKfKhRO8UU+JjpR3FsNADAQeUPSl3a36ll/dd902
JxaiUNWXciuhV6byWLadNDkQDTpS5eQka+qugVpOdKQ+q1tXFIaoM1ZtWa2EpVqV
BGz7QI2pXR4+EqZ6avS9oZGcJMKjkqZ8j0pLCnqXxYRtlTxg//bxeDcEmT73FD7C
GaBPDWzyGfiApsK3AhjXifUi1bX2JpXxo0qAO1tial3UnYLGYn9jAkMc1c8580HS
X5J8y01JkcjFcRfDfBOfVJi9XIejT8Gd9/eo8sMSSIq2NFrLLmP/U1BOlVwEF7Pa
9T6dMowaBQXJI4dQ0LJFaDtX58p+1i1FNmTsUEcAlHUjciq4ZobuqrFGic9K6dCz
esd9lC3XRtVSfke7PtFza8kX77s/cKBXOhdP9n9s/sVvEg8WGQlRGQnnkgGFaZBO
7GAcBeNzNVjlvwcC4LTNTmmWIk69HGGviIYZIMom3Zh8xNMvuxhyic18zuHi1jbg
Fewshhhr7tW/qQ/F/wukULl5Zy3V9XBNMzceUn7KDLLCGa9hXpQgWS5BPkqLDRFu
hJcUTnDGukFd/pTV9+G+2n3xNk3hgetITR7Dg64jZ6hQE+xCNnbQ/sy+HTucEHoM
tQBigeda0IZmJr/ZmKh4ZGLH/eKPRSPysEeTFnFsu2Kh/Iq7ByU+XcBUXVAkKyNP
WH5MRLC8Kjg512nAzyHCcp8+8eHctPbUB2SBppw/VyZuPl8HvjQbxkDME5UpbuAP
vm9xuVL6Cn3JArdxUSQmzms9+SPWxccHTzmBhsnh1P5x5NYym6x5mQCOE3Pp3chH
0Sm10TybFMlikW6u0M3x7CC+ZvzCMWvsuaXxeBCgfR+d2AUj3q3a0FrO423aV7kv
HheeE8S369yQrWoIAFVW53JZtnBKOrlZHCMR/GXua4R7Us3gSZ+nRYYX3IJmelqB
cQduLabTPVX4CI1MY/+PJnwpBf2xHXubGYz1PCQVM6n+NlNi6vMZcpt9+iCS/Z1K
dRpuKVmH5k4w/DC2WwNRgLKLapPUoYg9HwCCEhuARiIMUq8YN65oBAojFN7ZCXZ2
i3knzGRhVIAcP43UTdCJtQJPRl1UzWJo1US0HtGMuHUKy3z9kCayF03XABKM59XE
f+o7Q7ZYyz+u5np9h3wzExqAH7TCfKAx06vPecnJxcSHqpUObbM3xluvdM8fKaQj
xZjAvZQ9FKHz3R3cYClQ1kRfSCFTEq1PBcC4D1OXQQestoDkBCPzlTf+oBiZ06Vi
SkfwNoDw3zXWXPzRvn5RwTr2bM27NP9XTj2+AvtjzVPmP4vB16hBWUzFl/UH3aO5
TyQ9btkomdQPJRXvyxscAxS52wvrGli27h27Y8Q7CsN9CIeYqGaPVJ18UbVyGnDS
yR+sfu1/8QPBAtGRyhVobJJUjxkSnxhTkAq0bG0ASAB98gv5Pe1pVQxAE6hNCvg8
H4xj5KAgnKKXXKkH1HqvYtoVMdbwgeQiBo+esg8KrvnrWZ4c2+N8VZzMOpac3M3R
TRW+gc5V1O7VSWVAZtTzMqaapPN5U4LK7l1cPSH5m1KDc5lVeyu1w76wHV0bCNhl
D/6/II3ggLhEUd2PXEQie8Wz+/r3sRCDRUWq7Ylua9QdRPx6HuvCUg0psae6P8E4
QcC9HAhKptmDio5U9l7GEcq5cAi1ak5cxhW5T4l0YiCrsiZ1yui3sVxI2hq12fZo
Ek2/nKLkL0cNjoFK8f+ubtgkQRohVasPNGciWoC2ek3OBYbn8K/phYxbKsHanOfp
LfCHFjpp0YvSO9ix4M0Jn0dZJoW0caz82z6A8z3SubMXzYhih0DYWp/hWevovTp/
w0LGjk2jDNhqgCm3kG65Gm2e8iQ+BINul3K21q+QbgVTs7qAgnNSaFB320BCyUxD
BTvhwZLtS1qFx1RRokmfU9097/2XEXSNzvfqWuaWHI7lsEby33IiK64lWi7R+etp
VmYb7suzThZ6nQrKWaiXgFXjxmqE45e1fYXDAWMIo3A1tL2+TqyV4g1MAbV2LhpZ
grA6PTX7cWkkFDay5OYOq2OEq+QqDpvomXNEN0Nl8XB3X+umvRyB5qrrp8XG6Exw
DjKDpmMMrX6NySM5zl+MHlagXp7T6V06ZSFzuH/aZef55nfkY8VuV9yKCBdq/9C5
YI7wHFEn1sV8qh75FKFO8p+RuEHTjglK6oBTDKYmCnS+yuno/Zt8Bsbx94kQhnLI
r8pmI79hgKlcTsYYPqgt3N2UD65m9Mc/6YmDZmdOciyk/G/gdIBxprIck8WCYhBd
q1sBDX1v+g/lWMHl/fLfUUax8P/7SVhcmiRF/yxZcUiHosb/ZLtCSwmPMyZDUMib
7AMYwMlU+6g6mzHFZbNe9tPyoa+rlMTlIEafKiWdEKwu4ZZfncM7DwzeYuonPAhn
qHQ8t4RigY5ooeo+5wxGLuADv/L8WKvrTzz1nLDCJbJbHfeRfWZCh52Qt7YWqsmD
O+oYl9YmuKSP9uNeU+/J7ESGoGD3vuhdZgFF+VuGOYY5dJG6Ct3/O7RknOBcDK0j
J4QNvYRaCjyGp/x7UDBWfEc44qT/PRW1hv9A9UNdXB6njyIlh2ovUuWSuwPda/mG
Bvo8u/W6cLCJ01a+2HF2SY6+PyZXo79KaMfmaIe2JOcdoNU366xErQWzWdBE0IM/
Fj+rUHLxatn/vQYHFdsZx7W8zgLeILTKm5unVu0A0lq7g3oZ7nCz13smFnfXj4xC
N62QIOzqJC+TXui66i0kpXw/CTqEoz7FTxWuEZ3l5B0dfs3rNGk0sZzgfRj1UD94
ja0PJFNq4KqmqV/2T7atodkRciPzpe8OQ/iIj+OhUgMoJN52K6bLh7viyGPvmHVv
/DXT7RKpSn5Ka8Zi5KBl14dROCQDLPFbY2mleLZX556j0d5GruJyxA/8ZWyYd/IB
yQihITeDCpPJxW91GHGFyYH/l4rWpduH2VCj/sNQsdQUS6q9IH3T6Ye1GOsv/WXC
HMIe0w6xqn+7ruNG73nmOBRphGiNEPfFKOyV8MH5eWDDKCtpD76bL1ZTYYA3wg9m
CkMglx+pzuz/DjBm+UZztBwhM4Uc49GkqLkdKhndWVewDSGVdHqISY9E9mcwTBRi
T1ZozuJeOlbs9EWP+Ldukbs/G/v9Ml1XQad2OtxcNKiMlo1IQxJ0hOCnB65DbwfV
rOjQxBFK2IxyO5geVUstxmEFLwOK9pE80QO0wqhCKrkY05U18lRubCZ6N8EdpsiO
0ipgsy3Nn/y8ReAvnhQRkaTT9oHBgbE6puYYri1g4FOBZ7d6/9qolLBOJAvdQA20
W/+w69AOkM2lJYSY8+XPRIg1/7I+4vuU7WsxrjOfjzFzOZRnSn3TDpZTSN8Vw8gK
RvvYU//UEdyZDh+mAW3BvUVUesFUgyCZ7SQ/lCCHZ8y8PECVqXduLFouZkopc9tL
gCnFrHaM47CJ6j08SHVSXUS32ls2HKMnjDybqIOr+xzt8sRA/W/kin+pJZ0vvMbj
nJfOKsTsVmU5AgT4kQAe8GNVrZ5s//YsINR85KcI11z19YU86bLG+m9zTyIDOgPP
sgh/WwSxemTXOuTcidCRLqz2Corp8nMIscohaMZuOQpFESBj8jpmpKsowpmpoOhj
6Smoc0rl2Usu8MxfAgA9C9CHNqWs9j+YftM2X3TsOiDHkZVH5cOzvdYP0xWqnsPr
7bOogaEhClWbGYkP6EjCDgbUXZkiewDiPKUxCFZVzYeCPQQ/fjwCb3JSGJB8pQci
u6oc1Bt6+iQeajAjR+Ox7nbUnwKYFqTSTd1wpEIJcvPlVGgbY7QHO3VXHkR854Dt
`pragma protect end_protected
