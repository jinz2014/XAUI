// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HBdN+uWlKIOW7zgrmxUqFxdv3Zad20K6VWAFbKkQmenS6PRHAoWl9v8gJAPRLjjg
b1gey9MNxFIoP6wu+/0zrU6AeSh+N2FeU9GYbWinuxsHOYciRqW52D+mm0//DnZT
ZZrrngUmWgm0qRvfJMUufpGLxsv7F6UKICzgpvys3vM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
+6Wv1gaoyP1F4s1YqZ04lASkMUpN3lc1EBrDTguIeBbBjx7UVc/VeZJAF9aUMIW6
LR9jachS1Xj+TZx3iZVl3X03AJGubgashtsi/T8OuomOYi4cEyGZ7ptUv6CZR8oH
m3KwPrgbYWGmK0zZdWNgfqH4ypOQO7sx+VdqP+KsubrOAmAbQ8e3dlN000chd9Fc
WBDWezqafqdOmNPoz7lxGDCwl9CtlXvtJzU5x1fovcr7trVaFkiKDAdsO5dz+UwP
EbDNPHVNqwFeYwB4dDo6mi8T9eCKDP3cni2/SdD8M+VkZmkypd4NH/8KOgwBhZAM
x28BDU3UZowHb+0ibkB2KHVOncrIOwuMtiRuNLnT8Fl3LR6n7mx/E5n8NcKrPptv
nr9glmn6x1LEMTjEVpS0tPOqZ/1DzWAUi8gqbO7WKi4CmGbozOmdSJ6fj/dMscse
CJwnrBJcL2AY4TPbnQBWhl7Uv0Xa9KgIde/7YdUUdOiw09cxs3ptXnkJ6wGdKizA
Iv2L8b27nMY/jyl4D86GN+z+6oCAifEUL0CeqS5RSJtT76neonOF8OC1ymNG3KLU
DcbLs9Tnjzn0PbFHcdRfcCzBVdMwp63YM9rGTpy29MAguN8IiFNgZBk+ai57prjf
Gpwrb0SqFOexASVOHYmPn0kfbo8H3fEtw31Kq8vkNnRhgr4+FejgEEvaH3U8m1nI
M1ZxJ1wK6uZeKKnQMOtW8o7i8aazdmqNGFpgEU5zZLk3yy1F0/eCTbGCrsW+U1z3
oMnq/OGjir+DxRMUK4hE/SWSCJCQsOX6Uf9E7ZoVc5U1ds2jWjNCt9NXvpvMPVVT
MlleihYjXfnq48O9NX2zSxM7itUSPUAKLy8/t9lxzie/5UYAvq0Z4vC5h71dRJUU
wD+8p2CplyerR/9O8+qCG99QLSiBkVh9t37g1be5CD1kMe1/3eelXlKVMHKT+DHg
R9bHxWWtmFBXSzk28b2d2/GTnNXPiwnfAKKxcU5IqmL9IIIPSf6VglrvhPkX35DI
yIUD+tEjpPNOk9UD1o3NxbbnSTfxuspEA9LRLBEmKDOAFty2OTJp6dLYmDlIrTaQ
seNIfAzvymdWzTDPa/Nhq974jLO2yWVJaCjPoq7QVYebz/DIGUXpsiNdJHW1jync
J9xzakE3kk9txxqeRSGOJFma22KGwNDYTYpJD3hJ63kq7UaLeqa0piXAN4uc3ATn
RhBUFozs7SY7FltwC2XTnC0s51pRgMQWsVcGrE80uuFYxKYhVB0w2rhbTIgjKJ5M
Hm8UiVj9K46csKjUCaNhA+8tuSn+XC4g0pky2tOpaIUGY33/jchrJp2Bu58Llumt
2yVRWxWeRJpmXMBZYeFlim+3n8EXECfTbOyf6Rf7tCefMw7JpO5OF23eo1W8LaZT
QhK5Rxj9p+0udNf6W7hiibOxkhXG9yoQzu3rrAFwSLSHUoc/ERqni580Y+gnFftE
voWflNYLAQStmYzAmCR6QQ1dvvJKqaXwm6/qbXSN7us51U/BSamIqoH77dkbv1nG
GmyUEiZGyLiUTztWPUASHCp63/9EBnNoB5tKWyWEfWY7iTqoUmAA4J1f0nX/pexn
k6gNaLng3MXO3Bhq2qnALCFw/jhG60i1n0oevAyH58Xi7bFsHT7mE9oyhUyOm1sj
6A37F0NNXmCA+bIawjulc8iDrcg4wSBf4j/gOfTkjFXMPGBHrfJYJx585WU0r3iT
pPSyzXTfNpiEvMzcF3jZxtDSdKcsFnPseW2R4yZuwaLhpWXSLjC6rEMjiE65fvNw
vJMoraYeMbzl5gxHNP8LHt1CDV/b5DB4XuymxRQ1a2AB+RnYyEljEwvrk9SB/1A/
cqhrhfgFNdrDxqgtpEAXrISJMR4+VuC/iwFZkMe5fvHqugLGHqffype1tQSK89u7
z/136ArFqmCtNSDBCTEiDe5CZVNHZWiQMZDLSuajqh7bok+W2fKbig+a2If2ed8z
6bIZNQDyXQtT0dj2rB5f2WqnZ/WoUwtIFsyCJljisymN2ZQqBM6GLOXxNN+wajl/
B5KO0EH+xvI67L4dNHbzvqY5sdhY9QYRi6d9J5B1TOHHL46oSJcrrIBo3L9GTg3z
dCsI/4cV1EyO/cyJB5hffN3ikBNubOwHdte9IpxmBBvSUyt+IILPaJf++DBbUwff
+lRTauswAGAYbaDVlNrkZyj6xNnWOr9B3jZXueBQo9LVhjewGZbZQEVHNkEWNWE/
IXZ4n/iqnczz6qcI4Oqfoiya4vyukSS1NtLlWPdLzm3n1gaVZpet4CFs6ETilvzJ
3cHQchoIDT0qGh6V3iOKA0KDJkrh6msGdc14bAUpZg7SsajWzUDYmA2OMzXxm3dL
++p45djHgxT0G4BYI7rY/NSHOpGEGjVSX/lWf57aW6+yrszoN6GINuWa3Vnlq5dc
8Z1mRQsL8wsajx4c/SkCjGCUEHCGRnrEnlo+Jw6TtddIxlBI/UEjdCGNL3LRP9d9
cGcPSQ8k8J4duBspRi8UrU40idohKUp1yb422NGtXq2bELIxj+94jy6vKTjZ14pH
eGL1YVDo/T3qPbbys/eMuHqpGz2YaFSZwA2qEBXQvz9h8aq+ZlzM9BM2PxzRUcbA
kCrTMCYqVLjam/l4CZ/ma1K+GK9OE9Wd02s5jYE+C482DgIWvkwsEMjrpiGtPOny
r2n/69XNfQslbLqW/MNXz6WXZ4VLtvU1Ju5vl6E/kNKo+e4B0QPkOmXkGR9O0aIQ
OjgGE53rUQDM+GQ0dqqEIAB0XCCi8PfXwjEM7fb3wBVocIbbHNNiyjKfVLfPxNBy
HrLQ5L1z0RzG0er/yBBsJhEUCdQDsGzJjrqBntAyMWri7IdVHQeWJOkXGuzeq6WN
Uih9dZXAm2sZF84pen3f+Y8VtEWER2yu95q0xZkgowpDJiz8TcYH0lr2bqttg6vs
g1LgoGYkchWAS72OOVm/pEYjryFJANmaZeOZiAFYpkpJipNAibR38RAyeFGAEx+l
pM76oEIng9l5cNikMV2OG1/odglVYXJQvOXAXCXxhP7Zg+Y+fAfoZq28KGw+9GtZ
zqHsoaqDc8WNOk6oYbD1O+XC9oWcUXd8lhonRJZvxAWdj9Hrr5S7q7xAqh7g+nkg
G0lCUc6eq3yTEbCxqfDNCaMWuUX//9+5ih7fWXuZtFFLPomoWz9w8/GijZfkSaYf
jz/JqZrtZMOmCyYk1KR0z2Q9ABSBx2fukaKfWs7hFEU2gK8H+nA02TEMoKlDPyqV
9YWsff5Bj4tKOKde6fq5kJd0Yl2fSiSZcsK/SJoXA7s601M9jjjz0H0y9uPpvjGR
Zd9+OgKvT7Z058jVqUPEJV6Z/dVGgMUOyFw/l+lTzKtMOypYUuUADYXXozbV4jbe
MlYb5uQ8KBWEOFtVIt5RDxy1kynS0cD+mpeQsLsk/oenj6pEtFtea4X8IgMILXOH
NoqVKfuFM4pVYUT9NfZfHG/UUchyVSfRzzyKoINxZcy4TrVUX1X713jqu4OryNwl
SCYbjLxOb90c+Ef3kuQR/pl1jBOxAEBG9h7FeO/wPD9iM+ffVl8QJfKjZH6+ByM8
kFGji1MDw5LGKQ3klknAh83TFIvRV8EPvTF9kYWTox7BYmAlCyPwm0peAEzHk/XG
vRzRMvt9aH/3n5Rt1+ttFRU/pteDXLlDLmSEjLHj/PlfKCRRyhy/e22X+FGIeDBP
3FYsF3zhbK8xZb11Ks63U5Vaudwf99vvH+11mF2aOdQ4kE0y7vqEM0Tc/YkrsBq6
7+2xRA3yznsieQDYTOYaIcAdkYTMhb8QiOhyrK2OnymKGoSbAYZUmnyJqhZ8L5Jz
REE2DRWLcIfktRvmfoZyFoiZLPKdz9+wqgw4T1TnGusi0PFWDpL5MBAiXzeWnZXw
II1zCMR154x7aNlZhueHaNssuEt2/+/b5gT5bS4WNMiejXPecG09cJUMShFJ31+e
2mdS0HoIAVg7jf8zHcz77Ih/OEoWHJjz4jPPCau/9MpNDTqSYmMH6KUoOwrWWQbn
qwJ9Sd5eSQTXPUi/pr4h/7t2N5qWM/TuqmsE1mGueNT+Yc4/lMmlCAwcZ9jaap8H
04wK5RBndpg5xwvYAZghlw5hCZ869LhgV2PRYaxafnNceMNCtguyu1VghXVwi64e
3HlgtHNVy+yxXDYheb1KRD7epxGARaalYGyzAUQI2j5TTFzuzCIn6SxehpugrWUo
eOLHBNbe90kDZ1NamVXBtT85aR2WUyt+AZ4c7XbYh/PxT8zwEmA8kpB0pxuvQEmC
vJpebdjfdnTjWanZzFO61xOaFyfyxRxvFjkDd92sZeQOPzDZ18XFUahuRuGd+fRz
8w0znS5NR2FBHcL6rr1yPYWMdiTfS8Od9+SpSiRT3GDQg10JBoOeWE3xdSfweFwQ
wrgVThLlkNljzcBAIdiRBCAV0SShYaN2r6+iadcrZSSdYGK9qkG/dogDg72sCN+Y
pAeiS+usny7NnkAdtWr4vTndFrk6azIFgmsneLJlNDp38avrPZAOSMHtw9kv+DQ7
kfXFf1r7vFFSdntx5HfXo7k8XXUxjTcRTiGjxLjKILRakgKGe1bSoHAyr2r+cmQi
wiP02QvEDL/hnSTTcJCArZgG2/DMdjARsKCbLxm7RmQglB+RLedcbWvZnpGdEmi+
4gBPdsdcnYFyUaaXFIM7CugB6o2F97iUuQd0BtB+s2wbrfmvb0Iv9Y+Lbev+wJJR
966460vcpghfgheyyHJ77nWIibuc62ZeaCnI6WMDydtc5iXiLzxJSzqDh5eP6pxJ
hvau7q9nwSjgjshsU0+14dKvRKqH7ILhkwnORT/T+muBd3zFxR7UjgamFa/XbFAk
RDDuYHLo7EuKgEyKnSGQLysumM/veO/z4mfOs6a9KU9L0R6aXkqh5nWbqEIwnwlq
TZS7sxlXduC9ArG5IMI0A23MBmpMKsQpaLAXi+SgaY9BZckijtPsTy30INzvyppV
NP/RzkyE0BthhMAfOFB0+Mm1g58yLIutP6fArHugAYF8LZT9o0Y6ahT+6M/6VKuS
ldIZXxw3SMIz3qwQOl7kX3g9Kqfnyen4rJjLHo0nhpXIiicPdmvBEsguutrNOp3I
vHBBcF4X9FfttSMmHJLXr0VTNU3rpZhzogSQXvGNmWjotUcxZfLyLTVdylXmEDSQ
IIx13lHc1W02Q1z3Yh86JVfS0fySrq4FcdyHamZtLb+1i3WZPdQknhgJHrXg1VN2
YO17GiuQjKoCTikQSJOH4xIU/peO4UejdBSy2nUqgzGleDzkTjVFo5f9DOBG14qm
KKEIHmW8VezeoyfIop5DJIQVr9Jm5zCZne7Jjr3zdl5dLi8gf1zSJZX+tBlNtTQ7
37h6A7Jes5assyJ9ZmWhY7H2uu34H5TgV2CbpkNQG/1JovBA8BKhUCXLkxy9FDG4
sCiR7gmbeHc++oOtAxxMrTIr5cm72rPhc0Td5SpopdlFuyXoC7XvNXPSh4nYMxU8
TQt4yDs2sH4K49yL0Jkcdjf6TUmVwldFPSjYO1uke7ZmnGPOjH/wVJEJyVSXorud
twwSg67VzEq45wneg6sPR3zW00gu4pO2x+OS5MyymlKc8AXZdq2yvwq3eBOrHJl4
fdNB8ywIHwvtdnWr6WklUUjW94Ky+bmWxOgxkHW6T/W09BepwkdRSu3hVWPCX/KC
YdhsdkyIWpovuQigMBtn3FZYtuJjRxl3l17lorXgnIevzoiHoabqeH5vBYDmp8ce
q/68sBbQKsXU+l0Id8wp0pptdtwllKd7nc+EiXvzu9excT96udXT2+xaSPjD2TnK
a+vZocXtDiaCE3CozGenhHPipHFU1/NsJkkWBRfMkCkYz3enmAb4sPQ8ikYSjLYN
Jz1HgW+FFiulkETddXfqdjaHYNXh0xz924+S1IoQPIGF1fuyXqy7W3or2492zCPR
2ylBz6QQ0LqSqZTpvq5rVS6LxdtmbRLqFVaiJqHDw0gbL9obSx4TKDHBc2fxfINV
IvBwZtYEDnUkxae6SIktEqA9l/nWtKx/MB00wuc3Hji+4v8jIwVlmwxaEak85tzL
Dq5YV3odoh+g70wpgVxVOtRXPe8bqtVb5LZ80TjQZG3sUJQMmx5dUAzQ2LmX1mDV
BwOwJA3AqVRT+H6kj+dQ2U3+GMltxrClYvEi0AGzjaik3hXLUScExfnVMxrKakmw
aXN9uMDdoyFSW8S84pfIAOj7hYnVqF6zZQYkTU0OJpdD4QMU2MK/eyRPpEWNayiK
UcDEMxt4fAakxacr+mPL6ufTaEuacfggbMetKHe5zNgBPNbxcYXmBiM/ZLjBqmks
BCFP5WgR0oOgVcUZxZN4MLLvIgAPTDQVK7PP0bxMDJPK3jhIDCAkH/geNAltXC/s
F/3xiG1b/VrYuMM+ij8lRwh1uUxfH+WeRGa7xyLqSBAtlvcqSh0R8nlOHkqp6BYc
Au3TJjBBecJHOT+izqMiRsI6uZr8wCMKwerPR96Nn166CsLZIOPYrSgaf0iPeYdo
5s1JJfZ48Mdcm5QmQNjaAlLYt3osoX5cw/Z9VpiIrHSQWrpzvkXAmNvNIt05rkAY
UK5k6thkHN8ECbmcgwyTcvxIwDByzsx+T8PzfjeZQnuyRoojh50Hw5a+P2D8SSOv
WoX7qPHVNXZdrorOVusCQhw3Vie23MJfx/KRYlK1+OaSsmq43HXdCNeyHsNabtn3
pFqMjAb0g9Ti6NLUaFjOJZ9ZX26j3zwPa8pHhbc3pxBeCp3rGYsNpy1jY5UYvgPX
oTwmZTxGn97wCA5VTFlyt1SI4pFzlJauNHROufceLLmEzp8rZlXB/8wWHvVcUTfD
ozaEr8ZOh/fpoL8IdqXmWwd8k82DRF8OTgvzPCg6XKJ+3o28kD+Zlhc00Gs/TpeD
uQ05uv+zxBb5wC8l5HtJQfwjQ9SvCMDcOCO+/LQbGQIY/V8DPBOEwwm945GFPA7S
zPpWS2yTPy9EFP6ug7zTD1CUfWta8CF3LAsimiH5SMWOQ0Fre8BaEzns9kW2q1QT
sXQ0o5dWNSLXozmyZ9kFUgXy7/0u8r0y0YcNtNoaYErpMD4sYsoZHUseRQkxP+on
nMOSpT5YHt6WGI762xZ1lagYCgFB8iYTJEuUYSG0tI5FfF3yCM1lLxdFl/I96uhl
3cOe6DYc0Uz7gMW573lh9ce+4XWatCdLmEa93vOHFXnrE2wNi5mRenwf4bOmsCSv
VndkX28+udbSz2t2VFXfxafxJaSoIHH7aJKQsVh/P0fZtDsY8RIYOso4inSOZX2Q
7XCPd9M31dIhMrDYMaCMVBeYaNhiYjF8ZUoUcFjeVFWncvFQxAZjhXrZFwRpQS4I
3UFi4PgB3yXnXFm+0ZRIEUx4/yR8+tqw6K8rzGzekO9sccWZ/p8iBO+Uzti276zx
eK7r0fdgVvs4QxuEBPDuFpMA0lZNBAfgaasYNSujxH8JqXPKiWICnODJfaq3A72T
uUY1wQCPhefgvS3J110LYkZkySYUmx1USVDtwa96B94Ewo+k0Z2V1yUjlFDWyNT4
92nstp+hkeDogV3YAXH43bnAzcfcluU1mgN8ILiCuo6viX4xFtytu0Pd0siaFr2E
ODnjBe3PIZoHvnCIZ9EpAcFglV/5WnD3QsbvwhdM7WWZK/lpGtBdXZ4dA2Mnl2RF
xUs+4Xc1kg1P4UCUFB0og9VbmvF0510+peyGdACiFoE=
`pragma protect end_protected
