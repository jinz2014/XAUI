// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Big3VSHR7oUuVOC8nRvdzt8YcM/q3rXUYVSoY+rNvb1O6TQ0kRGxc6T14SmQl/Lk
24yYzcIVrBvQvQqrCvZoOvzlc/dMXVL8eFthLBp9alYtClRrZXLpHgXGv/Ci5fOR
ODTjs77tRkKuf3fjp9lcFBiSxS1VHY4rSLxIrqaSLCA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5072)
ll0SXj0lhgeBZG0HAUZhkkGPg1VcqqJ/L0EgwiEjUx+rUuqbh9tSu2YWVJ8BlB/p
t7UHEN0gCLxn9mzbPDsCA4my/RmW5vsNuzf26k8TXRAOhJa4Z/+ZmHEEf7+xamfX
UpqrtME5BWNpFNkZsWFCFjLj9FbJ5xO/+TaxGtGEhq27TMVZpdwLiNMK5jxxzn2p
ccy/k4FqkfzBkls6l3kk8CQjmdXYOrf1M0n8HM3tcrdvNLupeRS5oTUX3uhNmYAU
0KQQOhnRe9af4hiQX9LyreSDpOG/JEJoxsGWAjf9GuQn3iBLsZ+TAlczFgIScXHh
lG/3GXCWGaP8/hAnscCaXK2IEXcdvWCB2EdEHbxupMCBeW/AEBqznvQEfZF2VnTd
T5pv9EOof5fOmJvMqIu5E3zTCkWYS34F38nBV9kv/BZPB2UpsPoewcYVoOlv+FH6
ZdU9wba+8m0u3Taw7Faz2qlQvcOeLy8V7SdBoEeRpLGG/BbC86oX0hAwNH9InbhV
gmBwUEfA1RtJXfrha1Gth0eQKAt/b87fixdS4DrZdR/wptYZjKWiIWmm3dfbzVZq
PATWBgxZ12zracFz6AaVyQXRVsRMHFfy8zVXLK+yrB+uz9TENTWrm7xBly00Tsfm
AuL6IKvHTdP5GFl30Bzp7b5sFrevgaO89qi0hBrM9YUzyrbhoHB3JCcS8HZ9/CwF
EYaOAuL8kWBwygc0cl3MUaJ8EXjVbqUa5Qmdeg18zFgKRETuRsBStRVnSnIbcP/r
kpnjeKuu2fbV+giECDRnnpoWTU7xz2HbQQcOIdpp7sV8ULCztV+gTmyshbWVCu4X
0Q2uxeEqW/NGbehOqrKSVhYhttkzkJhZ6gbLXrj3CxR67qsU3gsuPqXlEMwsa3lc
nBhH6+1T4UuAwtziMoXal8l58Yfko/lykp+bstXWwbKtq3uiqPQI0njWNtzAuf2l
0a5f8jAcmLOQGkP0xfLFQx0idXNWB9pCa6wRI90leTBMLMCk9nX2fXddKIoN6cww
qJ/rCsvmEpB4nBMadAxxfXd0SUerCVIGG4IlEPGyJFSGjTQR99XR4tJgq1GgFCCp
VBhd5/W5/cIEc/rjrAGsBNdEE0hKIA514vpBQOpRGmj+SLMF3HcBCLcrOB+9G6Lz
5/hWblP6ppEnbZxIv23vKBPOyaPd/Corh9fp+n0PScYT9gtSuEa25ot5R8lpaED/
yhFDZ6ouGPemdS89FJnnlAGEikwImk63bKB8hcKpHRxZlMZxkd8/zmnsiPvJB4u3
6pwh4zFnsiugImQ0iB4KpEx6t7vC9RGvIs+TNDlEzHskz/mnnmELm76zXpS1rzHT
skjxuSxleGyrX2MKaaPDZ6ST7kOoS07neANfzZRkVGJJIn70q9QHXn/YbK8tqngz
+xWUzF+CeTzu+F1aXg+ph8oyuhGAf4EWmdapnA8iQjZckxeU3DvqS6MCjChKO4fH
7TuX7qfrXcxBaQEMusEwEDhX+BwgIIRsuAqQ3mT6LaVBV+kD+7uYLND9ZPO1ar+q
Can9mCH2W7qEKtt/RM966F/4+46slr0qqn/m1gevd3+SjTRd95vcXOnObXUlHXbj
qhjkD+Av1en34qVfSZa7ozlBQcHhI0loQma8lRBj4URZvQTpmdITgpH4krhIPR0G
2rS3zdNfSvvRcVw7SgWpQVy9o5HIMhHARMnoA/9o9uIBrV/F7Y2pCiLdwj5OvEew
IKGkHahZWk5AcGcieutRievoOCHPJkbO+bSwZuyExdU1GCHJaUBmyEtYj/HTy5/y
yrBcNcovKAB2bydzEWcbeAB79TmQDYjgBn1TlFp8shgbObg364V+ymQEPwRSDarB
LXtDtsHkq1Id0w0LahPM3R/OpipQSAl2RNQHQScPfQhbuSnq4DLgmeHyPkbsFMiC
bwKz9oaE3bjY/qZsDdRC0HSctRrhJzIGFNjgjD/MqH8Mh/aj9RStq12NeKcjDGES
0koOJ6+jvYlJ6wnkvNJZsWxvRk9B7NCOHmqCD5zvUuHj+HliSRolxdY5HbSg82RY
pVNB0zhad8JrNsrn6GtX4BSr0IbBAJcFEX9BfAc0/rb3W4/sCBn9p7AAiTuxbJjr
xZL3KcPsr5eENPjcjkZYIPqs5nwDW2/Rpyt0ZZvQC2EH279LajUkfM1KjCzkWiAK
NYbfRtOBbUP3dj0FKk1Ovr7NQacR8z9IK716E2Y7h15wak/1L30aCEkRwNGHJ53N
YBAFeZXu6qksqyLHcKQidYtKHt1fW7Di9Z//PV05dPB5kbirm6nVfCrOddXE7nUA
Hhi/QC+KMarcXcsqSuUlOTjyurEqEsECFf6Qa8Ple9Jnwjb7xW+hMqTXvnP6U/aF
FyplsWe1sSE1ocn13eqbToYBvpqm4vGgr3CRbCL3NFYsh1YGi08SqAZkEUHlzaNG
CGNRKqHrgs6FwoJ8EjZBzxrtx1f9KXKGAbBuTb28u9wnANVnRzaduLbV/XMPupN5
0F9CeidyXlvW5QuK5dn7WrMwuCqHOpXJyj+AENxP5UjbWffn5q+ch88/U9d4S+YX
X17ygaAd0ZyA3paKR8Svguso60W9j/Gbq/E78q08U4gYVQ58+3dnpDWPknaZLVXI
1Rd2KV2FN8kor849gAsKsbU3lVLRRiFv9QrnarjRHeLSpxfwuhpRwQaAc790VPo8
qYC55TuNMd6w++tkClB3muDsQzM5PPTq1tmwZA3h65LpHY/lPskywhkH3TFPgcee
0koG4BADJJ1zl5UMNUe+dnkfVvLiLPw6TIiN/O+XNKHc5vighMvawJIAnSDlg0pN
DyZb3m39e/wNLacuvGaEuKGtGFkGlP7FOxkLz16hbdjMLSyZ6M9NTkiCl4r8NXpb
lIOe8V+5MT4zBvZrk7GJnVU+pcCCvlCfy1LKzFBj9rmJUiWfgEKbW81zgpb3z1/Z
w3fTnWF6meK1fsWhtnplWAI/bJfHcRo5yPjtsRNPIkUJrbez4dvdKnS7Jj9mySt1
vTBoptRoe1jEcstMnX8CEdwXEUm6iSYiddEoNusBPBIxf0z72UnCnlmUKACl+Ks5
Dz3WRIRaCd7IUN0MZE8j6rXRxoOf++1xXnscS57jKEHhbmYzRL659PbcqWm9rNNZ
mhcaT1/NyJ8hKPkozzmzK2UKzDqaSNQ89fO+0xWs4hBH/ilE0IcrUb3OPPJ/b5IX
gpbGsFVNC9fgfckB89Ot1mlFxLJ4AA2aHudxMHgAdpZ8PdiL4pmvh63pwhvctvGD
2ElG73qchq0SqTLueyvP3j8UdK7xNqMdp/dbkD84KB5hu9c+X8Wap0WYVfGnsZKi
/LTgVh0dnX8Ct6e6CnwmHnaELRtd/K66HpYnKpmemzRM+BSHzb2/4HFSsuraME63
qzLWHv5id3nFtdQb6mCxCOlUtXGSql87/gXQayak4ovb9NcojGA17vxkFKDjA7mc
M+qHWt5R+n6WC+GnP1Pbw6WwsnMy2XHl32JqRJzmVM/ROlgxdlYpqo1DTLGYCmgL
Y5gZL6BLE5+Xhgz64UjRpgNwMpY3p2HDPulX66CXigjgYcx4X+NMawdE/FFuClz8
he0OvQ0URcamwCvwe1FyC3K1XtxM5ukkCyUPIn9MOUDEqkYOUqy1Y/h7CHXVBUBS
cbH9GF4UEHuWgRJzWWF8cpFRC9+sKJMqx574eicZAJKAzF7ml0omzn/7Cuyqlg2t
73UYRv9Bn0RPMqKUHoaWOTuS7sCjenYFRgn0tpLX410MmXvjtSgv4873DkhiHI7T
ZVxP1b0DdvCnV5PAvgSXwqnmXU+OV+DyRKcBc1Th6im6IeVvt4/sudWruuFoq/8y
QGr6+QZYydo1Fh/djT0JUe+5hD2XOqTn7CWf4E2Icv4SsxD+mtV2PGq8AfKYEDwn
Mj0YPjwb4xoZf9bncl7u3JLqxzefn2OzehFhqG+xgCFd0k7iAzQY4+i17+4OVaLo
rqlm5SXeYwtCDo898RCudtf/9s/r+OvjfFzf2tAAYwZzJAlsSsvITG0WI5+t2cua
enQfmqtLc4brwnnRi6dwfQScBVKrLfTSSrHaqx8SSpzTGTnZCzAlmihfmge+ba2D
eHkzImmmBycVOa69gsNXlCI/8il3FqwSsZsBWbmkoFjCSbfYlWL5FbSEe8a7QANR
6eiMQiFPjN8qp8g5PDmh3zo2WVDoVyAPHAc2M/gd9snQP+KGqZZagyR+xUJVhmOo
gKR1dzH84EA4OFwJVnckBKva0iK6/vg5GVJhEUXxjtNKiFPdcWw71op7Vhr12jy2
BXYH02pdyj0S9ZhVmW1aPdzEZN08/uqXAHMzogn9WcdViTB2D2A7Z0puedam+TmY
vfX2JZJM426UnH+bDVCBgzxtQlJsGqxUpaVpXJCALH93MNaa6wh3WVOV9zqnMlw6
LvpJd1KNAqO9b1apuZzBvSxRyconmLWkCzdXQiJT6vgpVAZpc7Aijl4BWWEBfXeg
RQGxojupfAwalf8+b1y73+CJ0NTa7uakrrJjc43/yBn47JwFzXmlryfz47Setojb
51VZAk1pSSWTPKT7UR+hssWKfper0cLtnzB1rfUoUlV8N69VY3njtnZglwnIpcMH
sKAAe9KV5yrfrhXIcHuDMsyhdlh+zxsCY5hepylfkHeZA3UF8fblhC0bgOTSThVY
1nk3CspriyCTWJzY0eeAlCUEghZSrL0sBlxf9+UzsED2tuEfr23Ht7raWdVmc0QD
OC7s62IQF+FRrw3NcoqIcsZU1tAC1E7sdhBLvK1YGuMj67+uHIm7ZQXMv7nsA886
jm06Nz1cPnyqRJ1FlFNqrnKNizQdzyZldl8z2N0KYkFQTbosAkUdX9P93jlCYlHa
i8LEEkNHXRC4oXhhDqFtiyeyjWkBEW3KZYlDYnGvJAKBiV5qpSVMLEdkQwtd235D
wK/nM8CxAuI2KxezYjCL7IWVIpmUcU+cS4FS0Ky3CFCk12DEbGSzJZGk4QhNycqa
WRQLEjVzbx1Yud3zJODSBRIvsQ0cxMiCgG0mkXtp9AahZLlJKXEVxrFChS4tCkIk
UAhOzpjFLEQJyGW/azseMhqGYqG8vaoD8b2YhBDnv6+ADiaCtehdzizH85s5e1Sl
cQa5oDFBCwDULbJsZfU4QOKycSO23ZArOMAmBS9n+/GMWWVhez3vVKZMtGrayyJx
cdlxSqYnvTEpcuQUD2GYPyj+jT0KyLi3Bgm6UcD7TtdHMmlPcIfX6dm20GKii9OI
WNxofpWY+zoeaImluUvYpzbLy6WUZim0ROGvkOg7vwMyNt9kNeRLrrtSkAJtt9TY
Xn1MNgAW9s4ySLIj9aYoUDIVl8ZwYMOk1XdQkobfjaHtHY1OfMn99pugWgCvfbmL
aMl1WXPLrgKFJMwzqMjRs0DGdQC19bxsEiB303YWl1TKNMcZBgyGsAr1XYPKbc8n
GCivbJqSgyEpF/7QTjr5lMS35nWDFCFl9htSBTLm/YbPNU6fBARic/D5w9eReepv
i9YixxgsDEyLVPAj/fhignCMIvZzaNQkpes3ILnIs8h5i1oqIu8XvDYM4nI0wD7v
1fCJgWEG2oMPmOVoomquSBelwAXm6ZBK1YeVLFmEGYMoEuEFwYsCJHSBvbBCEBBd
zAO/Xp0NkidG4rGPdVoFKPXTEphdsK0M9bEgvBozfTt8+T+Iq9WN05hVdIpexQGX
c84tJhc/hnynzGWzl4x2gccWgay54PSAkSTOXG9bEDjmAXM7nVpSXnkIPr4AMNAb
R6RkBnd2R5YNUHsAg2IOoMb6UO2w/JMo+tP8VjOaUtRoIUH/SMEk1poblB4ImXLa
D8My1fe61pk/Gtlx0PN5IecxDSPhtlapNbijWA0Xety+wmI6GxopmyoMapZNxTrb
nlEQJqPynz/ODkh81A/COISQq1qWmY+Q4hDzaQBAt/WEMWzbJEHoPTPTkDS8Gr/u
9dXSwezN/IMuuLWbGw4pKWLUJ4SxOG47IV0oOLNXDGhgn7tqw7z6ZMOKGmfsU57X
W+s78pienJ6DiWHpXKUiWlVTB5rkZquPbDM8dExqixqJ/caN5ITvvHpL9+ppSdDH
0gqWKR2b6qWm6MPJDCFIMcBTHvv0YoGjplrj7C6TCQTt16JoyUnzK0uxukHpl6gB
jay3DMxDZOWN+aoYC+DCa2x2ZKUGr8WWVJJCnmvrlPPSCNOMFAjSAqzqUuQOKCtH
DQO86huE+b14FJ44AVD7tKv16Hv74pGQ6f88yQCkcinRjMCBaCbAns4+iemnD54a
Hanpwmi+SfxZxtHASp6DWUgZTz11QrR5Xa7e2i32tqB+rfM68+fcPwZzR8FACHL0
GAkLD8bKmPM/u0kGqUvKvXXpCWnk1SdtV2VLlwy/DUfT61YLK5x7DTaj1QzQmyzW
EmKICgAiw3uxtk9SxJXB0Cwy+hL8ZtD3ikbfFGVRvPWZ67XXjNthNIgTYZzUNXrf
nt5Bk6g2KrtlgQL6OLdJAS9GM/StaOtqZJgKUgSVhsECEWKWxlVd38zgxRd/bncN
cC9+J8Ti/A0mkLLi6N3yVd24YdqxS0voAb3m2wLJasERJSisuNR9euOBCt73laWO
vIFTqnSJhaOwY4g0lPKBvs3ohsN1JJMPWlr/Sv0FEJukr+xtotnLO96XHONWDE/0
vKoToGwoLJRbKF0RViRNxkW3IBFu4K4bai9K1uMzCsnNdS0xJIEhm80lIM1wRzky
GxjFHuDWi/RF5KEvRHDdKlUpVV81pFFKhKUXQpxPZuU=
`pragma protect end_protected
