// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kHOBK+ubeI9EnSemuTTj84nSD65P4yXxTyUX+SOqastltCb1BLZxIG0XTmJXR0w3
WUxNFOuHCJKK5yQJ0BJeOexjXou8Ic3ikV8Cr3P3fcT2tTUnfcBeo5mdIdvybYi/
vbyp8TsfBbzoBVu0/XHunV7FVcbapWCDlJ4OfgRFGIE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 178576)
IjqLvAMZkGcUxXmqxVzIODCcw9MrAWpirJTPSMFV843IuJCa90PguCNZMyjgZe3L
SND63HTH5zV2AxfE61SvttKTAON1IWi4iOAkMI4WfOapbS5mclpth2YykqyjIMsR
XosFZQ8mqNb1QvvXg2LQgbcgrz7D6rDSxyoyEho8OZ4BtXbu2YUgFnA5ybq3K1b0
lOJQvkdvEEGDHAKbQksq4g0El0hgB6J647oiuUBooNV5cYRDNqMp1c4EcXkluUD3
+aAz2CD6OvqU9DE+6NGxD0RakSNYyPzGMjhS6LkNKRe+W2AYfRiTVLZAnrNUxsLe
7o3+lTyGpRaruRtAXwnKdN/9+j+Beuo7ztLp4/SIMvZWSmRwFE+v+5Ynm53Pnosk
8pakNUKixLEMNhyDhzQvCzgoG5O2HaLu+Asc6egYJc4G4I9jXlIb05Cha8bgh6+q
KbU4qDwblPy4OglerCjmtrjUSXnr174Al0a/ZI3sX2BQJSM1c0vaIMB6rB8BaQhm
TEqeQ8ISXvkV3yMi54Yy7ELrcqB9mWf8nboth+hZD4urB7V9/Lp/qPh2LZmk65Ks
splcp7H7j9LD9THuoEkQOlqqaKwVT91HmChrJNmKvHUse7laVKttrBM0Etiv1L/b
wm6dw2V8kVSfeG6VQu/wgiteVyRMZdVHGyJ/3MxcXjrx/r39GbPHSlpXaSQQksgi
4bqfpxN9uVXh3D8gl6Pp3FvLxeBsJ52kbSerjzdYGyGJLlNEOspBZE/XzBLf2AkK
4TcJ351xCiZiF4sfaRzHJnOrFBsUkDTNfUuM96BPqWAM10hKtTICDWCOmEKOd8JC
1GDGD2SBErDqUAbXaeiFYqCF8vPqhHy6TBkBeOeJE2xUSBTzQe4vu3j/RWlqglQg
YXxT8TOqssp+Z0GfPY07LDHabdOx7cHtgRELNxuK/x/HIYXbzBNE+WajtLpkG2S/
6MlKpvq2pfQa14dKD0AJBDFPelXPZcLCL8HM7YnZmZg7YS52zUScSyu/0ETZkjHB
i41P8ev/pw8L/pxhMKZfJ2g3k1WFgS9eEAWq9n07Fsqp/rd9Gofxo7hAN3ktFGFV
Gz0kDjrgE8fIyE5WcNS5sXaQMGPSk6ha/JhXieQLrtbI3x77+hS7nQZJnIYFQ4of
qokls1XNS5RZw/7OcYPh5JyIv6k0Uy7fwUyWELJ/5/d+H+eoLwZ+EwvEaeXjhoeu
HGgqU0htB8E/fkvaMcU1oVN5LpFbS9ot7wAORyQpgEoDbWF+Pmqwqj/HZStxg/Eq
MTwyDYA0ayl1KY4a3UA3bZmAI3jfYA9bjHPfVZ5ks+4/zUpu4hV6ogh3qJG+RcdP
UCCtg57QndBkwVKFxtualIVTycMK5dz/pmHjM7+DgqBTgH3C7F0RVP47qdoJHgfs
2SiZVX8EjqB9HVimp+65yx3Jhan9falmG2drWdAV5ttHqGwEAtZv4G3GJ0EgZVJz
g2JEUefK+CX2VDJYHoUSExb5GYdJrpfWIYwNJlZKnbV5GqkMvydmlDbhFjssTHSc
LqUGQGzGiRa2aSG4eNmilSyZTL0lQvKn1yOOmgNWhow+s0it3vzeAWIc1fx7GTNb
3jBgC+j0vJodN5E501FBKNd9Qsc0/X+tx1hDhyABoBo5UmAMGFYMj+M1WgtQPR35
CUNZLP/c5h76SWpLgydt53dVYiuERVSxsI0epOnPwC2U4cI64C48AvWktIUHwD6Z
NSubAqAD76p+eSSKQEgt+CDTqItBwwZOXCneISgxKgL/HSMlAXfnvH/5OBJfrdGV
TUEpl95u3EdfocaYhqewcLFFm6P06O/WGqYW8gLGEOJPDiCKvsmIqT3nVYTQVFS3
KrG+9tGCH/XWtIhoekI+1f+tMjb/Hg8iptIUNwn5+aa53tgE31ALmwB2UKAMCNK0
kIXGIvu5K7LbUOOfwVu4HGh3QuEf66r8d5RPB4An6T6Uci8YnUusu1KSvos55ahG
Sy0I3UwUtSst/uuTy4riILOtGi9/9AgLntZxc2cNRMTB+ZEnrvohUIm8FYfSyJj0
KMFexuvGdK9asYwfznCGwFr0Y6HC+qwsWh+M+4Ykb6TrcLNgNoShYgrAZ04imQY0
XpVDnn05qVTqLLCOitE/QsdW+n9nIDNtOQC9s21fxemw/5kMrXtvn5Tep3KJlcLw
V08tNR7cgM3tqkAjfqn8foX0DXo9xcGQntEtVWqzeiBCAm/L2vWEzOYdIyczhzZG
tekqbnDBVjgaqIG00G2EMjtm2XkLSrEDJkZAZ4gzhSzNJEhlnFSPMaml22IOd1el
aecdVH3NhemBy04J8NtGR8IFyWVUc/P5elupo2VEFImx49eoDYmeZkoYCfqXz25t
gBtI09qydFAfL0Ou6SbMoDUChCoFJ0yA00+gbjwOKXs2o0ckl97laYu6sd7Utefz
KWZatVSxt0/F7GAfoCbx0vW/+bKErjldwjAqrh9ZrMtIrOQqEZJJrJqCAcG9kYg5
gHZWO6B4cB/7yjm2kpLBDhmUDajdIojCV2rQkJeDFxwH079G2+36i6Qe4WfRcYvw
R3AD/OlJJaTSOxPJ1gM/1ps5edd0lNA7QB0AK+vQZpVkmD4JGHr+bkEUaVQgUn/v
rLpmAZP2mnpNr1NC3eZ0+opYdf//eimgon46jFVKkfNFrC7Rkk3giC+9yJsGxKmT
rZ5gYLIxOaSRwxC9czsqzmZDsoU2MvreqAp7uISHHhL8JCEyl5Xs2XoCFTxNR7BR
9MX3rmt5ot4N9OVHwJyJWJpVTEA2XyCevt/VdkNXoAyi+wCkUms268KlXYu52tWC
aVZw//4ZINbS7w/GpRhJPVzWwau9XU+tay+cReVz8vbxDVRmy4uPzFOi4kskLnVm
MKsoAHdW4oJcM+nyTSgSKekTutm3HtgR1b+qNoEp1EkndoLzP2+P117xxEo10wFg
HhMJc17N0OFQQsvRzL/1+ltQkqDAlGPsBacoB6UxyZCzFqxcnMu3ymc/82+8lN1v
Rgk14898sf4IjXXK5D2AQ8BwFIcgvfgH+fegelF9PYCyBrLfHhMja+9R0qpFZKJ9
80yAroue1XZ6xORhc+rBABRGVzomImg9j8rEBk4kPAPdJrXhNzOeeFxiYn6PlhPr
MOlYYOsFpyUn5cGDagKNt7YtKKxy5wT+8yloo4wmtNvvpwR3CPP1f4eFS64LDfjd
LXllyP1A11W8xq67aO+ySeKnFeiemiqf7/2OYL5XK2zdCQfvWUSXbrem0Cp8VmHw
YVS+yg660jZ5XBUBIwXiBXdAkLrfR2mQeBB7t++E3gi59WBs/numeyD6trJeZE9d
GWOtP3jDwdj26fy7CtIuDUl8gKw9WucBzGyAXYwHBB0eWULTzNf3TM9i3PR3tWbZ
xg9GEZtjD3cLrDWRf0QUZuUWtGYpbf3fb0y81zunHMpOXs+3l6TaJjMqw0uCyx4q
dpY/jjt9+fxjJMFIUiw0PfV9fJYf0IR76YMpCgecztP+S+MHg9KIqC4iMohHSJur
W+PY7m0odTMYRSxk2eP5Xkw8W+0qmtbi8L85fHFi6F4IRO+w9XsCT7L8fyXH3DDq
TujGSqPUQPgZdrMLmgoKrH+ReXK8oTqwjaQamv8EH6DjZhdjfejVO2Gg/NtynBFo
SlNOSQTYE06ZqXCfwDDe+YqBC3mmvmSmyeIFiID5ntxGKbvy3rt8uUtw3ScuDqNa
eHBDPQL2xH/xw+80CEVzQPt0WoRIkEpuADkj41+UlE0PixqOQTJ7adWx9/WMfw/F
az0vaUvfnwkqqaMEkrg8q/S0BDDEKYEB0tduIh1/8LXYw+Xqxhm2Ody7YQz0dP1X
kYCeU2Bu1mArD1lcT84gkjSYXKia5ATrUYk9E0oxOV0tqyDopqCrRPtX3G2ZbZpf
up3bnPfI7Md0Rcq+BHdrbEWK4GkynN5BXVItPcyGElvnPxX9AgzfOL0Q8/DTlJOd
8SOeiBYuHTNSgrLyaGN/V3Xtr+PGswXN25+NPA7e9xEt5TBx11j7dmcIZJKPhW3c
CEa+udP0fM//BnG5cTnmg2j5xYTy7YqDuv2ZNbH0ecirS2jD0c+R9cMiWu6h55Ja
uF8LQpcw3ieRIOn4PNC4TeO9y/4PzNSNbYa1iqj2pbQrj51k1zHyYQVb4NOyP6nR
8ozySwljRFpHApEmDylT02dV3lPSRqou15lUVR0fC3U2cPnmugyFMYb+YY3h55Bc
l+88kLAUSaE5UD9HENOH/OmTRpC5jREI8qd8QQ6sNme9X+oQZb6MNJRfA6nP4t+B
VLSlvWBPJm4mDXGe7qwMVfw9DlxmsmoKhkkZsERtxTiy5GwefDuevzP1mQmjVn9T
mezWjVdcI9Mx/L7Gqvmhbg75XHaFN+CXb+qO6kV0+wRFgZ1DNF9K/zc+dJ/k7Sav
xHCCaDGQjBCAUXQq5pjLu8BVpMzCeZSPMa3RI1xYMOShpB5gwSZPf0309B1VNL6w
0Z7Q6hiXW2mGWZi9XvDgJnc+JZNngXOvD4efjRunWFFI01qELQ52LSyS38H9nW8P
oVWwvKvJ9MAgyApp6lqlbQM0+bKhMO0bylpxc/7hbzyAc6fHrANYi3K9h8DYv6Fy
UkTFNXcVO2BR8DhYhV1hvoJcmbPAxHKZDT0BckkyBtii+krmP5TPklUuOI1GcJw/
H0vFENGClGEbbUMfJqWAcO+7g8nsvQViFYCfR0utXc8w3i8SQlF5PUBXTO/gvy+T
U23MGo6p1WaWgqbx6DY/EeSRwKfqSXIp9VYPPiLXnFePTGcZz/HUSeIZAIm0+qWW
d+VgqpHjxOxeMd/Ol3xObPLbkbtwzy9lavjKzztuNef9zFp43JhTrwjtjggfui5h
nsCTj/OYH5B7xam3aIkQGk20wqixPaXrdcB+knHQDF3VzHg3B9FzuvyR/CDMWOqn
ol8pvFW7xhDhL4QMZEf7A6/KorgrjbPy4iTq1rx2weR3eK95j6IhTiaYPy+rsyl/
SpPOW73p19nUFr+BuFTGqi/d9VZNS9gNEU/tmHZ9WeS/T19VKT5zB3bq2iL4Zfg8
Mu3+hvtWsCt5bgWrn0nwFjv3SukiAh83lNhK/BxzPPBHQiFG24Ha/tuFfCSQCIEY
KXEDDDZe5KW+qHH7baXQsCTb8BLBBCE6WWcVIlJVfNHMN7m0su8239TlyshcZ/kg
KFCdrcMjnNKhBDk+qFySJqo0MAXyDQMyo4wjRVzGy8dJpIBoTV2htEoqmuP4ZuZp
bPK/kgVbeQ8lt9TucaeNdJd8QbkX6BYkuidSQBJV//KuRVqD8PTOagm8rLTmEs0F
HesQQRfF7er3PFfSU78odPx4ffAfTTwPEAq4uyX+4iV4/GFLgbOBfZs7uaXIse5X
p2Djl00jXIvx4rMh1P6T+6tPuKqRn1rqUdsOz/KDVbUb4CDPfno07AR9xzYXxd9W
suuN4Irou8AzDgs7+16QcsUCa+Mx52c4B4BXGMDX0fh9wucUinTOEPCniW7b4C5F
dqNm0pMrdhE47CchNw+Wd9ySxD4CHu0jaFV2fafmD0KQ2bJegtuJHMhrLsqOY7MT
rYw/7OegFiYI27dkDgXPnAxE+G+RUHqwZEowkm8IzILlpjm7DIfUn0Sh+FuVBqiR
Y8okZZlyNj6jD9ygwxoe9ytyHFQiFWUjG5BLLwTG/LWwl00xlkXJ8AL+cnUWFLxM
Vl8JNjQdC/3RMEjM/w/6DLwj7J7tcSMz22i6ce6HilJyeddio2FhMmcjINK46F70
EmUipOr+HYrjSipV/9IIDLyU2bJVcDQBf2663jEt2/hf7wH0rIUA0R6Ke5BdNxZ3
0yDyD5qc80Vr6DEpDkDxcKzXzpxIOqfw0822RL3I0fXQH+ZfFopp7m4Z8lbi7kMh
7tOEF1RGA4kZDhvOXJ6TqF0vWRbN9FYjBwhX7/rhcjcSZM66iTXdzkAm6XnLCQNp
fWj62Lc6s8FLwo6/OLRiHC0YPKldXI6ZLldBEwFFpAHDoReB9Gy/7WuDV/f9zlGC
hmt/4zrA003mkHInHMZrq/LWfG3UXv+q8Mnq/QnyrBGbK6PoesRPPWiSDz7ybJ0d
e8DWgp5+l1btEZonhoVsgG5KTocVmXzvalWoCl70ueNaq+bru7Wpafs6qSOL/Xdr
kfPRCF1yKU+8xRhO+oDuJMKnDqwRS4/bSXxquoOdaGK87SzHKtjmcCGDzwlHQYHu
aRI5IuEBMNiMA/NABhV2nsrz3IaSrFv6/W41YR3p8sNV/MiE6zmCW6g58GOYdxqP
fPKvbeYO4yybv7GjtJym8nOzPX1giXwBqTEewBWDhuN0UJPjyCrJwo5SZTIOiwpw
sXXw550pKuici7bw1TI8QLXxoA14t6Pz8wMs8FeMwAR10xomcRKtXY0E0QvOt3J0
EOf2zMseUkiafqILF+79OD7OhlsEGwqWD/dokVL1PXaeN+VSRmLfeNRV2gYVqI4u
f6m/6BB0kSumUULL8p2+UN4vMIzzcESQUwX31BzbSXb/zv5Hcogvo0fKi1NLCkWV
eN8LSup8EoT+2FfVf9yqzPyH9ahbC+rjmSVbaRkRLCKlUEf5Q+USvathLO6f4fwE
Or9V24ZCDgy0y/lCsAYWTNA2skIhnRFYDEeg1ER/MBZsTOUGHn9fa3oVltz2qT9Q
IR7dN29DGzVD0U/1y6tpCQ2Cqr7S9PnsoSFssLTbfg+iWw48Z0Fw9//BzRpOlMvX
ZEW/93HbrhDzC35OVTjXW/kk5MwTDadlWNwHIDB1cDukWcLwl0/tBf7JOOoh0csi
yiiVtnLji5iUviIzsfPR3PUA8tPAzw1/XAPrgTjw/MHIacK3qpNmJvz1qMMoJfYT
eZfgAQZZX1i7ptdfCNh9YNA2qx3CHkoPhDj/6H24yWDEuB+xjLfPF3iUML/MVpPn
zRZKgcMvseLHR9snMiy7ZZA/GNnZeZX9RA3kdkjMbKsA3TTd0rZePbeEdqoBxEbL
2qIgS78jn+vZ/OKdoQEtdDpTM1kxOGmekVtvy0ha3Pd/a1KMrQqt1KjJXQJEGPWR
qQdaqBf4rsyMgKlukfpTl07kqXzRQguA4jOJ8T6xwv52YLkFnqUKp4EZU5/ApNeN
Br+p8AxSk2y/7QoGvmIAU3mp/FsAPOSsLiyFIPagrl+v67/Mvi2VxaUafUGpqccl
NoVb58q0B2a/Hzn+JkNz2zYQIa8DApqtJyg+PEMR67jRdS8c+TGCOiTpYFKuOAH/
HQs2G044kj89f9gPCpHzZhFjU62CqsWjcrCKTbKePxnTl2HLMx8gB76BIh5v8vvZ
mrjCDk67krmXLpWbVNCNYRevxKUDqFQw/2L7v2Szt3GMaNr+2IMQGZ+cfs6sYP6S
1HP00YqWsnKBZvqJCSEQRRZwokwavT9EFVl4baNAysq+TzIeWZ1ASKQ62vHS3hcW
9+5929+0JDSb4YWNhMzSs6BiwVoBFQJj6qXFsLW+LtOuq5fIZ7TO7wC6BDSfawlD
kUd9wxGPeaLCAC/dHkht+TApJRLzqNacx9DweNqG2G6XnViio8yaktm/d02sPqMk
YZ22/KbXavPzlWVBui/KEuJFq+E9u3mpP4SL4jmepLC6b7QhfmpbvQHwiWHlPeqj
WnpR/Ktt//VktXZXyRk/TZ6H5D9aWFy6TyRRhasPWScg/vuTdLLUYeBXDIuCXjTU
JocahmVG6iL6euuPJKgTFN9bGZbIvb3L7rSzQmbtxXc9H6vOBbEeMTS356+wmmnN
EfrA0brX5Fy/0z0T/sVwitNrCEUymfZgXhZDNG4nN811YhuBKtGOB4d+prb6vWRW
+DQ3O2hIRhei/TSo56spuYtOUAXikvERQEy4I8FoSHUAKfWn7rowUwBOUXeHyZgu
nADgnb/60x+749NpYOiKzKAGTGRC/Zb9aiGuSGucuf8tl2W1tTE9Ln5v6EXSa8N7
P9/WEIn1EEBifejaCM0LLN+Atvhd/Ntv5YlWNUzbSqzQEbknZe4bLlKtb8S9vK3a
99V5QwQ8BsShLqVzWd87fpol1myVhVKIOU5NXSRfm7hBiK+hgm07+wDIDrb4yauw
uSkrG7vD16AA5qLM3mc23t6jCFj3DuwlBrLBrbQXOKzNVhyf0LsFUptZ44ubILl7
yDlNdSDf0yC8Iz86OGsFQj3QDWh6v0ZcTLFCAePpInHbbwrO4hoI0/IkcjYI06HF
Tp5kfXWiY3f/zCaduN2om6iwop6o03oIwRRajoEovxtldonAqNgU4Ovp5YBK+zLx
/qtm3wxwqq+PvTMn72l8Zr0LHuxOgGoQG6K1DHfZVZC/elp0D8gsbJS6m0cQgodT
uAWAo+4c1Eqz9gmADEC0gCnfrlQbsfqH0isrlvU4LnLGni6UyV30/58vjgHzqSV4
QT8+aRAam9tssK9dBRXIYPjYPlRDSIBaDgH7TAP68Z9An06kiIuR2SYk0Y612e2p
dtQenPrYY4+gxKzulqQHKGF5RLYF/eArvCeIX4jNDUDiQ7d1rOui+AOQzkECuz78
mvm7Pi90RV72N7d8roBeQ9bNjprKnabDwCiFFsNiVI2qNHvbTsgWd2Hp5JAufcBh
EFs/ik04hZB5NqxgvTgqTSwq8xGQb0ZdZsiI40gV7fCFyvZzdmuxCSC8I/MSPuLp
cR0F9i7ysXKcFDyuzqbUB12u3MK7+KK0uBF8p3e9Rkj3BdyR5ts+EpJGYsNswOoU
ZP+2c394anl6FwC5G1NVw+APuID1A+GXXOqdo24EFo7AoxjOifwyvODRPoAbW8FS
C7AihdjLs1Ldvtibb3UJ0KHF03BkHOKAd+bTMmVFTaqwbXJHUybz4Z+03uIwxHy+
ohp1azY/meXeZ+l/NPqx5SxcQV1aBju8yO/Z1BnDlohqZgQKnPinsJ0QpMNhxVwK
JAjjOjPfC5VniaV/6z7PI2uKTWGGmU+dAndshDco2FFlbV7cgdsWefe0kLOjnNWC
ln7xN5xKRJ2VnfkSgatkzcZmdRHcK19XCnvypd3DCyVNozVFkED+BnWPJzZHLXz8
9wllkMIP9UHumd/TClbvsG2xU48c4UuXO/pOHmy/sp4uOGHAhGoazJ9NJKrSUWkv
OyF6Zi7/Fr5WUSOu0X7ZbJL3GFZ4yY/5hrnr6dDkjPvPtOeaJlJRFvCZ4jqEOD2T
YuDi4XsODSr/BywQ/y2sOcQxyk+DALXebtQ8LK2+4Abd1BOSihWbxRvAQi0LRZJ1
9CMY1Nd7D6Hb14AXJy/Qm0ESwGgLjToqYi/BFjZb4lW65cOM462OyHQDHsSDwt2/
R6AeH69OtlZj9rGI7YV6SQOrbYyJkBIx4Pb9ieeADuJSiRdoYVwK535RpPwRd7kp
0/Yk20QDNwb96XR5+kephCKVFXhrRSdC40oKM+IDw9EnAgBTeVD371wZrYpZQ2ZZ
amjOcYcFUFVRH1rhtApgd6A0S9PWV2KYVNvkFMtLCfHEtzG2hBFkAZtih2TIi8v7
IAw18/+xqhGUfxt5e4WDbc1F2LvwT7oPzAG9DjP3+ZlXliQP9z/SHdg8WOBe9+G4
enlLIMYqw1vaMwvWwJ2ho8CGkGYAPSWJJSTyu/Z5dPNKt7odxu6z7T+Rx8DAT4o6
4VNkEHCOYzYXDgkp5SYlsGMLaRstoJKGwaVBLaITvGaAgaq0YajTyRTdr2hdUTkU
xMjhLTUxfaZ8krWrpugZRM3s66flNSD1KaXplerLj2Fb77hehl2OwmavQawGil/u
n5rL+XbBjv7Nex6S3CHfYeE8QCaN/mItYSPdTemjudngXmLkHlGibXVkszh4mACI
tBXGMpIeA3EynCorUtGJ2QD1JdZJZIAbaPtlwCldn2VFcvoj9vqbIXBbkddZ6Y4a
+oomZF75cyGbXqtgaKL3t4jhv+xQ863T43oMFdEjOg4oSh4WSmG9cno63DF5/Pt7
DRZAh5EZQsd7YrUfNPJyIpJUTGIxZaP7Upt9wmHsIjQeCLDpwE7Wj/gp9QcqP1kU
zR91Wagt7lFLohyatJNrye7BFpvbwr+v9HaIw98zryq1sO8t6E6jmFBSJEGDKf16
TNkSkpOQmKwyAKXLT/p2RPaY6erHtnGhcEAU3lZ9+4tiNXhLyozRkeYGKoEawGed
9hARktC4jyeSefoR2p0c9zYB56OC7zq8/kV2CDGxUkPNaJ5jkPVeTvUimz+OK7Bx
OmMcYDyOaEawP3KTfIT9F8rgAoOR6rBJJXoiNb7ctTjMYrG5XCX7Hd1ITysnCRk9
5nHFa+YkVki1FIxSh6x/ivQyLs6irmIaDgndsXDZMG+DKlZUsKxcOTZ6cos2s20l
dDjNYCpwUu9o0NN21KQz1UebTBYiXH+gJu+t/GLxGD8mFZFJTBLV0MrAhWh04RlO
+2VbOi9Hi+iqMyQYr/eKFJuGSvG2zXsoAJweDAgLvReEekXLuPiqs/bjHFh8IsXS
vm74uq9WeAXRrAbwj967m0zqpnAoUJdelrFDfO3YgaWLf4FKyyqguAFSW+jn4Qps
X5x5tlcGPJQ8+XT4hkFxzuDzNNnrzdEMjgZZ9nhiVPx6J4RIYY9gc9tgFj4UfTC1
LULHJYh53hjqj7d7Ml56wwpg/39gOzrLnSUnhjfu+qoYbr5VhubhMx34EZL0UEoW
gLT2C3Dyf1BU1FfvBcBB16P2CnjdLAZ5+Xqbs5TBQFn948k202Ild5aj2qn2WjFE
NhrGAJLpxv0fkHv2YwCEfmA3jRpDcawVCkv9oaHUHZ3e+Kxi3cnL43QgRLAil7XO
hcCm5PkJ5hXIftufsEf8QNP4afHzIh3BbTNafEJlC237kSinw+L3Vr8yI+jO8sEp
vq3dhxIulFoLdVrWOUUUf4P0UNslPB/sgnAx3m1DiRJ30UNkp2LL2QYcZC27GeVu
rykJmhCtAT4tiP//iYG7EaHA34xXloBoGQA+Y4hr1VuGPkBdqiwSb6C5p2ttNW5O
pPG/HLg8dCz3PJ8YA7uPjTUwZ4sps0pHe4JtXK75QrHpMCxDVq4JmBxjgA2kaieZ
8/XNawO6i1bGuj1iYvoXssFje1WHBr2p3qnsIdzmjVNHRPHYdLu/0OcfUYv3kNe4
1ydACX8J3l2mIZi1bmZh+arR1Hl2lbMkADT4gK+o93mO21+xjrCNcKvpMjWrKDG8
ajR2kOhblE1qe1XiBhEUYMDZz9INRjPqhqmU6gLV09Vf8U95EWtwBODFqzAwFYyA
XVM1oOeR6GyjgIEXxPidXup0lCiPWHYYY+rPymZFVqMe0eNWxA3dlg6oiZqj4m1y
nU1dsSG/blmmtTfCw9MZjGPLQg8erUb0bqRQXU3zB3PZpTjdE0oWWoVC2uz80kro
zHTW7ncsU3sfOmCIx06E3u5adO8Tak/Ti/+QeaAwZtOotFBEj91miqCJe3h8hTXx
RO+I1E7ytib1x0rcSn+qxBkn741gmZ54reZcEBP8Ai26VrXzVyTU1vwC5TN11o6w
wwDD+dvpr0iICwODf2EvODUPwaiclwzfgmQPStiSg31rNS7eQnq0syxIRSeZybzw
g/uF13EhIQm8or8n7uIrw6P6cROmKqL3hRIC+AvXIW5HJS3tj3YumtbkQEde4dDG
elerH+CbKZuegBmAr5cesZF2HAYzBowy/w/FMWhqYoOJTHPIfWt+Vo4ektukBfXI
E2cWmtk6A2Vr8tfWAwqmdmYJ6g13dexXAKomx3Ot8ahaFwgTtiiapbkpaQqBnoQL
qWU8MTE5ApvL+0nV5NHS+8JrD7lZcCwmdoypZ1bAHfhyF8GT0IWuQvaWLKWRc6k6
P6ho3JHuSZGBqsDHOM81Gm6H3s37Y2kwFmf6DLGicGs76foA6S8vQbol/XiHmKj1
uLNvzCSH9KMv54B8rul8SxY46H1uHGFcEmieBxfR3FttufCpt3rIKERFy2VquoXB
SeHCTJPzDxsB6E9YG7locuXHrwFbv3l1+WWQeAD+1U/lhXHvlaBwC/vD3At9qevh
sTYVJk/sA4s18KlKNPCNQZxKncuqSLMnFUzW8ncxe+wlJ+HtULUDPoITvMEUpP0g
9yzn/0qJGonHbqM9nzVNikh9aPcwpi3q46uP7soM6umXAt8cOiIRaxraiO/kTKZb
w8cGZFjW9DROC6vRl4Kjii9pDZHxkdnjIH6hTKTqHzaQ6uqgJfl9h3S3jPwq+ffI
AwN9ks2Zex7cWuBVsfvM82UGDyFBwLUxP5lp7tqwaJKArIyDTf5LvJNR4bbyiRIG
79nMmmFBcDMVsqx6zivpBiIFUtboVtm8aHWa5thT5F3BYm6zFNtgPOQ77eQzjau6
Tl+CUYo/lucgzLJYfEiQUlT0+lkxviTvphptYyILouRWbzqaHjZjmCDxzkYMafh+
+1zFeRlLexL+ODa6pd+fKtH5WzXvXkiQfI1hNH823pOSlsInFkt8TpHM4dvHStsi
E3FEeVi+NvZ23oNBVugDP7hXfs/IQPXyhhavg3ewaT+8F+x1mZZIGGTcTwqObKCu
L74An2LNiaT9Qg/oPKp7rd4ysvxKiHdvWjykGhMRCc1cqrLonaTPDA8k3ad0YirY
o5PNasmuN77tx2u3/eVaYz4NsFqGTV6qFp2DuJ5LjUrRYiIkn6V2KFDwe+vpX3+s
D3A+RuSgConLrdl0xgeluNkcbCx6pfubMquCQ7AwBPJrKSbgGauGkpSbVUzXCtSN
V5f7j1i8ApzvB0dEw5G1/QJZ2nwFoRrOo1IMPGQEpuoQjX5Ml6dX9QcJfAiXTWJE
rMRom98hXqc9NIy4sWXqruFHDs3ZyMU97b46fec9D150CwuFztSoJyvEEsegBQh+
VGK9no83tt1Q1oEo3B/8DTisrRo6ARwlqyYmLzj9r7hCcrHRs21qQX/LCy372AOZ
Y1GgXWt7+RJ1xu8rKwPxsksdsqT0PRPC5Q5e/jvohMtJnejnXWBSylnl0MG5dU9m
vDVpizATxitwnS9xELh3oWEj0KE3aYp0OVGlQDGhzX+9pKcA7HXLoxFXJfUKrEzL
bv/Ad+5/lIRAB7uNFG5NsNXlsxboLGmzrRgRe90ErpQ3BhejgyHwht5oheeqnXDq
sDLrT5TG/UX9Xab6URmkL4zD732bttEVY05fwwitvE5v0U5IaFD7fIkeaqgCkl0F
/gry6cVipkIdeuCnBXUICppewYNBEv2yBUh2e8Q09w4i7Kk7EpKmk45qJcW5a32F
rx+F9XyBf/CoTRihzjHeWLCUOgldGZSta5hqI2T4xss01zcszXeL/EVIpiXYN5cL
cl3SapvWBZ3Nb0+p8V9mHTPMbKIRyD70veg9jboysaah0+XhdTHubxtxHfZykvG/
TnOdHYRIdYPkQnp5rQ4/Z2YqXUpb5nfH8NczFfwIgNEZ5K00e6iMTc8MwVLj/niv
tgJpv700EqEcC2TckACboMUcU2DHcScf6iu/2+a7v1bjuWwByxtWhOhFAc3nbQCa
x6RAO56to5tZdWvK+pqHv54mShNQD/6GJ0ZsdAPVg/0OKoUWst0XzyBQwN/eBP/K
0xQkHRSGCyIeSK6xEvBWmKqbkJLWh/+9txolfPakRLUQIwPwpCn5Qu/qu5+yByEZ
ezfz/ZhPvB4VadsirxV6DTTd+FYVnHVTZbz6KFVy6sPwl4hWPbIoy665OKa94ZHI
70O0d0XVSWepxRNva9Zks8XBmasd+/N13p0qVh6Z69lAcREy+id7MEvSYnRsj/pu
1EqnnXWAdDoTNMv4PQfqOfF1VLUsd3PEa7x0p2tI439lzlUyg3wRFF9F/3xes6g4
/FzhPAtLyfiM0Jtq58sdqsrZcR6DUZigQ0sm552p8idkr0+is4GQULCvglFW2gez
rCXhWqMORAAie53ACQR4xbT4cihDjqv+duNpgBxaH/Zsou0sV34mvQ/hG2m7gJsy
CpHKgrXDJonrbRx0XlUKwKxuH6f4gYYsvpUASMTcjSmvR6r/uoR7FclxEc2XR+ZT
Le6sujXs4jr9pJH7W5jlbPrYvd6GWR1bsAD3qwdTNLB7EOPL6JYoDW6ldMQnEgkk
2CDNCm01r/M85fObYv9S4kjvBTLy3ElMecTQaXxtMvILQM7R/F4PeVSxyCseqO9h
ljXnQWScXZfZCzTS3uwlT7QrrpEGc+SyNvScGvMle0sUJLAJ31MC+1lYysuoGG3p
p5S86XWjkhr6o/4iQOK1qDkIhluHg0am1mVHmfHAWX6fsv8xItDb6M3lvJvp07TG
EPqlhphHXe/kYSFQQCQAe6XWzg7XxjzjtbdytRkyCoxCWf18BH8uPi4z/XTGSD5X
+Q2fxjZkN02D75J9/mjhwd8KL6gYtxTlf6cXcvElXt9dwXshksfFfyrW3o4w47+j
ZDC4GXToBZssd/eyCwynxCIQDW2m0IW1it46A/RWW42u0vUD3jVSoADZs71YmzcF
hBmNLmppRNEJGhkd23lvXfCFUUiLOVMtn6vN5GDSQrfx9fLn2HsGGcvDMaBFTFUb
azL0Wo5ogmjCxD0ck+i4fUqcQa1+HUjV0HLm9Wb+CfjhOXMRwWQPlJTnPTslpRQS
LBVsXkfSycfLrjPJ/r48i61YAQL9lZbd49BQh+1gdnJpYigsDloLKdmP20i5qzTm
IpGK2BJ3dJvZj7lBcB5/gdWLk5Xc6vsmRY+YQmXpMXCv6OO79/F0xINbCAyQEDE5
IiwBTJVk6Vk7h/isApZiw0EvGNwizeQ/uGT1Vw0KogczFXIwokXnlSrqVuPqoP4m
QH9inmXmK00e7ePWx2jIO/okI+63CIuyNSP7f76KFJrpjIyrDGi6BVEr2hyn5kIu
jGAKlH+F72TlWP74Sr4LKC7/EmiW8wc2gL1grPq7bK79f25S4noS7oWomvWGftLI
MQjt1xbncIdK4/3iunT72oKf7f+A6zwMCtDOtqUvnLJyV/D5tuE2a33igg1zqzPK
o8h8aDRwkXrYZM2BpzenQNk6kqnL9vuSf4Yuoo0Q0CbdI6lzkYqIXrCuEWlPVvp7
E6PWnDRa4M71t4mUICmQeL5PuyEQ6K/bfxHkJsW9QQY5T+p3nlpvZJTjR6oNmQQo
GNaaM5FldYmuOqHu/zznY7ayFv/iCnP01csU3hScYiSaZ3Po68vOcHOwkk2Rx+XX
InmQHkl0eJRSa9j60YfFt0xR+wnZ01rhPinaD9q4H6G4xpuQuum2zVH/E9ej/wAd
/UiAV+5/TbYGKriF9wZkWb9GfULrQ4p2pRS0Msiz7Yn8q+uUGnRYKg/M8ysQ2B95
BIcnPpv9nJRLFA7BVXf9HAx3D3c6bGFiOb5W3fbyPbLcAOlCbm+exTbd46h9SETM
cy8yM7e0uhGEZ/esP+2DCiRirmfBt8JNuXj/N2DZ88PwZO504S7Iqj5Yw1qv8sDa
eugA9pnKCNQ5DfqzDXy6fMFKUjR76e2n5wZ1Z0BkQvSaiO+pvQyVstM36AnBwTkT
l5njs1wFsQKO19RuBonoJD0iEg403VbkkAZkasRfqGKZjHtA3qhRDoLMZzEYEQuV
B/W5nHC4Ipb1j6i6Gon+VoDjUlSEv/7vLsx+6d+fF/5E3LeKApFzQVi+/GI7s8iq
K8MKRChYeXhqni75uxDWP2d0+PR6o3qIZUCeU3PtVNfSFf4t3Ud3+uFk0cOsr2pa
7X46PcVR/uESI0z5Ps/RtjwOhELxT2yyzSK+TgcAdTvLP/6HQmB59WRhiN5Uj9qg
aW32gn9XlubM2SxG+9GXZ7mcYJZsy7gWKDfE/Hz+IXVqJ7lqVuB3yhAbJx8d4z6q
fKDy/vDq6IdEx0lwWjufihtKEERR3BS2ualwTKvm0vGTon9M7a3j6etVJLNY+E1Y
q3ZJdsgQA3uNin4inmIIfVYnFIWvaZ4fsfT7RCTpEkNaUP7SiR64+il3uDR6EYIM
Qvyn4+lmOVa3vqSIt4V42KyJ5/Lhx+6tNx8B7llVo8yrcQTKLPHL9KYGrV5ZTmlK
6+VG9HyHpPZ1RGjLdWy6rJczmzSzjTrCp71afyfenRnyvGEwkCy9N/eVTKjEnFig
OKUZ+6rXPdPBt0adfbhIAqXwBaOQ/8N0ncVz7eTy7h17jGbau1lzoazuFldSRX/v
cIZ/NixSiwqb7p0RuNxakVHUWIm1NqMJrM0BkIB0qkVOApVSW6lnwICUt0HN/S4i
GzsmGhFlUhmFtKC+2XsjRAnfE6FplZ69SVzAtHvomMLV0Rb4Ypcc4Z1Xmt9VofwH
IxKO7ADDbvQjFtEN+eUgAW0kT6WvgkSo/dVuocsbmgRl2puSdkHd47hu8HSoMVRJ
yOIU3Kn+ZRfwcPQhY7bO7aFA5UrI+1hqXAW0Q6JjqtNwLCce6nc1r9IFBxT8Lan2
SzJYyrJWSuCSJ7UhaQDFJu+9AKXyd8YATac2ZxsogcpNxUD0TWBsThOfiL/AaU5m
S7Si1SryU+X85rjNx2r3WG+RVrQE1i4tQYjQGaChyUwOOAG7avm412lk9+93mAmw
hz/Ut2I5nDKJTkx4wKWa3ipR8zF41re0AlD3PFciWOvNkOYeAJuBQr2rJb52l0+M
LI7E38n+OUt1MXn/JHxkhFQGbe13lmXETh94VT4jMVgwYO1k1XngEEb97CmcTicF
ia71Pl5XVli7/XAc330mXW/1EHMU7ZSMgNoJ+boD0DaoiHmhPN6T1kzapN3pOAF8
Wy6klbBSPDDchgkkXzK3s/EN5njLafQgqcimUG+bksaD1WZZ/o/6Ecnynj8g9xyX
2F8ujAsgRUo8j2bEsgZdzMCEKoi2RMKwVwo096/Yot7k3GgaVNoWz71NMopMYM3K
Gbxi5G+zEaqWjMt7F4Mz6zQEulo4850RyZ5eTt2Mn78MkAOCJm2kfDXwxp9zwDz0
BDKmb76sb6pZvZiVPJeGXz7SWTkWs+bhJHV1oRum7dep3pjbuvWJ6r+9jNctMuT3
Wof61bM9wlfOxFyFiZ7TsuRReLJUx38842SoBFU+v8UrQh6uv55TJHurpxtKL0bZ
qTVfvrowz4pOmqL7sLgFRYzYdHmFpHurjfPX8335YImuVRp7Am/r4CbYvsVdAcze
6+EAqvtSQfdInRCXTOpagN5ynRaw8oLKkJFvZx3aE4iV6k+1Rw/2eEG2IlsWRAaY
Pdnd3j7syWW2hegWZZ48JZY6VAlabWgpM1DOAXj2d8uHSHJW4oNmiOUOqTYq845L
4GhNwNsbsJa7Tg4hMuHwsfFeO1I+8Rh2HVgrL5JMaGYIHGNGtQfLc4KnV6cbCt53
gqHc1E5ftGyLVoQXLULnPHgHgLndMGzhP5zhs/kpED9w5Ez4joHjR841+9f4sgqO
RqaAKdLYSKgyDCckreQY1euBpSnoFb+ms0YnAu0+89ZBVyuZfrbvWaXlIeMrVHAB
6aqhTX0MtveyyYXZO1YMgr5CfTsPoZA5NmNFHw19MfCaMiv92PuKXFpZIt+BBgmR
60EJj+JVr9BOayu41bl/84ulNpG+kLrvdWMdjLgDp4b6UfSbFSqZArxKP4olD7iY
/Vgq6oVPzpYl6dJtaf22j6yvuw9Us6Onb1F7H/p53CX+T2Ww+USq5oHuSp8ns+gW
9bqPkJiS40vLDcKurMBrrYthlUWnbA+bX1Z9H6/nVPNe5mUaaYZFdswxAdpTDcFH
454h1uCQHr2dH6CNO7mU+bRfczjBiLcOE13UExjEhdI7iaVIH3RCmx0miavsWv0c
49zwPuqu60uR7QaAm56BMP5z4sdGIE+lbOAOCBVCKOOXrU9OLAmoRCzNxi92eXlU
JHVe9PlI991jfk5deC+E4TlM9AdpzDQGwrMKGDvipfi28QlEEFuEkJQJqdxWpf+x
Hsc1BnncebrERrZyQBb6Id7/a3Wmi78ZN7hGM6UJ7DFrv8w7MeZeKysiXtD/VTIo
Nzuisf4C52agWW8ygk0EDJVcEMEBZ+/OioPdPnbB7ewoMnrKLKYkPxGCnxqDFbD3
UUO1ujrbmh7O2D5KXKiAku6CWR3p6weAnHGyOMREhGtN5xOSdHxvpatUuc5Pihe3
MiZOQXp3r65WnTUM7jknXJnGSWHsgxqx0doJXb3yoD9wBC1cH95baLEIZNym1QVV
lL5vtaXD5fdAPFAhnZ60yp/kteXEaV387dxMA8fwa9ksYGcYMhrC4Tst3H71O51K
v25pEJDokuNEqF3WzPhtG9YcXX9xCPbxPI56ORFrtdjnIjwfHHPGCRm4uvKyJjWf
Hdn7fgKrsBQUw0sB9jcaoAyfJyPTlmwDqjbg+h33Uw8NpE0sVc+Fcl82m4RqtYaD
s9tJ5Phy0VEo/HMo0dcyehyIVe5vsr607V6bbp2rwABau5c0/YB6cKRTDZh/zmjI
9fHUxPLUV3uCfDpTFaGDDsYOnr0tDGRXbVHFikrRhNrL7ZRzKl7gLMJTXbtOpXtB
aWfEAYptD7qx0O90iIE9IFI1ClXAIQ2ogpGQonRdZWo5h74XE5pe5iC23mH1HXHv
gnHGn0ytcz/n2Xv83Qtt0EvKRFj8MahI+hLkqzdTroNbfYBytVoJlw5t3XPNhrJ5
HHrA/UtTAh+sjo1jss2iajbhgUinRK+BxZyPd7sKP70vkX2usjUtEY48Pl1705nI
iFWC1fy2rtBv1BxoAGKc4jCaaGCdaP0zra/l4T/A7dAvY9BO3iNpl6ZC5HNo5lng
3uAwrh0l9CunTJVzNeNyfjJgnRZy5VU+6TIn8UbxUZdbEjlCIhEx5NPohHD6q/y/
R+ER+vhvlt+LnKMeIXorsV0PYxqrBj4rhC6n2IpcMHMjuWc05gJT7d6Obgq/4PIF
EZqLX6hqkflJsLnpOhaG25PImv3H6y34uQQH+ZIdE9Pepvg018DtpT4CNgqhpCpW
U33nE9WBG40+hWXj+BKt336dmFt0otKCUbdsJ84aQmAv1YLWIp7V3JetrtRcIpRn
WlsyyisTa4YZjsPSa8mWTKEOBN7/TlVJf4eZcAPzaHW1H/VDSHaHn6XScfR4wJ7w
i2dMXwYT/tPAdih463zGzIWh3ieQenlChtyarRfF8oZcCuiwHIF2ae1bTC+mIcuM
4PIP4BbNWVGHeYq4ZFF+51kplvxEFQn3hO+6NRXDulycbMHPWEVmpPOlLYrHJF5W
qAtt5uXTv64EfysKNZoU8PtC7NXoL/OiM4Fmw/9hatax1MK47+wCYARMzjTPVlf9
QXELGfwQcZ4W0cK4UVvvWs/vICvqAIgPHQmC2N8PyUBo1lRS/SENWFdK3wqahA2V
Q27tZ7ayG3YMR72I3K95C5X7GTa2MaCIwfIo8AkZAdb1dc5U2WX57GmRv5SDe9OM
EX1/NQUNPlNhjhV/P2jil4ncvwriBSzA9MR/AOkpsslQh/WlVZEF/M90GEc0ny1g
7/uGR9plTSjW1naW+7fFSVyf//drvwfUc3H/VszbrZsqSmJH7VeYi3CREOhFwB6t
J71lMmaC7+htf+SZ2+8fPzz5k/dFrKG1JNNb7MkTzep4QNcmVY4oAP85xl1iNd9g
yEKtTBG0Cfyl+nuGqaPIJqejQ30ZekyEcZhAUMX5cyKdyfKDQB6nRG05JVgZfni3
k4bTrCELF7CTY5Hj1xu7z7+/iH5wzuRUjtsq5RDhLZTvaWXRhpJruMBgOvZw1tUX
QpLLtE96JDpBFY1yZ77nWSNbIzs0yT5w5wVwb6mBFTyEycVwhhBuvgabTDcVbLt6
hFkJGAPeBEGJxeuTE6AGTbrMwWPdQLNVbnq5JD/SoghD984KeBrvnwHmtVPz3N/G
R1UBG8CGWD8rSkoW4OUtdIT+vfWUeoEP4Gcbq5XY6VYX1Q5Px/MSTQro5CyIwrE4
pnB8jzPDi8D7WmPYxkzQIdmODcge+cBuSQ3u87RT5rjg9qr3ZD7cmX09movJdeGh
bbK7woBYphvGCLKRgTs4TNfIyCpMKoFAVak6ZQcnW1kigXswG6XNgWROYO6iDxm9
teVi8VKH6MGJbWWs5aKqb0E3teuuUzi5GCuOSBCiO65fo1l0n0RSBZTflmJCbUmA
UytNL/iDMBci/jddYOcshkPDr5VP5RppBbdglG8MP0wGk0KBpSVRk7ikqjr3Iy77
e5nY/+7l3XfzChAGFR9M7SZCOT8ou5pqJcBS9zgrlqkxVa/SSKFk08YrhZwcsX56
JxIR4/S5SwjsMTc8mA9jQvK3yHNRGFZjBczDqXqLPcq0MQu3Fi3JYtuc+w9G+UUm
yOXpuR4ZhLzQWVirK1SezSMQes/fYzm50x32EF+8Hxgw05Nc8NhEFVP1X4olhlPm
fLUUp85FCKp/3tN1s+Cyi3pu7A3tdSdI3cErJgusLtKKIuXqukCbWU+BWpHvtaYS
BRhr06PeJwYFxNJtPPZNpIa2lA0WlRxyMwcuN1IOEPHIsrkHqhYONRMK8V3RUFNg
TB71x/RD/lyFcDqYrA+A3xmfOIF4IKJlShktfmgH4yh+didNUehckCRQexD9KTYF
z5mmHnQOmkwYVzIBby/FBUzU1xqtr1VZkNcDg1Ap21Wz2Wz1v8WXSiCqAHOpcF4w
ber6TJnqdSIlBsZfzcr3ccYvj2HQ/e0DEgFkUJ2UeTZNEe/DtR59OMUjN7cP6tAz
GltVn/ODyV/ekwBF0YInWa3OV/CgUTnn+uvRgd6/J5Vgx47iIXLHGhJpFjw7O681
mz5HXzWuiY6viCOZnFTLnhlVUbrwkLmDpUTNPqe3Qomm6160yyOvUqj5NdVc1USF
rNAVGD/mhWhhFk1887gbGzlmXqtN1bvk6CYRoKcJTZQ8eTwg6c81bG44viiG4GKl
WaWTIhtgC5u2/hevW9+fhMFEIooorNYyEajv3ZsAuRBMW7DUSkEVaVzD0464FlhC
XlF1uHJlBVtzFDboaEbIZ789/yyNNS1aqgQyZh9bPYGNcsWccN3uQCcmXm7bzVKQ
2WkgzwMpY7zFhQjQsnQI3xnuy8AxU2jGSTVSz06+Hi6oGsJQPnx2NOI4ymS3VHyi
p+2hjjRW96OCW7shqPXEeMC9HF4klbVPcGrbm4j/ZLpj4c4J0A/tmJ34yuyl9mHc
r2l8p+Rzut6oxiLexVWUgWtszFfINKtoHPocCKOylF9gZ7CT35iDiR3DB4DaACcM
JZe7KyJdWuQglgyjtJBlUFau9Mn9dvQANA8hhwbj9XvY58jrQ/SfITFLmmyPZ0dm
GXuf9dTJ4WGO1bbnfcEj+mKDkkHgbrqLwZQ5B5JuV7VjyEq+lJFMiZdKPgxYnTDV
YBtt0+lbvAkUQuRb13p+4W4Nrp9ldtC0FyZc2q/3/66w1psc3w4mHyxkdXSQMzPM
RApn+df+O0NyqdyA46P9JkdjtbpaKPSR4SVtCHZlsii5xDbOGkji9FsZzW1WTGrZ
zS586/cRhC95Po3WhHq5llE2yJwIMQKw5mgjcpVYRzJlkG0PKbfyR8hm4Q3ip90X
VmPvaQdZx2CvNC8z8SE3ceTenWgFmNRyjZX9/V7H94F7J1lphNit1e3zMZDvKVqD
uKPwV0qTpRbX4rIWcImFCP/OLEIoVqcJJra+Fj+ht06x6jx9v9VvCCEvFFpc29Dd
E6C69mAsNiFvZ7SkGuX7Uwc0qpvJcba5fQyfWVYF2pDTLol9rouvoF/pO52DkdaP
hu4yqEVrEhklM5CZ5Om36KTUzGft2Q7e8xrtkVZ9/EGKgFnl5L7CKD85FWW6JuT3
oZjZPkwZBdHSipSomaaA0oYBavjBRSi49jLHh8AJ75UwjXX1uPACAZzaIK4Zq22g
jawW5kcBpbeNdM+OahPVTM93AudBWNmOcCUIT/LiJSavvxes2IkSphoMqgpAG7kH
Cu+GVUr4ygT6ApQQ8ri2QotVChQSu8eZt1PxXdndmoXMfxPAq7rijbgyM9suHZyq
2AtSuTGztHIt8sR7sbnibpv1tSDYSDPAVZkJ1eVclcYbBHCE2bgvnrpoYQ7lpuQV
uODVsbh35O4BOo81+pPIddH+Bya34JpdKKWD2/lpYL1d7quHCcJE7cC2p4693L2/
X8pfLsQZYqavKtkwFy3/9kubxK/C8nOnEFuj7l3xFoGaPV0+7aDr4G5j7eCBsvaF
81BBWgUXtadayTynV4BdIAFZIt7K0TKXrMFGow64teyFki3ZBE78EZSU1+ZdOdJw
23jk4JaNIc+xltlIDXQxPv0NgXBZAOqLu/gKYXkcmjv6TdmVVeu7vochP8HjUDHR
LLI7sx0azQxOhAhK6qVrOB6lNUot5uSe9UrIHYStE9o8+wal3a4YLgqzsjfrASYM
3P81Ypebg+6biFpNT2CMl4Zh6btyJSY+1y7Uo62pMUpF92tUv97pxjQjGWlLrviQ
fMa87m0NMwXvsPhS5YgnTCeiBjjbkcFXywvMHC/KBA8XRfa7kXcC4lg1URrx84xD
wRC5+1d1sW2UXElr1NpiWttktTtg3Gtmcqch3zdIJwO66DJNpiYvuu+R3knCuYJ2
G4XniN2FCTWYZl6SWB3U5KYAdqwh9hAmW96nad2wsOv/tuLN+U1/IBmxS8jvOJNF
BDTLRjMGE2wpBhLCdvvmg+pwri3htdtfMrxZrbgHl5WpbjIjWEASx75+OlK1/iuP
sUxhDhaVjJdqEZikg7fadEoFj2pK2+KVCde1INNpnpxHIHT3Rm/0/94L2vEoUxN9
wvw4s5DsAkK22xs6xnTTVDIlifb32MJlY2Iqyfbc/AmxFqA6fLDDcL9h2P6uFz/2
71tWjcM4ECW27nGcwxnMQy+ZQukFH2poM9Ov7KT1O4bqW+y4QSEKsdYFFhMaXP0L
h0hxySoJVmcVsSpT09QbgRFtH64naDFYFEYyRWfJ1s9P18u8jNA0wcyqzyBmKO8n
nhXYzNII2y29En9E0TC22AdCvDaAymwGPZ2QD1z/oRr7qRtcCtXDLZYVozghFjc2
ed3MoMLRyGwtDzZ1keHxf4A1PvYOU0n5g7HCWn0AO7vKvmuFktVyDxq0KOyQjN2N
W5qCUBsEC3Gg/HtrgejFBKxa9ELFRlvGXCeS3WCVgA5ZeTF1A23y40igDyVbiSmr
y0GeAbVYvNqQ9Ij9jOrEIfED2RQ7AjF1okGa7yYxbf9jycwQsIQLg+RsLYRK9TuQ
427bc1oD4mUROSZ/jt4lQtE0oHj9DFyneN6gOame/vOkAgcmIzJvA3FuRqvicc2L
Cy9TbUcJ2JJKGd6yDhGIqt9pRhcC7Tz0o4ZyLEFFcL0Xi1syeZ7Vyv6yZ5epMCT0
/0BVwNXQxV3HYeYtSfj2crwn0dqH/rghMAsMZop1zEkV3Xrovd+NZ5Q9EJSvdhjC
CuMKjiRqdWRe2j7+fYoPuuXMhRtvyV0yc6i5FS+0awg8RCiD05I9+WhRsEkuzz4H
3kXiYt0o7AO/qbDWwfaoVdvy2ovW8Lc5OtM6FS0hPiXq3+be8h2MMm/BSuMRDs0u
8llFwrihMscc3PcZkrtZjrjoFW6Dhgncw3N0cyvYV+fSWGw1ko8SO5bhHaRogrpT
rKU8OdbK6oyiwgV84L3+bHlXZubh70RqEob4ZYFi6jHg+/dC63qTOcoFv9FMEmQS
dZjV9jkiazRQfJ4fom5pOU924BT04OxMtOYLwM1Ey5Fw5/m5bTmkyFX7WRDHrtqu
tjLRX78eS2IBtSFu+2202arokTxFIlSUzraWvLLAX3i7rNV4NSq1Vp124SIO5/8N
sfKuUk2HG5mJbzHjmPVkeZpWr4+VKI9KkvZsFuIoLkR8P4H1h1QttkbnuzlJ4Tqi
fC4h4L/YOxjwBBCwAirBmWQR3FMtwJji8r5iy3nuDFPLUTNWeDVKRYopIeMe73dJ
Xv4I4/Enxie2KZ0A8h28yf5yIq4s6DlwgUKunwXck2dRt1iS/ufskyBUVNs15mm2
yfyf4K3kNpoB3BlwRVe7MZ4MvU4twceRXL+yGhXTeN/IjcWe5uyzsUHKz1/1Kb/n
W4ArHT0h5FUvpXr7CxH2UJghJi4RM+Ef93Vv1k4dgzjjrhC0RPX1QpEy0FqSOeV7
Irl/K5rXW27w5Ldhm+HAT0K8SHz6xtWJMdZp5mGthTOWKGozFO1vTShY2oXgBe0C
Ii2B77IvycvORo9eAsPzAtT2zt8kzdj4FM4DfR2XtVUcGF2VtcSoxo4YyasGhSxk
kXiB+p+O9bsQQtLbF2ZFuW3H2m/t+R0bFawSEnn7/prfJctNV3EDFDAJeg/G+K+s
ZgGyngk0QjD5qQTDIw4DwCW/flatLBav842I39STtfHse+34g2gS7iY0V/VK1Wvv
TDJbSopfQqrHg/Ww2+DjsHRKkGLUaOMKf9q/qzJdRSj1/2B+OaWEN5tCyHMCYO+6
laVVNcGzwMotr3jcUq9BUH2bCfAo8bZYTPgLpMqhem7luKlB+A9Uf5QsxFWo8YLn
yXnmSyYUf8a12c542dfhUFmXwqrQ74e/B5GVodkuSLyj0yYW+Yp8yvTGyX6kF21d
vLy5slyZZ9SPxKZOjF83Xy+5JQOr1A1epsze87JhJ7FrQIMucGQVJQjNSMLuYVv0
k0RgzeJEK+gbSw8UBVjl2QHePcj1yophHHrL20dfsB/72SUyAVKWcvNy6tiVJeO8
mH/XEfim5MosjKcwJ9Azuu4QsYP1tBYm0r4w25AQjZ1csLrWXECS227NeDSBNMUW
RvZoYLJ1LMz1LbJdrz2/dqHTTIs6mQXQoQagbqyc8srxEmcM9+vSxuBSxbQGC/1u
e7dlq/P/VtN3MvUQ3Q6BqHQd9KYFTTpusbgSLJy2Go6dPDGUGczXaslm0Qs39mNp
10Ikz8d50FDfmQ16i9gUIaBszO9IsRy7KbX4L5+4uSCTdMytZiJUPTaU1gA47XfY
wuFuxnrxvjbzV2Il9ZguvSPLAEuVDGdvOhfTrHIRmEslBe/BGrXE5T9G9FdmZ9d0
7JRHj80eLB3Ud0ZkzbxnnsFf5Lc6W+j4joLYF7i731muHQQbfN23/w+1zUVcz4F1
sFEtfANCdl/XivuylLAwEsg5TroqKNpxnMh6gWjiJO8UAXhh1MsNkVrdvQdH95rB
uuHWqZ74A0RNHCDmSuz0nyHjNXpy552mxArI1tUS3TYVvOg2Vi+ddWTqOUfXzki/
u9SWQIaYUhS88N9ZbhzeRdyDo+Ry5ZlgGQ06zmkRavDoEAdF+uqZdIWpi8E82KVi
WYQPeap3ahUICV25mDyYWpmDM0mYK5AjVtt1rNC4+8S0nyFaiu18dSxmAL+Cug1i
9WYjGSu7wszxyOSKA4UreFd+weGmdl0soDKycxrevnZ9nf/wUEVg14y9pNvHrA6n
C9xryOxeNOK/YsQPqgCFSuKR2/a0hi0YUTq+k/4lLoGR7EoDhvTXG1be321Kea1W
vNgGU7ZVvLnIYQA1fazG5PC9bkBCT5oK5L6OMEJC/EPWONRIzg2Ll0MVVCFeSfeB
wCiB03Ch6du3Dx37tyX5Gb1/eDEE4YhibHrf15oiOLNX5jB8qX3uz2oHk+sOodW4
myLvR2IJGiYy6Jui0XQJRj/MKXyWsetLqDMrMLFZ1016N12NzGeuH90WYQ+zAIgH
n61u9rfVzvLTpKLvA57NHhiMUGrUyk3vG2Bwxyv12mKdgtG43w1Kp36WUhNHfh8S
6uV2543rhG4PQgNZGkIMWbNvJJh8eM60ZmYYzxlOfOcfq1fJC+rUKg12fn22GzTO
X9Ru7ObtSyen9OE27P1RnDZZVF26scHd7AbLvrGw1Urh6LoHni/Dz/9NLQIoyJEU
I1D4BFAsfv5VNFWRdMTUWxN5LyedNyt2GRa0TTo2z9W5L3eP5H8mQ/wT6eKLQTXf
6Eehjqma7ImfSgUnFYNm+ZE85vJOTqz+dzxOf1CNjIUcG/6+29riSLcRx6Msdvmr
7qd0LuIcqdUoSvnJEcOFNaEX4QtBakbOLpmVmzVCelta/9g3Iuk0VH3qhdx2kcdV
Y6R15GN0LY1WPpNQ62KAXyq6KJCRkviIEQQ+N57UhvIXA/bG6H52uIsPbaUxVFlh
rYFIi/m2T2Whk54Qja6fTS24428lNbH8VKIx8iHtSgispb150TCUanvT2oOF/CgL
vsj6u8rb90J8aU2fUcLnT1Y+5n/wTMfPlVyE7qcuFANze0mjoar+xojVxejZ+737
uk2yWdLn35JNMEdyGtaYkabX8PApUBKzw/k05xkurQQCmFamjhW6b7CVbv3ff3ib
wfjMA+6flRvk9t4KGZklu/C7RKzBmrOrWlJ6qslI6HRYX8mfDgW7if9k/NQ4IEto
3cOOhUzdpiApYVWVke54qJtiM6StTy/Ek9WAEG0WZtKS79OqD5sDwpHcfjvtKgdp
7Yznk+46nmIIiQeJaGgnyu6cZtCy2/xSPGtBgeXbGVXHj9fUO55zKW7WmyYmlyPD
a/a7EFwTr9S3lUwRKdGunj2BaH0s8kTSBpNUqb/Lj+Dczpwnd+jKgCP6G5l9TGd2
lhCbLar9Pl95J4qs/Y393JryADxS65cc7NsgA9Ut50hpadHD1GVNxf4Bg7SqROOf
+Cy5oJTi6rWt68ZOjASO2Uk+IYNcg4hm68sQbQgVrZWOvooTk6IDtS9rG0d8vQ8h
/pMWvn8nsniWwVWqApJ8YfU3TsCMAK3V0N5tDvYx82mTBaRNxMI1GUBUSm59ei0W
4P8DWImoQ6rEC/W66fp8Duv/Nq0BEiUzB+rQ8+KZBLEmLE1OHwXQHz+jEYI0yIFC
zb30txQIWnFN+A5LXOwIj2UoqkMDN/J5wXuaTHcNtO2I3iTdNZ/948rFDtg4+g0V
O1C2Y9Rt07FjtlFRQ79R7UZZhTkv//NEFRo/YsAqnOy2zSkIeB2lpwrUSUvYgZLq
3EtVKQfpmAArjZnH0RtrNmsEHSAFH2U6TEPtjYgY4F9xBTuG6ZEGI+5GrwOuEEqB
EjadJpkFKHtpdKItUfwoBzhVUuuOOwXMMpBNnv1oOeb1sMa5iYSeR5H1oMtt5VWV
kc9pD8Iylpo3y3rBWM7LGc4lfpvZpt0WNnsLSphYbyDEwvaI6sjaXnKKFUE1Xdt8
dG/EjxwHVkEF1dVKoywdOWLzUPupMUDIfHXp9BPvQ1krX7QZLDUzk6ZcYNnya7j7
hG+IoANpdr+PO7klAmnDHE8iIBSGiMOZtFU6P5rufD15nnFRNW3BRV25PjezUSKj
II7gQvbDJRRtF1loP3im0EDEqrkpsReMhT+ov7nMR+yZ9LNlCmmxbRnWCqNU6GUg
IKuPugUqDnP1hZXlTU9BWlhKGkgILQlkmPk3z0a6HDDKJRiF0nXzKDRo/tsrYdH8
2y9XZHZEOhDFZUQQqit0cDGaX0zvzYNA8wIbj41x17NYjGXhpTmAZ4hkvjlxMCeP
egbm3Pf6rhtkSjpMZMuPp/3AiWyzf9e5NDyajz2ULJjP6hh4LCrzKZvpSe6ahReZ
8WNbshsdf6USmQY4Ac878AEeJCrPWxZ1BmMJZHNfi2nOwiyW3xiLA8YntDB/jwAj
yaLQRHjUTXJsXxCQH+xNk1QogmlcA6qfDpG2rflvzqXkmGqX8/eeVn54c0Il5I5D
/bIMDNUpuNYgXlPS/RF3NIIitfGUWDJxRhbFJlYnAGKdRySIt5XSROAIhbrnnW4h
w7Eb2E1Xmt/O/dDFtB5uE5A/eojE9OvUnXfrKGiEUYRfdWht5cqBVLHTJGyXjcPA
iy7Wh4c5T6TTWoz2Saj/GYdR4ua10MOGs3mm7qoZVg/iFzXLcDYPcxcZ221khVEl
LV5AOu2J8tdo3WhPFv4UwJSyZo6J0vY7HB4yJjkuPiPaUmoHVDK89yypKOZxqrAJ
u9qoxNURZIp1xNLmQwUx+WDDVBLfaSz9y6dMODgJ8zZfli+ziy9eTCW5V4MuYQ2C
3UxbIlp2JMuMWoz9y5BzwDjxuPXQXwX2e7bgKc8b7b3M8D1+oP9la24Y6qc/Nlfg
zX7svqpul2FzWW7WgNsU0w7kcnG9JJLJ8UYdoBC86bUWEjPsyv8H7cLdkWw1p0EZ
J+K4IWyUIvxLN8AgBEBRBxKAFfBbcN9HcOaRCegEt4eNZP1NinxljX3JodCL9qsv
KpRYvu7T+7mx4H99rnwoe2oIbhN5+jMLN9xSOsc+BVU9vAmLIop1xQ8DShZoHXRf
maWLYIg+e67pK5DubWqv/kG7tP9mUuhizTNYRnfURPBL9GrFMBNJcV/GB00+Ke3N
zr2hQ5+txNXhH1xPKygz6IJEeEOIo4hJZPCJKUS905rSTZMrYksYpYU0VnOeqofz
Dk+QmRWNOO6Ea7lR07OHmLP1a8HCcATy4e7PJa5tlZf243u8Uf3JPis5S4Nn8RX4
hQ86zh+k4DQndowBCibAwq8u08glv7LxtR1Dk8CCKLUyc9tp9yHXewmo1lz/6VzL
YwDEIiURPuIO8yQggFH5kz4CPkcmTkC+CI/3/Kzz6i5TWsNvmCju8q9Ye2U7RjKY
tpvh/ZN45qCubRJQ48yOiSQyBIX0EIeUpR5GZBicseD4IlcjA/q4ixS2gbAiyck4
RptbEA+Pgutq3tYbRMhH7xhI3WoUMFpHvWe5NKO7UZMX9AjYXmgAhbSI5OfAptxT
jzeCA/EHKUDLDSjEJituFyHoYO0nZ27U7sbUBM7tEwgszR5N9VqncguRNKb+kUat
DvcCxSfQKBwfJHNtx7g0rbRsxfVNeN1JLbP0DDE8tqYS6hynKLFNitRhVRX1ajJH
ZVGZ6t7Kl8Z4YKk1SU3RLYBpp6wG7p/UeUVZZlyPMH1XT3l/ADOXXk6T21qbrLNB
aHoXkmhHINLd3wBmLYD0Sa556NImC+PWxX/LrXPWwj9AiJYPX2UuXJSVWnwgsfee
DGBRuX5fwyw60Sfxg4tUTKpxadC7wdED8mXklw1lEEwLYoAPflvXeXG7+y1YFnTj
CxhwmX/Pz61ZLuE2QdP6W0YSbSgkL4wfNccNRjPsgKB67bLh73we2sw39628YIHW
NyZHTKyD5GK+QLQiGGY2tCdn0lDWK1bwNAbN/PdsEhtcIl3mAZH/k1sAhzAxlZwJ
rpeHqORknzL4O5saQhCjhpM7FJFQTzYJEOKFLzhP1gFcMIkRWH+FDUzyZ2Yz2v/9
kr1I/sF0IX+98oZhqBL4skheKHgjFlyYCdskl63HNwl7LjRXYWliM50m1r0bhktU
tC1ii1/llk5gVtq8U13B4sdTZiJSh1gVYe5csFgvmlFLbaRNxPu84H3ALMtl0qid
/ZteT5QBCCcMtOLg/+EyiEEF3nGnxgsJlaE+ITbR+QvPlM2Gq9PnPaIe9A2LI/TG
Aq82lU54iDJhXwHh0UiI1uTsbxOjJiA1WxVoeyzg+mbS0++cyz2C9JeMuezjg6Bu
gaW92xXWnAGGdcu/Aeugbxuq3zI8yX76CEVRGOZR6FylRjWbF+E7WQyTpkgo15EF
ktP89iaMjLK0ZbPou1Lycvu0uWwzZmSTGBlhmGcuUXmuRtmXG1B8gG6PTCzEZF5c
7uUqdLBkD2VQ+5Ivtv48XmpSfHoIvTgGIPJ0txK7aO833xmaeZSE6bOHol0yd3Vm
xt8YKu1v2r2igVmt7yQK/qRORKrac58lnencSloZoHLBA+hb8qIAOxXooq0MUB1Y
+ftLw9CV+Z8yOlOcJXXQA3aA4gPO3tNHv3OGa6km7zM7P74N5bVdpK0koRGcefc2
4O/ssllBJf/88fb3hY3vRpTTDuPKtWdWwOae4HC1L+dV6TWEAKgyjobsdOGHics0
zKjuMUZrlLCmd0Fjj+TA8AAhZ5ejhRJbbaioRmhAp2VhH7aR5k3khBzScwUo23pJ
+J2dMqbsDTgzBcVLxlyPgcuF7UmH5Qi27yXuu66vgEMq7XmQ1rcAVSTi/yio/Gdc
1XmKFuF5EwrrcBykKBGCUaz+6wxE7ZtVXkUEF7opyqpTcd4lXWlKDJAF40chVise
t+J+BIhJpbLisfEMHNq7qqXgOQ1D49e1KrgbPRohsdLfs93adSe7GaCck2wCnNfS
8MkvOHLX9Lu5xJW3rHZjOY9cAyldUiD74vFtR3/CtyYuKCdPGSjWLPwdOwF7T5CR
oMUsRnvbz1uw5IwGTFWHjzN+RkTVSG0imptwxah398GcI5jXdzz8eYebgpsz3vjf
QEsCxB4/U4xMWBvpWotBubx7lw2GRj9A4fmXogk8bYjBoUDY1PpTDoBW0XMEoch1
eKz6aihzSMUahrKHc30AK0cDTWWBs6k/MckFiw0uzvK2q5zOMBrIL5oLUF+DgaWU
qhQkf+ZHgQEdal+QhCnh7VNqG8ssXnVTVKbBI9jk2bEJa7F08wnJtOH+PFcFIIsJ
1zC60+lu4mBq7S5UGMK8VS4sqrOyCV8G8Q+Z/UuZowTaA5R7bvuU4S0Ip2ADOWV/
ad3ihTGP/pZBJR43Cyp1Va0KOsvfrC/RJdBHD8YV82p4Ea6QtNB/58xQD6/jATuE
1PeMEwfIj3IvAUGbsDUNBgAsaufcqEfEX1K2p+t1RXyoG1+cSf0jgdWNKSKSsat5
tQgB/TZxxDtWulGe9D8zl/ifBZACXy3FLjsx4ZJJtZlEKp9Nl+0MSSFCMn1SXsaQ
0BAKPqUU9I50qtZ4j6q9cuee23cgJsoRiDjXBCvlyqFVi0XJuujNOWfoYOqIcfxq
TaH9nYgfGcqd0SwD79G3nIRFtLsz7RPjPvPpf55UTQ78QGbnvSylww/Tadi0ILf0
iRLLk69a5YlF/TzkBTWdFAmYWw7FZl861k1zY0e0xdBdQggfD5mDzb9UTj1hMdY3
C5ihwl06ivbLze2s9ODH6tp72nsx4OUwJFBuTs0+YzWJ5wH6WkxJpUrv86BdbIFl
MQ+FwuN9CTLZvdN13hhUEJGU7YQQg0DknSjK9kK//Ilv/e+znRBo0CKOHU3mv57e
tsm/h2GyDDfJAdr5Iq5DygIEpW3YeG86ssncnJBRQxbvlNBiT2dt6/MG8MF1pvC5
INq+cgWHtIVnPfXnDOXEo2DOVzwhZuRdmkWpDudCPNlgh675ywIH1YQxCGotYXuB
OwL7VNBLZjkNKHRqiuAb0qrTK2hO5erpHNKqLyVlkUHXmjKV2NFWwjLQ2K6rnuE1
4HhxJsHcGpDhNENT0NjnTpnCjwI0ZhI0je/+SUDTe2xI9I+L5M4A8/AvKSXrRovs
NyIHYM3fGVXXZkZSJFQLnZob9/pZ2BWioGmH+YEAValM3FXvroJET60DnwTFJ0eH
uDVNXS/c2Hc0fDrIZRrUZKQBhKlH0AelTnxpiJTAvsIpmtCdVwW9f4nC41t0juxf
EVTF5iNONWZdLZ2OIfXx3RI8QZ8cj6PkbVxow+v7igqSl7LdZMXwULYUpaX4emeE
evosoLhcNBqi45Vu8GxP8fCBlaoul97cZpUw8VdkiZgIkJ8gicVjFFnlflvn5jFC
cEMcvqGZqvCtx6+Uaeib147ZDU/cA2YfqdedOblCskE52FIyTRQy0rjd7/fg+QQc
t2obdADdBPgK/iFhqDh+tWSMLlSkL29Q9M9fVB58STWujugXK7fsdHyvgs8r8vTb
LKf7KuNnMuVtIRxy9EaHurUjP4ofR38d0qtOngc9Ka5vfg8y82RswRERW9NY8mBS
h5oi8BUpC0mOGpgxH7XgaQoP9cReIf/6iSurHqAaRSK6Uh2svLy9TD3JOCQg+MnP
N41B06jRUY5rGZCHBOaC/ItbGpBYH5J/5F/pIt4pOxny7kW4hcLn1pM3alOyWhsv
B2PiNx4PDBRpdqjMG0ED6ICvxt6VCO8aPASjZYkE/DWbQ/N+7OSJKu81gZRJlbWc
5uKHwwhq1EP30WlopW+eQ0ceGwgLHcYUO5Xsig08XUrsUzmihpHYS8xfwpMXGxME
oYKNdPMFi9NdPTkNtKWZ/UxDmiRUG1gHNaik2LdbrGZePR5bkNHHMEVeQvaIkq8K
cJMJLBLTPxRVMp2+Ym8h16h9P9zQI3b0lITAIWpZYAGJ+6hj2G8cpHdW7YH/J4wG
Ja1Q4nIn/mk0rkuDmLyU+HA/glu8JmGYNNCAQYY0QTIru5AQsBsLBmLuI3IhC3QZ
MycslfaVlcLod2R2Uvtm/8mAeCO67Gqq4HmeqKP9/AyjcRupDDJXKOw6VvnjyFwV
zKQtNJF+vfRBLGvFEAk8y17O/AIB9pG8aTf/Ylz0P3BOHnCXIEaP9Q+Svahn4fYX
/59urnjWAdXvm4bgqRXN6fU30OJC4YxZveqgIpq7/U0ba/onn32IRiS1lXTT92qa
NOR47BjhVZOTwPi5Tx7kdFbJwKZqTU9pM7TDmgGr8fMCbD7oNrgESrz6BlyJ492U
pxkfCc54RqPH0HdcovgRGzDi+johlujiiZrFGpFYL69fzP6L36rIhQs+G1jG1DLZ
4zNrAktEm31AlaUUNIED1Oy+RY/g7nsK8QAkh25EWyZL1ybx/xs3gcvfGgcRhnOZ
hZwfJsz7H4DNKpX2d2NklmNxN7H//9CRwi+gfjaquC1YkNHBSoM8leHiPmnS3/17
fW9+GPC3dzs5niMoQ9lxH8OcjmTWIYvyVEjvwoUNu9ZzR8QAF3+iyGgSZKJ04CK+
Hp2JFaw48Gxhz4vOIW821tjNuPBiOVpeHE2o9BkOs6NG3OQFadmLeT8sH0tgubPX
LPVcQYxnAsdjCX1E431pmafdrXBZqs+0AUrbesQ12gx4UizZFPjFDwB1SXD5zSow
A2t2FQAFlwK10Ss2Osm8vIf/0dXVdjvcgNV/pX3cx6Agcqp1zIQUXqdyiqOIeMFe
AaHEVXBuHaMxr30/CwICvG6PJ9UHpg2GOeknW43rOpiRa3UpphYdF6df6vIvqlQM
BIdSsVQOVBINN4KRX8Ha58sRCoL65DYVKr8NWUOV5y7AI2iDRfk39Hr/uYbbri8r
vVYRBg5yfj4mNoEvnht2d4NVtZv5FGIfEyKmQqeXm3QHk7wgO6pa7CS6cc8nEP09
HsZvgZJdHlDJQP5b6aNV4YybHRR52IHX5H3+T3wnXGmQG5j7QtKPlzUw8Pit4eMT
YFUxhJSiflj5ITQVe8bzr/Kbe6KImsxdcAz0ap0F7MClOWLGP8TNNk92fars0cZ9
zW7QTikX0ZPNwNSB3jzxZbZD+Z97rsRjcuEqeEFbE/HmAqRLLmfhx8iA6VmQaOAW
rRGJOO/1fO7wszjiAXnK9Z4nrFNOIwpdXqRnGbtcfJvv1ksvI8h6xyzYmRxNs3zd
R8l81rrBJi0+N4Q2qJacNfHrWxbEZcy+GOFwKBHFeSra2ZU0nBszcaAXWpWIGbXe
tztLM9ICyxRvCOIM/R3s902LuqgJxTG5Mbj7bPBKtum+sImcgWNb16eNLVRSB4cn
3YHighjPiGYCtQjEQrhKGgrWqH/AE1TZUzbWnHaKPOinCCtcCB+y8/y3ooHz9jzN
bg+oKWNqlYw00xmW7wLBS4j+xVroq2rebrYhJgckqO2XoQlkpshTL973DPZTBaIF
kyILmQV+NXLwkKVS48ZYfJqEwRXXh+NcVPbXvr+jJ00zIeFtCp4NyMDFdKy1XbZV
D3IyrpgJLnpyQeqaDGriNr9sWavKoJbMx/Kvpj+ROU1e12/1n9oA7/y/OP9qJoa+
/dSQ5AVWcqSbvxYQk3ad+2FzkI4FzBZAxOHlQmPfwOVy37pHc3lofO9AhbGS9mTH
pHvFi0GAWtW7drdA95bkb0UYjvQSC4M5so9D2EgIph1WSif6q9a9xRDSHqGR+gJ7
rDN/Cn3Ij8xEloQEGSnXYsnC7Gia3F14McHNPpo8KvZpTJyP3kBdvo/sU8YmQ3o+
I4vkIhd1GH3mP1UMZqVCbdPDHA0SMZ04p/cSt5d5jsro8ZAPVy2bdmP29hSB7WrH
g8LHrVASgS5DJljNmf6crKyjhqTGIAgu7iqK2/NoxS1C947H0EmwKnFgv//6OngA
opN6+bpzekyP7pcd4ojSxAmZSxMcuPD5Uy5j31aHqnQia/YSggvaQ3fwXVO0xWVZ
L7yThm1GzQvgubTf7ztP/G3JNqW4Xop71DS9dCL/qvqrPeSjreC5HxAz2yZ2Fqtu
BjCvh4VHn9sHKMYmF2UXGFQlFF8l4u0vvt5OJWYsFW+KTFzmm22inGAAsSSwEYwy
CHXIgY6qVKJRt39gDlvoha/TWlx1yx5gHzh+3jruXHoAM4ZVcqyB1kVwzTSKBv2R
4ZwxPU6jJgIIXqsR0R1pJj4DmCua05h2H/At+uhzZuk/B3fehOK3aFiN/vxUHo21
TKFqrC93C4Qa6vr0QFuMNI4QVMzSu2GMVUyFdSCTGgTHb13U1XO1D2nw8F3537/x
IklJmsKlDfNvPiUN4azwzh0w1+SaByW21ftok2bRy3eErXx+LkEi3eavFR4mMCc9
M8zG4fCvHYT5w35cG6xz9QFGCsvG5YacWcQjPSgB0KFklYf6WAJJmw4gK4GlrxbF
mE7UeJ83ufkVpmQLO7Q3Bxcs1SWWs8WhKIb20I6r5cpYCn+Ke0FVt437IEiwwusp
YptVdWSAcSmaeyiT0lyHsyQu/CR6toLLy2CzhPu17/W17WG383kMgx7ZyPTBIjYC
/lqPKRdyFifO92i0rRePkmG2xZXeskA8Osjd8SYaDVdONDgDDcSx7XiiYPYyRCVz
lnNE+e/41AW9V7X7QxfVsssTYiddzGRqFw0Qc5fHgnS37URMDucvTEqydMsmMLnc
y3xKlz/UGukUkr0F7SeVulrUUn5+OhQQjdExdk/gcNosCf2oYCM/McOwnWQqC3Aj
ivRM3AqGZG2/kafvYgrEnLm8i2CYw0KILB7c7OzCwSPjpk8o7oIbpUSa34/ChIc1
YDDwYeoRgs1tnYUjQ54DaImSZh9qV4jGGPWkm9ntCYMLBLM0m7dWmcGx5I1hJUrv
Nioc2ZagW48wt9HDLLe2rmZJZhG+6lk4OcFK8JyVr80P68g96cuvTFyvDZ59piFM
LukWTX0nuDB/fPargJgIeqQGK2XKJ6RwFwJRFp6bqFSalmG4x6Tlb6aq6wKMVdg/
PilXDdUlV22zivku6sS93CtbEskMhEqhJ3NSR64aVQ+4vIsmgkd1FAXtC8F1PvYD
IvsPZWyZvkghPvikX9i0MoihdsGrHhH/RQ2A8T7xPVI/22Eo8ArjsJ1HFBrrgvuo
USO5ydVreUkDGUtyltn/HpPbIy1X3y9tFkf5seb8OqwmOezEBwIeKYHzSpqAMy9h
F7w+91hnSqRRB7/8+D5yN+SR5vi7djGdXd4oEGglfxwlUiRupEYS6A1bRxbNKm7I
Z3fy4s1fGvM4tB8Tj/BbHsxqTOv+RSk2Z12UfULqtkJDS48KZWz1u+FCTSMMd/DU
KPADnlj/vgl0D6d4mwdmj6dl9Ukq2HMqJiUZwbaS6sTl+I6ix6eIIY0h8lECMWtF
1rDgHbBDUSbSi1zRqgDnKs8pTP+dMhogx7cqnAHAodn/XvYNr/nkILURTK9ac5jJ
n2noktVKRCFEeMELeGDdIQD1b1XS9g2cMKn2m0ubHWPW2GulrNcGrMqqzcoOLhMv
lcsFqRkZ2ExwWljN3uWHvxxNpm9ADFCmxQXui1IzA3bem7R84138OOAZ/yCXNflc
6KR5TZJsBLQFPB81nKSYjiztXMj0rREXGSsaCkGNqwn6YxAeyUd13CC6f7msjgwi
o7A1cHYrkXsshDH7jDdtk72dyqiVaSc188yau09nBMW40fBikb3QIcuwLeGMRPLi
pL8KYoLyyjc65RiLlW/UVeRhzzXQbi4KIt3cfQxfQcDoOP0Y5o6G3nhMBOSS9I9f
Y78JmqMMFBfDol20y0SdZ/MdUAkMzdbtLCKR659d2ri633JR56jFuq0lTaTdlWMq
EytQbJehfVIEJRQvIWi0JJ+10roGsvnwo7mWh5evUotfOyfOnSZh0LBxfNmXouAn
mqAR4DOVeTralIo3Gu3kEh5FMF19uBFe5ns8XQkopVXBFKNt8xPxOm//o+DH4u3v
zYcd4UqYd9oyv5se8l7WZkzNVrwaZUlK+9P13fHTiKkriReIO4ogQXJeWXHoa+5y
XT4KtMp936ISLESBBhP+coEgHGrQkvRUocZ90YqLGFSF8+K3YPMM+KMM9n4yIlGK
TH/1AckVJO/hVQiB8guLV7/ynWcTCa1xlVAtjPzel1ktS9sP9215mDM5HaX29IbU
m3Zw98+6eFq2XRWDKcISJobDhkay6QFYM51yewso8aTOtt6K6Gty9NzSUUqShj/Y
cwvxJ1aPoLlwQD3wzRSVIoxjuYQ6mdNtOVG8zNiSxQX6yco6TlY178kivrcagzMM
LXgQDlB+BThB6E/kieYsCC1FBBC0Qum8RCdj33M+JDh7ANjw+twcjGl1kTOa4Z0m
lgP1ORnngbsKFSuuvb1NaRtEmfMTpEA+j0L1LajyrT4h4sSJXOC/kHrb+/AFlCMF
o8yOVoQpjA57JYT5/frMxo1Ax4kvAYLg0F4eBUhuHR2CXIQmySVFDYgCIVrvTOEJ
vpC9XPZdiu8s4ed3PyErpY+FBM5vIn/pM5HMht0IKeI2+7EpE09U/2VJYSoZRv7z
ZxVSEkIC3mlimm4eSZdJLge0+HBDiTTJ327SqFKFeYImmpd1mreY+9Cs9vpyIicq
j8Kui0NGxcL0PtKXavLfFNiwjWYJq/czL4AWUSMuy4pGkKkvh52SNXyHO8DSkFJA
2JlILZY1T9pHlo+SsJAn+VSQW1S7k7XNLXDXJs86xbUZhVggbKtuyXMUjBJOCRpD
hl9z4AUkULCUw+FYilPj2Wf7GLTKlopB8TTOGPyGu1L9a26ACSR0XEIyt3mRJGMC
RZ81QLBksJO2f+7mhojRZS+xhP9XdXoakfU1XHlzSmkuzB7YBKgi5vKWxe2pO/bi
7Pg6WMu4qB1XRiLP5MaxC+ZZ5Qcq95qJtuBYtuyR2MxkLEJV+r1XbNSLDeOmO76r
ilsFnkOjLEzUpGPqkO7VKKih6Rfw9i+L+hj78ELKUZ43uJRfXpDqv4xdQ+yONsNe
EzSyFiF1PVx9m2m6mUVORLFGne7wnqP6Z5YVtyRWKuPeGs+xtjPER5PJ5DYBcXEt
Ce6eRWHm29LDn8KoxLWjNu6oOiDUZAH05M2GZKGe+gowiF3cjaAk3RNmsMqz8m+Z
5G85nObx+Xw+n48DtzhKOrsbzNIkbOd92lB5SPXYYxKBurvk/2E6g8MZojYRP0pB
hdRDjyN15QJ/ujihlsUB9LOJ7Lb7FH2Z6FJYSimgxREiHj65CHJiLv11czwqm+qp
9yjKeQKIhf/Qzy0JpsIeqaw5GXxuROfQGJ5wHwwg2os1BmxEzXXT9Y8/j/hZmGWa
fbjs0oarPMdQ+OLb7ZZxDZTkSHvJHJC3O3YNNWrAsY3Z1QrqB+T5MU57/HQloq9R
6QNiDn8fqNUAjm/5loZSPVcIJZJtRmHxNOv/aBLGxY1qYexVwNXf6nf9X/E4gVJZ
ouhMBOu6M4ahJyvT9718eEm4EjQZClH3j5OexHYk86JJ6JWPZFEvzOzHTVhM0Vku
H7/Npz73vU2lQ9eUjcOJ5lS++5nYy/4tkJzEFAlyuC7pXPcOAnie0VAaKg5cxlv2
5+IC9eb63RYrQLKJ07f3xSfT2CCcv2myCs8HwZhQttPuolFqWCX8L2iF3fPS/N8m
JCFxogOSX046+KaLbn3Vikja9wZe8Q+oBXXG3wLlGJhBa/+sZtGJ9cQHFheudsYe
lcCEOsv7JI02gaZ3U+b9ciT9GId6A/Au4PAaD9sxGPqu1j9Qq+rSwQx3GGvXvkWy
G8hDWXkJIqv7siaI8olat2a0HfxPkF1HloF0jlQV1YPHU9/HibUX8lgFlVURHIQY
bCaGfJiLzv8s0xjmuPUVQHqaQExlQkjZdBY1qH9gnYrDNBG156gjG9X88QQYCB6c
KjrgRE1wW5k01uwBK8fcfLElYAZinRNN9Q4n5mmXN91DGt7cjH7fHRwAHv6ufsAh
hd2sZu/2Kg6A7ZhjQYAPFQvGHgtU/K7HJXKAiW5IeBRJOzemJjiNXAhUqLOTlzLW
7wUhzY3VYUVH9Rt93CGfNaF6dFmuL71MqsHVUbzoFXMgLzsHpkyL4tZGSX0lK/34
ixsMpIzwAGRvtdmjzBrM5QaDWuhkBDfyD8FXtXSeC1zy+lVhqMurxsEY4Kwk08eS
7wgEj5hiBzcPs81Oit6LhSwpN5BovdI8/rhgtLThOvGREN4TqGGFS7HEuAPC6qYV
zGZDYox5bNOqhc4cbnZkhUTJq+B4Y7FhdRPaeBN4H4Wgn3ObE1FtBKOWZhBhKlwx
+xAitPYxKMvTLo+eES9NKu4IG8KN53k/F0uRza/Vz6Lx8eDCaqqLoruU/4kKCfEZ
lVY90JsaOnJLCcTbGuECxg+gH5yLXrF7R8SHxDp+aK15miedgNbhFvaEa1tAkIx4
9fNxGRDiVh1E6FeGgnlxit5FZtotqiHEOO61bd+qZLEguML2NoYoYjW7cbmNp4Xr
J0XQ2AHVgS6S9x/bGI0HPWbqsMYL6HO/sfm17+Jx0xuwHf7pwblYNH0yC1LVAfu1
SJ3VCALq34qIuZl8ZrIok/pdQfX+WGZAqWykCiJhkt8tk5EBI93gpYYqP/GSCy+C
C4498KK20+x61oUSwXh6nfAzoxPUIfrOcgmSVktCA1PGjANzgHlXHy8bKnubUlwr
g2iMw8w0Ej9VdRUwIIAj1G69x8UTWB+ntqxypX36Kvvko/+2XjW9jCOyB5ZiJhvq
ticRXdd6cYBVq83R5eU3Xf1KhwvdUIp2Hb/gTdvHeIHpexlrZE1W4r9WrIEVRkrC
ljY+G3voffsBhfaOF60Ot0v47+KeyKFSCAC+K4QsjZnRpI4lD3A3hMLpnPOvwzU+
CIaVb1d/nSUCK5W7zc37ZvY8iBmVakUYfYYbGBOp0qWH49vxAc+9YU+HvYyvPgja
10qNRNySOGwWeGL1avfpWNKYZayT5vgGI1h8RSh5kELKeRNnCtMmfGl5hKQteTcr
mnpmxoQPcuQ0yCvI3+NYh1FBO1Oz8is7BuDw4ZwKRkEfMRtNqXVbWfXHnU96Kmxz
ExbiVKtpAKNnJeVYG/MPV+lsFX65NmAHF1nLIHv6uDRftncakgFjAZmlTe757Swp
1LQLgrGeSCMhh5w/fmHAEGwlsFqQl9eONmS1L21oeBkpXwA5H8QXAXi8g8rUOqnF
M94agj6W6+di5vGxjOSb7PmPELYyvqEnAYOJUDTkALaSJ3IXdm+Jq3UVeiglzAth
pTHDNHwzkkEWRI6XgAIvwawsJuctUlm/9hOcB8lPoR780h9HgJgd4EvlQa2s6SsC
0MxI9UxDK/Qf0MboJGvOkqV5P2Blq/+CWahKlwHX3GtVNgIt2DDKy1vwkwJdUBXW
Ty9kufk+K+7FtCSbyXwkjuNU0wQ4LXqpTKlhN+St8BStlP/9YiyM9dnUACcHWXsZ
fxNvkYjbpy8Dz3EOT8h5dB5Gwq5/hCg8xIdkKKR2YO2EiUaXuZmQsT6oSKej1Sv5
vbWyRToIk9ftYVr57veFrhoN9VvAUVt0OGlgeIR5sx2kp3F35CNqXM0NPIFdq3zE
Kh+mVLX2b1MNkT0O/DcbOrZ3Ia177j6QnF+IwPPpFqLFApjwUFfzBm60C1H/jROG
WzkVRKnerPAO+GCXSvYlZIKNNeDVm0RYwgrn9GHtTilne3J9GuKhYO2luhmDcD29
DoxvZziCaU8pP/80j9CoQ9iavWdo7j9uv3FukvTvlPQ0ktr0/j/OTnSOxvEYox8B
HgkTmqHhSda2SyFZlrr61+gHg1SkGgD5Ph8b5wg47qCyMt0E++gkAaMa1fNPt7Ci
0y0Zo5C4jBu1NV5Mmxa8mHB8PMRJY0kLAp6QfLOMfLZih8F2pWsy6eNnsztfEPg7
u1ySVl9Bkw1ZsN6XEdwQok09gg6C4j03RUGHoLV5h7JGA+QcCg2h/0YHzTRwTo/Y
cxOOrAl4NH+KimteMeIqgPKMOKYrQ9E1h2XYFrH+odIfRx09qBf1RhDeDqDvlq/L
TLOVl88mFYgsGxXZfhxYRpY7ZvBxu3vTZ/+dmVi2B0upC/QOG6H/gp0UZEtES+Xu
J1dFof6jTdKMaJLOGR8Uq497xOVVwRs3o8ezbdIY1YoqePkryn3P8UEQ2tjJQL7Q
xfw2fNxsggtL+/mmlaicuEm5kK7lJ2i3HE/s6/uFOpdAkn7sBNv7qtOpPxLIh9BA
XMfeBGDEwvrSQL343MPMittI0FYA3t3Rha6snxHofQWLtCW+VzwuM3t7GPo8TyLr
Bco59Qc+/Vt54ad8TdawTVMu2QH906cTKtVLrgV7Lhho/IIFYCYfdYxbEewkaXYM
dALju+F4X6wdP1R2JAJB2qqeZyZb9oT/DfQYDMR2/paFKltr8lXbiDeDyXjkukkY
u9hS7fc0ZdVv5pDdzGg7WS+eYW4IgLRB6pExdRyj0Qbdr2nuPtefZ4wVnz0eh7/G
b/NY2Nt0ONzqc3AFntsv/qfGLYm93y54AnWCQsnCTYhHryOvpb08mvoobShdQzYX
WZxcMZ0xy+AYaaXInFuCY68//+ZYPNHw6Gk1SqlsqdvPKxPsHto1xPK0ZfGplsrj
nwqsfCTqM3RUi5m+xapQV39O3aOffW7gAcpYVhOOyOwc6H8FBtYRsKactSaZ/Vey
11Ng97fE0pzS+1HQazr90U+DWJUQMt/DWIfY4dwno1Ofo+O6ChJh0/ylwNFFPnFy
CQUJb4LNsIOI4SiMEBu/zFPCw0iC4i3cWLy2ZXc6x1OdYVqvzuS+Bf8OHDOfVa4G
fP93+5PGm5s8vPuxy9YlAb8Al4vHwCzbyKjNqrA6OXCECa7ctKH0lGexr1PsWTjx
OLw2CyOGCaTvE/9LHSJXgKjg26n1UPxWCcunFCjNuxf6vbcDNX7ppBo5w5AjE7JL
rCg/3tSh1rvE1OmI9z+3dkNS9+UgVFunhj1wCDn6M7VqSH8guuZwTJ93Kti1wqyf
xaJueH/qCcpxvOsIFEw3gRrN/zt03geNfbSv9i5Q+br6qHzsKFanEN2xeOAkEN5T
JDjldjcbUgb1PLACvI2LWey4bnYfvVNIhE797bq+GsmHlQ/LU7R5OZTROdOyzkak
1Ku+9azDAkNC8DNX8qApss3zSOKr7/y0EUQZwKO+99VCs0ImR0qc6kPpPnRHpBG9
004gfmKiT/DTyFaU04VEFGvysfs37mKVI0k3Q73harInciAi3wa7eiCh1yRSa7F0
wECDmISBykjrhVuVRTLS6bhr3onLRmfxhf6jGgg29H05iVNo0//vxLrLLC/WVTjh
ksQ0sD5+q6TrgAtUdfpTjnyS/vWN95rpIyDRWzN3Vbxpn89A9K1KDWCxWchyk8ME
zLkP8qeor5JY2y9E1C1mhyDxFHzaN2mjKtoZOWEBizQH1X2h5CHS1EGCTfKw/0V5
VK3d7yHEAf9Ah2awLihYaap6hc5R3SIRCFhsmK1qQPix4cwrF6aM3dYlUWL0isH/
vAfyu+Ze3tIfGByQ/4VFG5r2xpXcgA6NCYWEbnzJeOMrViiWxcWVrTYgyJaXpQs/
tb/ndHEk3bbhFZe1BLYcm7glwEyDeJ7QnX4MHRoEZgE8H5iFMXgbZf4x+Q2ibJk7
CoMHXeU6Sj8daWAwhHdV156hLIVun5H82G1JQXnRqqog8zTfto3One5ZzQvjM+HW
Wc4SLD8UrSSPruuSwoI9+iK32SpTD5lVruA+ndcglsZFNt0y2DUUI7g3ufwwlbnU
nvKuFlh+M8l4Y3wcSqKBArAE/XRFm3a33vucM9N9A5TWKQi7U5MpL7FPm9CY1VSM
T9sU8Qn7Q11vWD9c9Z6Cbyi6enImEGw41aLli/VlJ9xydq569V8q/MTvGwdxaIsd
+IESkEQdT1oyW+w0socTMyHfnHf2URzJQ73qRJQ3qB9eElgl0gUim9hpXuFY/q2H
O1LkaPTPq/f0GlHVi5o7fjrtjGgMMN9ePgDuBrM/ROvfgViBSHNssIcsz5aV9IvL
s6BSq4XRxym1QA4cHZsTGgYEkoKtXZhUyZ9hc+++87KOEXaLLNd4Wbaznltzvpyc
32j4JBT7esFKJxLriNfXbnyok9594Or5uuNoa897CkxT+6/mgSa1z7Deup8veKPx
2Jwbur5KuDuBVyn+W+PclSzrzU38uDGqsOjnvfKM1dqahT8vtuGzNTWkDDRrLZcH
zl9gmuTgcUEcpPDMqeNIsjXU/byH/KkY5zmrlogOqMCwMxaPYVWqj5hbD9nZu33q
Kkn5gbu+p3yTrwrWd1ONTvoN4Hle2QntdVzNsA96We3dJKLT1Y21V4CHeWieFBDh
BJWzAYUOm8nO0KKGIFYH4xravtlymDGIO/DVwFrir4j2ldB5AMnnXqfW8M4ovDSz
23Ma0S8ADpUSzxFHUYc3FTf1OyY0odp5cZGJ8ZREHBaaXVD2xRmYAfCSPrKCAjhC
IRu0bHCcvDdSz4KqwEP4cGRMmhk/nXMoftnLUYpOGOmHNHGX3fDtlBrUBvQMQXpj
RgLSt2E2a8ier4Kj/9oV26BYebV/RZmHkNehBuH8L5qmp/NQouCwQVFU8iiVi9pO
en0xAR3p3hbUAm0qzralDjLogm9ebuKvOEOX5/E4XRdkqWTOOOXxx7wtXzhcjuLy
eCdskvuVhODO2N6Cy2SWcY3cos0bBSpS1qpYsqhOM7NORR6OQ4z0ox6EuofSAoFn
4f/Lq15GmnJVhztHNIvj/LNklS+qusJWLrerOb5tNFLw0+/lQuly6tqy/Gma6vCO
lo6ImecKYLi9KC82IDM9HreEdHD8MVvsci/Cx895rPBz5AyMP4UZNC7nc6FNLKVJ
t6pT4lzl7Sy5bZT29Y21AfPsCzI45F4aoGPpLc4hixmTKft8zwpwA5U5UPp1lssC
e3Eo8OJXhaNRUU5MjDiwgXJX3WjGOINBPakuOIA0ufde+WpWv/fDAjXu9VrnHkEF
xYmOuuz0keaARAjp5ObQX4rnioel/jwnvWNOPKc9QpRYKe+rCcQUb8QTI0uJaWlz
e4w4EHKCUJy1hoKI3zgoamJEH7DndyzlZL9d0UUzxFkBMxprGnSM5Fm+DzPDDqjF
wU71nWKJ6PHoUwrIie7T08BPW4Qt8zyZvAGvCvaGwDE2AQLPHPzzmvrxQL7F9VxB
reayHBempInKriv4sUR2wSNNkaGw8ok0BlTkBWozD3/OPNIgMlfMXgND5mmwagsd
MYDJ806Y+bXZ37qL/PtAktDxIui8LcfZqpqSaJC2+99PSfpqfMOldQFGDISk8M/M
ZuKfJ0n969ugdBcgT1+fOpR3bkomwpVjH/bRgo6jkvt6eFYI8kNvzsz4zoudz5yu
PCzbEVTTHWp16eJseC9IWpPV/ibS/9uhwOpIhx0XXDeGUZxA+mA1/ojKcx887lqB
iJ2LMvrvpEIwDrtyK/xy5JIiaoVa2EpMtQS9VtjUQ6wGxVd6R6NGesJ5DflIp39z
QAIEOC1VOhF/CCXVpw0TpahMMoDOFuz0Hd06sLBu/+miXkh2Wc/ZTQX6GVxyog15
TmH681/8ZMmWVSNVHeE2XaaAXgo5UD6KFFw/DEn2XvXbM6wed334HAbB877lSkVk
JnfbuUUkAT3V6RARu/MyqAi6WHYq4sbPlfRc1levDDmk0agAtOoyPL5LPTMUjpWw
hLEmldDCNP44bMuzKWsutVqAXTOOuf3b13FnHhNb+256dFdLSakgUoWzbXaWFH5b
oMoTnIOmwtcgph9N6fVTn+aPB6FCUp8/l+b24IAZls2T+FPkMSCMqQIUgOIqyR5b
BhzoDUS5VeigVCpghMMCUe2sguLAN9Tay0U9bLc+xWvG5wx/d+HBnKpMHPw8RwBF
zGzOYoij+7C4F5mRr2VU+DN3YDBln52Psf9D6aBtdXTH7I0hkJK3axK5IHnw3Vd9
v66tUVsFqOFGDwN8/5NZkAAZ0DwJZy0OjHrkuX8hfJ3X8RhI9BBD6tc+hWACVgPA
4yzPNBQPSkF7mFrmb3dAaW6uaC/9CGLMWYcQ16Ic4d8fi0wSdzWIbqwzSuc9b9jM
xwkatbPHHmTKYyO1zX4EyhgJqW1wgVsyW7/PaIJ11QiLctVw0wmlMmsppHaS7BR0
QE4IGa5nqw//x5rjtWVKgD4FoxDsFbhgOE1vlYAqjNW0LP3W1dn8IurTjWNpVOpz
QR6xXCsGO+1PJtrjtt33Y1D4WXuFTC9WmiDjEC+WDr3t2ZObl0m0hQYrY1RsZubL
zMzP3U9KzXcj1/Ia9PQ3fK36PQsPJF844spaKaW7eHbHFlNvxsrmvbWCzRP4H2X4
27rIU2JOBOb55CCN5t3t5PCgHJjd+CqLkFjqLcR6dEb51Y8Xarb1cnXtx77m3TQ9
kMhAY3f6a3oDyi2+vj2l+D1p9+xMOHxNNo3HCfMUsSGF8+clszuiDj9Xh7k2rAWG
bm7P0lRUYa6Qg24vMs3iYf7lqklGwLQA3+h2amfcCe9KvbosCwgR/2MGo9ftx40n
ouPsbLiHC5cLQwbv3wK7WA/MgiLfLUxZmQ2gMMGYRdtTMnIpPLJlYMaNf6aMvYl+
e7beiMTX1Asb/LFwuFP3DgQg6x+BcRLI/NSc9y+8dbrfenjnQ6+zxzKgOstiXucD
6XFK+vIeRvdhk2g79y1s9CPpCEAQk6xdq9Accc7oHv9jP24kBJ5ULLdSnvY30Nrx
RwDXE79X4uodHqfeVRxm9V3bYBZEh2CK3aR0l9fZdENHgKPNJxfnLjBYDwcwWEMZ
Fzk/4mXDwAUbjGbmTvUgX6lgcqKwQJhFF6xNEDqHTCu4zxGkEkiMZtLAvXiXAcwS
/AfOAc8eq74fNW/WT9cX9SqNMLYTA7Nj11Q0zAIismYSCXBpwD439WxKpiMYiwgo
GeDn/tze8ni4ytJ9yMrZ/JPF+lSpHoyJDlqBeiS8qrQRPvXJfdY/RK81VxwEwJLp
xu0Ao7FYR64GbO38XyjRAYQ12joXbxjWi1+W34KfLnnM9EOS5rlE+Jny8OKwz/xr
ui9u6dzlmxF73rE7VjJgfG0CnhEPOlEa5ADO1a2dYe192YB/o6HdW55vHMoIhc0J
17SXivxQi6SHqAqvlFbNV2G0xiwySJgb9EavTalLRdKc8oU1S+3EZ86KpN2FijPA
c5/FwmRigcM+QyM6nk4OeRWceloT8CHQ9iZFh/0CQso+/xxpfXzVUlaeWQNbzYRR
K7Hzq218Ne6Y1umZWEE50njD3C22w0FH3bmayhReLvg0qWNO32f1hakWg9BP8SrH
kXBlHVwNcqXwiHo6FNGH+YKQJ+YlHwD743np+aFzhm7u3QGWf9sUTxHbcwfNDa6h
h89+cFyJzKf1u1jYtId60o2010BKwN+v/HemDcYHvTcNeYz0WaGYbKvSKmiTo3CB
V6RQga1JY8rMde0d6lMhD+oWuMvqDOEfVrq/tjNMqtbX/Ifb7ZeHUrLo1vZHrW3b
8/jP0VE6NEJeIjtJQK2FXeHe4dL5ddDu/vhsOIRTtCQvSdwRHaKDb8QHj7J9WHiw
WS9dOrbuQfwvMKwhiG3B6ilinU8CKqg+Jjp3y4YdAzS4yezQX7LT1cBucmUTZYA2
jk9vkbFzIuxfcya+40RVz6lPI76nxe3ctMDhjvgMc5rRQfvIP/MJRP1gjuN2XSqE
h72+TME6U4f4ScXtLH7al8BvNwb5HSYcplfKGt+nAfFi7GgzSg3tL84SUlHXutJh
LhEQDfxz82xjIABigZqpSB21acp69hY3qkn3wEqX/YF9fZUnTpoKiRxUMxhWOuQk
+TGUcuat4C6ClyTo5EK1FwFLcHwDvw6/HzqKv4UahBGZmrAchOySMxUqTqE00PWc
ftjAoYQBKYjzZqy4w2Yz0UwboKnL2bxFXnqIXtLFC941svzNu69GtvZPu5xNz5nW
/7Zmd5La8Ov19axG2DnhrNs/OQFBENxpTGaNs9khTqBMYiEoVjveRSd1nFh1Xk2c
Gc52v+OfRpdRFS+S/tWIt78asmg2evbQqVv+SZ186itLV9C5xANVUpM8MGNjtXkE
vAfXGPwCxHTnSVqjN1HB5/6Bg7/jqpMjvqFM+Jq2FeikyDZeCGZSlXvi/N9g6iiz
ZSyphQBl2Qz83vGI4AfAMgcw5L6YOBGjYCABKJHfIjCJVyz5wMgVwAdOvY/+0m2g
tRh9XJQBrBTKlecqoHujYu9t9T3aLr/lem7WkEb+DyFRWR6Eu+0bTYmsmXkadXZ9
Q7hWGOPD8cXzuEPrtIKkm/YnfgNU3rh5uqzpWCoCtna2FuyMvfKIWmypnOJfy+Ag
/aATW2x6Jesv8hRHeoXIJb0dks8M5NoBgZAGCHFAz2O68Z5raJmtOZyYn+c4HKT+
KIDBWGoHo53zWeQv3cZ1p/I/kNVZ3pRxZIimE33sY6JR49XeF5KRtXI1pMJHuoa/
mOK/aVVAm8trsPSqz/WQMSaj1eO/DZ4jUr0LNfiiWfaH+c9FWz4LCz5/8Dlt0UmG
5Lu4axjimV08lF7yL9n6pAf3AmaEfvUXugujXbocmiAxWfFu2QTITyt0umH1qCQl
a8hBmtTR+VSgRaYIGCwCWxx4k2ZC1iBgR7bcCqyzOAOoiLQTBOmx6GpZUESpWs6Z
x9uqiNBtgEoh5FAP0G0roAl6bos6szQqxJ+zMZvkIPh2r4/P5Wb8V89sKErcmctH
s5lH7WDItAgdW1vliujEwa/TvZbSIvHhEZ2d/N1IHTDHMVMxRBk+2XYn7IFjc3No
yAusM9FUZz/sRDp5If/VDddmo12krA8DTtcUavwo9NGJ/21sUxcszvMfNuwXc4xh
PnR5XGrZG7zzKsKr8ZLvkYwdotOx9605sh2ENbjn5sNiDl1nG8I8n9mt4WCkApm5
/YQfM9KE8A2AqqyclBc+nHg4oreTXmx5e2vyiW9gT90Y1pE8KoZs1OWcYsIXvW+d
Lv9gKZTqCry3lqRXU4kBD+msMO+0aXyZ3JFTy7/BPR8cxer4oyLhdht8b1bsDMyf
nKnmk79huZ+BZ90Jl/foAS7bHEHWdHle1JF55J2R/f0DzvjeQQ6XSfy0Nxt+iwFz
HJ9dYgjCTo9/7WcbSn0PYJK2PfkEELjUyiuV0OmyGMUAAPIYNMElL+C0jRXYVzky
OB93WvBznv4Aw1oZMhHwRfJzBg3p6UwXZ2/8Qz7sNLwNTnt7sf7KgeeJGFkU9kxW
YWDJQAJmxs/EPzxlQW7Xc6yZJShFOtrNRDKodvhar4uktO+uQW+fFXP1FHQfcYcq
BEXc/y+MwpINhwZIEp3Vm6giqe2unf858Upi2CsAxlVunfE0GWAI9a3tN8PFBvL0
dI0N+qu6QXZSeQ9M9Im5/GO2065GaXRCmuZrles+FL7ER/ILdWxO3ja6LHLfqKJ0
46A8Wlyzv4JuZ5b7Fe21LJenNahNEyhhQ8beFe1icHxxmYrLPJHMvFMJevJQCqhB
PRXLzVAmaRiSS6/Aq+neAhVN1U1J4zMENn2+z/DoejPUCL28wLIk5cVQ0e++h57A
w45FclFzjzx6gVJucfrrsiGl3RKC+Q9Fyd85qVn8EJjSm5PBgRdx9jZpC04+UKAN
QtW9kj8/vOLF7qu+fjhjEkoxf5B4fXrNu9tGLdPGX7eC9fENysccl5/2RLo7OI8G
fd7Y+TmueA9+xnWmjxvrxoOy3eeoIT5+50RyEDBVnYr6Wy95yUAUiqCHmycg6s0s
EP0AGi68/6pMVZwasO8vsUDf+udoGKLSYr1eRnH0wjohxacLop+qik/L8UErWUZ7
xEaFXCJKob59PBg3oWiq8i8SiwpAgh4yia8+9E5EO40Aqq2hebNqdMdccLRYhEBb
CDdLx4A2D/QK1wFOytKaXXZFolF8p2FcyaJwIUdh+MmSmYZe2mONrNYHDWVz4xzt
M58zAQ7Wy4+NiZ+ws2QVbFwlWCWsZqDknQ6E5IFhajpQduG8s5m1Tv3F9A07VnSW
f9hZpEXPkxW4ExNjfk2DYVygoSUThUjsWrpBh5ZjVBTx1szPgCOJBtAUciGnvTbn
n9M2vQCQE8j7ITla6eFQbK3eTYb4LUnYg12OiTW+/JLkL/lv3io3YPJ01Zla9Rug
UZEMoad2VLp5sB4GidFs2SeGz8tAYqVS3iLh96C6IpL48mT80GR5HU1hRB95Os1/
QlOZWUnOTrWcTAEK9JUO3X5zKpTjxJgTZN74fYZS3p6ih1ft3o7I/1335bb/g8nq
0pE54DwjPyFLoCJ8IEdcWkHzEKT3Hzob9KpTuYy1UiQRufTN680DXsrzQnKBByzY
rSjrYFectkibLYibZUCfDKs27PmwsRme09MotU20wnT1/3hH8ZpvVfDCr6Gt3dER
AmQYKkw+uozcYRTsLbshFpveHCWlvJSqamaeyY3Z/ZbQOVlESJdM58WJeEU+Y8Fg
+L+el1FEiqiCpiBY7p333uCj8iOLqw1gWizhBVfT91X5Ny3dr906FHsa+a+Vs3YL
JcVxD/OBzQJFCKszewzp3JIYj4G0Vqloc3nzMtogeJrqwgVWCkyrkwi+X+TB4jan
zN1/3NGbxatfrjcM+cN6GYBNVDJrQG/mAoS3Ciinrgnjf6Rucu3ZxpJi+WPBf3eQ
MexQ3r1bXcQ/IDDuUDH8JT4CJ9tu4Mc/J1OEzKw3TmbUYX/cGY7VuQyS0FxN2bbj
/szrrnsnPcWSHlJMzzkh+5PLm8Npa3EHBDfr8evn1XZhB7ADjdmxRIuWJjQaYkPK
rZCPD2mymhk6SF9tFspKoqv6yeYbGz4r2MupPXWqPWx9EicRUhXb9f6vBMYjhmR3
MGC5wO9jvlK5qJ8MNeVFd1BGTIH9Opbis3TCFLs5xI9AcYPa1ersvdoOymAfil+G
ovCcr4CL+63ix63NovcfCdGwwTA5sW2pejxQDHVckw9LOJT263ygBiS/jTXFdWTz
8iYsQzhzM9pxwfPCnkFxJOw/6a4jjolpdTOR41FpwsrAC/jg5PUVB0VZoVBPmDkW
wnMcwsj0BKa/K0l9Log7ppWvvbTZBbaoSLRM1bfbpAFrVZG2DF9GNmW6HAG8gLjX
UCAWt968Usn/7RldI8bVLFb2/orqEnyHSMj+1PtxNGYUDNYQYLxRcMsyPS18B9TW
Qf6Okh3bSSd/QGNJt0HgmYFZFx7ygV+DolYH3SVZ6vtXoGu0a5bqjRVk1MznyyfL
yKMITW40NeBOTd4CgaZaVNNOVUaCB2T/Cbi8xGSC8/CVrmh74JTQ6ZT4FUudYmrq
4I5GiQF+TRfyUL7cQVq7TWXhJEQb4Fh0DLlqoBc+zMOz3Ls/YThS/wMY0pNOZadS
roBtKkrTU5fVT/HW0do4hrKuxP8M2w+D/9YGq6Dx5JMpYvmjKMkeo7+HSh3YGgFa
Fu31yP5hjy9MDjEHAGya85t1meXQFJAjYEg9xMIWfXCLZk3fFoZRWMsiIvBOE3Mm
3OVZieE+LkV/sEiDKHJlNXNvrTVZZPtCPk2f/cJeHXv8K8oCv8d2xQmVJ968WZMI
rzVOFHPcTpiNguWzYRyY0Cr+w/K89m/SbDxje5cnZjtR99M3ipsnZ7Wb3+jo3ccf
2qW+qQdoG0UXA4XfH2Z7fZCXzNLdeIf4sM6TQrY/WRbjbe7RgoDfm8SNEBy1W+8C
fNYEqvgeDsPPDfUERD6HcOGDE7yp1/dQm7fSvDxt21ZIPSWU5uSaoqd1zAufDQkV
1FJvcygZ3/UN5wxzttY6GhX6ohIcDRHJ2j9/nM8X9yFkQex0sGcE/B75L5rBb5xt
gwDP8ppOhk7fMofbQygbWXo8J6B0gJVwVxX74agBZAn6QQYwJqSEY6JLwd6pPoYV
COxz48OkJfPKoPJhY1qp8SiihPPXvDpF5TVkXTl4SrlTrIdpxP/55k/wuzj3IK+L
xoF4VkPyXlQdPiKBNV9uXTvo4+HxKTls4Z6MlT5zTWIvGBJJJ6nY6UnOPbWRthTH
ObKWSxPOUiEmNtgVhCDQ/dZzZC8G0wFatjy+urO136xWLwOqpSmtcYQ+FRdlTAfm
L9zsB8jRlLzfyCKYO4JA8tfsG7JTpNfoeHFDq6919wsLZQcSdfsCPDi8/cmJNJXY
JikETrkJQ1pZbORhxj5IgEcx5qvvP382cTgahrfgsP7EQ5rUFryBwTR+OM9l4Ycx
1YKEsVQoMrQ1SjePL8zN2s7WFkzaGCJlFk8Q6GF7r+B+b6Gr6FxZG0kH9kSbQmrL
C+pPs440PW7IGm402L7/MVnyrDQlwg8LzrHYMXyrsv0b/d0vtZkZYd1p+eq575O8
948ZMJZx0r6yFGnbV7+PgROZUYc9FFQME10ErzxZYbODdW30COnsISxAOGpqNRLW
eKy43GN0f586EM7ngdjFsOlubGOGKSD3fkyRmkZ6RI2HiH1v6jsurV4qFA9C/mLA
Kr9w5CTjDKcHSo/WDz0TitFZgw7p/r0sk72teAdOEU0CLEdW+viFfvoFtEqygZAc
Iuxlvz+hG/lq+fQjvDLjFdKDqCPg3W5lFl3ggp9lWz+gSXQa2SAx+V1BqNbjvB3q
VWFUkW1GFcdZ03P/cHi9+x5DGr82Npbvi0qwiBqFSEeFuMR1mJOgmuwnBA6c/X6/
XmfKuggZTGD7dzQZ6N/lh5/IM7IxtgvZEJ/yHK8h2y4Vrb0CFbmD6eDDJPpSXXnA
o1DPeY5SYBDSJVQfcJFFIwMu8E/BwVpWKC4KAOEB6hD3Vwt7JPhc/TX4tJKVmEtg
KJxCZtTa0Vtiqt5ndsG6USlnUryk2roWqeK+/Y3l8BpipbBQa8lrybVslLhY1DMM
JWtfeclM6NUT66igFBDJ08s5joVu4HPUWfPmlWTUCkeVBZ8bQBvOori9lm23Q7ss
5fYVwVKXTa/DSrQsjJyL4RqvP+lfn81ugD5w5LR1cfs1yrebt2CiJ6gwv186ynM0
fdPt8Gmak0D4ktSmYSLD4NOV1rXmxetGI7a1qiKWHWTcO3SPpi9bxeNzl8NhQN1h
3iQonjpYicEtxOQmbhICUYjb9XYdSiUhuTSg9mBjyph4slEWV9RJnUbFqPGtp/48
CGrmOFRcpLZyr1vPiPXABeawkrFiXAPpyWBBlZC8h3MwItCAQp0uJPMuSRyFIDhW
qjbr05KrW/xQfQMGS+SikYoJLHOjRIlkOI4I78ErVSElGD4GNzN1q1+GCd2siyC3
dmhxESG1+dTOKvY6p//O+UzbWN17lXOfuWKQDs0o76SX5hRTF1hxuVzuLItnbegb
RG9qHfMB7okQNY05uENyNBOXoqRceFEQ20VOJkql6E91tylhlb17l1LmjTjxLoGs
GC9enE9v8wA5Lrv/A09QZ7ImnXLHvq7npFUQZm9KXStBNtLIZ6CjaiTPPwrso2/t
X25ZZLwXRT9hW4l/EvGI+dpdqvNBH206b/6rL8QCSurTbAxshEd94sip4E1MZqnn
/7JS1Ir1JI9x2p2+8mRi8jf4mcNYwOL8fNu9qLsT3s2fr6NPVhEhlk3mBNrVApq+
6c4lrOpuOoqvAzhYwobMmjPCGBnBA0qevTL/Mz+yYClmGxsibUjFdbNvxk7SQr0j
zevgfwkuW301eiRLS11UcxDHh/yKKJdXG+sth26xQeqrmzbaLt9GX3bqZx0qUrrk
qva5AgfmXIBM9pgF+cVfbngZbOQWozpKcSRATZCydhWvzZhhttQ4gs96w1/oEDle
zNC8jRNHE8ZBLPykaVgLTMFbX6vl0/K8Df2DVzuCb9nSJVCPhovwSusDVxdkCnFs
tw7LGRev/RlTNyc2l0L1GlJzf/Tl9jL5SL/vIdu0NfQSktNuhEZY2PijfgmnLOTX
0sc9z24HyHorMM+Kg+3ZubpXhrr0WcwrH32Dd+qku4HcxEoyxrBwj35rjRRRD4Qc
+GT8pArVlwx5m+b6oSl2kEah6QWMHdc3eBmJKrXAnSeQaWIjgi+Xg1ub7FbGlbwa
V690h/EC7Zi7lgMK5Tg+klpImlcz8NWNQWMjEVp9a2b8JXyZRwpYFZexcbpDM1PF
0oGQbq6nUnU7LSWJ7kKPax6aGGCRbhJ91WrtX1d6xmD6FUUNDfqSlxn7OfRfZ/J+
VMCgLf0/sQoXe4brVBvwjjfG2eowaO8C6y5VTXi1p1ZvEMesBu9bCXF4WsQBQQgP
j4YInJJ6iC/PFSXVCFEY6i52B+9XZkBKirf0JWTSkYZfMO+NhTjmBz70t5WA28X6
fVZE0QwzV9bMwNq/gbRSIw8o6N/1FlcOYfWsEwr67C2fQwVY495BgRcOzhrQkWv2
A48gHJguf5S7Cv9YoWY1JK2CF6tNQXb8De+9ynFGSQMmcMyakFT2pHkenjOu6l1t
HLy4XDzXzRo6/6pJbA2rWcLsO3pM3c7MavFyol8kS3xb7zUtVKtPQs4N9uPzmQTL
ZlJHpC8pb2lKowtqJE+PGiowqvx8td3akxkknlBtfBeOgnycKeUpgMR+MX2J7rma
zK4kNGW98VC7EDJmdE7it0bzy639FwUa1M/xVVQUofTAlhrsi0emigwUPboztzhV
miEm5DIVCD8YoFgtV2q4jF0vATL5lrspJrIbQcd8R+uW3gkSHugoWqrKJ9+IpUnV
zyfkkKjoL1SIzKvFQY+PkaQIC688qUNbqxhpcR/TzfmYYphuY2uNxrS2GTQujf/h
B729kTYooKFv5OLa0u3uXALWT7W52esRNfAvyVVQPlsedU62k6ScdCVuVynq35lE
tfMd0+1nX5DCh61C1szfmYpDdEDojrcbPefsINdIsCsB3CZhwSi7fo0hciPaMQDq
xtKQaaEM+UwzXNpDzR3oXkEC4w3WRqeOjc6ZJot4uG+oy6we1IMcY6kmGZjRNWMZ
r2yMGOj1WTWFdFjTOnjqN5ARN86K+84Yu4js+ENX/ho5ZhTRwBd1T/DoB+PB29kz
qa/PCUPE29qbuHH5wXVeBx/SuMVVTU58DKnPxEimUcXBPa8+/iKLGWL6FcsaSrcl
s5P8BjMk1i13VeY87VdfakeKlTfbTkcEyrlu8CDIsonDOZYKs01gUwPho6aS8d0E
55BMydkuhD48GgJRSDkVHwacKv0ujGb/CukpaDvFL+l4pQLWh4kXKb1unRjnHg6G
dMmZ5a4MCdQs43+xBiGtl7EeC6Q3LMVfCd28bYrs/mVS0gpU5nc1H5DKrD5LfWIR
ajcdUNaPQoKh9Lwria9lG8XHhIMg2kGPXJDIxAIpckj/ZLTW4ahMN66B9c22C+WP
bU7Uum1GRbzMDcLu0SExmEVkfgBCUkbYL86TvJPJWJJ+yEAAZ+E6hnBGwGEMDmfa
tt+vpt5gOuOFAzhNew7kiqGiqq3eN/0OkRwGnirA3hJcOvCrw6Ze1R0qaz7fljSX
BqP1CajwB3R0+Hy4uW+rX+RM7PP/x19iElxypY5Rxs/fDJVMgd+1t7Re7qOm/7pI
Iv1GG7wHjn8MqHa9LC05pW9p6nVCPXNrfQOADMh9VyxwuuNOkynY7uIhqSgUW2Sg
iYVyDrTI+60HhY5yWdGmq9Oflv5kQlHD3zTeshDmJTCnDm+1uNi3BVfLCMRejGRs
qzUQ+/hhgeV5kIz8p0JZBdlbmP7MOtKfchE6A8q5Kl544yErMWwAimtqVJKO/bo/
EzLX3LjY0uZXULm6km+03UXDagYZo1rWgArr0LBQQN7udrH0KOeUT7IF/gQfuG5+
nMkWng0tnnLdLpseE/l2o50BXDeDXDj7yZYzetjbXujAqYMqjkhQ1hjThwPh6RL2
G6WFPoOGgWrMhpsGgxhqyjkblS9NH9+R5JOSYrVd4j1HOKjnd5OXbUSS5jp147ov
zUp5/YyJTkAn1uaBzHG5OhjHaFkkhXDr3vqkmYU3yN7JycnwXwLMOT8u/mce+dRc
DBqPoWDoYaogGQpYK7zTojzGL6Ymfj0W0RdiHTrkTSOW6LSn3FKYRxbyQHzw4IBZ
a2HhJxsnPBMFla7RTSgonye3qnqWp0eSUdQDY4kiA/hz84Q15OWLmliBbQMwYsc+
uT9F7bJA/C1s3QAgb+Ho0zX7bNtfinAI+k17a0WQinUErqL+6ewqpo7+GaL9Z4EX
7HZrfHULsuntu7/KNLu51Jbr3E7onA07Fi1xHY7sxC66oqaK4mTAb4nCHH8vOCC/
Q4bMhOq3kaOyCcZP8f4aRukr2BAkZf0zoZZJtbGj+otG/54qA2yorj5W+WRY7sss
VjqSeYOsADP4x4iqm/Jw+yLwYmxnub13jv4iT0W4fhNM18YsHpLRvDoZ6rGY4GT/
OEFdQHKfBh5zwrIZtMpxGPM71igDddGhBNvA17CVjf9N0iOYup/jRfxZB5c+2ra0
C3cilhuRFJ97MdI+Wh8D/o1bgPn3nJzZ5lnggPFvYCg7goEifjWFvlRDOlPouwTl
7hlvA2wN2zZCVvUBnpeNwO4C4uXE/WE+7AuBLynrjtlHlh80qhw/Pyp7KTne1GAT
bqWs4+o+l3nyhsLCWRUc5IKXuAoTsGNUGxt5piJZGBPrn3oXlWyHInnA7oStoUQ7
4DR12M4b+96wmqA9Yd5kHOzJ3jGNreir6Dl1TfevFUeUSDRElhdkXklcZBFXpdlP
+F5hZPa8gMYjN8z6d9OFiWSghn7VlEJIZa2Je70J3lLRRhyiGSspsF6ZmCoeUD9i
1hHclFRVDMQ7uCZOFLRMFvugV/PWtZsgUUGo0HVHRYQJW+DmYoYBe3gc1JY3LQKj
eMSzaHXwXOZV1sfXUCDoSn+3U2edj5pKwCXWj4mIVosNmGOUPYWIby6fupGl5P9W
YT+/nqbT4iva5ljbPegsqMyVvR5xrzBdsl8418i6PvuvQeacCV8rCilxvnhkey7k
9tJVLq2jGBgc31ObOrIRmWKkiigrcCpBBaxhK2gWqBtT5oXol0R/1VH4AmuQXCF2
rTQSjQFq9jNf9B5M1eoIALlr3IrPwnrZ45PYKjhPUVJXKzczpbaF7MvmfhjCjPUf
hnHzdPezS8+PkgBMKd7kUUBdKe3z/sp2EpVAnK/b3DxBoQO9xjBxmMuDLA3TtknC
ifBZf/x5lmwUuISjUxpit2K2fetlTKDoaaNRz6duQuaNdaLra851f67ZyMj//Hw1
nafXSFi2uwH3zsqvBKDek00wXQCTUJixCQnmpgCNbpMx7t6UHFC6zqbE+xir60o8
59yaNP1w8XMnxbv8tQVwkyfua5f8sPQ+zfWS6HMMY3D2d9lDPbisGduC+mJDjngu
OQph782uaRDWqHW5mhWG6avtltVqGRR7YUQwYw5lbscJskC+NWZ8uIMUgilqe01V
lyk9HjjlikM7b9lAHbAhInimQGYTAAmy7nXnRMDAMikB3V8xr4Asg+vdtEBi6VpP
zTVoY83tF7bmKNnN0i4I+XrtY9iTpIcIkOSg5S2EN4Lzyz+MhHytQBhEsDqMUGKw
ghl5r2zJg273v089bRUYniu4NUrxsq6tRIYxEvGGlVyZqEezBB/u4fYsyffac6C6
kqy/ZJjhaIHfz/doCwtkKlFe8q5AkX3O3XfIAzM1D0BWaOTDklub8vCPQjZ3uzXE
kaNeIB5tBVCS3HXFF2jvVsnCdDXlrmBDqBcKDkTQEEHRFQ/78lTob11XjabfUxki
0bzr7hrGxk1vPQKiBUIIRtxDw4zPLSzhO0n5Zj4GuYkpLKLAgSOibCCBPJxpGmLo
+A5X/Sv7pZ2r3sLIFwFkoMMa/2FX5fI3YRLi8xtSBOLYC7rttJt19VSRhRnVePit
vFdGXlTsGgQqIK33Ly3HAKe+z9J+WLPB/+AoRhOuPgUXqDBV8Ww7mtg8JWtafAGw
47Jap05jwDk7d88WOSO3b8n2mC1rWgI+Q5aN6chV9FL6TsFmLqtf3hYNQntXgI2y
po4SEh8474iVVcXamyBPhhyn5Oq0Ay1Odh+ucFInboEx4+DMOzn/8HsyssH2O1w0
njIgrGd1sNKClIWhoVDayKMvgdJXOnTzv2r33MD0jMWYs1pqY4Z2Cu/B6lVyoOSg
v24b9SQmznXQG7OQrtjwWVnX+OxTbK+lTcx0YZ8I8GMBMGbRKzGQag7trQOZVHLF
nV21jCMQ09MXGB3XtopWqlPxzK5sdZJ9DCf0wnL09YJpz+w+DaPPjzvk/DnCCUpY
4o33cG9Nl2c0j/Ef9R2bixfvdnAHKzjW422h2xfjJ17Dg52ADd++CndBf+gqROUl
LJ2rcFOIyImNTMR3d8c9zKAjKVA9E58xcUvd0x6P3GacuQF/C9nb92vOY59h4+IO
/wPWQoQgK2oSj55L4S/p7P+bvMN9fzWwdNKyZNplRt0IfSqhYB8MbhHoZaqnyhCd
OHIGS5n9sCbZEy1NMOgfMLPdZT1ISAoeXZkwAycqdkiVqTQ562Np5+1/7xF//wnO
tlOlD1Y/xjXWPHJRzaRVjTDyN2umcptujfnyRaCJcJImAHVHnl8w39zLncU8vJWz
NtgylYP068aZS4UTwBBGbDMO2mnSnYM21jCEs0YgiEnjnGL40YYdMoCfnIjfytGc
OayJFfkYcQHyLs2QguMufBFPCC/Q6h//9cm8T79mfAOs2AayBRNj7FQTEpe396k1
UkLzyZ+22NgLLtWfD6lkqOv8VKQSNOW1QeOYWEWL9ch07Zx02lQQOEEqpFBVNwOh
HG5zgPQVTu4Wr12EYveLWeGHQbuYPy4/DshBSA+YqpQ++oBqg4jtvBtlxhpv1CvA
oe3Q5uQ4JcCFi3vnyS8Mg7cPh18zK3bnPQsvZrcQFBStL2xm74I3NyjWYej+bzFq
JViCXZPEtca7Le6bTTG4zuCO1eB9wUCqfVEtpd3CxRy3NhCpgr54i+drZPda0UOn
CHaB7Dd+KVrWBEiDpqeVQ5tTkZ1IMPiwC81OAnx40mO8eFp+cfYbFCWwtJPcEQxu
BUZTwrjkxpQ5G9O0N50pBOK2fBRivZwFdV815EnMSNgwKqHrvBiyPgunsgqHKMKw
U0fuLyjRMsQ1Yu6Kk4PKTPnB3JWZ7z2KQOwUkEpKgFs+8MWnqZ/FTIHVh8V/sONW
TkDVHCkGcjOQkt3FkMCb2Wke5n2Or9ExovJA9k2xuPEYVyrkkkvg9YGJsmwSvdDT
bBym2HAQNOc1FjAXvb3G+lEbBheJkvVzs7vXER6sKRlAYBWguDwcUy67CUixnnOa
FmFdAzh0642yEHju3oK9praos6NlAJBtQlBJ+EKlmcY5ZYL/0i+i4F30kv1a7b/D
nzTnILdiydaEDGCsUmhWuqoiBGQbbpvWmR81VG7vtyVf0clO7+dKMxHG2HQPwnTr
g99kCOsLRNKEzz5sv0W+d8P3w9MUSIhu5GbeV6T9fVgnih8kLyJDVinwov7hNJ3q
ed6ZSp4A9s0RvahhUoD7WYwKyhtPc+GcaR/ONApkLzk9jVRguwGt6wg9cPUvcyXu
jjRLe7YXFrOr75ngV7NKYGkrWUa5gRISgq2P7vTOdZ/DHg4RfYld3je2EPS8ZZOl
Ulw6zjxU1QiSdKkb943lt/SgD6yMV/xynED2n1dzFzcCMdqvNKq9aefGYXKleGZt
AT/jV2aLmXL1lQ9N+Ns3s70BBIOqWY1OVGrMiVFC9IelXiWBmlXrU4VFHXWCwd3W
t+K5LNjRnTDMwL3UmG0/kvhUM1whFIZ7d5fLEGUW1bULJgb7NcIrq9u1XYaZvJVo
jGPF06pY6U/7Qtonqc5Q8BUhRlLMdSncXSvipHZtLAZza1FN+Klj3xa/nU2PTTZW
JBLQjxl8/VUFwWbmXgLNqJ5P66dSI3TbMQkrEbqe8RcRwAzlEy7JeSgUvUvPWrvL
1QdxBeALyBl1ASBCyurnn9D2+fhQDvPBRTu78V2v7CSA4go1BLW+swvUhZRN91dC
bt2T6Ds4NkbQ4DIt6TOiiUdOoUEL7leB6ebYrQ8dCgOdYADySX6FzQ8hF+Mb8ldg
CVaexVTJoyEhsJMIolMifF2kclIu10KMSmDgts2eRnZTA3jyV0szO+7eIvxuxeOG
Yot0y5rD74cCyXGqarP94N4NELPDYUvd4G7e7Z4jwre6EgX8yBElRzSxkD5sD+A4
8Q1BlQwnq6LC3oQT/9VOuawmfqSdGPZqjp2iN4cWJQHW+ZBIeMJYKEBV46YjPHP6
tQyxAU4iMu1lGfjjHkhF5MwolzZIYtOnXqJ29mDEwJ872I8Qs2NA0pO5HVA8cGNC
MTu4Hf6Nr6wsClYmmA1U4GI/N9vGVUH5espheIEXzHv4Dj8oLrTgEftvDa9wky9l
w4ebD2NfzFV133KNJ0t3wxXBv36dQfjCTTqf3F41LlKbqEPhmQKA0BUGEz7a00vI
f+LMYyJDhPGCXb0oyLTFoD+V08QCqt//WmFFr6DRST1vNa09jnJiDHt4m2OcKHaB
f5fGkLERa4bYey6ioVgkz8TAd8qLgwIee+gLATFPyYMaWQ4lj02hFbXkW7S5rRNt
2g81cU5JmJW9UPtm8a30C/p9ZkW38RDbf1qqRaOHwaXHhSzZFbBkLkpNi8hFQJP3
ccu1xJYm5DKLmgqbeRj2AeCC6dvgJI/2cCmDJ2rhUdnSYln0jsL1rFQ43aa+nomL
nD4shByEztJ7waFx4ykaEl+/hpwe8Yent84nAiXsxuAlvYVeqOmS1PpYPSQdgOSj
GVBkfMNEQVDQq2TXyoqp7LSbVeKhrMeXe0pvz0+gaJIEQrDEDxTXsGvmlefx5vW+
F1IgqOeBexTfNflnSYSfvFXIQgeq7XaIIQvUgBD5SN1FiDqaFnFK3ATj5ovvY3Rh
xQj/q5V/6806u5hGQ43VD7YvOChKkgzEjLbuMd9sW15SNP3+iWiILcozGwEnbsqy
FENPm6orLxIG1Ef8i9SeMHO3seCV1Y0R3ayVIlU8j0HGModvZbw655MoWQSxiAm6
zfRErD0HJPvObSPZWHGTkm80zHEkLZ0KhyRfGdC57oKVHtDYzHmqimyYL726VPrk
tNS4t9AIhIpXT3uGtgP5yrF5eJQ8Uy5Ap3btBn/49ieR0rzUoc+xTtUrxZGTsjXY
+lP4cLiFQ+hAossjiXkzZiIcC3E56QBCX0Hf4P0wqQJWZNo0ZVZhRuyCcJsjIxhr
JAFLMph8uhUKyI+kmxVdHvILFvVE/ji9EIQQyp2Oq8fEwyBFdxjkhYGa21bPwCed
5iH8YwulUkZ8x2pU4v/Yhn+/vaU/OnaEv3+y/B9nt6r66AHkLn/TeyCjIcgoVdeM
pGpAorJA/c3H/i+e+z8LSzFOx1RqJJz4BudtIszrlLPJ+DHgdwkR+iXKR5CmUMYj
aEGShMnwXTan/lvDJo4l47FhSkyfUkqI0XCDduBQTfoX0M7CFPSSktrvFUUDuiTT
Oe/psv/Col3dIdUqv7cH2P/otgBUbl2EwX6XXl8gy59A0H/E2V80Hwx27Ha6kraz
fzITwd4NJK/SXVlyQauZddn3tNLHc7Ju9NHht4Z5LmLlW2a3FFzsIkZxZt7/QNwe
KAV4eYCVuFKo1KhMONslLd2a3w4INEWL3/NxmxmvUBTABWr9ONYm6kdXlxaP62Ns
NvKO0J9l7vun5r081LZr9/UZ7YLkmVrp+I+1DYR2aChUjFVwOjYHsZ9nQBIvk1RE
OKot2E4tkbcJhMASfkK//n+tVr6yCw2BzMSVrl5IyPql6wBDAfQ9j9rN3V3YupZG
RJ9nbauIfJEFZkTRrBeY5P9nrOZjzMBRcRiLwfRR1Y67UuibEn40wD/XaP5c7Gto
M76W0pkQHLH6zgj90UHAqOSsk42kzEZP7+ZFIZFki66V59zl8GlUZ/XwWclITl56
14zAUtBB2OH3gleqgG9Lfa6nTDKn2DFT9NyJ1A6eha5TjaUT6ssjhnzxcloKDd+p
oLsNbFvwdbeJqxQ1w9fiVOG4QrlsQsfejf9gN30F71Z38Zj6PUC/qOmWTR++5vnr
hfUB4joN8C/U9skWxoERI3z9C8jksbyFA7MRqp0jpPseUOxOILDRENGU7QTf1ms2
A5dqW2L9dpLZFnNAcSOSvfqwpxGV6PCtZdTaceIAAUTyDFiA9AgaCazEah4Zs4O8
mko2JZrYO1gwaosv8zs43IFh9dvBp0evhmcgOVIlINF1zzkD/jXXpo+8pp7oBJyB
P4LqcJ480rudB9Vkb/G5dMJpHpkQUt06WWe6EYkks1wOHQI7EaH75v9HrYraBGH9
hHhjTPnKWQfvNFGO0CMBO9WaL36pImPvqI9YrLM6wFRP1IxiXIgjsAKHFtRK5O2j
VCZTNcIfI+QJAW3oMalE1g7MJAEscPr0m8xzTz9OwafcvcZxZhMqQ8p+PQnUSRV/
HBjNX/XCkz3FUvyGZ+Z2UGphIVAlRma8T/NhSpP1tbFcOw99NgpuoizQObEUKdV3
17n1AbufQq8ZEEN81u7DFn6Kv6nO3G9H9EWULXUiB4MG46pRNzm2TgSBXltAKTPJ
bicRJDuWedaVlFtm4g/9SqxeJCg6lDIMdjNPSlNrmBuPAvXFvZcwXWK1dxPswvAO
MuWHCLykvOcVo0drQHphM8Bq3vDFYIaIAJQTUmIXf0e2AKPX/ZfVCNJwKkfCZuRV
tOAix7bmNyyrL5uIHWsN8dudlwJatTdl3vNoAPwpaO3YEiT1VCJ2EmdA72fJEyaK
9xX1MWTdGCtGVWux5zbC8Csf2ulyUCwK1TDoC9SbHfWsHRRNNgzWySlG4FBtvJaZ
eBEvMIF34+u8odSmDHFRIX61mZSnUPTX7kqU3QzCFpwu0cGT8Ndiysv0hFYChQCm
GA4FCEL41w7p5pT8gn+NGNV1hOZ/lAVEBecAS0uckHe5fgSiFxwI1x0v1rdlB/Tz
lcVnSEhDN0FlzyNZUcL4oO8FrV88p4ljsgFfRPp74qAATxHskRny0k68rUIat9+I
ZuoC7/WRXKQ0/gYZ9JGLeR9DIjdUXvZ/W0sgWpSz8h30PlCMZvSgCEydeXxa3cdU
u/Uvz/10vcUqVSRSF6je64MUoCyvzMVps46EBczT8WK10cv4iS36CZHFkrK6jkG2
stWrD3C8PRkJgzPDbjFG7IXtEWwW2LXYNboeuvNW9beBjYsjSvHXihRUxfmpcRce
1XQkeSbu0eomrzTfvy03QUY7/Qc2t6EfA3qRa6wlcaX/6bygwIVC2LZy57rPY9mS
r2/so2HR4wJQuLw5WimFofXHBvlTiOOmHxSEzHBV4oxVkTFqkZolo2vAs8p2jS2m
NqMETUwA3g7cFa1iWxahhPa4kHJaSfSRMjl2Td7V7oZclNlTsNf5C/37WDIkLHgs
Dlxxhhr1MljSC5xBr+u4srRQcmSP1qOQbjHre/mV8orBVfPg6XKZPupTdHM0cYGZ
PW0yCFqZ/70WmZMO0okrI18/LogyxELnbo6ikKRtV1pTlnFyFTx3LYXHNjgSujjp
zED1ql+quWT6SjknRIdVSCkT/t0v3Z8UZZLdxmbolTFX/Vmi+UHfmpEpsZQPouH1
HfaXsUN5y6vZcF5NctjZlUe0Y0QIj/ezcAvMDY1QRM6MWmGEBBMJnVmLzAiWTIXo
+wV7IGiruDusWFKwlCCI+1EvzuQdgy6aEiqOeNLCM1kMYFOzusBfwWfc+hx5qgN3
OZTpMKGzqdj5rO9XWf/gQRKoNS7oHsFrDo38TqWP8GTYstX8yQykcTRtM/4Iq+9z
/OKmbkzpHyJTnCtQk6gvXbFqOaauCHnlAsBw8XY/+rqHYon5pn8GgpR0IDMKQtl2
TVhYKCEYjSfaJpRsllwdP58aMm+L8GMb99RbJIHhuAJDUGYUMplwYG5LkSWam470
kwrqfjVRhcLaSBNdarTtcxqGBHn2dcLVf2uPaCX/YazaBOAtHyZER8mADLFvCfPN
oZelDX8ah0cfQFCb9GUsJ6b5ucO1UEuJO8wxVymzOVC+CNL2BCZuu+DUINVZz5+D
jcjGv56Rg9j15DfISUjc2PjQ4TrIty/hl6bFgUrI/0ccKKEVEweSudzr5mEuZyFh
Waq/P+Xn+Xe9fh3uOyhRM4OF9TjmREqhXKm1bK9mltj61jKGFgU1Rq4vF8H4tIJm
+yROHzMFmxvSaLPPdmfmi+cKV3YlpYjsFx4JStCsRpB6c4KGPRLg/dSXt06eytTx
c+UDqYGF8MmMW0lj0ac9nAxhJ1r0EWisIU7IdWZaozkMpzbIHcF1zvxQ69IHGp3a
FdHN1xbFlC48XQNv8wxtYGpKJLhZmvYxshR6eN0ZXsdR1BPfwM8D07cqEolTzRmG
hOFOHUIgZFldhRXLqrkaSPJdeIBnV+9MtvIgFpja0r16J31xBU8a4XHlVBVB7Fx4
LcL3j+MjYUjdYDLAzixhylaWu4IoM+iTTG+9GEuW4BrMIpur2xgl4LSlExTToHOE
e6FTP8gUdcpcBOphHDrjcGoE1+nE51MVn5eetER0883E/0NjW4ny9jF0AK33Kfo7
BdpJoH0qEPk+BIdk+tJrNAggltpqPev0k3Gzm85K3TLRsxiKnYSqTUIFfqHOfjrl
I40yISvGItVsUuVo9LgtKYusy9OvxgoqhDrItMlqK2hEJ098PI6vx6LsolnFTTdZ
iOS3ztjHwyMDkdgJCkkOtNuQwrkFLwxezf53cGhMovc+rNWid9ykqKn56XJ5+LeO
a5QhQu4/6Nkupypw4qEriqK0Ln1d4mv7tGCKNsZMdqrRVCzkJ03QaF19oFcSSUVe
ddDGC8zdkvSYitvWYHwdNTTK+x2gfubmDHAqLMqVS3bgsx20VoHH/gmZCEZEVgQY
/fQzL6U7etaSSoDKce5MB1VCIMCGLL9rtXK4ttmMyYOmc4MKFm1KpPCSCvUcW3q7
Faz6L3zW0prqhTJh1kQ4O41e8NVgld39A1gACHuJ36VbFtxxViBtkiMLkT90Y0on
/ZySifNSa39jBHcRD9DyFgQcA9vXJ5drO9i+efts7k5Y6ukgsDwZkK24NpPaSCxB
h6xCSfseBXrqj7FDCUGkPuABYCScZmQWrvcrw4CaM1mCALWQ+j1BQa/SRf3vijCc
qMjGDA412mBY7LdMvgsfLgoGk6nl1xO9bIPb/nt/CpNjtCKXt/qCD9O6SD6AW2cV
PeO0aN5mFpzQU8GWcAstnInJTJIRABnPU2W1GKjRnoiabLx73YIyAISOzOivgcAQ
yFmsXSVG2j5xqv07xi+2YuneTQvqedHlkzhFbATxc3AKHh8a5rwLuE9bU/5CScCF
c+knvkaHfYmN62rZIK2k3TUqiucSSPTTDTT8hIS10DHmh4DlLqeQjdg572QHZzdF
TnVYGHoYoE2xRjfNx6sbFXBzCQONfRzTDr3Bd8x9nDxev9AbZfKzVInENwPmVtZF
EyrTkRhz7w3c8L849CT4FmMmWLl5yUIJ/y6afmLW3GvVOiucW44u5Alo4xfy0Sdw
JenEvBf5/v3QHmKdAzPIl2t+ZKm6sdRH5x4bVs1JphkfGaP4/cgpdJ2xbrWmSgMQ
Ljsl+LgiXZxSZebDLfCvq9P8yGhW6ck3nvDra97ZxajmWygoQzuFj/oMv8ReB/Dw
C5uGdLvzhBAm5HSkET4nptKae72MwQWbqT4AV/6gcHZZnAE6Tiv3U7sw/iEBaLQw
docDvygHZNWEJY1tzJawi+OuWQj8m/xYFEbHma3Z8UkywJqXSAXSmwQcewQv7Tr/
xVW2JVg0q2m0Nt3FEMewf0L2CJYw1lBcHty23N9TXs+GA+0kTbECm7t0HNBlnxUN
m1jn7ZCL8ey/kE3FdMEhlPm20I/gV3SNc8L+sHOdL/K303gG3SFlMxTkJxkrahzO
UHhxfl/UvOh9zk9cag0vPtekuRE72xbrVOYMsaInUHG89CR1+3JTZXthJGtx17y4
Y3Np7Kwv7iqDA6U8u57illpGA+rp0xFJYxs/2EVAFK7lZcy5taZhtKDnJeB8y+6D
tfXtPbNkWEwsBK+iJ46X2MKaI5MYrkCBkNAwW3cM1PBNQAiQmjkmm1M0NZxSYM6/
rlJBLDZpNg9JiZlsYFRS7rfoX3fWZ+kVRuXLUD5WEh5GqCmQT1aYwYQPsR/HTGjR
Klb2qjAJsiZA+3E1avxNPqwk/6piOrnMlY70GsCc8PL3peO0YfYDlzN79CQlGxE2
iwxY24k8IGDSx6CviRLZD+1G1IppzXR24O7qQ1/MZP4pQOuEr6LnONUnNKFVrXml
7Eg/WvDfsRq82ks0kPHlnsRjOMZjLGkDhb3KiIxNIEF4CPCtH1bZJ8lBwmxvLsKH
ygQSGuPySGIWhJ+YtGFAvdbP/FzpLz9FFj2H9hgHy7S+LYjV03bDhzbDF2qR/yu9
mKi6wBilaQ2wSKklvFBgWZvx7PK9SKCEtM6VU3johW0q2KM67N7t/USiEN2Rs5/p
9dT3kny8EMEIvh98ZqW8JXepHZc5qS3lEOwOmNTRi7ys2bA/wnKKaeGxWNA+SSa+
ULIEbMwCIAjHSEECWmx1uN2Pf5EIZHyQukEDa//x331ueZZ0Pqk9pVZZ6iidceJy
XZA/KiU9xYyiyK111VbxLf7XCxLuR5VPN6x7PAilRgy65VMvCfkjCjRv/Z7zUMnJ
hhn6QkHebNVaQRn1hFFOUTBRtZVJcs8wndl33WYdJcVyXCD121DADBpigQkoS9l6
mQkgwukTSrpCPJLUEGv8PIsDSjHu/gdwIxLJCogugrmOHTI138wfCzvZiogq9U8i
/7A7Fi3KoAzHnbYloZcooyW4ea/25Kq8chs1kUe+rqxVVPOAGxl/pwO9oL2D4pvv
rvNlpKzASuEdCDcNK76PloM4yAxyr40uVgnGLwd+fW45F+pgruIPQQPLpnBOu3kr
ZBM5wN2zZ+ZAqQdCfpF0u8ifImO0fv37KyOAoJR3fxclYuUwsAbt8oDTdumMDcBW
a5CSPKqwUYUMS/FGawIcn7eqQDYzZs8vX5L7kEvMNu7L6RKd4Zxt25zQVVCcEcCc
YmKjLuGlLU831V8yTQ38YvqkRojovhK1ObLRaW4KZUTn8ReQCKa8eEQ222w0YyWk
rXW0x9YuylTodL5GFIQMns4Whr8Xw9QgtWWLpHFwLuyOfI7Qn+radjUvhz1LTvYQ
1Z7R8o/MWEqVlQf0mzODv6vTgF9J/zfwIYTiz8eMJIrsvAx1K58nkcSeYl5fmUn1
3VJF/g+VrRdzMGp32Qh9NgkKhsaSl+fyX8sewwyB3/1H6+/wyIJC59eP4w5Wswxn
cU7mufmWMY3RJqnt0XVIzNZ8nh0A7dyuJAS99J2XZp58XgtrvgSCA6R1OZ+sUEkb
xVlrvIfy+iEW2IgZc/PgFMMsuZunf41DH6RzqCQg+W1OGWziHbKAFepPIoIk9D5L
iSycfO60Q/1MT+jtfl3KxLj6AcCLI6MYwpIxJ7rL9+G61UZbYoYMoZ6lVCMDGHSP
ifmEsIRdIbGVHXX6Mst0Hy2PsjJpIAwfeA84c2XOUa8nFeUp0YLfuTPSJV7HlZ9x
uFTRag9BglAji9MaqV/SdaxLM5Q6x7Oq4v0S4RHs6wBlJ5t+vnWpGNkR9xOdjoW2
xMEXokdPLwR0eXTurXYHEzWEyPB3+RRynGGohJWWQ6qt/0HB5KozdUFLqTuOXQhn
pnSoXet1OM1HSeOT+lWC/V8Um9dl3o33J5HEJwt4OP1ik14DMx0kVQWJKyHHcn3p
wwUbYmSc3h4W2tSb95vcrCSsh07uRhBx2BsAzhwz2V3gKZ0uDbX9Zf3PZ5T41XYu
TuLKTnKBRFz4kBLFii4UK+OYYd6wsaUXVkSDhafFXPyNHcovcTE0IqjAU2ml1ZWF
LDZk+4eZmSQ7InKO6C/zH8dWyXn0870WAugZCL+i52DzoHKnzj4VS+XYsSFWrK+8
j23/kAsCSRGNxFh3JprvaP8tX1qPRF2DkpzoqfR8BT1J8MXDynsNdNOz1v0QS/m9
Kw14v+jaQet1mhcTvsRSnRtXr8k68gfYtN3mUD/WRP/CYdXrhsMDrTWVnjDK0ofR
Ai2bsDZlSk8pyM8AxYLne+xfsD0+WqWKP1F8Ch8JZyueBKBLk3KFHKF82Eu5qQu1
jO6YyY+HPi/nrAGx1jmCBwDF7MNcJbxlb+D+igxfp2uUte6FiPEVY7oqWZh0//tu
3uqjcqlO8HnRADqQKifL/E/zMQGB+tTzQmSS12NcFUhnMVGSks5BMrHohFqc4McO
4gOswCUvk/QnxoXHFobeguyYLIDeGO9KDDcaU1KzWAGepBhS5LOcJnFuN1yTzwc5
c+koZu2mrfKmB3NnDSEaJ1YZwCAPS+oZhjbAGy0rtMcD+aPwtpOBAj8LXBhKz/8Z
hlFsuUh/rtWlHH6pxf+W2I3YZVzRMuKiSK0a3LrWoAw3K72MWfgPR4muupdzZnOE
cqDLlF39Am75K+bTWMoqyD6nMVhlbDyDUm5Fnek9YANxTqfGqyGQl6fJP0hsaV+L
MnHo1VbzrC6gGCpuQ9qSB/OK+UqQ+PydpLtdl54GhlXYCCBXQvcI55O3HzZ+Nc9S
fXJ2q8FfJmUhvi1/Wb+Wnqg/uBL4CLXyCQCVlJcVUaQIykObntm/0QkLy9xzuOoc
7MIOqJ3wvKRZ6XzgAeMvQDQnt3I8FcEUIoUN+0X8FTKd0FlsAZL30DjRBvKg0/h7
BBSkXdWy9v0Kej6Pe/7IRTW3d2/JHiokShWWbkcrSlCAJXsN65G6QaLLxxUbTJTs
JKJfjYHgDN5ICo8iMtZPtzxZjohDmo7QfGxPNSyuCDVv9ltLFNHj6K9C5BNfB/oa
pzsgryNucuu9yOL247E92q+gigFKIO+CaY7sFpn2Mccr7Kl3ObN+gvVKiDiPteOd
7btQ3LZJBpGgGOKsVPwg6X7lN3TJwTo/EoWhVH4fH/qRYilHia9+tIdWMebR0btG
1oYcxHU1TRHdAQuQ83BgYyaqfr5pB6HmGAA+pa6oN/1dezjLTIWgX027yzb7jrlp
6JO1hu4GoEiuLeg5okDAolukNzcTMfK8xWUfKXvX/DvI1D80y33LbreBXXdO0FPm
jehfRFkBuSil8bHVdvonFBu9szBeZ7cd/s6HpIpCwUdSmqKIxT0l8P6jZFJEwLGK
QAAH9ApjNG/igSkvvw5cYpbYpR6a0+qmyczuAe/zt/ri299/sdpKCh/cjznCYvcP
JdKlQ7+YNJu3Ge/TDFJ+YmUFMspsPEuNfJ+Yb/rj15SIrK6NgehWVh0yd02tcWax
g1IlbQucruE2LIqOtcFqiHMnRnjyarMoMry8J0kXvv0mAjKv25hEhYsFUxBqaK3E
tQC16x7XidT4VwC4C6JQfIsi0rrBAfmP+k82g2zqhPj9vHEUmg+NB2GExVBHUApV
70pBPZ5H/nReJYV3ID9obv4ogMa/nYWjZ7Z1EAHiT59j2TMJBzCq5go9G4ruPDYX
Eh1iPy4QMhr357J+lRpsQurz9nsfGiIMiZN+0jkVF/EQy2hOzWUCfyqKeCrDkPXj
GXaqybCVGpsxj7WtCmLOsKVFrkj2OrwfPuqJiGYKfMMiri/WPwpsPmYoeJw76yi/
q0cG6F8ZcDKSIYEUD3CQcDcery2MyI0Bn1S3MOW97EYY/gqbM6IBx0BghMKpBajz
bqPr5RBXmwcHCsAP6T1FXuj8px6ZkHeOCzGHaLe/Pt+/MOANDhw0vg8A12Lb+5AH
pn1asyZjXQ2qY1VET6vGV/4xwz9RkwnYEEoyI8Aydwhe5qtgGJtd6cBXaHIuKBXf
z80D4XOAx5WccnhzPoOLVWTtoB0z5YCtylKpxwu5Sy8x3hVwPlsHWLnqB/APgBQ3
AYYlpcVdBpOBJZjmjASsjZQZ3HGWaj0brHVXuxTtMPB0nlQneUtW3mNh7bwj7U5Q
J1Qznma5h52YLppUe6haEYQY9otaOtbnCaw08RkRqQTJSa6ApsczKyiUmdx67ifd
E1B5iHx07ep/KUxk7uBTfZFFVe8fN40Tfp258zYmb0yMM8EK5AGESDrQ7Sy6dWvz
IBNo8ePTGKgkR4Y8N8cDEN/23+7jor1levTE1IHlT1HyURmXLZuf4xgXIEkykt8m
Bc8IuLNPp799Ls8wlVcmmtZV/5uvd7yp+gNlczRYNuoRDImFS3i7U0Sa+aKYViSl
D8gDBfTIrg2A1ib6BlFAFaDKagr3+RFCnEsod3I0/ceKQLr+BsdfTXprk1qDLFbI
akZv0/UGax5U6NxmWZrUWhFC1rCXSYeaZTnVHdzVRR544wOLeqq0nJvT3p+A400d
SUKqzkKOPJ5K0yE1RHL/2JRGmH3Uy7jZNDv2zB5UYEk8LAQWII314/30kniumJF5
JSm1D1uOMRUtGeQRiMWhT52cgYm5TA0W+lp3LtqggUv2eFpP9D7nJy4Rgr64ZRTS
27HFnUxsetZdQ/o0X2xygyhVuH/EQ1D0dfgnK5SSgdllo1HS59dV03zvpJezrO9i
rsCPSc6VCdQuZkq9yikHg2JWAIUAxksrSuNOVm0Ksam5Hjm2KuKTk1I1J04mHEDV
xUWLLbxbmkYV5/JHEPe9Mc8Q2ZU+kdWtSPtr4JjS9TOIeSGuHqicWRoklMiKu640
flm3dP8O69bbLkoEa6iHx8ifudN2I3OFcXz+IdzWr+RRKN4tBh+2FHi0H/6jn4zK
5dN7zB50TvOzSG3NCwcKqEE9AUai7VwoXByGSuk0MUEWcLq+YLkMZJ0DBi0VWPm2
7D0rFRUSf4vc+1yPPELEgufuIReE2KI81nt8sLJnYLT7ruE5qo8tvdtuCy+m/5Zq
89URmy7cYm25CXMaDDKkXmTbFTfKZG26jpOGqegAOOCwSdAdsot2psFgIq21nEAG
mykGTat017ChzLXbv9YdG1UVygoMKwmfx5dUe5cvB0o2woFQZwo65dWt5E2/VdvR
qcUBFkoDO8VyR1l/wSYyZLwPibLZShhwhzDyGJPoEE1tW9cB8gkZdorbFl7HzQdP
PXTT1Vtng6kUxQ5N3tn2/Ix0buZXP1Ckfo2/hbsxaKC3xjixUQbzrCDPPjwQwi3Y
8tpvEsJfetYzHlOP8CbxiFLNcr6iN/jmZqcJ0mE8kTqZzZFedwFK7fR9bLLH/XOe
XLglEu2ckXrchn0RyCXjM+rI1cGqWXkv7ysUOgB7gCbrf/KqbVIzEgMMXTWHnGjH
JxKIcQNaLDZ51RVUn/Z/2rF3V4LsgSn9oowNxetBrvvvq+FoVrZOw595H2umoyvo
d6EYGpPrHGaRguKGnuiEWTAE9qOpyRdqa972gRpFUHJWnT2N2KoMTSsL9531PF4E
whe1KO/EgmSdkqCgt7vXabREOivdDZ5b9ljR3tNeMljN/LXtOs1QjZhuJv2IhBSG
/8Ldw9LGBkym8EmbNLcHLovzSmIssm70O27NxXc6DW3PlkMi8nDAQBYOJBUE5oyk
iWyhSupAWrW6R9l5tehkkzZSe8llS2BNtoxekQZndnmtlI08Au/6RRdEfl7M5sAa
lOMwrz7Uyvklfk9yAZMFP1yumu3MucsdvEbeESjjoF6ataglPvXmihgpEFQ6Tfjw
LQgPdWYXKNqC9qc6CH+v5wK3JjJvWhl7yagbIT5oaKis6W2DdneQC5uTm8jXBRkg
md7KVOCI8D+Kv+iH3gyun2AYcmhp3atZsYvWdlFiqIpge+7tXiafFF+kYZzHaXjo
JkcZkDOKzYesZzRZE699rkteBos/cR6FmlQwA8+Ej02llrtP+3CrcvhOLTTlfBBU
/W14Omte5d1df8RBvvJphKAf/oz7t2C/l0jB6BPjQYrUN4CTy1fPobzWZm2heJOX
03Oiiuq5oqwEE2ZNbZR0wWt58d1PLJ1XgcWXcZJPi/bxXL5yax3NdGu/fRb+eEqi
S6pbIRtmiGEsrK6NCHMJpFriK9lOCUVlH0IaVEwl4ktej17G9h95CUKVwv8/KbKS
JnNSE4AQwX3ZmSQrsdmP78QEHdnmZNDxbKVqzbUTLC2oQcWnLn9GD5Lpm59OaURC
VXqvasl06+kKAqoxcD7VFpryRJCFVDxx4seHauMSv0tu0j+rkri3lZiZX64nTP/G
7bDue9toZYGqNN0S4c1ZuU6KOD9yNo/qhzHaVkb4g9Qu0hDQo6zIG1HBUbyCm+Li
hbLkP++WQOZCpgce7/ryGHgW7iRAN9NQoidmZ2zfuBCyrnJdL5XqZZTktXL/Mc/I
nyUnHQ4GrIm/gn2meuVxtQbLjgG6oowncL2cu3gc6YqyWpjf6dZIu5AOWQZUF7I3
bd7jFoN7xPqxzPsK7Z1NvmTieb4E9/xKDNbGLRXN2rpk2fP8ejTnJ2sZ77Mx65bf
102iiwCZDbCjIAiwgLqfxlOghq5g3PnavoSNdTZZQI8xURtbEcwySs5FomLgFynp
tILLcZJU42nLTLh+WEeZz9GfTxfvXhhf4CDJ1SkoDstGWisdsyxo0OgMCQKqXmqF
Q6I4B0xje8cAxGSw+MGE8n5hsRwSLiqbFNDNMSXnsryjVPGZxkbripVmrON8xAkP
GAOUEK1w4hPxoAdFzzOrbpLD9qlL5DzUj6pXy7NM1bJb1EbR6RMZcMr+Xv99e0KR
YyOdtwysX2kO2AKgJfC2EMDw+R4RaRE6/rumFSpO6lpTGqhFoEeeo8ahe1PYKBn8
aeIfX8mii97kWXBJDw4A29dY7uFcK5akNbu67H619qYvB6O/nH8L1jss9VCGF48H
ureigJ+JzhmqrWzx9Wv0T4XG1MrofFZKs+/lQh8/ENYmbz+2zdEI6beTpAdNSI6I
vzkIJWuCnAZyqOcJUYmPZ6Ll9hI/dCzfYIbioHQm5DvEWcOajsRPxv49PFY4yINw
2ZBs9U4W1NofeOc8NZkAj4hU7uD8izDPSx0JZbei+Ud18EEIcMILcAzC38WulZLv
zmh994qpWJftwoMTRtLw5wV6YFM7iGjoUfTidYLqJAKo2vFlPW+qsXslLiHnRbCk
YRSitOiBl4eJSfXO0KoO+rhyOkcGkrhT9LIxslBThKYiMh2rhQbW9Fa5xS7EW7jS
jdo4hWjumrIz7xlXKfO4jTfUBPpsKPB8zJhBsS1BBIBPhYse/BkgMRSOnUepGsUH
0a2CAIWoGDUWC2PNrxTc9WFWcloTriKzf06yAjbWtl6EWMuwnqrgRFW1vLeHmw+3
LlDZ/mU9DnllTqTUmrZMV7CTZ1HWSKFKxvboVzlwmrLUn1uBEJXARmUlBTSuTKEw
KR/U8NNS3G7Icob9ubgNXHue/VrKpOcDApRbpPkkzVhHTAyslr9DIHgqBadZtT7P
L387gKmNm9xSgVUsQUQh3OZuH7Sr7UouJNhoDHF3Z7fWjsHFb7TJtys9V+UEaDDc
Ux36+fDl3AIH6X9qZ08esLXH0A/qQHJBiqD8NSATJWQL+lIgNtP44we+FQP+yD/R
f+xRtbo2K6MxK+MDyjgZRqMBfXxfp25f93DPm/KlvcKtrYwLBeb4IaX/ubE8vCwe
+J7h3zIUBV3JtTo641fr+39LqRhtmTeELcWQVQbiLEzKkpFPXoJRYvrYYgrP76Jn
D66jpzp0icSsyJubU647h2JGH4AfwuZaHsK7+s+x33iX5GsM+KsJOY7ZE9OyU/KZ
efN8R5mQUefEoLBxtCCNZz8lRwBHjJ877wooUgWyJz42Gnw++2a46tbl36bck7SS
cHfA+HBtX1AIBpYXs8mWULEE4bQqOQrf/XfiecklwyoB0HNp9n+X2qYy3ILUuS/F
LXk+sXgq1S0AmzaSpfBTX53qe1Kwoq2DXiiXH0xt9xgUNSerV1LK54k/7Dpuc2uD
Iww7tBADR+lK0IvwRWMIrNcL/KMzcp5Ko0dU6yahGZ7BAJdK51H+ZcXxsl6RnYvR
aE5WQgNW6v++2fIwS0q2paaKkTYDuNq3OU/toyDbHQ/DriXZO1Uy7Wg9M6bysstf
mxGfWzp65oXmQcmaZXkf27SJ/tTEL6yVtluy6SVDSJeAXy+Wc6+zf6dEQRAbpRRB
esr8JyJbCNbpi264SxLuGaTVd+DFCyxOhSZMdW6BUpDnhHAyz+iBWbQUyaSIxSW5
ZKyR9Ic475qs4lv0ebONeNKSTu3WVQV49QIleWdO99Ff/EQoNWeDw/GuURXOcAEc
uSy524mG/K3SOZRKwv3YI40PHd1wUpb//mOGNHCCfD45lx4v/fjmUDen5cgCuIxD
xQVE47jZR+kJfquMgbgq+RSOcVfg7jdrnJm6FMs5/MuVWzW2Vr/hzlCu4BDzbRYs
Xz5nsLmYagF8fLB7KO1xsBEWf4v4z8eIQwxbrDc59ETStW+mFvZ6SwkwPsrxnGFz
asSeHM6cTGhohICJkRxrp/DPNvLiTNeJ96hR+DcF5v0OjnSaNjnrw6YdY1hn2V1f
jfMPquxs0oCQyNTgn7IVoJCV2FAK8on3l3ZL1IPprdtCmwQCeDgRHnuuKknMyC8r
xmoiM1diDe8Va06RgMCt7QiQT//PaS7hjeHJtZyMuYmHu5XN/TP6+KnrKMFpiztP
G6V2PTAvlxETclGpo7OJRhGa0zXIQr/vc7ZCZMvk63bgfuzYggXz6OfBSNRM6Zp6
hoZtDSWILTAFpMzqDj4tDAa2Ar5epNzBScXTLCC9c5iT55KwNaYgMdZOmqYKp6vj
3254rKofkPolDMY7zGjf+n9q7NE8XCWf/1yFZt+NsZVJrHLHvXSyhCNDW+3CAbKz
khpA6fmP+/9BLqN4KDYsI6yPGJ1NUCZgnAklpvVB+bdrLTPOItWPcfD/VadP43IM
Nukt4l+el8werXxutHhEdmzY+rt4T2ZWcBJA0gIp3UnDaEOVmAk9EwCMALvE7VQs
X7UlhZIaVZNRGzV7gbO7esocLYMWBe9em7K/KlJj0QfiEHk3+dsrBaIjvzG+NvtP
n6no8Q7+DsPTp6Cs0hV8yjvzmvYoguoagNHvpv0N+yQHInHCNI6Nx5hof5voAQMn
7IKxcbHL9fLrnPG8FwgYyhNB3IZiBzDi6k6moMNOyiWb4r/pJ5cABVIYSqm+yOdZ
MVqHPx1WdguI6SHnLNgDktJnxMDWYy1neOELYWquiuWNILJw8EltbW9R+ahhGFCZ
Mm5MFpCngrsl0jbMX8YkwHBPZjUc4pnjXQdDqVjESH937nhEBqPTA3TcrKCng6ZE
yiq7DLeCHHwiF14J91EXB6AuH86s5QWtpmploq3dQ+wC8fHIx3BpLq1jBffRdNN9
fpnEMdqNS8ULyIl+fVQpi/BUhkdTOxqoQ8NJopak86WBCgdy2W5qsX7ceqGWdjGa
ApTAfiyboX8kTFd5cFcrkqsK18m2YtVVurp1roT+N0NT7VBPDT0SoREgQQy9gyHr
QWFAkuRpC524Q7uyOp1RAgOHdYxxadfB1NNGeZdjzjLeQCA9+obGNpObe+RPIodF
4vM1QVl/EC21d52AwRkGO8PS6wX/F3eY1oFkonGJnGTCrNs3ej+lsTPKCc32qI/d
q1YG0H/QoA0zDp75iaKdCCj6fFAcSV5UiG/eaaVFTFw/JriKt4nX1PqxzLI8BDZH
HmhgIQHhpf5Ovg9ua/P3zMYQ6XEo76D9FdwXRix3vc/EEeSn/iW7Suix2M111bZM
vKKXirHnC6W4aCMPDpA+5pFvXjszANt5yPNqI7JXzJqhHqQeovg7BRBgftqX3EiU
nkvZiYfIFEopEhP3mtZshbeI4AGCMyTO4QlXOa1WD8ZtrIUsUiTvLTejeEw7YsNf
i9AXk3WLo/yIUaQxd1Tu+kd06ybknBpffdoUwhKcXqLWkGsJtuQP9sxDxFSfzOUR
cMhwOwCg/TlzYdWsp+rnt0iHSvzxMJPQA2/3lJGqdj2TavzTbRgyJI6hI6LjKHdg
ONtlzQ0MP+rUoHGmbvD1+c4Z6wtRlbvLECiiBpTn49sMdvWHMJ/J3xLH4h980OyZ
n7gv36zCXh4TtYPde/cWAL93fTBhe5IHMZAXGu4PmikUhXBZDGZCecm7G8e4Hq+V
RtO/ugfBozK1tSVzLM7qRaDdqCBYU+haKHVGudzwGmKDE7ACxxAeme6nPb5U3SV7
HRBL/oaX8P7zUJsW2KEw7JR9+FZWiUmSR2JDyA9Qy3hM9sQ/bQHNLrFi6i0wHJrI
Kww03d7rAmQaiwzXlcI6W2RPDd0EAQJdmViYkjNu7JjeBtvKoLMUnFJHjNHvB+gy
h6vFbcIESwhRgUlYOlm8WSuZ4O1U9phhzyKbMNaXDSsB00JlDXquoHZF9BUgAAG2
v1/mBkc2ETehnLrHIwMOnuVLx4G2DqXcv1rNnGUraIw13hAN2f9bdTnlsuxXQbQ4
pUHObezjfA4j0OwV0+ypPcCNgQM+yqrs5o0gEY4zcCYR3Qeo4eE7dFo8UHbDqk5Y
D+1JhOZLeOpOSPQ78EvXCIxu7X4tZmSMe3cVYw+hiooEQ7VbEnvE1N1he1zKgUVD
0I0GYOXOo/dm/7hxwBwuj8se7+fchtMTR3sB80aJCCQRjxTKXgvCEE/9zH3x6bnA
Ss0rQ+inH2Ag+h6g0CIzE0RtUnnMrCsQCOQieTSpCYW0k77zwek70MoB4Sblxxze
Y0Xif3d/Emwf1vkD8SfXDkTb/ML0mjueBLDzxIGEkOy25jbtIHbgg6Lr6ZLpuAIw
s/Ul4Hk6YdGjhXmwHC+WUKkK0SU5DOTqM6aQU6KNRzNR95bDQmRVczu2M4w02pNm
djyx2kbJ/A3FULDMGHFwRuhp4LMHp0tkkwqDs8NnlFfDYfTYUnHwZjXA6+5GU9do
8aTxMdhGCguGUu5qcqUrkwgiqYDxnBl/PKjtJrH0kbrHGHsRS5B2A3HZq7wyW5ZL
x/4Tzw7+Q8xhI7XKpz5MJbTMh/EvhrBSidyTQMB6HPvl/COOOvkOpvcL+7eXWyDE
OMnBjFTiAL/Dc311Gc0ywF1/sDryyAheVMCLZGn4yVrf4SVhUmpgCWwSx6uCFQvU
Tl/Lq2BGrrWyR+kDablLCiBoO3RiYbBMfWb+iIQvCzry8ljgbpveLj2IRNa7z23v
WBu2GpoGrC1mwXoU0qXBBUKXtOpucum5whnriFN3zOU6kEq96rF6QkfNM9uV3Cn8
FBfmc2z853QIRts9ifh54mHyi7LyrHNGIjFUjGsKUW5x6I3S89h2FlRLycQj+6nA
9m14Qq31l+wsm75rDCFKYngPQHkU1XDwmdukVjq7jNQjDByc3ZX67pJFGN6PTJCZ
7X01Iu/3NR4xtwfeZe709c8VcC+iTgH2QK7VjTEINowcsN3ZBVR1EyXFbRmcAR8c
arFWnhf6M8SA9JfGvMAK7wewTi0aF7NWS+c29zn9jIvoKgl4sQ9nJIRf5dKzCELy
NYFutN1RlSvPcEWw6xKR4WZGBpUPwl+xSbmNZvSes0cvL8zRoYWCFOKbWyN8z9Fl
caOEXO5IHBlBva5C2JY7PS3zDyasjgXo4oVUIjn76gDSran0ARAvdkiC8eyOu2s9
D4NyJ9wVcO499lXDPC+SPwGw/kDvdZ42jZJ9jMBs7+QfPu4k8atU+D0F3bVBCgpW
w5iRsQQyY6X/4qkQt/RqTX6Q2fRKUhpI40wVm/bW2i0LZM4hFgenXxEdB94rwWti
lFQZmPUT01j3boSywUCIn0yU4+nNJUKubVSeRCFQZMMuhY8ZYjI7TTAoTi9AywRZ
B51hGObthkq+9NaHfB4jEzk2O9q4FGJZ8MOPthtgSyDDeAT9ls6yUz/yb/81nKTH
ZbX90KDw+PDJN4ipdH5UM7V/JP2X0UGq/wDqWN7Drxm+k+NKAfQDO1vGH9WhZHDC
CbX2Qz4TaAAnPbXmmqauvZs5dWYTsWwTgwqK2RefnwP1CFonuRhLCS1PqBpMXCY2
MCcn6JdDmcHnFveCezBuy0NJ2s8rFeq9vNp8hudFj6cMR5eykl0lHIBbwMPXhITM
vxFvA5nrjMzUqM4tcp5U8o22P4/W8XXR7LKGb9qXbxwGygOp9NyxgDN73DdaGtC2
u/c7pzodQVF4GCQHAoKqKA1wG8z7YO99OmFgVAbyeQ40KFnt/J3tZ1G9890d+IZc
TAkcb9KebQyEsicP3kL8RwlSKQvxMe5RwXDqV2vrtyUBzvS7EoHnMJZmpEMYj+Um
qlNFTPLX/VToKL3XtsSX/DRBl3L/Jh1X5ICVRE394Qx7ELWRa1InbvtHC03BLcA2
WNvKMarnvUKLJSV2ds3XZ3svQmB4bhWQ72XayNrWJJEczzNlQcn507wyii8VB/vY
th1DxPBaR1YQo1lG/X+V3zC/NojZcjfPe5TpkF8DsPKoPMOS0RyQHUloATwChui8
/RTHUyAc7dl6AsiLVsxSHduovj6GXmhsJadQEwdAOCFa7LiTJvPxTUedj4gswHJm
yele/YGkEe2etR6A1/CzDmVv5voNYdjcCS9B7USfje19+YpfJhk13qqHln7TGO/L
EENE4wVndQL5RWUHVFjFscpqxvtw30ovndCoDVONuxbaeMGHaPQ9pIoX8gaPQ0An
Mb0MgBZevbnFmuMAXX4IiwBjdDLzqJCUA1itqPS2pbE6+dzpP0s5bmyZxNNpkE4e
1cy/hC69yEyoDCLIZMHS20fCt5e/AGfZ+PUhRlBuzROfUEvSSfMpl0/Y/Sn/mttn
zL3hoWTjjmcdB+L1ftQEKsZ9J7mZm0SmP8sBphGuItDGg/jOIOukJKIH9SEwc887
cGw/3QQVT96l0PC98kybil1mldAHBnq3cPoJ+/jT+pIHiNu7dzIlFzRtflLSN/i5
CFbjxMDaqiYtiX5xvukRwaRlbA+Tc3mmHkJQY/aEkGP0qbJo4AwAF86/gHOS1mRX
bfbEkZcj6rALFC9hKKWHHrHJCdBSuXXhK/txF8lM/jY84zZqzymrGFUY4IQZzRva
7TGUydazve3BUqHObwPVx2oLklDbYtyzV7m8gS9GNAov+WewLLR4+aliR17kLL/l
Q5iRe+tnpyrPOuu0UxTUYvuqX4OYxQQFfSPP3tWRlo9g5Y8SjLTUbmbhiRncIvde
zw1uaY06LpZU4/TSTCQ3Fvfi4ApB8CkYMigTvQ+qGfawJyeaHLmEBnt6+Z9v65Zb
e+UqwT9TTj9rMYUIgcKOxGUOm6v8h0m1aG/giVFRr5fKnFWfczd+XZY5tc2n9fdX
aVyPmeOJ1dxpKdj84NksUgjo0t8rKXkrxxRYUl3HbAw74zbb+I9dWTJBw38E/z38
MP4N8T+rn6XRP7pi88wDiTjk7IKT4uMSrndnuR7Fm47HIXHbXCdtwc+Ws7Ey0GyQ
euSuJs68ef6ZM09BiT+UBkYiKhhn7hP+YitliEKJFn1QJ1HwAxY9RRlw6p1EBGVt
C6rEUp94qbBSprWMVXWiAM6fL3AYBbUd+r2FQeKFKk3wabIVroJ/6whI5dymq/yz
rkTDgyXjsi4ZeRPvIDOAgJAzaptN9XAOEUrTx7SJWk0ThhSLUaMSnAAR9/O49qIw
plUTeFueKCKlS3X2wWCernVSBiW/H5VNdhEXnK6yJGiaALpT75V2UHtd5fZVgo22
Qpzqu+nh7sErFj7JS8V6kzzgo9jyAkTySlBXEWFcdOn9Ujn2hS1X3Y0+Kk2PBu0Q
Vtdas4AQOX3owDL0RvoikdpHL8ANLQSTmXnDm7ib06OfcpvQEkNbLS7TthK2p8oA
IjU7DnJj9nCDHPwS80mygN0U7NMifzPyO9QRAICFy9jnKZQ+CwD/ZNMD0McAQH8y
vCTOo95Vw1VIW+jSoIAEn9wzyceFcdEkiMTDd3prse8dkyNc6WGc/U/7HnXbwEQ5
SbEiUEBXDpN3JxuG9/E19Sx/a+s9z/B4nzNf/+vCfbPvaIfr8Olx9thspPh/BnTj
n+LCxNhVF3XuZMIwCeNBt77BLDwhxCaojfaqI95dKmA1hgIqwLGzA/5To4laJ2eq
fQYjC9Wyg6q3PIV5WdnZ7KexfFF58eoQ1VcUiyo35o85HCxCzypxBtz76T+NH8x9
rW1p8NOf5+ZgW2lKL3On2RRc8Hh2P1Clp6EngR2IL5J7cJXTmn2JN8UsptQJQV4a
iEMFWl9QT7eQB+K3C7SA3My5cjQpu2jhupabLIKmcEYFJ5edZTNOiJ8LHetixV1E
40YgaSFPBpipa6C1+CF1lVd4e3nz2KGkpmThimn0491+swZ4QpmufL1VWr3/0bt5
ONPFIdQmlAJHx3w8eKsjzFiQxd0A14u3M0wX8UnNZaAoC18/pDk/pxby14wyn7Ys
EO5LvDBJYZhUqwOZvu3kbs1DAtujE1wapQFBbT83s8ywxb3E+QU/phAQoTf1GXDQ
LzMokbeBwvoyMOJlxhYPNkh/YLpPiT87yAk7uH/0lehnSi0/OmG3iIulWdh32SWK
THbFabKbP4LXWgb12bGWLeqzUBNHR5HqtvBhgX9dCA5nyPHnjFEeaLmvjQiEhOo+
S/wu8l8oBK97wRfPOzfz4+ONUKCikFOb+JzPG6pn04f656vqGoUmsg4g++KG6xBr
pASfRjiTd4wKWoTG0TEZEqqm2zicBo1rch2NPNdgBuuGnRrm84f6WwrEKRMkdavi
ZF5m+SCcQXzCPNeSCkCBzYswlUL1lsyTE0sI/KTVk9FG1koQjwxXtPCwy5ySI28J
Bpa4YeCeUdqF46T8qcMwDjByJZ9TlJkYPS1sEklE8dLNw/PbqPxabFqd1mP47YZK
mC4+jcaWR6puhIQbLK8ltEpx47toME0bYOfU8p8HkS3w5rBH6w7dh7B8A8QGRK2n
2zPI1OCLEJSj0NQqRLBFR5DXEFQ2SQiQUKsw+AbbR8aSErJ3tzH/2e927R5exjoJ
OSjGfnUGjEhBVuZ4lXlURvhzOsRLEM6yjYajhwUquIdpaDALBkD2rN7SNHgnIRJQ
Y1uzMRlHE4BNJrZ8hnxgFA+3v9z2CAVP53ERFuBhzZE4gvmXW3wyD9N4Z+yxJj1H
L+sBdxFVKNeL4WGF5UFyyctA3omc12veGszEn44+kJZi4fqv7lsBJyj28/mL1vPX
z4M5HEywz2lpGGv14HCmBKSQJHRczskRA4RFw9Dvh8h5rfTO7HJOVpoRLzHz59ix
Uw5t4It1KTHtPyuyDh0fcScdv6yO2yG7vax7dGjcm7kO67tTIeThp94IhjqkAiha
yOz58NrzsXxkfWaP9dHgNttkkM1amMIsSbv0pUmU5eOBisd0K0kIgWiQDSi84cNC
01RBE+uX/SVf5PXWFc8RrXnSuK9GF7l+NbW5QNkNvM241UbluwJQ7SIvJ1djA74p
ustdrrFFrjjUucEljZcgCzM9SDPs71ZUL4uh6bG/JwU9KZ3ZsV06dlV4Hj/UM6bk
PlQ3cE8nEDGJFmm4Stb7MOCK6T2NVHRpo733XDbx9hFlnckRI3ptC+iJx98Vh8RU
vaU68Q+GSfO331Ia+H8bCRy8+UrCVAedQMk8Mv7C9rqhROQ7ZRXfFSiVLdEcPJbQ
QPk6o39OqlnHrX2zgT62Etx4pJI3eCDsovSxAaSTk9e7bzYarB+42MMZKHGhKOSc
Udty6yJrp6rvkpcmIqjJPOgh0/2qxXEKtW82Q9jKI65zOY8DcYJ3HKEbLynDFRpy
8Z9dLnBk8V9/fRmFXOz0uTii93GCha3ffPiH+Civx/dYBtzg/W2t1latxXYdpLr3
3kw5Pz0TbP01b8DO4+uh5DZhwgucQ6JJliw9fDJYxly9y24A7L7Rw7pmdbP6Cjwx
lYLfOtFT52O5aLa+4IVLjKcZivrlZIWH+s+pdC2xbKGfE2GH+QC+sQrMPZqJY5jd
aRYGwxUqcMe64VqVP2A6uq8YO4Ucfl2PtJO7nBOJsf/bsXUEAuR3xXg3+iizl55k
pe0dBXMAXdPRxMSLpUctOxEtqD0Xe6U7NjX49kmRuHhy3x4y23maBvpxF6mM6Ac7
Z3gAKSfJswvKZypEiclXjp+7HZckduy9HF0Vemgd48491yjuY2d8x+FVVZxm0MJn
U7C2YjIHuDYutSdpbnwoDpNPdTZzjERfY6k6Nuj3dMNfaXfVnP58l8xKEcV//6LG
IgnmvQJ4VLf9fL19fvt81UR3RXqX+bLmLVnvN8Zqxuh7kQPciC9NAVLTbxZNdqHC
vNWe83n85Edad4tF1J1q91qrrbu1Q50QXuaxs4+2dJr72ZsjdaGz0ZyFs1Jutb5k
ggu4WRlI0DXXJ7aQPh6ptM/j25RMExnNBoN5CzqSCZlOmOeU7W0N6zb8jE/CdTc9
M5wMp19g4MJF/eBqFiVY0GaCFJqYOJBulIzDNvJFpZzGIMmHbpFPWwMxSXQ5Rf59
reWJcprr4498q+mZeCHHQjqjwa4QTiAzBRDb9S3QfFJahiQuzdmgz6QwQC0f44BN
Ig1efXUNXpywz92vscS5wW/9/tUzjGK+Zya/cygM78pOcYfifqjqxCtJxYAnV/Si
Rj0m7Yw+WANkXKkAvHZDwU/1jLEezHgs1yClU9w0ttKSCKwhlnVnkRp8f3AgBxSp
XDYcft4EZLVmPVNS0FnnyS9KAPPRa6hXOxSdOTsvfTWHqJr61mUNl0hUHCy3PAx8
sN+5LRbwdnexe6rQIbcDVTH/paj7LYwTIb67E/pykcbXbsb9X/AdEdd3eGS5+dIW
lyzscXznGMdTQ+h4b+MssGcOwKAD2ESas5q+ZGwv0i2P7Yv/JKoWPKn1D9Z3+R1L
QKQeb75G9YrvrWQqvt59bFCRB3gr3xQJ7D8uOyQzUqCVZK/71nH0lHw8aLFv0AsD
jaqs+iTiEFIzv7ex/WxrX/g28IOiN0movtQ7SAjkEFB8ak72qjpVeBQCHCT4ln4n
KmlIhnDgNCzoBmNsFgEX26uLdHCEpCgSzHkYYfeBDQbuDiMUc2erKCWgUZzgQbdu
zS4KFX95s+Im+eVb5jB665oyhif6hAOWFr2RUa9fN4uQCJFf8Ocxwyjb48FjL2Qe
dZZHWhc9AGOlHNSfQs69np7nrb5YewAOl8o6fITyB2gKK9jdHdwuoNdIHXpO1BAJ
ZijECrQeibsHyoNjRGG3xhj/2mzMeW6MypWj3r8mjJP9ROwgDl2bsmhMstr1/tEe
P+WDNFYIRjClMzRU01YT/r4kRQKe6yspHI++CBXvSvl51TxPuzuwQDoK8/IrrKEH
yEVpBsWAW24rzJF55C6BrRKv70IbV4LFpgqg7c50I/vKJIpiOQHqc6CMvS3GUFBC
x7Zhx0FTv1QoW+FqifUHqoBEvX3uCmj2YNy1tabX82NdLfhfN0aQhQTaRcj+OOF+
loMFP3PHbyudNybbGlqV7xXdOageV5QsnLJGEhNU9ugsNq3ZULpR32zY7E6x6jUn
V/nzoBpViMOuChzQyUrhhWPHhN+neb7E3/1a5OxmYoTbyxXFZTV7UcmIUAkyHKt/
qAMSUnOlwnHZ5RhjQ1QtkJ8Ya/SNOhg8KVn63cvRvr0QQI37ongqMs3IdIIVn7Qr
rfGqIGsHVd7+YKVxhBaHZEbdjWBKG8PZPVfKJQ6ERPFuECB86hvEC5C//Dy7FlgY
Oyw7mI8ib7tCKT59RZZQZCIO6o4bb2CHVknAiG0DqCKyLm0kYYyxkcpc0WtA+laz
VdWGc6vRtYHVjEwuHDUf2N2Qg8iGc4C7oa1McnzD5lB8ujggd/aocVbyQ+wKCUBD
Id99XClAdA+FOwhebehzWVEVbw2B3rqujz7uJ+4hrDYfxdJNsqoBmX/zp6EGtcKf
UI6E9RXH3RDd5QMjdLEf/kNHp8bg98VZ4QDrPIVFbwKQDyrsl93ASeYYai5u8I1T
EljGrRukR/IqWtsWIEVeLHSuLPWqLbL/0IIPHpmYlBOO5KHI6cox9HGH6NYScbwM
JMel9NMLficDR5K3wcXpcH+vZdQAPVD9aP2SzOIT6h5kkeMC+ImKqinpAeYZhfge
kckAa1MwQFjG1B8buy1cMgbTCvT+Ciwu97ydxxvI0ICpFJrvRnajMamS5RIrfKW/
x0ro2kQYox5bhSuY6mXHWKCeD8iuknW6TwFH0lrRt4jDMeYxIx/aVmjjP2fJ2ttJ
lgmfbESLEZXEVie+o4s7Qvc91ujaKQ/wzUxdkAIfS+krrPJ/8/k76jzXEgAbQ2A6
sdr9ajcPnaTeYK3Za4ZBfsZclCfwQ1Sx8EOAGq2bDfetPjuUgwD/7IH7C6fX6w3p
yInYdLox+mivtgB8nJNyYzPyg9atXS+CcDkN0VFvNxwhi1PAhrCw+JUOZ+Il4wzq
hjraAvHje6ngPjnOKEebwseWYdDxiCPEJkFVjdhTKWhgEKjE8VT071V5j0L5mYF8
DDL4FftcSmapPOESfD5vUTxDDk6HL3J3GE8SLY2hBOTiV1Hu0X++olUsrd2Ki6l1
37XYtwQEDsqtSiyJtNZAiIzioQ7lIhSCX3Yd5MAUMsYeJZj/yaGK3Ark1g1TdD8P
SC97EWUaprc4KrSoqLE0/xXO5j9nR1IxKlijpGI7GTuuZQu/yvHh3MXqRIogUpCd
FlP3YPzUTum9s03p8ASkKXyICTVZ+xP4W6BNcthzFKSzmmFAVfunLvLA3UShwwP/
kqLzhR3mXcRpeTCmq9Fisn8IcUz8seW9xIbMHhhmlHH1JuvQrKFPP87Mf1QZfBKI
MOyO58mcTP5J8NU7Pl+UKlWF8NAxhI3N+WSsVcyjOndxGuD/dE44pjGN/FHFTmZa
a0cO0pCGBzPpYC5rT5iWZV1NdFCglRwLjAUgLHV1+cYRqZxcc0DhHiF1gqYSFO+g
/6h/A6f+qVLshpPZ0AkZPDqod58KqkmSgivF3cwapsEtzScro6/cE9QTj7rIN6lB
rfBq+R5k+2VRC8t0Amk3jqTxR2JzzYkBBiZ4YCUCQ/QWqEwNZhRJCdBJWBuCXRts
4Ap7/dJXZ/okRpR5WrLl1DhnPt81Syr61g8abdTo/egLUnHrEdYlEeDZfkzEMAeA
rmeVf8VIUwLN5PcnG+On+j1I6aDcK9s6RKhu7sWkXNnSvXysXrNQCtuA5Q3jJIyH
S4lMbtVRt++LjDr6GIojbfuqjl1wkqoADPlgvhbxfjKBKyFOUnJOaPrGIkdbZqnd
g8cree10y4K3GuDTUn4sPPofm1fQ9lRaLlnbmyKcE2PHea5pYJbfcBdz/a2ybccL
xNkwCwT1WCmsUs8yod6AZudjaNZMKfaUSRE9gm8bGqmaQGAHqz4P9am9odniqZgF
UCqTR7RDkiY4EZHPWNA15jViMtF3LF2MjtzRnIBU7p1UXomj8Z2dUGyMBbISuNAx
16vj3zC99pGJWIggm6CEZpJOnLRgj9u89xmPuFd3okfn49t1iBCQ1ctv/On4l9fa
PDd2zsOvzP8Vt9cFzr90WyNbjggCdvoFxiqoVCaa37rKM33h+HltmzhICW9y/Yly
sIV24m3Js8NtzuHvql6ls6y8swvZk5+JEPEPUPbQe7Twf8ttO1hWjdWOrHRc+Bul
35ERc+YNI8zhmKOBz3ONZyHnjOB1h0mL+byien3gWcsFKPwKueUlxnbSSvD20yPm
TH4n8SFXYMSe3tHp5Kc+1QOaRWsDlkRhRzEebyYU0/A1f/hXor5pajm73kcpu7Am
HFdwJ1E0gMc7tVqeBpOcFHhh/phlTBj8n2f2Krn80bDjOOc2ppC+1F6uaKuEHwkF
ursHlbPFjqFMNOVyDmeqHwo7QdvybdZz3PBEWvK0WWsSnd+kU9e/jKuisAvUZQYt
u+7aPUADdZ1Jf5zJ3v8h8jTvTmQ+gR9UJF2TZBrW71g32U2slziw8aWWWKxy6/A3
Vf2RHc6HK8UskwZRCL+1/THqvSbJ4Znxlhy6CHjH7z0SKvVFLcJHKDmrjwACvyCp
r5CFWFi7XjwwSD82eRxZWKLcA2CXzrGidnODma7jNYDjptO7qCLcMN4Si4bi1GCA
QmgTm76y6WaecRDZ+IlKxV9V6CP1YvH4Q4Hr8HTuiNSYnuz7JXWzM/sugM1z30Gk
7oBSMWlONMOJCHKrqzoOoUJDjJYWQMAFiLrP9l6peANS2GjNz1uSl19YJQzEKKlI
BPLxR3CypNt6sodUz+imvCQrTXehdoNnPDbKLQiptIUCYeguosa2edmdmhR38xaj
/9JNAf9jOpR/zSlCzhj4ONlBW2At7BgZ5DLLBGa1mWUqSLAkb1ltvUHSUZEyTlNd
CpVAUDp0575lyGzCcbH9gQBduJwJ4ZM7TEbi1iAnd5uHBnebEvuqA5rUjhDY3Pkl
lI2SOLn1g2WN98q24C340NuZkJrUmyhpPmBJrEabatY/vpOpir0+flYKg/VzDtOh
KxkZSXlBg8QPMqjvjeOThKcj3WoZKITQqULkjtfH4MQr/buN63wgY+NDiiZyxWgH
2fmkmtkRrDCoGcQhcZhM1ZYpGY6dU8KSuySRXI5+vDey+R4jEEArNvFUjhmC9E5s
tdFrIKHDgHhxXlazOyYANWTuUtZRw3V3r2pNCwPwNAf9lNbhI4MNyODarPlB79Fp
SHA7bqhmH/Htb/nQUsnv+ghIwVQeuxW1rDy37IJQhjutOsw3e0uioX8Wq8yHxMgh
ptoN86KhhVeHvluGwmCrvDScJGw2EkXLB5SSAEbserXxCtEGJw+I0FZvlPceJIeq
5gnSpt0ek8qKXjtUE80kxj8A9MkJTInLXWyoQgTFWUL/BTddjiosOIJm6ZxcPh6m
P+7e983W4BdTwSTXYSJtSuILiDcYLwX8G9xOGKPEOSDeDr9UaC1DTtvKhyCuyEhI
Yk7yJk5m/8aTm8v6Hq53B6/GMOegvMzjy6FM1PdbLGHr/kY59EugJB3aTRvria++
UbyC2WdYcfPKDv6ZCXTXI61yWA5Vc1R0mkL5uQHi0AVBZrARo6PUmo3p6iBXTxRv
MR+KbSJXkjaAZquaoAiTAaIrQoGFVZplFx4AkegDSjVdgnD3ZTdaiwn1llfaqyb7
D7DBziZ5qSpFvOYb7sAS6KUayPKLbCxXrPY4P3MJb/umTT+L39ts4GbpbcwsjmYn
C/38rgVT8lWxBKPXU0oG8oL2hziz6cjprj7FPRNZ7JdwTHv5lCgfac3Jvy90pPRO
ownY76t/9jxBhMW08dkt70NJyrYdaCNTI41kMdJ3Ku9qtTlePNp5901x2JpiM93x
/+GgWmQNJfrBEWdhG7VppQf9HVg3m0MQTws8Gv7D3CGmt1e05NUd3HYPzHOdBrUU
BU/1YUbyM27Sjt1sdSKmKrukkTISAn5aiUkvEW82/FNDzfPhF9y9ykF13nMCLRbs
eiIxhstnPSBIbIFSSM4BcMUlVUFjTbrVccYHCzTjB15q5pWovtI+rFisyq4b2oM9
FqHUlbiS3XVRM33vCHjxeeEKQPw9rSWsxvjPTuCsfxD5rMIoutrR0eu7D7xYf+cB
A1SghnJCCx+bLIj3LEuNQB0tpX81hR8cAZqa8LyA4I89AXHRfxN4zPq0ePKFNa5n
cssjNIZ+IyJIWc3g9qisGqvUtj5upB/b0K83HsUqwPdybA5dynQ+Wc2FMDhIVx2t
KNLut6AyxYOEHhIqWYoWNwOhvGDb+2Ejg+ovymMsuowbISvi2EeA7ZhCgzjcQXZq
2Zf6+ggTKckdX9hjOcEKlSolDf2gwPisAr62xnHMEKxVSxiLvm+NjLK+4jGQ+hgN
PVBOmkQmTvOiGr9jhc2xv5CRIKbR7xElgmcJp1uFtU2d6O7F+S0LlmzsqVx4lDlu
HPT0AB4ymYx/4FCasXBFCguXUWbmmKTFpw8AXxf5johqJahAmJ4Svjs7ED+7+OQU
HEUKX9FDS9NvWMFPlLfYpttzBp5ooW1wnLXlJdDTFgyblF0jnr+Mjo1UzpnQZ1KN
/paUzPa2cqYpZfdX40p2CnruDCG0yb7+S17FMrQfak6v03G5+9V3BY4WpUqAXwOX
B4WOWERbRO0uHrbk6KBBWp+2TkRccbwSBRAEWjaDiinkVK0EikVd8ZJS/Z3Zr8Np
Iof8SJD8ugHGU6c3A49aw7E4eZBjeBU+o8aCMnZ0kAhFrTwaDfnJ7eBFqTo/EY3l
uTed5IhnBITlEEwQrGkZq24X2d86C7bEhdDGh2IEIIsruzlpuDaLSTUny+7WCaRM
3PXBXsBAkyGkBJ8DkI1XuFIUoTUn0Qn3hAjIdo3QVhwjMOzmQtjfsh2Hxembh13f
EqWKzlw5EOio3JrhQFsTB+OKHAq7rFcyK/RyhpIXc9UoPxq4Cn0IkiC+7S2Dur4o
05comD9VtxEjxmPBCsOcfEf/a/19kxeUA/CKFR+ItTuxq+Y03AFmDIuMq2bXiO6+
WdMSEXsi+bUP9tQ5SummXtnFmv/hKsGIDCYlyn0yskmjsu/1zHlw3oczQQJLjdb7
Q8cedY4bOXtpfWsUyngNTyQcNfha1JHCdwvr2ov0pv9jziMs0vd2yUP4cA3pN+0V
lV711FTB93B2wist4toPBda0hvOMof/toTdSTEW2zDRCDJDg21YvHWQkXngUMPrZ
yB8b6H4BvumDbyUaQc1SzmOg6CBAcSker7uXVgxLI4gGzEW2fWwTjwlmzkm/MHOq
SfbqdBD4T1qIi3vRhHEAIcHBjwb9Ft+8MRfw0k3BAIGb+e9h/qm/AtWtGXKXHPqc
r7Rmwt8EwsTyAWbtS8mukckHBY61ZVYo32vLzFdEY5woEtz23fSEfwAKXWew3cNV
j4Kam+Oa8ChZFYkHZBzK8vSmKvYHGmg//1NB+NQ9CPMdvpYskSsSHi2gSpYsAVgQ
V7yDlA92xhCIcVZ274Yw+wHZBCDhouM5aHIShJRIqvtj3plq+gsQoHhS6YqgVQCI
KA0xZ8YFLNbV7OF7pub3RQH07PEniGeh6Q0IV3508F0SiSJYx+PK7CotVEEuT6BD
8AgC7vstxMbPYCLsl5vxO6yWSa2o9F/Mui+A4eW3SBCvPnkpr9d5B60y+tZG8sTD
PLjxxPwCDOfqa2MdZ2NkFpu2D7MTEAPN2HeD+azi8d+0YYjUgcdbN3kJ+flJ5d7f
coPJtvFmc9yt7HRpQYT40Ef81GGGrG9r+TF45PoK8uVqfE7QJtbym9WGmRs9s+nf
GLlbs8/ITjVE0t07qTIlDg64UU7HDRH0miuqrhRcl3toxKP8zPMBocsXWFTbPS3Q
XhnoByumcpyCMv2ODmQwxLg6WT15zEU3/oo/5c0lZhNyWRCJ6H7o4ewcm+opAfz/
574lMg5fIEHe2wsoaDB86NbqQtv0cEShf+TxO0oI5IJLRPn6pXqRoljnJfHxFrxI
02fyVwNfAlBVmQBaigdxl0RGKrae0ocS2ZH9CBdg0bX5+YgdW9pdgOb2GuUXnNzf
mbrT2ChRaghrjnK0P5l81bABove8Sjg9/1L6x2MRAKK+ylI4bAMahqeXXjKbXWdn
EbPVS5sD15I2N6E9WVwNA6KqGxcQ2cbQq5K22WZsdHrB1eR33JM5yljg7ksV9Suw
9GLdDOP7Ju7DPL9iKEiH8xJ8FjxCdtANTe9MCYA/D+uzPcFMb2tzo5Fx0ZRo0/81
YvPHsjvEL6mgmhMNRIS1BoPTn90M3O8mIr0/7g5/EKWUqUNwsUCjjeTFilWYE97N
jG1CWfBvmybWPuXCz4pCDreMXnvsZDX8462Ky47qaZVV+xRFkencPBunSiQIPhQk
Y29HNsJniaAWWT6IlkQr/i5jdxgzMfuchCieSUBLtgtt4kcdzL5dQ+uvUtWhRCh9
dMLfqTdG1HlDlncDuN9nNijdc3N+BJVyCBakKvx+suAKUYQRGQgxQrllZIw/+CZN
cr140H97UutjFtyUWiKDLmG6f3zyKkgzQYBtIA4IvRCBNQCby8kGR1YPRzLXF7XP
1XQNUQtFnGkfhGf5yCjRWqdIhSxpAx9MqY2Mkfifr6Jj1GBtFpxWTWX9po0TwmzN
NRdi5pyCpV/LcLKuR/xJtxJXt4HY65B+xwi0j6MIvgQY4aS1HmRCPQB2kNNI/JjW
145o6h2LtpBvNB99xbWTQnjbq9xZJhOmy4Z29lg6TOd7k26ck84tK/0QwpAv7KKn
+taA6EOxyOJp9ziKEvccAW3hBQsxiZDQl+1iCNCNe4Zlx1s8Wax2+rTlfjktjMo5
fI3JyyEOVy5wHw7yXprN/jHBZdlSd4IVCKZthZZcdIOsD6HHhYIyX/39RFJl2vAo
w5k0wHbFYNW4DWvuIcy0CRqIw0SC19Ytw1yPbEIFOUABtjpmMPyVgg40b1k20KxK
nEPdgTsmnDeEfhoIoA3wIhOAFujApTTk4RnVRv1yAKnlG/WcnHLya7kXsQ1S+7yA
Lqs35ukE7NtQUakhaCwIbaiE+CCZxHMmaXzTtXny4Vw2LY6eCagv9eFzomxO1DrK
xYIYrWk++dGoHpJayJ83i/Ihc0JX7e7ysHk3YYSlmZXrn7nYLZyBn4BKbIUjtH/L
EZv3WEp3jH/8hBIV14C/OcnGv3dKBzFaDJyS50aI6s07OWkqGtCXk+6oUlilSegD
9tkl67ggsFAGrPLf/hwn5CFWiVvTak6RD0oG8RaoO0/aY7eCLL4oclzcg3QLBBr0
49sCZnQxRQQf/MY8FoeuD35KccEc46dHnncoZy8FLlDFY3eKf3eghq+h3ojt/3tt
KEUjrvv7vpilspb8kzfHPRYd7kk/Hk57GZaXw93CBkU6Qke4UApe+Xbhm1PslVpw
KwUg4TDUqKA+f6EQ0ThMvfMToS3MD4wL6TPQsmjK+8mJBr/VUng16Ko/D+1hJ1oy
lNXzjEYsqafyho+P3ap90LZDtHdlU4QifStaET6ciMVG+qTxy7OzOMXhbPvZlc4V
t7VCVAELzfA9p2+T1UgcnaI4mFaWjDKk+mKJ0GKgtvZ5gHgmpgAB7xHVhDng35hx
Kabmtpv0ZkNUFzRqBQH+32zW8kV8/7n9cZrpFVuR/VM0f3beJcb2uN9Qiqs+0MVq
ELexKRGi1b96MllVekzrDDquP5wBBIKMZMamYo35eQoy2f9ouJmdS4xPV0xefIie
7ypFmE0ivnokilgMmjkNUvm2FdTr+Ar+t8Z/6Rx1uT23sqjkSThDs7/EU5aLphKM
jIa/or+Tl1XOS/hqLmh1RVqs3USfdMbcJeVCKt8oH5oX1y8T/Jtq270fiq9HuTXc
CefWEmU3VCTHPO+bxmfxmUjvUHXbJUMqB3hisEenJjM1XUgBih5IqBv/5MvBoxpd
eNkklHP2Qm4nGmimFegNPM85hNcKyrumBAzHG6m24b7MVOsILMNAKucs4zNKBg44
twvT/VKl1Qt/k0CT/xdFBcKlx3Dy5mOY5WA0SsGcMStqPzPWMbcKDHT2R8mE97+8
wxC4IjJPo3q9+ITwVqk80dirklcedVdqgZuO7HqlnxT7V8te1hpkoHBvD0QGc+vJ
gxB25xK7pWdEZlO2tjwMVRWawKUHcrmq1CRP8yy29NDYIGATxnvyh4d3mJ2DiFEh
+n01QTQWQGRyzfR8gIMQ6sLYJdR9A22AEbekAiPmDDnw6G6iwxtyNBxsLuSstYDS
yzKey+mFcgCcgEbbyRtXROUx2GuF+ksD43XnoIQOIV/TrR5E1WmVKAFTG7P6U7lK
4lVzqOLWEzi5oUhrGybhVdEGKLLyFt7qXZto5Xy0WaaXz4fTm/ddPCbmnymamXcx
7LGE+QkCCQWa6qZp3ZCEleMPwpJnj/HDouw+Yll15iV62lvUoZt+Yz4KURqz0hkQ
XnfkJRaOXNipZAj491UMdeGGfkhyoLeFVpuzMQ6+3pBSkR/6DAqvHY/QNZw8Jcz4
aN2F4vv0CwSvYSyAq3x0YYi4+fBMBkUJii2joJw5s/JnYOAI9O3uqdZ+6YA3UseU
onVbZzAxejHBFBsP6O1hfPI4OUh/fTR2bjUVGIikg0CArJ7cUe6WYIn1gdn5rBFs
j9KXmLu8UHDis/WsaOyQpc1EF9hqLiBP/zFFlpKFa3qM0/+dpcYPSsgzlhQCQJi+
N8olTABeWGvVCLVDuKrTp/40scyXm3ulqCc4a+LrrDX1v/fFe3NiufLWeHVWs6/F
8+4LSB6Lm6oUH+DwywfVguZ3yDFz9a/ayrxCYbxk9v3Ie3iHIraG7twlIxMfB8Tl
IrEoa9gk8QI0mDuS4W+dGuUga0iQSqi1SqL4mVIRF8eHXF2+MANofQcOEkEU2+UQ
iqDSdUvqDxCiscadH+c4YtW6kTEHwM2+KAYLWCT5YzvneVFyAoNNLaH2bHi9De2S
EwL0Ay/YaXT+Dgk/b4l/yOGhUZ8hy+mLdCTtRGhS0ZMTCMxHLSRhROLtXqaPMGto
ZROduf0V/WJ39pid2qpHNe7UJ9t93Tc+I/9DmdZfKVw7EPDXFuKhpoNd5j816y1l
CLaK0UJQpkJzPNwUnYLZrHi9dCkOGNi6BKixbZyQGQzoZPZX7+tw0GiqjKFfgxTz
eokK0o0xQlwN1prZiUZmvoNqiBpq3KAJP74xA2iMn2xusGSKHntZhD/fL6119nAc
eACMHPl3jFdUTKI6le6KQVzK2hRM9dYnU2VpdGoyOSkhoyQriZIgwA0NEGNN2mVB
u27xCkf3MvzyYuhWZB91cEHQkLJsv4iPhqf8kGDOiLorBzrwrWxtmRa7K1UN49h2
DtSK+VxNtMHVWSrZy7Y6cJvP7EiofNCp9sIQdsMw8dkwzdSdQcN5t2/TnVrw8Bwp
r6RN74vJhUm3X2/G5Mr0fZrysDPQHY1On9vjUGHYljnJ7wZQI/SV2Jtt3j8Ljdcg
vpljIvl9ls/3LG0BzdiCsk5c0DfRoT6ZMEWiqn/LE/X1zHmaloBVXEr3qj88tB7M
+tCJrqOAdlQnLYSTDu58Mt0q2vpKKJ446yjEgoWYvQypbxMtiLoqro7BDV09/NtO
N2ITbhu32d7IjGc/2AIF+nUK0KHm1ottW4FM+LJynjB9KraCe744wGJz4KszaYYR
jrEHcUfORrnf1yrh2ivKVKmJqmTMpzVUWtljvZW0s2yEZxuSVAc86jjYSzDcFxt6
OPcdjDSLYGQpbjbqjXoRJvLOMjo46Q8JjsE4Md0+aaZScRWga1Y/67mt0nUvoZJv
RGtC/GMUdkTp14x9i0WPbdmOWpYloPCxdEnMnyfx7pTjZyAmPvk+n0sYY6BnoQef
gLZevX7PG5iqoTLRhPAfA0sSJ4XQVlJUsHemWoLROpJWL8w5BF4TfaRviTnfAu6+
yHe4RKVe3EkloexR+LYDUxXpgoydWLnHWuW7DgxqHCKwmVFN0OF3jeTBiGTc8hRz
GjBv7m0wlnINsF9i4loAleRWuuDChcNRfFkQzpOHPnzGnh+YnHMG7QmtKI9AVG/D
xev30RNjKboApptmWnTqOUp655KlWT3p3g3qJ8oJiHMPYVBgx7ggTMuQZcVSfmx7
5Y5Jy6WTY3EjyGM+grVnXihDEPUTXFvdwPe5IWfSH7QLX9i0TM/Zwqlzo6Ato4hs
cmCw4knoDep9cpYvfI/TQcR+ycdwAvEgQiWKueEW/DAEyJnbRZkGQmsb0AuLOkhy
0fPwCbS9S8i9CvKjYluqqXV1LSxfcVZ4/0RYDDYpkgeREE5oE2fVIEJmPQRRvZN3
cp+7D3LF9M44hvRzGFjmwbhySEtLdlg0Mu9AZAnHR7A5VDJ7QvHJ1uo4HfM2HzAg
faNClox7EVBAvyOYiXkgnAs9dKl9tM67iVZDpfF1yDSpSXruG8g0Vsy8U+VpQqCW
W+z/2dKme1evr1PKdzRhaoU4HMN2lbg3BhN98KzqTImECkMFL8mRi/gt0+Oj3X22
iA0PLPIiUoa3KZ/7D+EiSPULSC7+4TFpkdQrFiM0NA9Jy1oZmddmFAX/CNj5k38E
xo8UXrMBz61gfnY1u3eI5fcqIrVJ7ThTJ6N1aCtbfhaAeg51J1Bw5Le6X8VFLXOO
7VgwMqjnLLj0T0Cahp2Xu+OnO3INTrZ1j9n6ZPfZJ1/ha/9Ehnqt9NOns9OklccS
1BMnXz5bc8OtWWDkWuPnSZg6lToWltXQFvG1oPp+C7YkeusaOaO1AJrN0IymMAzP
uO63cIhO5/3NzwoptghIofGSmQT9pa4paYkJVvdT3ndAFLL+AXqLS9VcgP4s9Dcs
EKqrELSh4jeAUU8pKxVcrZ2rgyxNFBikjuTf7DSXqDZhJyxqCLJK08Y/QjQ8GvWe
5USRnahS0yNmZN/HkWhim6QmbritglH+32GuUvR4+95NU4oD5vo+niRwFMm1+6kG
vclFcBtTi1rHHckuDPTUg7xBAL/e6Ur6ywBJk2Ew8x6cdx9PDtR49wzl2b80+Yte
VxtzmVZ8ljGMZ+57OUwhxnIZ0X3bqLjNHNVhTCUIOPJ8HAIlz1pF6+JEMtv0o7l5
dKQrZT+VIV4wqI3jy/Ok9WhMDWay33zAG0lPWuOIueM8/15i4y+5+diJQdkSF4Ct
4R6Fw9IVqSQpltIdIr67pfhC7eZhDEUGccXOsK8MHAKCjJajsGuq95QJLLCgWPxZ
/Dd6WjbxWPxvIsj1g1vdvmPGPxRVFPVuIfektEsvwI7d+dD6nVuzpqDtTOxDwK33
p91bhlGV0ZiJJm75yNIvrTg77L6YU77H/A1hd2W1C97C2DLL9BxKDyHd2kncesdt
EpR+kTeSZb3hJ0RU8YjQEyilawNS5xERTKv4uGGlkNaeRKWC30cI2qnRTz/NnUUG
aoBpAxvMKgTrjZ652RxvNyhz/x/G9bX0BbhWJSF2Izf5H4/1xKDxZ3L3v4+dtcZD
Nul7zb7KoOb6XE3gAu2h54lXYoAKN5ahMuhe/AfXQERz5oibHRucTqRyx1fY/dCF
XGY85jXLeE7EZgbTANehRfTQ0BvJsPuZQ+yCmmw1fFUYLTvGYpxCRPt3E8lX22AS
XcJQsiEr4GoxBkjlrwBPULZD0vyCPAjJ73MlbBHequPoorxm0YiNpIBqyak7aL/k
m8kTJOjdcXmgCd3kwFglegXkKsyysjFHCg/fwjpAQy4kprhyO+WrhoVVCRjGBXMH
oF2obfYKMIg3iq1G6SgAHbo/dyjPDRHu/CwZpXk/QjNdJlh6PsLJdZgDQ6k1zc4r
IcWb0iRAx3Nl9kAJdmulQRP0TEK1PlXHRSJXYnGckVImKm97j4USesrJywoour3O
T10NafU9SegaU/twYAT+WTWgcqswwjoRX1YnF6qqI0qyrdY56ZdMPkF0i1OeeTdg
E3Gs/wArzpJIbuCEnoaUjkxxitBowqsBiI2ZUc94TQp7mvHPMszejXDgnU5CJ+we
+2kWnzPBp//eS1pIOo8lWnQnzT98wNrQjGJd3JKFWxqj88I/x8j9RPjr+pvYCxwX
VnJhy4WVvD7W+ByFjIeVBXW/O87T3aQOMeaQX1H6RfaSQ6qNGggsh2YJpJM9h61y
b/IEkEw0uOLCXaeg7r/T+RkGs+ZoGOaL1Yv+JRWEyOh5lMBtCeiqGsb2EuZ1jbSo
10oQE0n+UP1ylhqgJHiC8tH+AIr+kPgjVNhL5LqDQhEoFS4eZIQ48cGskOsTm2DE
g1nFXBW2Wo5rUSTngFZ3NVf66ZS7D8Khz+ffKzwrihyvuUNMaFCkikdt4Ch38Jka
/5YSTlwE0FugY90nsomEP0sUL9OxfqvG2kx4e/1FX8ys7aeGIfxGwHCwLV+dXXl+
2Sf46kJZrS5FjubWYHKVtS+wzcHEoQJglKP6zFvMhQ2osOQVXDu7YC8guKKeznrg
fpS+A8ZxR147KegjDKYz2mLvz0cmXNOEwesVY2RN2dEckSpraS2LDOO2s65vFefs
xhT9Bv1OpEwk/+hbHuZ2mGzdgxx0aodtIy4lQcg4iXPefA/9CtIzkuUHA9XQvVpM
TdC5P49yy1ZVZEoBJHlXiLoF4tiHclvYktGbThNpIJtjgeqJ+AJ6pAqgb7qI1lK/
H6xqp/qqdQKg1WDDrmovMowZoJ+GvK+anmsmDdwQRwBTP5oqNDdtmlU2AmBFkJLN
1gx4ry3l3W58uvSWdR1d33Mj0yWIJZe7JsOjSpNGGBg4BPo+PlO0ZkKsYT7ufUKT
0l1r/HgsWg+pWrVNV1wG5r1JEz5/wvuLDq/uUAg3FfFC+sgmEqugGoyxyY0E+1ji
ApCzLOY7lLwvqdrrDfcBH+XNvdJ1UpvpfwMMsaUpSaJ0JEnoZIsVOC6AJnWtiX/G
iY98/+SxMbYPuEnPIh9i1jTG0tHJNHJBKvHllg1lEtMWZeOYvn5SRRgxtCKM255Y
czOJFeVmuhrb08IPXgK1MnUqByDV5yTX25NDyH7aDri2Pvx6nZPVefd7QSWqWZHK
MTEbj1FEtbe1zAGJ9B5vtlUS5ZF/C71BEfguJd8WxqO0svYc/lWrXvBs6dKg3/kd
F5r2Jfx50Z4/AW3eIQSLjnI78ZoEF+u1wauvyTT+7RzZI7oKgwyC7Z/SClvuhw4M
4ydqYJsjMXuzJog2I1onmSAuhGRKY+gu5/ZE2xqToXtb6czZrT72K2vvSdb7DbI2
Y7cSQjNOSkubgCsrp3tkoF1ny1g0tj3mtqk4vzNGV3I0T7Rt67MuizY2a0bPBoGO
+JYmG81HlabXhB2vpRZYX7aOB3ZBBC8alYUXh+EG8gvJuk3IqkV5sWn9kmLeecS5
5JfsoJhK0cUY3Lnhk3kQr3rQ5YoAat9C5wzApkcdNQ+Np4j09S+jo8kQxKuczy7z
aVIkagRl8nBcG5FJtfqKYWOQo+Wa0m0gd2TKrcQ/WrgLqC2q2HF3d6iV38jY6XBS
57H0H/LzFqSAZnEn9cyuvw7LJtWSML6adNlPjH74P1fkLj9LOH/iwdbpkmtzUdox
DHTJiqoMtgmTvv45TYIkj7FbnK7m3d6+Bk4H2TFytTZw3VJWR2jwGg2xtLsu/vKs
kf1muhjp15DMHEHEIlVuGEgIlod5in2ko45xuw8HDNzcydeLYEt4XAsjQbQof9/m
nPlL1fMypcFRiEDucfLhlA+zxExNf8X8i+dDOBb5IOrzX8Ryl+EG89suzvW/KqE2
XDH0cHHFwuDsbNP1dRZWkPqmA5RThpmWj+MU3NYV9CIOXm1SL0oA58KTU7NEephG
hggpMTnRco9qdTaDfsdhOgNdIuv4k8SvCSxw6t2aJwvL6tkNvRTYP4KD/Z2CM6Ei
zEkAGhdbyAOreaKWGetZA0SJ2YRu+NzNT8m84OT3JZpSKoI58IKaMRT6oj+Zaq4m
VbbL09JfYizHwNO+jioR1WzCuXh8W3RTGpP25xbJTYcQy3b6kZRyw1AbbXU/6vH/
8rRdKXfy+CVbtWZbNsUO6wuew/CW/BtnQarghZ/TsegLTyFhhfU99fPT09T72YZh
HWgfYNN5W3GJsHRnOW3xOoHWZb5aZhgMETR2x0JRgd2txfjUywrhS6PIx+aAz3SB
53moFYbzWOoSHfBnMgNTxFE0HkL6VA/Ow71E9Ejd3AKYTKz0HJrooUfMtrQN4Atd
2g++nu4/gBTfNJONkM/KS3Htf9C5wAif2uC83I84XofWfc7cf5sNNepzIkWRpERQ
Q5ghlE7CJkM8ONPUixYsl6bA5IDjoMiW7pQDj4q3up6mC5v2EIISPNiTCKDZdIAR
har4TLbXGSc1pUc6QpXTAN13k6MICcm9stfDJJgMsiWb7ij202PSPDRdDDj46Jzl
I7TclMjOStjyKuCACFeVE2B3Wn6qpEvRQtc0mzmrmF+4s3pBYN7tRmgtClv2RX8H
RvWEUjF2pm6kbiBU/z8oLknNr/Hm/cKvBFjbtyRYgub3J0/TuedSsSvdC0xOen5b
3A46zgUaZ6SXxFDZDcegbF95kqe+ewBTK07Rcl9EPrQIAgwaS4YxqV/X/ctY4+PA
WO+jOH7Uh7E5eCU98QTpTUXEoWbM17LNJq7RiH+WzgzYs5YeqMqicukt+NMW+xUH
Y4acP3bvY3TNlrs7ap6OEzkOBdLLEXwGghXr7ZuUuvx2908E+dpDNSbkwlkiSWq6
BX/IzOA4AVy4rYj2rzsuZVTiYS1bXf9/ZbT0YDVRc3r+UUJoMhCszfC5lPC+RRVw
WeTcpa+yDh0igZw/JI7fhh9V/iDGrZSe76D+j3bgK68KCo1vyyDonhh4wriOMwMs
bTIv10jvnWcifYncTZSc78J+w002iVLH19qCY67EVR1lWHlgt3JtJLZMeen34RpJ
wfYytCmIhkXXQyaq8M5/pgYnRIWJEEfPDYAQkVqpq9fKSgC8Wl+FBAn9f7LPcwnI
YB1tqR96SRQHfsIVfXuNsTVHwYIMH9k8H+ZVYeeAqR4lJn675GvoyPIFtC44LfS7
K3RnlFO5lBOODVffAVHaTELHBO6AjS8wqX+xxFAztpN1GpED+nH1mYBEdgWZfFFX
k6SThbQZ+2w5N0b2yyQg9ADVNqZo/k40CY2yQNvmdNdIGZUn7LTOwkvAa6bA93Ix
x1RpeZBWMYoK/680OVNYlW5LNg8Lc1hOgtQ91/i7r5zg+qLJpXUrUh+P/EdFN+uD
F0g+bEgytLUJc1E3JLlHeGxG6aGu3wINQ21TSESUdEjIEkPwxjjO0mEpqZMWgSvH
YHaiASOnCuu2mIwnBVr0oc1kIoFVpDgsIRpjb0eddZPXLKKJY83QoDZn0gVRxeLH
Nd6sNtGQUcqbEehOg0eHkoGWqF7c3VVz96BegBEsrluZmVh1JmYWcd9LP9XDiRWJ
D86Q2pwIbNGc+NfPR1HsuztGHQyDSa5EUp70iDxiakxNq5RHMZjuv16azrdP1Axa
OLlmy3SsPxyKOEnalU8QKz69Ink8JBYsteKeUqIMiA0rL+sRsuTfhFcjD4tQptFU
N+vDOTl5He7a4G+ghU5rWGtq8MeRrunUr4SkRyjXEw9Xd7MDWZpTrD4UaS9si2//
WfyiPkZokI5ZCiGFWC2G4LBAjyNdpwETsemZgqrSR3EzjHvs+hSayJigFjgYXqUK
wvwIMej2Esd78NqIq99bz0ALWGEKOgexMuYBe4yPVXyUyRP5H5ZA0biWc529I3RF
e3jS6poLJMu5f63v68Marrul7JrnsyDe/9hCPnrZpy4majnIICe+fdGvmctwiJkP
R4kRHoK4m7wDnMqh/EHbt1P29zHcZv5K6XH8Qo2SBmzlBbHNSJjHRMc63nWJwW0l
0yAY9cdIoeqiSpEEIbSfhWe5SdeuNHEG+F4qmZV/927EPSuQpGxsNL+8In7be7/S
lIcWWrpgOAWM1K4LDnlROoH71c9YZ8I8AZBZIgD02I2hczxN0P4YJ6Tjz44cj7PW
P03fDKGWxrx6vnA9CO4yeBymnb+EC3PquQvuasX3WtfegbZfJsQ8siRuf3WVw7Vf
t0TnqOZ75itwSAzDG6yAtt8/rjlwQeY91je8aThL3ClZMSdqqZJKCC/Gk1e1mva/
kuoZ6Q66KlV4g9foEi/EX5h8a6O0lEPt+g6WP0WA8zWT+CjjI2mVc8906ND0PBmN
RyQPuQtqwR1H/cPWICyZO0UDV7XCq79oI1P3zIwXOY7jqUSoaES9PyRLKaybRxB7
Yu2JA4H7hVCClB2+s2JaVuKL9NEpkubG4vYA+fhuApwSft833S38blKVi9Zm5TGq
HpoimiduKgAjDAdP5KAHsKlhqqQWY16tOxlWPD0O/k46/ILboUbym6RWH/FUWZfr
/ns9egVBszE2kVdDdczWqN+Xm2elo7keRQPlqJD+REPn8Ao6l6Da0DV4EypP9OaD
qEIlWVByV4j0uxrdax5W5siYpkM39veua1+2Fd0EousniKyCWx9A7ZlahDPxCcR1
eKxBI6IMKBJ1sMbbGgKTWFA1PrdcnGUr5v/miGWpRxRjSe8NiBLblPDBR8cn/NO+
AhhF7p1mLY25QPPVF+wJ7vaXshJtgnRINx41UD9j2eH1A14a1iBAXjzPkAxJnElT
9GQ79Mp8xWFFakutBSNjGR8HixRs+kmUnHNouFZaI9Kwdh5LKZWXtbeOcf3rIhtb
lg2RWQUERCc7cXTRHZuJmo31Q/qY4VRhlE0jgpLmMsl+hVZlsXWDze0po9GRHnGW
R/0vHdq1DenKbV6NvTngsT55fFHPp8Y6uWdwYJ7oZbllHDQ0SkU+rXMXtc3OC9hx
esp124z4lQd0DM5yQkDvNNMlbUwo7Fs2xOajutPqrRcApsq6kJ3j8DNqhyPTqO0/
fN1xtMmyxLJi/El2Er3P2WMtdx/kNB7f3ajGVp6k3Jy9eWoo7x7DVUvYUZFXhZZS
y+3tBjFmXJ54QQuAYe0qlWFqJ+kx2A8u/1Pz9jIXjIImedZcl1HEGS1f+M8wq8rn
sbd4YmnbCWr3foPdmQgAeN3Cx+c8D0Ewzjxg0xltN9UM0/eD4Q29NOwqeINqqcMs
Ma07OUHfjcDRY+WwhAMdJzfuMnlmDDjdVIwaZ8bIWa4sF5J9wDjS7w8pzRDX+zy7
lXt94O/Xe05ZDGhcF2Wi+I6jZb1AJcz9BWkdbL+Ei5vl7ShPklylc8jjwNd+6OIn
1OUnpq2RHpYXJTR2C1GERvc/mHZ/tJ/ozpEZ0mdSuS2boiJ5fw4m1oM73aYoshEC
Sn6GZoC9vTTbWsIlQhxfWYpA3+EfZqkEDcWfDJ//oMu47abJsSB6eOrzp4ipeuMS
syV+UiY6CKJ6W4TEe80mTrfmFaHlLHih+LEJ4fuiu1reheyJ9z7JW+r9PjaNGhJh
Hc1m/kpL6+59vo4fLNw+bPBuZ2a0IVLAHh5F67sRxHd5axcfqZwCqAdrxR00gKVa
8piyaip6sXy5S7C6W0JLIr+CpqXscrPd5P/6c1VrCHZzn4sSws1qtcwC2i47JF6h
EPfv0nAJxNgdd9a6mbC8NmcUgu9Cdj5gEb78CW8NARH2Sx9Pffw2bIvvcwGHWWjU
eQBa4CR7dR0Ma9P8eElnoMQryhFXIAOrm5LNJC55jqGjUAqfE8RZjpF88o/mBIER
MDSqHykv2V+jordqSqFhqpwCrT7txQ6Jxd64ttqF9Soc1Pgq5PmvrWKo862CNcBH
lYZiNlx4MqJ2EBKh+aNii3jW4GFizk+EBau/gbvfMhkhSfi/0jFz2Z6Md+laJOd4
UV44zSRMdn+ogXWZx2avh33uhzk+N5kNZLuiAdj8EX7YLyyvu61lIe6C2d3asvAm
nngtqSyitjhJy/uiu+MSruPRUcDox+OgmhVHxIfiUUk5SHmBiRijVHxUwt/W6AGl
wPzFDxMWxOk7rgjL0/oZs5Q+BtD2hclLX6UpLJBwvaPC/k4YhaNcelWMsCFvIhvy
PBwMUqA53LZ0ZVRGkBf/4PxCRmws45xM3olpdP7/CKzGN2uVn7EqM2jUI3zPbZqf
K6GkKADeTVudsdyIz0oQ548pg6uQSbqJRNyBVQsvUJOegLrreHNCGyoFplnAgj/Y
LCKiaGX/BMV1xIfB+imewRuPTIl6JeT5EUg/Uy1CF5eiT5L92ZQZNgQi+Sa6DuwC
yYEdpKzD4gcG8ymznO+YyrFHSpRqH3bYGRUJrrRYacxUjIV/H5LcJ05BFIELN2W1
b9wwIFGSBzREGH4SkHUSBKGk0ywROfYuQprZbAHr7qz9qvk6X2niuJtcdRABFjeq
sU+ke6w71TaoRiTycg7T8PhG0eR0eKxIWEj4KxxvvxZy5itWKHlU8D570KAWHqwz
TB6E2PICYRCr0xAfu2PRmSEtkUDvNFA/Uy7KE5EELVG3qjye+FEOEq6cTclyc+GS
dqD6ZvOUX+GbQqBR82CLcq+RzLtZgw8SRUTHrUtXWW2B5tRCpTP+WzT1Kyn93F2S
NMnYVX+jFSc8CtZKsQ8bC/smD8boOC1Rfv1QZqYkQKMNzVQgGaCNdn7oQ0G3OVJB
ZOmDequmcVCz2mBi+JXfySUWbGifJb00ZGbFcr1dT10shxsap2Co3ruv2SvMjkO8
LsrM2NsfRGcWRV8VPsAORqjTboyFntz8sNgnbLSxT/2j5hsWrPorSjqw7DwTmKiX
H7oekO38L60Z8cVCJPBqIkhgBlpksRURvI2rDvO0RKAu0nyKJDxQycoXMc2iMmZY
W1OwbHgbFveQt3L/LC4vEQwnGAc5TRQKFZpO/HSCMJqHKMaEBrNzXSL2VWuvhA4o
Apx7jBr5F9GD7tm0iA+RVTOfhyP/ET41fkw/sWKupc8csbVVk/ewKI3LJ22iMIC3
NU7r7Da6+TNyb5RJHF5r1NfnTJO1yvYFeGAmoujofBu5YaSs0kOT419Wx3N4YAje
ck2u5I6S8FENcv9A/f3eHHRbsJhd/7MeEiTHrwVczinGf7jDolVMnh3288delwoJ
0Y39DAAi/LoDjC2qCJc0HfL9zQUspBS7WW0KgME3iN3E2cFlubYrw1ouOpHq+q90
u3JRaDSrkId9dNW/Rp/NkZY940betTvkZ8cp5fVAoJqXQbaN/4u2V1sMvn94IHV1
DHJsiBhG7JAKPgZAajEy8l2bzECvR28+48wqxka6wtxnSUwmY6uQQW1huAp1dwU2
L0IgI580uPrUKQu5ZLQlbPrylRkq1ZKOjvetnK1ymy6axUyAhOz8q+MOSLefoNbL
bVU50PyXEXVbSlkoHIppIRy94FkwVdVjIdRUQagTO/aNSnwv567RL421Zk6CwO2+
o2jW+7JG+tAC/QIdSmqRkO2FOqqR92Rj2Ng7FpwNBE+oVg99UxJBe0/y4nz3AfqA
WNeg3E6XLb1iD986cqn8wXPb+4rwlE7S7KrTxX/J0GhkfMeBYnSJXW8chb8PWJKh
n/VX+1kMS/KLUwZ7qX6OFk3F2sKn6cQN8ZBC8vOl/5bTw4LrPZTgwWzPiBC5/CF7
8o+X4Ga/GkHvJg3FUcGhU1kYSKPLuRcOJ99Nh4K1L/LTsFuNVj59Wp8F2SBx83f5
R3FCzuEE+bcQAP/UhfptDE2SGquvLFKaOmUXgS3GtYHwcV4WUkC3SnXc6K/MPXKr
Uy2shHOjaiy3vUmtcrPYgU1aE1ztI4JIdmZuWvTjSTamiNUJxnYqCUAWujcA313z
jvbWfG/k+MXy9WLdcteS1unUp/MBexVHxX1lpOwpdu5cYmorw9gUwnaXF02iE0Sr
nylekrGfqAlbfIv25aThF8KVzZOr5ZwXgcG9hX8A/Pv6GJBlZkp0IQEiWhCXhbZ5
FL8xnCh1YYFzkywGS/re6aqxLDWmexjjsgsLvFxLSqk9YcHkqOca8Z8VSzXUvbTD
F7ywIKuPketQzYho4uNYcEvUnd4fUQxiQnwNUMsCs3ZYT4RBA5ctYGGsI9+Ygsu5
AAHe7q8iDOE1LFP8a+lXquEx1Aycv/JVEvWV6yJFkyQ3F+3ahjJzKt2yAoPF9AX+
9KHJ1sEXXJErDagtaqPJD95VTAtIkwlJFSa8vaNQ2GqDg1sas47YepZ+a9fSJYjp
PiMlq2F3s/1WDLKKR0gGbwg5k4K6L3HoSuIeBEkHWsdWuQTE+m1YBOYEFCZ1xSri
EfAZ29A9k1IGG83kPvm9cxPJ1Q/TENVRaTD9XqN48GgCIANlzRneDOuYaIcDhLnF
ILP9puM7KoAa9DG4o8oWZgIweQNlXwOqZDEriTTWfhp8ji5ruT6tRDk25QVp4yAq
jaERYHDEissLMO2vK8QXdX2bO0hzRjiLY4Wja5SnhGbWcIUXKGUlWqVZ5O+fk0YN
mqzyhi2WXPovsAzZ5k23sr6h6IX1ZoI4keXW9nUnI5npnxhAd6Taef+EA2qtRrKM
um+BB4dli8hCQtvKy0bA/Q2oIv2ZoqChnmfsNsKox9Mq7sNMFIqpai/Uv2hbrINX
J7EAkTjw66eW6V79pawgwnBeZLkc8bKqrMFIfhix0b+Rpkxyzbh2S22/a6eqT+jW
g/TKAQasIdaa8HjfMy1waBC6PMyLBDzEZS9lTvqnRowEDE/BogSmcS0FW/Rn6jb4
/KVj49dORuPGuhaM0r2v9eNisDK574ouLsU1m2mthVBR4BSrN+viD4bakuJwfxwr
7BbU9+rQhvIvSLFy2d2MDH6faIBMovmXhuJcIcGir19HmsEtGc6pF5MROMnyHSit
JnF5u1Jb5hbI00byP3tpoE+ppPpqxdgf92J6n1beYdofhP2HHsD9VHpbPAXvSlAH
W+/ZoepxI002i7+JT2SDVrpvh1HRI/zEZbHs1c+RnZ6mzW8DR+5EbOKpGcoGiK7+
KGbpgfLjnx85NO2zUO8TZqkZ+aZmWHUvcR7ZRWAsLoXH3AH9LE9oetAeC6eJt7+f
HUOZoS9Y6Wf8+JrYvVNW2t4r/gGAuHGEqNfi235rRBcsMn9DaQGChF+jexIVfUkj
YvgvVnZYdyz1sWCZSo1KDGdL2pArMC577TSQskqU+JfKrRhHc7Y6S1UDRPp1yulk
k8OaIast3kk8ByxzNhutydQjwG4rtN8jCIg2q7XVBJyciBIFtPCcp7kAWxihbWYP
Tgh8yvRjOS0feqS7crJRvV0fQMtzDdoNXrPZi1z0qkxyaigjHW5B8mP6bWH+7v13
2mYKN/yX1ns2qAW/rw1pYYnegywpMsz5Hp9a9gs5TxmiPEbtxLk+vCVoCsRbIeYI
+67kkrjbxktqJ5nVgW/E17v7VdC9lkvPXLeTegd/sXSrjIPgo57dj1mcH28xz4ZI
+x7FxlkHvihG9RBI1qv+sbsFVUJAmarRFsICIFjFLfayLHlLczDNPhcSgmfWO2pk
ViIk94Exjm1fxMGNBB+dFXRu82XyACDFbpwSNK3ksWjioOlAwBouoEG9Gg834C63
NY22v5XYbCXUpdgc5/IjDoqh5tvQ3pIKn7fsQQ4qp5R2wP8YAuv/kFJLSXQIDgJx
/lkn0u/BZsqCLa0HSYGU647a+ou60qGp1JM+v0tJIO7ufjvwG0xeryxJM+8wAQs+
x1uv/d4PXDNxTourV2bltm0YGUIy3uvTxIMIXMh3SgsMpw7Zwk+xsdWVHVn62v3a
4cLqkFHggGQZvik1fpkL6VEF6zAM24Edvng7gLvh/BCkbs017qedHyF0GwU4tIUi
8/LOrLR/yMLQGGQh4mzTq9tEenyIEE38ajPS+RsjFTe8xCfMgaH5wn/oE9oUJ2JM
0HPL8EF5xRuAoUhV8Lf36473rj29VhXrTpE7cUM/BmVtEbkfUk44idCrvxqRnXQJ
iZSSfR95oP7NPCdyBALtwT0YpghQrS8wlJQUr9338leq00ce5QQ+7yLvak3mtj3i
IjKN8AnOYGcqxoO+nRfEMR7f+f+o3aiG2ZhwxFs0auMQROrOboy6TbLeJlcjLhp6
NMnuVZoSmeaU98u2rU34rh4f7IgHqCERExPKs9woKNyULZPRhAJ4qo5qOV3u7Erk
2tN9r1JWw3WPxS4C6cqWx6BoiCcpeI+pZRzLrzHPyuxIRIGtofACldPRtRG5/vb2
0gZaPcBBHObKkzREaENe3tHVJbui6l0QdsVyKYjSgaQ85u/ojPl5lOwmcLE0fUTS
Hyqmd060NAo58ESX2yV9k50g3rNMksLYMIyaXaWyTEXjKuLZ/jeAUizQ0SdSPrB5
VzqRoLRN3T5SH4syhjSyUZOIu/27W0VIDwV8c8ihNVSC0val952sglUk6Wn8aGxq
+ubowafIW+AhHM9dwmsCchSuZQcmPDHeXGL12CIIx8Ldj5CrsxfVIzsnA7nudbgj
ltj5bMgqaUhT8n6gv3DongPUAYL7b87TGNXnsHQiJG60zB7e0KjvS1hJeEgrUku1
t5oeVcCVtNIwxYXJf/XvveHDEbpi476WAPuB19jfDl0hxM8wJCwk1skfcR3MaidH
sJv/RR/pIt/Qt0EEBtbgbEYxgSBFubX82/WWuCy35Ry0IE9I0NnNQmLgcTeGcasg
2Y4BdE0+TSlZyjQWLoFxLLILZgLQ6uqRggWkxaiEOT5/iSB2F6FzEb4S6YJJ65Bk
CkAMExTDUxvaUGJ53Uf6haIyQR9jjwAYQVd5o9/5XeK8hVJsD9aesU216mHFg/Jc
5QmqduoeUrXwsYBDLq84GBNZtVBttq7zunncfbcPxRj0aVwf7g6OO/Skok4DBHvL
DHArHtF7OZ66QSpLWChw+uEK22+q4a6GWyx0XXwHNoROiTX2HwY74kk4t+4hfWOc
WoQxRMpMGtu997EnYMPll5s1nYXXH3F9FFUzdg5AyNrhtuqetGAizBSa1kSH3yFx
KduCjClRSPSyu+sOkpzKIySnAKCuQ9degjgrdI8vkkw0opkslkfHG/I7gijAh9rM
55KVxchK/fSG8GK6YzvGihl6OvTzywhXsCz6G5+2lWGzM+zdFS0tS6Sc2mBef4F4
uhaQYo4y+ifbqRqZAt0On7/q9ri3YORIY3HbWU7hUMcVaZSU6FjfkstrQvIKmv0f
aTmcz81e03TWgH/SkKEltPNL1kivaVjf+QVdXA4+RxVzx8VilcaAkH67uouj1b6j
5VfO9+rwnxeOuQQ0pTFLbJb9yqx9MCMEPTVm83vHNTIxYNZjpmwSawiZT6Mwd8Hr
GsMPAbMkr4yFEbdhvZDAxT43eEYPf8KEiiXiaPPhrwq2K0gig59qz81clVLqIO+c
i7D5THpf3zobJwOHytb2ZRwA3T+y7ykT0QnrgMZNAUqLDWLWMMKIhXbihGBL4v2Z
+E2V+piEISNnz3qDfxeFx63p94B6mo2v69FlIBS7fClmikmENE7lQxVDn7/MVb91
E+DZSEffC9GR4QFPsffxPGQ4y2vfOQNjrwBCyuxNSw7NM/h4X8nRK0U7S3cnRjSS
9Qxny3XV6Kh8GanwgDNjfKGP9mM0dpXJswPclVnHwjgVZ+BEGXeOcct4Rah7IAGB
AGrI88ECiP+aiL5qKzmdYCPYU55+NmDAQmAzzJaFzGWuuUh7wOTQYLm10Y6dWG8S
oQRY2pyeIDRr/WhYoLt0W2PBBoWcXZXFtURZ019CFocvDExT5F8Vrq15EIpT1Ibh
eDaPH13ZSWEn9tsbGzgnypzvDijIWH5ztr9UmqI5mXCEvIwW5h3q1yzHDLTNVxv6
kuxwMWVLqzBMOOATONL3ok3vbB7I73dIRjVgfIunYHxlPOvgs+cgHwKtwdeQm8cH
YuBManjazUye0a0wRKSNBIaxwzganIOkSPKIq4+kR61oUoNkkvF+Ub7n9LOI6MGW
+p3iXR+ukFdGd9LaIY9uc0Wi5DPNZoSXKRhAvRE80BdyeOsVDXgXh+uzkQL8rE0u
Tbd7UxCPWCMq136/O+pwObB8pwkcCsHOMGaMTba7KfgAFY4jHf5pg2SL1WI5LwzL
cPChQ2DZnGCu2e4R8q/XULyJtObGAz6tA2lc9Ceze0rJcKBZrOf+Xd2dA/gHHqhS
D/RBTbABP8+NsHY1rl86YuBhDF2lsJhja/WVgOWK9fjtITuO5++AOeHb1tv8LgaO
h0vh5SX7gsQMIVNrIPJbPzAoPZhPJ8EftdWuo9g34JiCmiQ07Su8Jna581d5jaQY
Byoq5nlztkWD4qfyV57O9X/SgpFLpG7qFmj6nDNr2LhH7kFRDGZ176WHk1o7no76
A6l+uA8Df6F/oUtzj9etM+MQjhZDbaMtIefhEsN6JWtPcdUQT4n71bPXK1W7KalF
rGzDYgyLsn45yMg8dSXW5oYqL6RSaIBUcfO6UjFs+j3eGErGf9gRJqNsNi9CWAgW
WwTAV0DAgjH6Cqaicz3PnGxgYlz8ZvB8SY6eeXenKuqO5QHvrE+EJQEPHWZPie1a
as5SQXORBK7TlMSDaMvg6Or2BUIM+fH4at6ZsbqhKP3KPYrvVUk/Tg/Cc20ZNXe0
zTmPAyDY6mEofJhzFMRJ5gWXY107EbZd2hcACfRUcHd0IoVi5nye1MssTT8DQFgO
6b1OGrNwW6UUqMgknW8skPVCS30REgM103A+UUAdKaugdU8wiwR/O0D1RcEjxYo0
CfLEmWzWvFPu7/RksS6RRL//y603u5kNgRewZaVJi+m8Jxi2vEcqPIg97Xx/Gb38
QtT8GxnvhWBYHKFWBbsml9U7fy7RR42Dsy4P63glOChujRR8+Ldco3gv2d7RGZUB
bS/6fjTwdReJodFZGrlBAfwHFoe9Y8uzRMgUSirCiJFmH7s1Ip9/OqCHOx5hNPNA
67NthjvEd2YCsgH2GXN0a0THmWMf8rLnpH1v8pfQyVUlY7aTAX9jfrdQEXYs77mn
K+45wbM8f7YVE/vNWDJfglqUnNFLnrFx2DOuLEI3Ft2xGTIMwy1k5HO/QHVpiqU+
PMU0S7q8INCSQ7mKOv2np5XUSWYPXchW29O1HX53Sf7bBEdOW8skA1CLnmkDpavz
N4UJlxn9QzUY6fltNqoG4jt6GE32dPHAikv7QZz8t5FPyTeOaoB2fc5pnve7DfcB
AmCJtKpckyu6c5ctUpl9nrSzCTawprfMHMd6SOYAeOYwn7SSUfqCDhkPvUtYGgfB
zcxiuYcm4d5atgDX/iebObB2mniU9zjWWDCdwqGaWDqzOhnDTn6Imhyky7uTcxR8
eu7ewzb3qR9GAiLnJCPMTFbgiRREHi0bXTEqCFJxUmkXDnLVv0P4AC2ZYG5ObX5X
Sy5Xuuf/VBpmDNVaS35HJMQJApfV3S/Xidf15Dvfipgi1dUhqn6ORMPXBNEiStjd
8GgIJ1Ou79NSoTB6+FZiv0+8r+1IE5bh/9yTDDiIUW+0tDZx+U9T06AT1drDiB/2
TpfIwSf1V88fD0GrX1J6wE/a94kjbostIjL6gL0NcRQ7x/WfbfzjG90hOeWJW/uM
X6SRbu8sn4rJVxNHvsiYMtsKFPrTRRjL9R8ELKR+ucMSozE0nQswOaBw7dNmAGMJ
I1JPMnA9OqopkLztOQ6cqseXfPPZiIJuSdzNyHdy7jTTUxjQzR1MT5qXiU6NSZed
xFdc5scJ56u+c4dlUB18/YurJ+DDK3ybFId/QaXZn4L9lk0T2uchS8edUPIV4gxr
W1AGirdAuITENxAFgsmOQCZOPHliJAN3ZE0KbM3RmNWdjzUHnIO9jlQ8zy9rgOIZ
26n9ow/pLWyIXgKcPMlwaYfDZOInIt6ZbLQ2BLfnz9Cd7FpKOY8qp60L/I2QObii
rpXEy19fLel9l/8fmo9HZL5p1CmTB47EJs4dZ+8Jed/ntT3kI2Ckr+ZhHQsvjBWb
wk5mQ9PDn/ggLmB0z5csrZiM3ZxIUoNmbvzOs+T43f5s2HvrwB9N73SvKBrI2piS
zaddHbnsmy3h2DYOFMT3AfhhDfxdStIkkdknrEcidpwjeNos+Ir4uh4vh/44FAIW
O7xNIy5HP1nmvtL0epRBAZEb+sqwL+zftOWNrIAOIincHOS2/KXmM3gKy/BvbvcS
ASqwRLT9D8ha0K/EW/y5a9KXpGXAMa5R40riuoS0bqg6uKDMi3w2/uiMh4Kd0lSB
M61uRuXveJF24ylfghnIJP2dnulyRt10HguLjY5Q8nDha8K55WBX3qMSmrS3963f
ijIDgdUkUqc8E7YHmYtgaBrf1usR+cRM8BzFkbWueGq7CqQd89K87zLT+vQSewFY
EsHC7NgQ5bj4wNDz6eIrn+ABGWyrw6pAl9X6iGMbnuCz45lUx6csIcCOMkQ48jcx
ydn62PsUmVGdEUf/KBlCsCBHuDtYgLqREvGzuxwwp1In7V8konDRxaJNEbFLK9Zx
oETU3wsmbGgIQHFEt3ZuPTUDpoaa5zvu5dS0VbrK3lMZgYKnv054FAdhchfxaRED
G995fdx2x+kHxcM7Pm7+WFiaOeQQHxG5aGQ2WKbF94lW3Sk9f3wyjFRExFJnz285
nzu1v6u74X0Sd5J/Jw8B/ZTuxhPVDLXwuJWOr74br/7YGyXXRyMzoG+72QwNQEJJ
jLSXgGtRnrrjxi7GYk65Y9f1o1ICDdX1DuusHpBvL8MDrvYW2evwFmOJhhiUttg7
ZZ/wLR92kahG/K/Exyrkm0kU2jq73nk6H9RHVJCTUPVJM0vvXu3cKVjJNKfWiFUx
jybYR4tRvag3dISTc7UagMRYbAr2Cm5IroVU0Ugee5p0zTJ76nJVrmT4D95Yk0bs
AfyFQJ+eA4McSWRi+MiKz8PCbQLzTy44w9xZJzmELMDN+InVZy6Pgv/V/45zYt7w
kc4GMZkrLAVBSofPh3+/m6HkR9MbaFzOL7Q+/V7+YHd3NFDSeWCH0wyo+0dYGQkk
5P22O5Re8Y6UccJXFUq51wLCEoHWVV9YlhOxQR0O7oXsyDagF8OkIWamhDoXzHqb
hY83LiBkmXQC+7t9ScrI1oKBYFOPw1gDhc3Bnc8+EiINNqj8jCJzA3C7qvAQWF+S
M7bfilppoWfvh/S2TZuWgmNTpO72p/OTOi3jRPQPpj1PgVD7/nUK4lngbARlkpQV
ffoqmslzlhdikVzV7U2RUrhMVYThavBYiVk/vTB/gbtudt2+XT4y+oWGgAt5Mwki
WEjy+fMVxhde6tQr8bGc1EsqGUGYuu+Ef0jCiucuU8dljFiSANW7QQ9wFx0RudId
wdwVF0FUghJvlEguA1bvOnAtDJUwKlLfoN/B+YxrBpIRQBAEXjy+aOB9jdznHH0p
YxA7oJIZeWWLrTFe5+85SERiAzS4NvqCSZQcf/KklNkxqo0iAODES4mW3szM23t6
r31DS8CxCSvMTfeS1eb0QFC19Im/+VEpKrgR1VG8Yf93vci7aSrN9e0e5mORLfiJ
HwHigA72mKwMxWHUdn8XS7yXrrc3gH39ded/3cqD6j9wr4SUs+c5Uv713YskJOE3
A0jSLTrdXTfBiHyKyYXEE7mCDQd7+CMn0E6mw4h/k547GO8py9TVTbd7AHtsxnZN
WO1Xv0UhmRJ14eLQKa6HnPhF6xMqNKDBAeyw9G6wHLMKqSjtoVyT61jNTrRieKaB
EYRtDpU6cx89g04wxpTtsr7AzQLbpG0mb53SjKWjw9Ga2OUy7aIOMKfq2JR9AXIE
O3xd9nZyqCIya2EYxA4vxPy73wH7Ascdtz9hKGp54h5jztlqnvUXVB4eUMHPqdWi
mh0MvYXrctGuEzcwgLbDdHtwmCX6Dhg7Ab5g9hZ2wxOUFPntBPXQa5TNBQtjk8LA
SvyEmfiNF5kdU8gddAKPQxH96ToUWAQwfeGk9o9TsQAUNAOeOiYyQ51vIq6B3F1M
TkjCCW4j8h2Fh124FcU6t7vkJ+T4UB3347c6Fyku0kpXCcid2GtOIOaodrFHJfiK
LrjCtp+UokjzT7vOC6yeQ03czaXywTAHC5syZ9wt8bH6C1V82jMYuWTT6iLXN/W5
emluDBkKLhJAyAV+CoMzQnwmajtR67kK5ulTxd3RPoMwr/R/12niRB/2Hd9WNclr
3nIKe7Tw6MguaI5oEUiWY/oYWMrx1t0uGJo5nhjzfRNcGhlm7v4b0QvzB9oCiwkC
J/8xSF+dj/BTbTDVKaaLgylv2QO/TAMY3rE7jx5fGPFZZc24VH7J4+hS1IKZwa2Y
YlX2otKIsC2s0HgxfeMIzPaDbRZYW5lfcGpmUGYdAKtZbLHp8j+Gz4bkSWAVcAPs
Doqugnt8oZ9XZKkygCqjciks8QNoac4GTzxauqzCYc4hB9yBQNURSoA7FvK1MCB0
gAu2Q19QSoYPRIhJVsfF17BBTs65YGe2Q3u2eLM3+bSIUYKs+EKQ0vIMDNdU4OkY
jodQP3j3IbSakLUsXfgYbL6uTQvri1fLztO6hGxUsIJ7BJBwiRmL/X1pR+jG9r1y
SdQhESwstIEgT9919+MSwUg3tuhGDmJzAn1aPxZc1y2GkF0N3eoflm3u3osM1Qqk
0UwoKR8yqOWjjCKZeNsPq35rQfGPnvAdPmvigsdoUV5/s3zNwH8zr1OAqVCYlyyz
czA126u+Hdev/47OOT3lzxXV77VAzEUUeezD0Q4wonK+HU0mEYx9CYAgre1Snhm8
30dQ4e2fVCU2iTMz9D62OQA6DQMYnJIln+VS+mz8iLKS2/VCoS+AWVA+0HyEoVKG
LGTWKNxNSp6FGYVJ1G+I08diPxF8ZUAPWD3O2LAIXTKZItGsgBlLkTtWpHzExgRh
OZJ7ETqZgTcsGzkWTXJDt1sHiMdGG21CDAAxmp0ahoERu6SoxYnouhRVv1zmFDUJ
EiSc3I1k5wZbg6JD3ZDGLbnlljllP3ua3GQrj99S/6kcffj2uGv0UG6I29sPadLj
WC0Zchnp7SOkAjISw757DqwL3Blef4xn4BX57AcXzG/nJVDB2eKIyocM64fo7zCK
mYCzxgotsYYuuREE4KKnHYehDzxDzdgTMMLqGj8GMCyG5nXEPnA1GOmPxtUm5N/0
yslgCfNNZxUp6MoBy9UDoQuvFGG/MrGiqm32561aOlk7MXViC0VML8dULhdlOv3z
dUrt1foklhypCjjGKOM7jLmfpU+UAYuXuEZ8oY6ga6mBp3xhrmTBAKG4Oo7qUDyi
bN17vHvwlyH78d5Ibn8cgQ6LTWwHkIMICFWfL/Pr90EQp/74FJKUXZupnqaXI/kc
+dJZUtyhk/DrKqCQ+2zCq3sG6njyC1Z3hjH+/A5OthxonU1Y8m/BJ6t7fobn42UC
fkhFIryPGic2SNQZA6uOpnxcUd/+uCMkFGomxMA2UBXUDNRgQIh2VwATdOqsYgWt
FSWdimIKtxO3EIgY58WghOQryh/8XiBtCNIjaWwHussDsHzIOlGszYQxnOrYwPod
Ee76ouL2irs6p/Qday1w/ek9ZUinvjQuYlGVjX15SSXMfDk3JeF33DxkeIWMbzMQ
UfY6vuK0neS9wc8N9jUW+sVe57bBBuxOKGBmpoIFlvFuoJjqNlVySx/iBh/KfFgb
F3j2d0FDn/Nf2qZ3lEXxJJT916Cu7VSJui3qmp5PW0ASM4tV/uiIZ3JJ5OrBCeFa
cbLtoaVvWFeTk6SeNQTBKR1Gk6Sj/abV6OlklxHRYNlurEKfbcd/AraZoH2ntUVR
2zclnWcMxtqG1pCcX62fPBZWnUr2D+IH7t8HNSEsuInZDuEs1GaVT2rjfozu+Dvo
rxLCnQQHcalyA4J4pl5AnV0QQFhv/U6D44/mKjJ+idS6Q4Xc5GbFZ+Re0u1cJ5zy
OuDPYpdSXAeytv+c3AGxKJT4g6VtDGZJNqTot0t7DdqNFBG26wuHf9FageaExZVZ
NEWIh1RHyBN/niVDvBQFu8t2Rwv/+Je3mfdZpZ69sK6OiLQHituy4yq3WhDF146G
oEA6vk5UlNnvo2bj8dar/YviW7OA9SLnIyeUSfD0d6f6zgHDTYHqzX4Ho7orpxN2
eIOg0aKGV+XjaRzwQfxQnIfLnMvyBbHUPuouE8fE+m2Gp2LBlyzgMFFoAdPI/5mL
WrkYMVx4SCpe3tYVx8vLOemR2TNuunVtfMgXC0+7gWZsQHE+mir2AL13OQYPvAHY
WTI0HcyNt17m0TuNOF5dCt76wHq//HVlduDpVvh7wkynSTt8mfakYRtUS+4Y8pzo
fwHsCpVZ+DGNPODnMaEp/Pse+URP870WGgKZ8TfY73IalqFTEYrIRML+WSOFnJuF
SjRXgRBIW+4StLeHm/h+PxJ3usdThuHEJaS11B8Rudy5TCNOQvg0ScTVWNjJpaDQ
Vh2yIWMKl4LrCPpzO+o15SVaqqn/loDGfwLWQDmtLgpHNDiOlquKSNRt8AqppBWp
UIgPMErERhDwSYOEYJPfEfM3QnqJuyEEE7zABcono7dk+FAYdDPVOplp3ylLsRG/
7+Aelm8bBkMtVoD4x65e9Mpep5uhMN9upcsLdnI+5AcyvbybCWUxWHQqnDToMsYV
TlGK/Pd4jTe16HtirFiOa1R4ghHDFR2f+W8Q4LKTHAW7F0jnkR3/mG3gTLlcNZcG
ugj49DfCiB5xLAdmBihVxbWOFmqag2CoixxuWORTqYtobHU84CUiLfbk2k+0j7fa
cq5xFw+IS39TGCIRkG3jOi/hU+/iMP7SAG2sRsQCTgaTQbKX8N+0jRKeTzCkse8c
c5w+ZvtSZcPBs8+l69HzGvQxZRF98T5idu6MoBojqYfFTUFd9abG80et+Bx7F2Xj
ehRyP0veJdJa/fJ8XuMGWu1RSIxc8QRLjvvBv/bHcIJJvSuF6gsnz1Uqy/yADnLW
yZhW88iWUFciau2POUHNhPTwbYX1NGt+I2RN3XQCCHKTBY3YE+VHVYYG2CfJWUVB
hjv6sYzoXJC8A8ZMfvcPBUWwmEvPJ4AltMmk0myTxX2+rygqFdCHzKC0XRD2C4Dm
TPF6Qe38eOBQy8VXlHDCMxrmVw2mN/fShvRNuxW0V/j4ADQpp/wTuP4fApzW08Fa
4LsWyyI69tpJtEbBeUSM8NQ+iW891naAdJ0aa/JqV4sQGOgASTDxcoQ2kIopSPSb
iUdSFdyB3O6HfGUtMJEXAiGLpb5/TpZ2XfXH97kRFYF1oQ6J/zo/4F+ckAZrau/+
4/qxOgJJPi6XkM8HC2cuNm7sByrvfAGKaAYhlKcyC7BSnNn4JnPhsVkAqdhFRZif
jy0R2u23thEK6AT36aKF8NQic6fOECwfOexthIEeJqIFsyv+COGcbmvbUDjpJjWb
IANqXgq5NDjDXxRUU1YjNyAPwSRUxra3Q9dYR/RSpL3YeiAZgIrov/9SVoJhrFg2
jW1s+hUi/XjJijaxQMm+4HGMc6xAdPW4W+QmygsC5slj7m4kz0Gm82545UOJJPjm
MKsKzU+opdsRFlqNZq6p6Ti8VQc0kIiVfOcWah132vOi10UynfxqdwUZWFklfDbJ
FTH6GEUBG1ViIFv6wED4Te3DYgHi2GkZHrq1uiZWOMI8NE7DhsG566wvTzqDu67w
ZO6qRHvUJRUR+5B4iWUBOuHzSlZFwCckSh7QDUaF78iplcQXlyUt8JtnrvAe9kem
iq0VmdYQRFm6KXvSOrDMz96gUmLdd0Imryhl4xODmULZ2rNWFySMD+62P7oDlJhd
iPOouKPjEIBbVMNw99Vkqr/hREb9RduRoG9PxnH3ia50+5UH/X9gjUBfyqdWtm2s
CvlMi/rHl7Dl9+qoGaey+dfMhCFZI5hfb65gxc9AMeVWcFyHdcSL5UHwVmPhasYx
qi7j2JBeSGAs7NNCNSE3aL4owV0HE3AXrgQyDd0svYBbRQVj7+JsZuXAUAYmCjPI
DX6Jy75321Y7pgu+Qfl5RVEuvp56C4PT9myByKLRy1cUpDQOOJwB0Mgby8UfXMab
NWiOTNaLyJ03n5XXiDdUogWyQyXzQI3BjHqafu3/IgSEGVO5eKe/NLHWL/B/eKGx
xhcmwZg1c5sY4GBzufFi8Sv/t9Wmw0dHVdfJbpY1j/dCd3fxtJn3vQNDSDxpr+yg
3pm8fbSDBSZLGK0i3yixi4PiwQN4UM2phcqUcwISz+M4SC5LTQ3J7AZO2mSudz8G
O0uJeoFua5O4enmOcAaApLIPmC2fcpnrDiIxV/l4kSQkLgLCSIaoWkHQIX5tWMsm
nZiBm65aDvbO78wps0E47CHwU30vdA85bRXiLSRoX2H0yRMhjiWCEon5jR1hKzYR
+vld4hERBkDu7zYJ8Dnr9o6T1OlEJdmdgmCy6sLhUJSs2wdZOEKKbK9Cs+QsKkQm
yiSzegL9Rd8qLOHcj73eWgFQsAx5rXxwB2SJKazaNZ/CMEFDK5oRW6Ydbt0+D3k1
Yr/pxLkx52FJJ78/d0Zk/8WkDB1ZOLq7Cp3R8/iUYB0Y0LYIItGg9hBnRR9NyF9b
IFHMNiej02KgaXM+8K9tj9ybzlcXgv5Gtl+nwbpsmt4w9iJYwIr7QRtDrEaCP2vS
Q/RGoUF0e7mmQK8HlI9nR8fUlAj16PtpSAat44Ued092H4UhMzoQ0QtOIhlDEdGB
f0bh8MFGHE6YrFtVUhRO0Y4GqrdPFu2CefYcTWXMwqwKx1BuycMQDVj+CoFaXLR8
ogqwzMWhfxQD8h0uP7X0MOyiD7lc5lmPaeXn0i4CYSQTijZBQdwR20JK9QNTbo3n
tjOmiFsA0OSHU6gSGsqKlhXm/8ucwnodMcZBqZKElBTebpspKbGEF2kW0xfGH0fJ
u9VywN8gbdV+nrEgDU7p5efPUwDY2wMzGvxzNXJV+N+FzwpYX0iC1F+LoZo8uKUi
xWrdUETfyxGyobPaHB9nBfQRdkPe+Uovvg1NUZWpf7P7mGXE+820ly74+0Yj728c
SAnPrR0SrXtccJy6Ij28Owc/haBmnBhK5HBu/r2fb1Sse6EclqbAaycOWlnREY0x
dU8t8g9gCAsR/rl2vFLqVCF463B6rCszShTj++XFukQ8XABgC9YIDDUE3BB+tU/q
M9lzZHXG88A90lqeK7HjyiMkU1g5BG5YQwR3paga9ele9nlSwrCxVybHdec3nnM2
D+I1qSChz0Ik6Op+e5aMTtz4geJu6DlQK2p11GGDtWvOar2Fr/dLv2QdGY8m5ooN
u6VGgPj5EVl1DZ/5PM43W4+E+/GOF2RXv34HkXDk6P66uSZg5utuo+PW1JWyLWkg
wWm5CPj/FwPyNNpouXENxcVvusV5Sf8ZJIw9aYznLrbWpkjWA2lKokLwt51iq/0F
FJVSyNStxrtUBAkCfcCLnOCYCUo+diwTdqzongJtFeEt3bpgykUS4/kXrftOwkSq
AbK4uN1pEKTpnwhQUCIrMZc99FNYwfa9boxEJCfuZrSCmlmiEw3t8FwnmOl15QSv
FuMz4NICT+jg63WXoP0VvbsSOSJNtDYFBMjeaLwu2o0WGCa0c7EMaVBe1XV2zDXK
8aT21z44qaSVsbVeXW4RkuehoggKyik/Hyif/rOxsUOjyrrQECZobVp9YtBC6r8j
Cj8yU1qgdz5C710NjCYQKj4vWhIeU4rwiZEtuYScBCzobnJ/NjoUod81uqcu+EPC
mOiiubDAMs1VcSXMjySVNiqf/6siCU1sQOj7vaGQJojOuRdZsIZFRtmquJAVYJmt
Wcf1jqpD6jLXeCf7O621sbc+ZmsmnNC2ONHUgqqQWEpru+OV4kJeJ+z7kXxXohnw
v6CxI74FbA+NO/WivnBj8EgIutANIXt1g4w0V1bUUAI2YBUxuLHGdeokopNrlqQd
xkpdWQQQ6+bSTSBGAR88SneMOzmWpVs4EsZsNGi672E4IZk3qi/ZOGoyAQlgIEG4
Q8OoEQq2OmiPoFAo9RbXwq//msGx9bFCBCqXGIBOuEFJ9N5F6/wPtI9FAeu32urh
9Y5PE6j/VRoHmdYnVGkecqEJZcIZho8zorG7ONv8YBt3qF78qAO5aVX7NKXEJqhX
biWH/YBM7WLqv1QUBfmjeyvAMHelBkA7c318LkOS5zNUaWJfRW5jE66ZEdpYWgoB
234KUPshq2uXWiu4/w2OKzblqQ05raSGTwx6V2hNIT+F3obW1YSXDedoP0Ek+S4w
2ZBAVTasASm/wGhfvGOs8NSsmq/XzYVOco1f3eXjI3pSHM8A+GVJaUqd9ICUEh7e
kWgjczEOuiYiwmkvrwjS4B+ha+XeefyxqyLdoskxc31nKwEGi+FBR/P1v20FEzBF
g3Ber5QNkSehZn4gnwDu2VR82o0P2CCZgj/ERJacndxXpbdyaamdycv9SIPTGyyv
xbpc26+1HKaODrSUZuQWQfAEsBxeMAgevBldjHt2ttH7w86v9dcGNbFEchYbpfi0
t5Hpqy521R9103+zaghlEMUWT3vFs4v0FXut+0Nm1TIFyVWT9OvAckno3tapGQoC
61EpIIze6M7v63iCq4oEVz+YokFwu+E0Q1rb4OnNYlVgl1357li0AMRtFF4SHFh5
dWWFqDN2wc/Pkw+WtS12ywI3Wg6aAdSwJWXlQBPdbkbr84K+uXqoDqKKKHnsf2n8
YFWMGDiArhBUarGAcTMVH+hOldCjXQbJMLepuUy9UEfdi63fnv8RRnWd4mUUa7WS
05aw5yQB+fepDUmyzHfOqZA7CDdNaPzEmf6RDuRxjEc7hssHpbFDmSOZ6fc2JWqf
AnxJhNEKehA8d0rWM9UsZouonlsOC7K74ZB29Ka004zzctXS7P/KLKpHMaBZ8MUO
3iw5p/cuilgbOTx2KIeFQrxWRk4r3dcNs3qa3Snon/rWacmokrTY5YV7iIJwb5wm
POddY//O2/p7rP92AahT7myl/FpLJoPW/PTyeXDas6SPvjpL/N/T3OSk8anpoTLb
KVLZ8h4i6wlXUPivLeldqihkiWrpOzOY41EyqWffRwWwDkN+3z9BkmfRiSzQJVK/
E9U438/U+vhp4QhXJ8MyOaNn1zRPXDF833s3gCZSB2TDIhK0M73yYnytYCfKy76B
x45ESR4MwBD344U19tDB/qorIdPuPinQhJlxWCS5UQe7IMjRg75PWTwdrI7osMHl
YwFbMHaBLTpyHEFTLY69a8m5CCVSbhiIzt5gu8Bn1cpNcSOMLELP0k1z5KS6tsmV
1+nyIIuxcmTOQUrAj+70D9b1zSSx861zUMXp35wRGxkIryUzdQhl8OhVMtQFe5m5
X+XjwHz2OqdE8Md8Udo3GEmLQo8spLFCdW2pMUT3q/UJurtkkO5s460Dk6+SNJak
UOZG4k4xHvkpQTRAq5ERiOltIenRRcyX6Q2d0E2k5ReNvZSG3qPeoCYRYU705SzF
/ejXhYdZr/UJjvwyTImBskhe6+5tMgndkW7R/MgH5Xbm8pfitbBOA0JKiTMhd9la
h0YKFjJ97ptq1khQCjGz7YgAkTOW/nfk+qGf9ZRWWGV1jiwF3my9xyjQnYjtPIAl
AfZDfRw9mLT98P1fYFF0rMEtwVSTnDrvndbHTe3YD+93S5NVwc4l75CdRohmRtNV
J6HpJMcf+12+r+4npNr3eAfY11c5C+JeUM4vVWc2R2bBUXKqgIZCufKQtNkH64KR
xZooZ2t0/ItbAxe+TeIoTHdlhkUZUTaxN1VGNjsIxzxMmOLy8VnDIrNaSYQ82uQn
aOds2TNNZQbgbet2N5JgxrhLgR+NWikjPWD1NLMkyz8gccSxZCUNNtgqraw1zN/6
3QiGa6K8MRN8Y4D+suRFQB/3vWIE8ka96Q0ONnN0ua92zF6ZhCDoTLn9TZYGaN9k
1Ba7lvlsiEVs8f6e5xqgzQzOXwugTmPgyJ0bwUfaf8UyvXaH4UqQnlaousipk0zL
7KchDpQUTYe00mYopX9ND38wIWIWI9mhXjWRPghgwdh9sVZFyxV2ts2sVWVC9sql
U3pVos9rVXMntEdR/KXr/2WBn7AuXYFYn7KbVANxFpJQmOHieYuyr/ydwhXU6wI9
VkAT4uUmX6o5dnaPZb8h594JshfqKU2Qis4+c5rlB20TMtqX6Wj04WqxOotskoIp
6IKwWyWlj1CL4QyCrNHsr0ecJYVMPx7GWazrfYQrp9MhxhXTg0DB2zAD5kHYON2q
GsdoCfEWm9F/Dl6lhZpih/3pPQngKB00NS6WrP9gtzGTSTnreDrsYaO+6tXo4TwM
X8VSBVvEECgw678hfHk8BbeeyYhQeDRTth32k9ruPJvhqVQPcqIy948NrDeEGsDD
ZhmLILyvrPrreCYLoLWd+Opqi7G2tCnIVK/oshGmA7Amvti3zbBveiBX04ZXJkD5
JfE6v9za/TaObcMX98OsbkZb97efbQ5wA3la8Lcb2/7rle7RIgS02dduLuf8mp20
AZ/hOGnDPXL0yh/D4UuVXbAipwF7viJ0W91/s5imTxRp5fOwEo6zeDJo+8ObkSXS
RBeX/tOEiqc1fBSwxXXnMDsx42M4Hj+BaCXDY99flMqWQ0viTSxKLNPzAMXPSU0R
hAwdG/5lMO/zRBAveEpDqcV1KazSxnQ49D2BnS3cGby/WiA71OBoSf8RKMNdpmHK
Bk18bmHMrsq1ptnGru2zwpoFx1Dnh/Kmb/Bpl5qcAJf/QmLToEeuk5go1MtB/s0u
1LUgLKR+WWHrP+3v802njmEaaoF+AWYx6HbxBtIOhDoo5FeoGggT4w0mtPFDtoOj
ZAjOqBua4PxKwswWjk/YPMyGHMSXtdb6CYLPMgCulv0JlkVHKKGESAsj+lFhvHF3
Im3gty+kwoE+4Opt/oF9j6wYMAHPiyPDPCw8oCGccOICafPfQCDMMVaE00f/z62a
wwCO0R8j/LjYcppdYBmWBiW4PArezeqB0qwFvp5e+HYeRLFLWNRAN5C4zihMeVjW
wtuB/AhSb8//mhxdanRsV41/pPuWURQgi46QY6GxkqhBabT8pLuX48ApQhJnWNJn
K/NZEUdDmdHQChVIcFCf5PYva9bwrrPt3eZIykYrSAqnUbiVxlSSe5mVAEk8IOV4
CAnQrvxqhKKtc7uPcKjLrnXooififftb+bbIlFtotC7deyVwcxKGoOfo6Qxfnzqq
lyCEIDYrE9Xxmu6pKEGCBjb8xZZOrVcVD1jl1NJKzHNtIblIAiSWzGYCm1m+MK4j
Ff5Bguj8pMRjsKjYIxO8RVtfmKfhKzNFAu0/FhOiJIta6qxlY5qDlk04od3KGmV+
GiKrit2E+20Yr60BhJusvIF/bjUrYitaXYjBP2RQke6ahouwGd20SdnLHr0wyQ7V
ut1WTKZJAWDcjGF7tTLQN8Bk4nN1D1VRAyZh5F54Z3MpzQ3VMla9veh2o9+i5BAb
YeRDZWcWyF8cmwXzpuFTB8UaZCSpk+gXJoCrKSs71ROfWZHY0VZC3KjimiDaSn01
J4IDDNR3MIbr11Twm7VH3z8sh2xArkRQ05M5kzNkZN8VyVhgTO7zFv6zkWsRl8Oc
uCRLZ9/LiAW9RhV1XhYz1zcWdOm+O23B4lqPyJTkDpFV8IXXyZLWMIPdwdh92qe5
6arAgcUu4+udoP64gCPT8LXiU6oYdWx/KDjd3jW51Ahk1YSoCRASUHt8wJwXk2AK
pN09ZSy0JCOW7AZGJJO+4h/RJTSJYPpIg/353IGlbEBF3rWsSUy+96x0q0PMPkul
0MKcL2VCjAAr7TpdtGyf/7Y9YjEj4aq9vZxjs8BQvnmpfdfSv4VPtrlw5sgfcZmi
5NaTXtkp7fx5wqefhBpvkegob3EnJGpxBPIUFn3x2RePUDv4heBK6QkunMan0Gbf
2rez5tEm5qPoSb1ZYM1lKbDuXUVYtgt/8B52qrkN9IvyhzUMC9m4Hv/q/b+6IkGm
KhRj7IZV47foDRT69O+zMSSTCQDLSSb/0UiBO5RT0/7+L0Wr3F+eX7HsMSVbLryo
FH2zRrVYFGnD8Mbb93MeFOqsK7c7tgS3btm5iiC0KybHYPnopWOYjqRnrJn/IKhm
Fi/XCzQ8PUiCvT7CZ7eNpmWDxNE+XgO+szlhPGs+CEEkdI2glGffi3FVwgYw35G5
yKOMTLOp/A67bEDaxA7yO9v9RCElV42+PdR/8lCoFOUQh0nZNFzyerLNfG8Ndjr+
2ST+2Cwf2K0zeX9rDlhySqBMoS07/tRU+nfn4jdG/1adKdXCg0U4Q8OmkgTYJqHi
toqeThV73WoF1JcCcROwJPHxwMUhgO52KiKsQ+2INPfhJSsjEQVYU9iFT6CeT4gg
/y6mLghdrDhATEmvPxZ7k/NErqTSN0bRWzs8CuXNHLztnQiN7jBAsFjAPhjDlkKC
3XK2rOu9JhjZy1s7KpIzr2FsslfI8yaehVU5dZ6Sc9GbsRiH1Yo6kGSjMV7HeqMA
wlsuBsAU7KWfpp4obzxOSu42p8ufSIOThNuNDyMAn8UMxz6A/tESgUwbmkTaMSyR
VQIjoyI5lMJyvOVbllKDJ1vpcAyo/JdMnxM/MgppI0lWgC5b/hLXITcMkim9/Gwn
FWwXJSdZlflNXMP6l7dBVAT//TqdFhn8rSA2FpKagRfuidUATSPIPn3aFrv3yDWg
Fp3uR94sm1N505yIRmtxQ/rD5Fo3d+9hrM/TyV7YBtHZhyr2rzOZyItXqT4+VTs0
g2qM29hoJhpBtBh1UOiIhp1hvkEICgbXewRVDuuyIBb+UOOhSNNyaUp+LkieGpPn
Zpa0/gkSuhLp/IcpSWPXKv6WirIeL89g7or+PD2VOY921TXPBkvaDuFVCiO43vg1
827R1mMOlj06FoGc0cbbxKAF4Hj2FOeZRa+GG6KO7TnlRu2KtRfrEeFEaM8hyoFt
kA9mc9+M4EgZCcFYrVR3QTgTqTUMExk/0QLUZMBfE3SQb23u7IzyFx74pR1ShT3/
KBuELSHGEClJJAGcGQQ9Vy4jzgXmDS/emgnylmQNcf6Zm2XhDhN5Di4FO5B59mIF
jYotaI+f8Gl7Y4FpwjJvrFz8jN1n1GV5nVKFZUaWh551a9mQPUdXq5zgJncpuqma
qOThRoqFFVfOSwKeCOY/NRobK8P7ka1gcOH+FIBOaMD+w6y17olNwABMOMmHVjSQ
6d2qZs/Bjz8cW+iXusEsbwkY9vf0vLB7v+t7H3mGsoT1tgn2hipiBrJOATRcbzN1
Cf2jih9saOtMfOzlhCJgU+kq+JmRHpHUuytMYgn/nZ/iEXxHpZCLoDCP8qIQIAma
RG5Z3K7OFi/iF7t7jEFFyTIQ8OTGVeynd8mYh20NhHL/2GBDQYYu0mqwKop/04bq
CELjbqdnQ8jAVAcHnqXnwyJMwI8qnsHfL0avolbk00+LvTcFV+A9hS8HgEXQuepG
HtaFYThfyiG9RDrzzgI+4xYos9l4wVUn2xcQireGp7uE7iCM+VwPwqmAaw5r6MN9
GN76vsShHRDLnXKdhNqlRYgqO9vtUQ0CM9AW8CZyINYfPnPa0RhzCy8Pc2IBmuDF
+3ok9OUaWTl2ACv+Nzw6r0smnQJsRDVrD0h4tIHpzbEy9cNm8QP6Fd+juQnqdbX2
0gx2EwWZ4120o8ZgLoO0qn/svlMBuXpkP6NRiRcOF544d17ua5l+WUMAocElJMg5
2Yed8ajG8Z46k0C4uPwhTAeG1Eqp447KkoGDNP5DF8mFgQn/KNi9iDgGMegYDZrD
0E9vDlMUB/C80vF48ZMibIYyzxRy/r6WrOISUDc2x6yeAte2+Ljk78b3Xwp2MYVC
0OC2++HnkS+OS7MLetr6+LLKyf+apcu6wG1DBHrJhokg0ZNc9DiBFXncOnh+0BtO
K+e/X3VEiZLG3PMnxvmbsOSbB3mqLAFEr9sFroCSvk/ZINe01FmKu0vqzhx5akIN
HLOaTjbA2FO+0q8i25m8+X6KWafVBI/ErqqAd1/4RAVl7Hc1JCTw0Gsks/OXkvzG
iiq4nR60Lvk4dqAfoziAZM2uwwWjALQ8cLW8lMhbB+rDPxpuVqIyaT76HsBZJgDc
HpmERiWloCCA988gH3C5+BiNbIFQ4MTIDySZFKHrZ6FrGQ2h3gj//TdJgr1DypEQ
kj0ZyBSOT3JBnUPii9+6SMv8vtiUR8FzvxqTVS0j/hWWoU0RF+cwzgGmKI6xQMXz
eibP+ZsoyxbvQe+9PWcd9q9NwgnBZ8jx0BY0FyacPtgYi3Mt2Lhh4AMergeR49np
n2eFFZh4oJjL3Zx8iUsevRC9KRfvXMp1HY0/0+6fOytExST0lGnHkFzxbwSgocwY
VaNtx366gpq658irtzymjAS20Nv8QgVSjVZGzxEaAb2josPIhfsKnAi3nuQTzPCG
mmyl4ss8pQBaJ5NG0b+Z0f8JGOf8dm3OUZMQAQOG2ozvemqEsuRMSFEQYAKcFink
6xE+1Iv2rUeTIWCInOscLDHHwuSWyglqvEMqfefzWHhx4rN0AzY3G3koO1cA2jCh
MUuAXUdHxiVDK0h6Y3fv2tRaTXXdF4FOMrPmaBQYsus8f48020qnx5nzWqZTuzpi
CLEEvvlyHXIXVtL0LEfwm9MzUiO7Urmz9y0Yjc5NBoUx7zIacOSoqA5rZ3QYsGBd
dGNP7SV6KtwXLR85QcuNABfErCTvtVK7i2jHksYOxGtDaWK+hVX9FEQwg/xf0pld
/AQtjsvgA+dVSGYovCuoqYVG7VpukwAk8Q3IH4ajH38BoBMtP45fUv6b6fgzU9cr
yEHej6ftEdSqJIkV/Itaoir2X4ZrYq2+A4tYpXxgmay0MAQjevwNs7Wdg2FfeI7B
HuYcLMpS98PJ7v67INdaYfv2UTNzd9eZhs2vtNYPZDoEW/wxLqrPUNTMu7e4ulz0
V5o/oyRjiD3CXG7QUikwMMHGR2AM+LBQLxnE6N0h+8xddVAdbs01TaDsTnpgBbtp
7/YC44Uy7vPAw1Ro+YKJj3Y2xZSQKMQyd6ISVEsD6ucMfok6785+0vAbPWZDIMYM
P312oZzfudF/FWiro8fx0cZMNudUdoPFWVlk1+XK5atyVl720zCb3VJYoEs0ozTY
D0erGqmzG/NQPjrIxGgAF6lr6c53cpCERSBNRbwOkXjA1cb3PpQGBvIulNgT7YjA
5n/+kkTqTkk4223aqhSn/ciu5VaLNy4YL8FmLeUOFKVHe7GuTMB8bWrZv2GD73ec
IQaZ9n54HxfeCyvA7XOEjnBA8PXQn9uOJ3fJLZdK01xjXlWOE2wOrrIuE+EbXj2X
VPHbd1LGXOu+U60l7i+IaOVpqYWFu5U/XswndtWrp33r6jMm7XigjqsLsmv2Ddjd
RIbr+z9pg5dnNNIx/jL87PNG6l02kNtC//qZ82v7mXLBNuAEBZdk5Bo4224LeciV
ChwdabAM7122Coh97VGf/uTDLa1/369mn+gM8VB7Spegjs6F+DMyDz/xOpnSFx/p
GhGShJhmRd24Oo+9T3hGGrxdnSX4zuAvrsuBM99OGJYC7bU2pt3vtfAEnqg8Uw7L
+5ZpTES7Vu8JQGsR1bNLIpkeq1B+99L05fhMvCx3o/4fUzSMS41R/If1MowaI3XG
JHHWGgomXKgS2rejWzbN0MQ9VdTxum/NObbTJaAhHug3Y6BdmH9vDhB3NWlZU8rY
CWtSzQmn0fKrGUSb2N3ofDbrm390kZLEDLbSmdrHuHBfngkhaP4YjdEb1M75DHqo
DWyq4YtpCbVzXfN7ttFQ/W/NSYs7T/bP7PaWffzX/1UZaQuUWhAdpC31mc7RBke5
G+k+wz/sVTRtNcu6zixvEigQ2x82wOztO7heqfNgUTX19sKz1U51tYI3jiZIn6/P
hhukJb94jGGslS1u1HWQtrhQmJh52Fmxt+Ky5zWkK+SjDLLJjfEqHJXhcz/RIeFW
MaWSVVJFP0NzFD5N59txd6TyIxt0IzRMIPN7xqrLWUDukFppMizDyT0HZeReupUB
pJdsnUqAQrx+x1HKRJ+on94znfXcbydihf8hkMN4TbKNiwjEwwKaBlJGlt8It5Af
pjX3ZatPYKKzVA0qkmrP7Kl8IFtkMiFo7iFxpzrdn4b/He8+8s4RFTi/pU9jn0x3
XmVIIomZ4rDvfMBFgmGasg+n0umesDRqwmFtpIvcjtquMsDmgGb77FuCt2EuxFyJ
ncx+2GkIoU0ldUSwZ97xrPrnd038aQuRucY/RlrSHiXmG7wHaMI2AHXmvOneA5wn
EAPKMhwCWK0Pbx9eXqBbfLSLA25mFbUOX8W8y4Z8A6dSMcDxBWqOqKT+CtMGEqp0
suMzYIW1XLFSvD1PHC08yCAOl9pJ0/1jDYDgQ8Jnei8WHlHbL7ieyMjf5Za3bhmb
eBM/NjKvMu+hkAfUUzL5PDA7H56WTvH25M6bHfYFyrTJk5+ZuoPKlqfMDB6GSBG0
owhA56MAhmkz5aU9aXMklTPaceBNu1y7XDN4ZDbbNd1HWwR67Bg66Ko6nLrYelZq
/2HrSMdtus4TFKbpiwWPrSc0QbqYY1yWySvWwIYg549Zcr6JeX+FEt+/+Dbt3lQ6
WDMFTx0FooyG06P4IlfUclvK1tJoXwcbY6FPxV/XpouBhjKujmrxnLpte1G/V3CK
dY8y14/f+91s9Bv6afxPdynQt8lMJCmnUuFYNuTBUw6IGZaZaTrSsqDQ3aOcd/Xu
lfntZrBKRaUrTcBXhNAytua+QPvQl/qbU8ko2z/56baUlAJi/IUqvd/NfmJ3Qqw1
1QG3812HZfqusmNKfV0VZjsqCPyoMyGANWlbBDZ1ily2e7ljqEbIe2s93cY31Wui
evEEEsgmXIiAu9Ft5RKdiKiuaK9PPlzNGkedF00afVjG5QKYlwQOSeokkYKZhDFo
W92XZsWtFWcmrebhlMkLVmFX1qmgruA3iZ84xepo8F2dqKkOkIwwBOaTPBNpaKw+
N/WC+Ts7Sa3QxZdX6afkDSeX6trolOryVE9IseTBGLJ+GGu143Hzx96BZzI7toe7
5r0lGf8XPv5JOFo01L0LfbHASFaM8W0mKXBdkXgddVFnJN6M5PN/SmAdGOLYJ038
hWT1rrJtlpunLJxKdOoHyzbfu8FnQs1yAeKiaz+0Wpcg7ZDGx3s7r7hNtX/eOazW
oDFh2gl4EIt/2487T+W9lMh5OZLC4PLgc0y7b2YLUo+WSiAq+0i9BaiOXSiUtrpG
h5TWL/0/u1FBySrPR39pROo2/iH2H4T1ylOJPz0fhVckYls9VPK7UvgUD2DvPb1c
Ixpzp7896BZahbS68jp9e4aD9pjvr00ssISuwx+RSiMtrup71qIhgDJ9TYXjE7e2
Rtx2M2YSpawOfdMaXrulQYHzTIMae3cZJDfAP7ntoOgiuNRN7z2cDSyyf/lqLyBu
SnI+f/TQELXrYIQXa7sg0swsYVw1DUndMlGAUHCVL00o8YdNBBFHeQyRyMZOX1xu
BeI8Ayt2IpTqEgaAARYi0lFe8fwYdHP5thoKMsFv+pdSkNEzdTBMWaqoUyiWHjzK
1Swljd+PD5WcYap7DkMiUEJHfOR6MaTbXoutIWGLSsmBbrre3kCF7KrxoBsYhpKb
6VLy47Cq7fW/OVmiJ5i1T7F67u7lWK6l+Q7PMZQwhJ/0gF49bqlYp8Mrl0DqLRkZ
JhFcmTXmW16JMYaO63l588zFwYqUV2yyhyQ8vGxwCrqhpbic5RgopCQKlnkOqiK2
ocJFgOjUrYLLRRdXMGEdkKQVzeDb0vplnu8mgquv7Ua0fqb2XWg5/dmWri8PDjBu
4lp1MviU2E51emBqY5h4+Xnnf24UjmwO4T4GY/i+A75kca9KDjliog1RWe6xOgy4
ir0WGHzQ+E7ZX8s39F6pTovlw4vLRMVScmUyZPEmtlFoldzQzUyHimI27qUC/EJN
99UVS7e9CdWMAKZUoA6vs1szmleFgRXaTZaxGn7AA/pLGoWOCjQylgtuL2yLLlH1
LpYj6q+P6iXpelRHMdhQCDJ2bAy1UY/CCMqKlChpR3FbXspVU/PvwgVQGFd0KP2m
HnK65SwomHYCrv8VpjPsBO3D/o4useLjpcfMRMO1W6aUrM5kdJuiLwpzoKrsRw5N
5vmNvMexwOkeRAJKJ55ha30mKLZKQd5eUhqpnBJ/CKjEvEIndpT+Sxv95wPW43Zd
U4ea+Z1Rj5zYObKvcqjkkDsyoFp47rFvDiY2Ztcwwh93MyeUP72Jt58NCQWhFslm
YdYp0CgBHIOk5dLkdlyIufsiAOKKu99Q7vKCCoi9rOXIhHRyMzMRooyZeTcJxo9A
nSIMbAQQs0YWj+6qt2HaU6FTi8f2YemcSflqCOu3Q+wfZ0C2aBtXgWE+rABjVzGH
M+0JE1fNMUEhxtXvAPyR2ou/6R7ROjBmm94HVwb1sT38J0DlUIpWmlQhuR2uLey6
3WQABc8WN46i3Tr3clFeHBtyOJaLlGdDX+5wDDZ9GXrSaluJJQSK1id8PUulJSA2
pCgXtWSGntgT96oEt1fQY0r8ZHXRQGMlJWAeU4zdh/ZRxPe8EQYAidLxdhwC01Ri
1ZjOE2f7I42sRebE21YEEjYdmZMybx2ZcO393RjbQJtQKtuGFzA+O1Du9cBAsu+d
0yRWSxf/RqmSBVfrSOFuNLYRQmEdYX0R60RjPEG/gGkRpuvNTcm/ZKRX3ESJnsSP
gwdVmQGRipQxsIXog29BQqDZrjSDBGnzkoqPDfMLhPs6Cf1NqZEvRcqKMC8mWLgR
5m/nUdAo6SpDHVRWXAwy2z2gBGKnzmEo2Q5FA3KTNIHLsJyRFXFCKza441a4tvAv
hcpuZkEn42x6KOsYCe7yZczYDgGvD0b5AGIV3DdsfiN8/Zk2+ZKcSm9MXNUV3LLW
Jl/R/tpyqw5kIAGNiyO6a33vnDyWbOoSD9rIVwAt0K4CMlLC/s+abq9ySHQvCVzm
6FZubIdBX8mpUzH8wDQm4rb2TGbnzH9/QGnt9wk+i62/8lEXvm1QtfrrFXcAB5Xk
FqRP2WGe3GPbMQVJNCuTRdZ81t4oln6Vz84TGke+W825O5copFv1IMMvqmPKAtTH
ovmIkSeb+1XNgPeeONavT9i4gxQKEucjfC3rr9rfKyTgv6qURlMVCyG0hOcmOv9D
pv+j5ggXbEnLi8jSNnoHWLezMVIEoERSCmC9f1DFgC4FkNyApKwqaBo+MAzLY2yP
rCCSqFt2ecIyiA7Ub4XgMfREi/fTwwqxXasgGx+30ZTpSNbLGVUf0iAgi/oZQj/x
oEspP+gIeadQEa3B8da9Oz/pbGcPToK4MmVnh0o79cnLh4Ow/Z1EgIPF6oAEnSi7
4EvD8/zgkb9CUEFnZzTyqcgJUSbmuLe9rYNe12rsAo4L6d/EXmnBYnQUZ/pIRSPe
EnCk7XfWDfFmrS9VFP1YwxxfSbyaj4Jq7FkrcBxeCOOlxwrkyGdUbAigpsE4F88W
DkHAZWz1EhdFL3XEYY0I1DsTMO5Wi+X8CEU33fyBmRUi2pTladHwG7aW0NygYHMy
TgWN0gvwziiJXDQDNkyel1eNnBWe6fHwrPIeZfbGrRGXJLYr2+3/ghBjPo5YO2Bn
pcavMT7e7VJOV1S9SvfwAxuQ2m5fA1VnBsfuAJgOc6YqjW3/X/aD/nywSN/PSNAY
ad9RviTRQV8HShCppvdkf1DifTg8nnuK934tYI/et8grsjl4hp/tO9aPW5+8EFig
ZI0ClDGO1reACgYcs0JCzv/U2kN1s8Xwt7ZTH3eKENUjz2ZI/HmZDCgEIc/QaJW6
zGzMVyhZ4sqfN3ge4IWWqL0yZaOxkHspzqRgbXmM9CrLx11QV4k1Jk0RY/EPpkHP
heupr/h5zMg+DQLJJM1seQsi673ITE1JHQe0+m+2WCexWJAuI6M81DHgDhHtb+vC
+5SBafndaoO3qV9X4l1SuhazRQPjAQp2I5Lclv4/4ebzfRXt4N+IwDwp8oOzdZzn
DHCYl2iF6azTy+a0ymqcVzjaKvNF/SQGVcKrR/nG3RTYtHjV2cOulzlBOigJGras
PmiFWHUKqBC6htVz98fZvQKjGw1goBaUWvFC+hn6J7IspfhosV1XymTAJq0stEsx
IL7jxe1Q08ZmCT4ETDDQx2587Bc8oULMDsswllDqDKagelvlJ+c6H7f1taJb2zum
V1gyOe2L05T0lAcu1Ghb3RQOUm/Z5IHxCdK7QvXUR5m9MqGAT7LxgZaRiaQmslsZ
8P9gkiVASlYLR9UrP6+JQDI9ytLfyOa2vAzt386Fa01WTuQX3QO5+zibDPHaBMQS
96I709qfSpwHnGbRy9EWdWRBVHP2kNAsuodAM3HgEF03cgnFnOJERsIqZTt05Ziv
nIC+RIllTnEPzNTZ8eSXFxcQrBZKkyFHYA+jWPHATbeiXY41JLwVFBZ6kFserHiS
uF4CHN3agUGpm5DMeEJjBFJo/XrayIBAWkCLfFWkGxIn8YNqC6dRVV2XrlhoQEWi
/ibh8Y0Q+FMuZy+Pz6s+Z+ioG4eIk93XrxYdDiCKRZ3zVt1Zju8oxipi1ralCXDH
xAuMnAbSayf4gYdWQq22cqSzbmxdkUWxiqU5Bs8zg3LU9PgyeoDO1ZBs97O4IfJr
86eG8sz78fdibYtP9QrS3w+/oMtkWpDHNP61iAL2ksNbR5YRRF8dCmX/3bG57+8s
SdXSVdJR8CfE3es9M6oPTdfiRGXpRhK935mAAOA1awCroSyasxMrBOQz3orDVy7M
IfjM9DVHAhGKm5Nys5qTg0teXxCs9LHZ/w1a9V0Y1ikczd8ANzKD3e3n0E8j6k3Y
tz4kVCPH3wBh9w0memSwtXHgaIUX45X1AzC5A9e8/1qAxzBZwxaGojmNoYkwOqRr
fHRI4TdeNpifJLDKHJqMlvVJjlvceaPLhlf/Qn0EexK1UotBQKGmXbTnqKltrWDv
WEVrf83906L8DnRygeol5GLA1cYJTIQPGVORVuz9CnFreyJ3wZbjdGZxEeXiLJlV
VJPuDJNXeAkHuABWmhzD8UDjW90OjOQnVhzYtrix+GM1AV8BJdOfNahUdohPE4ns
CwErZxIngk2DpMsltAgEbTULsVSP5624Zd37hym88f5v7GRL1KoveSQ+vquPldFd
uprEUcmOS41et0Lf6JOul0XtxdQHvAZWnkCv80gR/7cYoL82aUNdYjzoFf4eU9Ey
jSqmxaCD7muhFANsfij0h3y4kWVO7RenjJ3NFewe2cbh1YFwq9rrccOcOWOeDxtK
EoY+bwLukSUHAz2koheeVTUFHul240cF0A//n68hkqNNwqf8EqzJe4Tmvythgl1Z
puJ6rqFzpSKtZ/VFEWY6Z2cRlvfLVbHqObORO1Ekh6nlADNnRF81W6e6lc/CZin+
Y+QK7Nh/LkQdM42hbAYHG8RdC4JDkfpmVyOyd245hSrRVmIDasT+AD/8AvGuUd3X
f8oC2UfrnU1Eyzyr9TsJNLaz2VUQOZxXIJ57brG03hAjm/GeS0L10+92ILghVf8Y
dvv7kWzLPdGKJ4VDH+E1+xKwyAQlmN3aa1/S8vmb0I8U55cYIq7odBlWzwZuD2BY
UvSFWTCZryZ9MPO5eqj74AEEsqPRz61YIlbyzVwuCxVlIb9HLDX282fI/+JDxhen
+fhdoFqRpeXZDV4z/lUDdXONfW8F9ZPZF8qdJriGjzsLzWI9wgm1uYPW/zOloQ6V
+RwiVwtnD77EXrBLQ6f7GN/DTyY98hAsG46UrXqvU4qUBjuhYrZtMfhN1Et1ZTF3
pxHhaLaba9oOcyGN3JS3/IRyAbCNjQ5bgAaA2ETU6pvTvq4FSaouEQ9FfcvDK7qd
OXl09PUmkRhOEHlZtcTxiFMO457TkY0+0k5YbiJu6fX5CNdsDkPLHyB+AuRZJywD
WLYcg75X7CEWK0hxpCBXqICX5UI1dRdZk16nb3J51aqUdxOj61HGYxigmqpvum4d
K0sv6fYQorVuVGTPXiP/mVoEBzVMU5bPJy52za3iUZ2zYb18BTaaOt/pM58onGqf
EmuvDNgw1uVaYvdIrXaYdL3K0KIhhPbITJus30GnAk6nDr8O6oxW2gutXzTAFRjL
6hb8LAdV+k0hY+hmHF5eLu3GlNmW8NJe+A4uJOAdkK8br7G3trA7L+Fqm5MewAi8
8bK3LVbNgPykHKrO3gVYFTIEmNBKiTO6tiwIdPKv85Qsmry0Rmg4uFu50RFubkSR
8Y9TPOXgab50isDnVYOQ2/X0j4LtR8fj55nuHVkthxZCtgRzfn+i+IbMUvu8jsKB
p6DA6qIvAjOJ5Ip5tSP0z6BrQmd12dmQgrD8wjJEM4g59tBZRzAovnAQbiL3AkM4
bPrJYP2IGXc56SRrHZOE1F/o6XGVaWkRtmVwYfm9fyzMwoLKMnrcxfG+dslRrrHe
TYIaZLrJ2iXyUMH+cg9Nn4dT7+GcFzcIuL5P1fPdhhQubKWdegHe/s1esZTMLpgt
AOwQpoRCYVQfE6ie/h4JD2de+Hk6HPGTukgtkzICO4vnV7/t6rwx/u/56bg3ayAl
Dc/E71jlccOUXe+Euu+wTAmkhxldcP5FiNiDf7bgkahTZFsa38hMTFzonr/OsHRC
dZ5GrgTxc2HrK0ZdUfnCTs9aG3FpdJcCoF//omlRXCrA8/j/NlEC+ER//dx9+F1L
u+A4WWLoFP+WHKG+rEc7i+sUGYgGj7yJfM+jFvSU8WMSLhase+lELJJqD0wTsnoH
2f3V+NNpC6iXNjZbx/DTvV8/YZsiRgiF+6NuNLe/212qIGtAydsE4UxX0237QQfG
Rv5qjuir+njCsuktRiUkd85RMIyzWA7H1quO3Ym1x3rJDWOSmHErc9Q/fgQ9yXRn
d870OLO9bRR29mhQnCnaQTq9q6sZX9fIxfVRYVgW75DycCZ2rUmVeiBh6SqVnoQb
IIEXWuIKMeJceOBWJVmDah55bcRMQuDuhY0R+IkIT7JAV9VWKvUmFeaI2EbBaFUM
mNxO25oFepyRtsIPtlIjcLGhFcs3RPum+rqulBGoJuUlC4H/2qHGMqGvLiSVmRW4
XKMewzdT1SWftKytm9gEVFT2BPYRdLtZSjaMVwUid3S+Aql6dB1pwxezDz19kvmr
rk0zV2v1ENkIA1efORrjp2Lwhh/EIQ8Fe0ElD2tbJNckYuEEUW0CuxLCWA1sbYV6
cP7kNRg76DGEnnAB0C55R3mtoHcdxpp8d7y1tx3Rxjpih1RIzZRsGWyQr5gJ4V/q
D997yJTosJVQqJuL+nDSpvjbC5nH0woAh7uecByZPqcmrSDhAz1ZxtdtV31tJjF4
hvJudOU5ZaM8+bUIVuu5DBdXVFH990Y3KjD/t81uSP7WGRWGF2x9472nTt+6DdC6
0fdUUiatFdmthcNRbNib46M/ty0IL1kLuATeT9pMx62C/pfq2E1cYgelcSqTlrE/
1Ig51jyc33cRTqTFw9U0cIb0R5m6hQTn5k2stXodb+CE98ZzzTvHIblHZu01ytqF
u2ylLeWOj+KI+F+g8Oj4KJXuHtnrxOUflo2GSgQTLNUaUdWfv+LufEjHT/jwK4I9
pFaqgukRkmFdbdFj6HTDse60FYdpVG+DZekbOB2QDFru106Td+6NGS3CV4M2Px4P
6uzUoyWHUPebfvm/dSY26bQxl+R6MAMiqa45wIj19E3rCjEFqTTAUcS1nFxWTxHH
+kQevFby5VTi/uoaJoM+z7dwzabgIbRSOlxkJ1ylCAHq3IPmeF7S9IFfTeahD+Jh
Ie+A2Pv1P2MJyhyTTp9JQhIASnq70rDe01AnaVePi9surQPTgFwq/0+w9jxptNWc
OWlMdn7t2MjKBPgxZceTiGWTvRN9/dchr/jgvS19vSKXDnSqz/qxEBf3ssZHYPs/
qOPLd9g85K3xRlw+auEZqN9VZ+BoO8csTpdtZuCilZUhZLdkNVPGt9VkHOYeyPLJ
AwFlJoe7UApqy1fvjS+NAydDSqiDE+euLFc0B6hcuKQtwPu3Ikdz2HN3yEG/Bvf9
mzvR0MO5HfzHBbjwLrpADwfE2a9WsJ4Gg6T2KY2/lkofOBC9IGp4pJ7/dM5afGbQ
fQ7R4V1FEepnZeWtkM44enoJIKgK7DID/acL3naKWfLzHIk9dxJD3Awpp1nsJTN+
ZUPrAnqucAC0Ne3xWqEe+VzVmJgEJuOQMPH3Cm+AN8CI7UDOcvsU+CDp/VBjPAi6
RxdbN/P3x58jfMTaTr69yKz4VbHomoHJNLo1XiYDHq6wjYhT0gow45IQ5QCo4y8Q
fgl9FcwonDDkyRZfq2mUkPkXv8js079bVz1n00tKoktz0mdKjM6DZm6w/RiVF6yl
dRsoTkkzGGYh84dLA7hJVEYtzTk3qurd6hw9YeP5yS0u2FOcTc/Mh9xJar1rerBg
ksvvp+rKhtKBFVnkksmoIyeZgAsXsiY9j9pWmOi4jPjsZaeQtuHt41YFN4FJb/7G
fLZP4tb/M373juqZ7Ov5wOlD3CU74a2/0MSkZDjfKJhyGfoJIRLckxnWpUEd12PD
mr6sJV0jnbamJK0V01HRffIMgai8v8kbx35t9iib50CTMV/CXFwTw2C0yMXDcy/y
CB/yLeaOg4SHs4RWU0PmPmT/2MAiAu09f3jSUGPvjuAnUnQKwTJwIXLYYHHsTlQO
5SBMisFC6uFBH+bbsesmAq408pBduOZZcfMBl0MK5hrgC0z61b7ORgqR9Jqqz2j5
bHbu52AUl0Zgxxys1+ycI44FfqKY9eKs3m7OHR+hK2kbsZvd8EnWkUuwPLHhoq6p
bhmQSLRTuGxTisWY4Z/tZcWbOH4x+fKGjvO4U8a5loXsxyoGZWjJlalhJ4v8qUcQ
Leh8mR2hOozQM00DwdaDyyFbiSeozB1yhVQX6exZqhzTgmKknwOsMat6MMcV44lp
sjEIYDzBhCc7nvgOaWml9OYpL60PbGw1GnxTIgykmqyRqGZzcN68lR55T00CDrrY
DxSX7f2+pv7N5nyD1qdsCK85uOBd3kUOZn5BHLwKF5IY7xHGagcHroHhLKI1rgrk
Y81a+jYd6nLlzVLQavgoDl2GLkh/fqQ27czNLikD+RO0ghb9HpUnao7XZaeqVUVq
F+A5ukGuG8V87dMWrUs6S1GZ8upKwegBvXULA/hjQIMWsM18jzez5Ay4GTNm3XoU
6nHNcLlieTKELboz3BxQiPKxWiG16INpCnTogT+9oz2QEQHThazBFDWGe1wxVIi9
x4bYEjMhgqrZsv6sRev+977Rz2ODJDCu99aX/muWeZ1Lxs+E2baWRTpfE7l/oy3H
1VWhPSjD1197pnASdE5wdhBQm9IO2aYL7yvLCCqCKSxHojg7gE6OdcN/94gfwdF+
ujFsEHd0jvHrj7pft3a2RBdLhNUAvW0Y3e7XpFpFd5AeDNgqISdsN0tRbTWFZ2zV
hCpwzJnQfDuM9PWPPL8fK1XAcirxAVwNyR9TkUba8qX7CGz/xoJ9moeDYOn63Ba1
9xTCoHC1H0fYmRXIfVlxRfhdEJE3bZgIyMA34R/AAOguUoYZ8wMvVv8ewsDzBTlL
3I7+zZMYgjL+O87Z+5/9kbS96dk7SgDiPohffdm0asnLDWN17Ya/psPdbQQHMFZM
j9YVFqWNNX6jY6+NI8DhaAPUUT0T8YnMgDj/0ZrEuaT1XMBA8IzivxFsJ2K5Loq9
nBEpM/aujQSdhT2ezLN6syFixuHmeKXQIxoThTdbI3bSzhp/nK83EjGb/ONbnANL
wNDS7Fy8l6QYhnOXzEN2o0LtQQHGVDsV4AfEXQ1bBeoIMYLc//WbeHoJASmpQpZ4
zWTF/B10BHM9UoflIsyz6wzmsxtyXpTayRl/G8T9EZPK4DhV5o+j4lnDznsj9FR4
4RYDFcPWJ+/JY9okppq3En7TDyF4eyOIVxjpgvvlWkLNL3m+wkQs88I+D2fkCIna
qhtcrmKmK1EaGU15QoSv+lo2pzCWDxMG3hQHfuoQqUq0pAKd+UumgadtYfEVrjlt
7eiad/Jd9OVBQT0mbNRYxLfv4UzzdWLlXkJ+bsZDcYGMzBS632JNSgzPvyyVzihp
m77HXVuh/4qRd+FcLk22c/25YBxirYarX+lAqC6HOJZr79KVyO/XfWymaQn6tTPe
/PNfG4Xhx46U9aIDuW6/7dTj4WdJUvDWoJh2HOxs4eU38qGdFKRrWRLwlVrzu5wF
FByDZiqSUCNnrWeqk9ugcnBqtC7JCZEglqWS1AtOGRfzVwh35z6opXiyGww+0SGn
bEBjXDA2jtG0wrBtY5eA7tkk0TXnqtTrIpnU29/zgIHYGf8xjy6yr0hiI9ZT98ls
JiiyN21xpP0t2oPlTdD8Pnr20xtX04WZLJMxaoLvuDhrETn2ZOZm258JGgHIfjS2
yaxf96se68zUdRJ4CDFIhov+4kmQQTp1rJ7WslSPBiNndpcithc3meuVkZKYjl+u
64gjwsC0cSbxM1wQRM/qKaokeywCEQaJhwwnfPEpITS9LRpNh2lxoB8Calf5jBK+
JafAGiRVmlZy/thJJ+NMdjZem2uY7EC6aN43On6fJIrzlzP6c3j9m0YiQ5bdOaIp
7W308CfVkp1Su8KEdIs+6fqnlwOEKCJ+fapKtxIQR0mfRA24LdrC2tY1Ygf+JCLg
afSfAtu/TXEkKJtE2ITYYn7sj4T9EYclrtak1ri3WPn9uLg2+xQd4N1UNSDpr5OS
suvv+i1z2Gib/FIKUIQYzJbBepXP4rc5Ue6epj5Sb6wnOnMbyT5MwJQUwt/TUBR7
ADefBpUE+QZb+iv2bS79S+yeoFvkNt9bjDceO9TPYf7Fbd0SppevlugVp/ljNUFt
MCA4aCtEe/21YTyR2B4yo1R1Ne+vmFMXyHK2+x+vMugbcS8GE0oUVzVaQaAx4O7C
a96GZwuiWhy9JYwplAwtI//u2QlcdNhiOVA9qaNQUF6Rah+pYVCa/CVt006JB6sd
MHCAFisUCMr5ga1xWWNKftyrCx0MO/m7SKdTDkCoPaHnqa4IVTsBoJ79WtpA0hss
z/Erqh4EUZ+6RslEKUNXp8q0QWOVPRRmcU7+f/53/JvzBZDuP+7cA4/4G8RaGr1H
0ZsJxMNUxsWN+qTgfnvDRSj8AokctghZTCGA26W5kxISGPMeNnvwLTpvDuL0AKZU
QIfl6JAzVhDY5T2Mpe9K86Ij8G801o+gkRx7aKq8O8uAbKh2KWP5nwffpqT2kqEM
60icv4nmSDpQLbanoAHTniV46P10GkZJ1Eenw81GNXFQf8EkwZjy4rRjcRHpbj+H
+F64/0Pc4a0UnpkqMRhoPWQMR8glu3wDtLKtd0ukGKGo+9DMCT/p0OEYLbuDoim/
v6BuR6EDDm2cWu6xUHfPVbA2pKuYl01lgaMno17yREyywaLoxXcamHZDkx9Q/yF9
VgwpDH/9BuFRE6+gswLAUQ2W/K3/jaa7zGP4jQ3XjtQCX3ZjRCz9eqdx+G6YYHqe
Ao6s10nj/4eQcsRBTEtQ5ifeZLKGOQVQ4fE90uDdYnzFKPXDRLtz31ZWcMJvmKh5
TtV8EqI188xPYdDOHdhkJcNH4YkBnY612DaErPnWwXuPK7m6izrFJTcQi6eTYtZP
dSM+x3gcA355JlEG9zFQK9hAEcGjYI5EI43OZgW/d+1KJ5ivfLYvTCOZnRjrImCM
hOHlH0KMpxn5dWL13DwvmDBxNtLTSYAmcXCulYAfgIPOUGt3ge43XxSduPzE95cm
2VQePe2Wnbkg+8PLHWF5XLquSL2hDbvbLqr9acaKOz9lkiQeDJo8gIx/2UU1EBMJ
DTtN1UevasiXWy1nj62yHVdMVauRZFhgjGqEomVCrUMuqzmnSrc12ajDBnr/uEOp
i7V3fW12wQSWsE2Brk3VxXUUNJSmQmTLAkNwNm/kUh52YBAVJDNRr+YtIFbPW+i2
2NknDHjwkV/0ImJ20kGQONHU/0V2EcJKRWs+Je7mMhVfqmxPfTfTMF7mpqnBMvp8
6Sud5REBqnKA8aqqP85VT8fMyoK2d8Q0LmEjlxPYVRw5ktjv1nl/taKWSCplHWIY
7ibJ5NadCviRDR3gsTjvFe7vopuo72JV1tgIhRSdAH77+PA9VE70pMojI2BXy9RA
7/TtVpjv1IDOz/nQftlNyAZxsANylbWSubY1fb0a3EIcBO6TqvpB2IHoxUp+bFNa
kX9EWy6mUEZUOQW6+1eLmizMjGyvG3bdo8rKZ+vPx5OvltDn8vsYKzfLBEGvbx9s
092/vkLqJn1MmRStJ38X2/BrnV2elxyXMhjTGZO1/cLKsxMMBfLL7tFfxt+4nlxS
w5R2SCJxvnQeBdKDlHrGI8W4FonMhtqx47c0xSBxL4SHGBZXSZGiSCBt0pwMKKBN
T8ocPHT1rBfrV36FVPnbrQeMyEVtMG+hUOJMxl3x8akHKQEOvmM+TPgd+LZmBRWp
rZ7P92mR+kSHZzay+dop41tLUczasQXhH7PH+Iv9Idq0AiKJS1kNSUhXdg89836n
UIgaw5QqwYAvYqO5Xsgdwgly+SOJn1UXR92dNteFuQefCz68IIdWZBrbhUYxWI7+
aNHZCJIipH15/Ibj4D8t73wp3bc5TNbbBElWErfPZB2aneQLXfklL0ZJVrWcsF70
bl1PEx9b9xk+6F9FRQBKNw7hotBESg6SUBKW7Z9ON/k4IRy0+afs2KLTPNTh8bry
rzl8l3mY6QarlGBKiyy/7y4yXI9N0DIrNSTiDkWRiIGYXDRTUc9Mm6MrwjLuuqTN
6JFrKvMIYW2M4SU4rDxbnBps3JiA5WA1PK/+TXPvQPlLHPggeGDKK7kPN9mCdurV
OpK1wHnC7uPT43Ijll0pLEHdbcXTI8e36DRRi09XVaaEBZNmN/xsjeMLtQ6IGqXD
Rca5uMKN9ru+MmEwyDIAbykechSaEgCTmcZWrsjUkcj8l/NG1ux8XOo/X8wXfOlv
A0Q/qV+BUkl7pFJNGm0ICWLDdrhBs5vtos3V7fzRFbQQqA4mUk2JQwN9svUFq2u8
gxDuo1ZlgXDTWOZOHI3lIbCzp6kg/wiCrrDU2vGklYK9uODdhfpAuNNPf9dCGhX+
oJ1+jptwo9v3oVIxiCS5DRmRoNH6ngydJvj90rLDPDPMc9FPgoPIgYC2fSBJIWq+
g8pdnfqhKgpvpYtoNn+Ivp4PWSt1fY2UAHZrku62vjBfFNbB5aqsacu+sTxjCXUO
wdU9ScIVGiRZ65MsI0gVgcsivcu9rdd7+UaZrSv7z5ZYdRYzxrAPHA93AhYsNaeG
F9mj6f1T5n2tbmqFHOCwvtWPphEHnsbMDadwJIlP5jCoH9HYy1jTZdhgo6jRKE1V
ym0tjpeYUzqte5EwEOfbLfbQS7MsKNuZcAZQlwrf9qLXw5LM5NexsndSxFZm/D3w
aYEYt5eRZ6+AylheGgs7P1aKzL40DcWuHiRzs1ud2YQrUNShhkarWk852kWXgwZJ
UvWWsNrpRsXe6ItyJVcTtgVVZu0xYZznyYjm/SLl8R4rOtdXHucwO0eSFhjxBqx5
hncP0Yc9XTzBaF699mGMy6IE9smUdWVMzdsmzPsIy/GdMVEi6Qo0Zp9jE6YGnsTa
qNNhCIXILE/CjRVP9qQPXzOMecMuCarjJDWKqdrTLVEYUaVxwZGhd212EmbOQNzn
fhC6H+stn7MIY/EDq7m+fXOtAP/ZHZmgeR7dkO9OLpKaoJrMWN/XpetQurYrboWP
lvGPXN7J+9pF+GGja/Fg0mtGlQK8DRs5Iu8CD/wzG2HjcrRX0yyoNjtnHqS7a7b5
83ASEVoDzhesMhI5RN2kc9+JhcnF5AvPH7KDFXMcPkE+uv7zWzIi7JHc8fYwDbkh
7ph5/XQ8knGQXEfOCBK/QS6Mi/XBpDz84orSH0K6IoNOiM9bn2z5gDDYMZvnSaun
rierKevxzrC07A1Rqy+NXF5ZGFZzBegAfD3W2SAAC/cgW77CYrp5tf39a5Tae1P6
teJJ3QCHO9wq9dlwyZRhXDjVDrb54wwdGjUh90khxaaxOQknKnshfKDfJkRLVHPA
e53Lfl73tsy7sfWqMG+gMsUBUFEPtfEUHgWRm5wQDa0PsOO6wN2DrcRXN35lS1sd
T7kGjg0hTJT5kTzTolfR8ipNRxNr2jV9oO84VXWG2wFcX8pyzBmmIuM9FHjvO/jh
eDL4IBysq2jg5Mc4e8h25th752vr0PxqqkPNJS7ViGM5/lH8cSqBeiV0CM4NRI//
iBaRUpW2eiZJQpiOYDEEt2f+C7YXqJLpBGjB3NMmA8DAoX1/gXIAmct6+BYwLcpP
P/oAPjbrwtloGNKRBNK0FTeudaqxF++/gp6LjJ1o8z3jrx/DUUrPKxuZerPaP+7b
uGTBHkTO+RijCEEQvlh0nzM4X8eNgNZNaOvlPXV2VrP+z68JJNLp8J1WgOlpshXt
58Ljhg+37b8CBl3KpRbXptR6HcZM7M/m561oDToSvR0j66h861oxUmVfj4xPEwNf
IDxluDffyeOL3AbXuofSnnY5KKFrZqanzBGOt/8hN/3kJaz90BXbBO1w0aaHvPd0
5Kwu59mtPsfLpDhpJtHhI08kIgUJ8Av+eiqJmE6MGkWVUFz3xBtAkI6unrOfzSY7
fJyGgFsIaY2DubLZit10UJedvz92wWLxRzHWCVyABml//e2LI7CSgBs3ld5qAS8B
+WCpD8TOdrkGhaCHvwbg4fzKQluieN/xn20Ahm373Hg9l2usOn8CLyabJWLqVXIa
zTUijceYMIRXmSETLvsRS7nirH22P6VCEwhU+moyqv71YLQzPa5aC/b61AxgpSc2
EDKe6qijU0ZBoxnS8EHmdaqrHxS0ajjNFaPZQWMmkVYx3e0jOwNq2eveXplu7i7Z
9q2L4bQsb7lZy6K4z/Vm+IKZw5iqDw9llb302FkWCYcYLrwQILY8MZvdVTA3/gbD
AoXJJ9Ks478TlYu5lSv/WAYq/Pp4589u01lMXUD371LK3KG1zflR3XOBdklfpDvT
erNXYJnBi79tjFaw43//a48hE6O3CPepP0idZ34S7OJzeKo6dkKzaUDSNkd4UfuR
PFbdgIto7ftKto/auh6z2+tUvwrafTiPbKQdBA3zEbDpMwSDmQflcazy0T/7kWI5
cpmqq/KbsM0IKKKPecaWK5O+8PORldxq8qbOp43f8C2ON7FAozQMQq+T9ye2F3DY
iyxpuXQHQ+aK5kMNIaSP/KpC1Mm4aBLbn9tffOeF2zDlkjZmylTUoZ5aEVg+aa7w
D9bvU/VWpIokX+/fiLTsGNDYKaNmArh/F7tVxPNWII3jGWiLaDr687i15t3FD7eb
PQ91/9FZOH3vxBjqQZU+r0mDfqJBSOS8fbgccueXmaRCSx0ham8v73+7IUc3Mqoj
D4AZhjwwKh4rndUx06EjZbfZB0UyRwcQbzlwToFFmQlS3cGDXpMIAy4bqNniX3+l
83c168CMLmEvXHYucDYGF9wmTYF+WDAx1HWpSBen1Uk/MSce2T/aAGW6zBzYYHJT
vuRykDf/zs9d3bVn4M/RvxViCiW0GznPq4nyY5rYyb1IqgGI09sriUyHOeqnmakS
Jelqi8Bs5qn9S78dbJEdX7QKl9uxNoDgw0StDNb/VoG+ffIM6WydMQaBla3qWsdc
N0qvM9JlPDyuwGEn3MuWTiasU9fdkCtIsG6Wp1Sw6hprJq0NwhlygjusS+ZSBXQE
vI1PIUSgy9QE2fDPje54HWRvHi9VpOkqEqMkVYZgnjcnuA3d5TPhmHm4TUupjIs9
8vWeyas53+48F4icS4xYWOWJ310YRpquyHXSau12fCHFirfyPChWZZFeIXyx+2Ij
RJbkblkyUb+yy55N2Vb+omk8wfwM1FLBB00kGMJNAPxgNaQ7jteyrp3M/fGPEAW7
voHuX6YLkcUOEAF/lIZnLlRrUof0+1BJjelCpB2su3u/bTs2V2E+IMXiQ0/2IeT5
0xG+uQNIUnzgqTcu6X6lgRetSgdDn2mKBIL+EBuEc3xquHKJf0pybdcVQ4mo1uM1
FMmfY1B9vN6FiYgRVcYECv3K1ctKVvEpvP7Ev2wsnxLX9ER4TMdrHCu+CyL/mO2f
WCsVS7t74ce/NEer6fBmsmGs2t25n+EGIOAjdt7VNS5g8+rccrJn+hPvN/yazKxL
r46PGOzTD7UbmU9UjadmN5vM+PNvYhJbiLGcIigPjqv6k3l3m8FCerz0woEfPp34
WIOXp6Z7oNJB2yC68bXoH9Xc+b799HcsvJf90fP/9KU7NPJmglUrdSH7/PLRTwn4
lxnRar0nt3rdkpNpcHo4hLSQ4UngpiTg9qw3OG0ndkmUHF7IW9rBawAt7HEFBdC6
9rPIGUOCtiCkek8SrK9I3hF4wmhzzp+QA79WGmv/baDv37erjq2iIcB4OWmZRv/i
D4JS1vAPKLTyWR7B0FT7ib80GAvTxHM9tggya+OdIJ/ki3uvFiCTrb9ctd0Vap8B
zBvlUgzIpWz7rg0vf2JO/nYsRv8Q4A14m8NiTESC+Od71/l6sgdCZEYKN5FJmB5c
FrWbQjIe1yemOaGhi/LkQ2aNN6L0e1O3yAerhXwpRamQsCD0TmpfsLzK2d9/xVnJ
EZfZaGjIpjjZETb6snzvSIoToH7wRRwVMnCjcH3kegBvyVk4VFKFLzrJ+/Tt+P4A
Yi2dYtPEQcXSeGSLel6UAz0GaNmKO/jZMUOdVgNnBBqV0F8mDKNwa9b1zlVzA6tD
MoA59/BC0j0JRKmFOW/QwJECGL7rwSffkkCsd9ikg5lpribhYGvBLt3vjk/RqhwT
2v3jrReQKcscK4/U6KgwLxZU33JrK9APLCXRbWS5OHGMi8JBVIhzXXAY7FMpawcU
ZLcW3RwiNrH1wCDRH8LutncaxQDHgXxO3E5Fum1w86GN2KPY7o9AVKgOAuVnYbs1
NKyltyXpOFxmlyyVk1Yg4YJs65SZZQkOhPljLOJNFyfSKZFu4VjoDU9YkSLi5eWr
HyEbiIt4fRBOVOyybsBlAYTk9gK1ktHrCtS8JhvZXQj5O6eRHzncMCRjNsQTCLpv
gWQhWeKhWHsuYdE0so1KYHE+uvwu6RD0xumwP8swb/bxNKa0RMEyyTsqqqgw0Gnx
BBs2MpeOhXyFN3ifGp2mAEPBbhAUm8+RulBZxxEJet2lkE6iYkenzCGgfpLEMO9M
+VyaK8USJrx1Ojqj/scPQ0iwWIe7NCdSZYDFV16PRRX+yDpoA9Oql2S9d9sgiOpl
afHHWkmtBgc4rt+fi/l/edFZn4HjEekNKJLjF3mY2yz2zF8e8EEMD7ovCNbxU1gW
RNaITBt9ITAM12j5Vnh1LUruvBu203nZZCJ/Za6S0+TH9ldAZVGh2j4u5dzd43No
sDkXFQ55e+qt6CLH0kr9cJpWiOmOQ1xYGfT/JQWL2MzG/v1vWcnQC5QDLAHpA5J0
eM+4iu4+xlMa80/rB7P9wk5jwVH290qhMWUglzsG/GIFPTU7XSk8nEpObtW0Yzwy
Ud3vS3xhXWFhSR35iOqezkUg1IsZ0PaPDyDmKDnbHSfB6ZDyicPlMAcdVLV9VO04
FK4QwkWqiGaJ38O9k/0SF1IGyqzOjR1W41nvUXY3BC+gkjZR/MPItlRDplDemYnF
94ghKcjoO2/iYoGSPq4tJiGuqiva7XpVu0vwhbgZIS2L1Bpsc48iipDWpByd1Mlu
h2P5RTGpCL7nBiZtc+I3NllNif4u76g8aUd5PqjUsohqONxwACM4pDRoxiEAAKdk
WVS7pQyI+IjK5x7oJBTzu1GJfdHnhd2BCDVD1L9Zb0TUHgPgJMsA3HGROgciogxm
r3AIVnKK8F824619F87RxD8ILcNj+6JdPMrpksjEXa05BQ3Zm1HzikgPGCv+jvIB
GiTGOOTW2PE0TT2/ysojygJ2HfWs2nWVYNLd0PZx/zobUldxcPhdCiqDVdCfGHJt
TiGBJz618rMhcTUnHnidDLe8t2AiPBWHiofvoczV5VtPaftpfGAApfPLAR+uRhd+
EMOXnUhdeLMh1UTQI/iSRlqSclw45czrQGadlgbc973gF8RHv+phSf9rGzEtc7Oo
jGGfaIPyExMcyy2S+Q5h+iFK45dIVf09MRpz4npIRpkeZ2EExwT8MaKbkX8sYzeF
KJ1eQDHI5n5WzHjmlaQn0EXK4sGR0toSSO0MWDBsk3D/R4X8V9RfQeyWvh3Q8aIj
RVM/gsvwU6RaktzHiqfmHoz5Ct7+eadsP8/hdl7eQqyRuZtRIVjCbU2Id3JBHYtZ
J9yGhNfjTsQsMRuFd+Ywu2OC/uiKBsm+TOD6Ye3uD3OKnFrFLDklDtSST7NszUxu
ltZUiNsvau5VTq5pJNUlpNqVtt7g7Orb5MKEeC4oz2ykZQO+2gnbE/M/OJadSz1J
79z+GbG/WIChGV7WFYvSiG5G5oQ8eezPDzKZPwQJM7UKH0m63HKdYHn6lbKlbTrA
KyeeyHlBvbgsE8YDrKPmTd6f2R/oEJnM4UV4fu8SOZyLKnx01t6tXg4xre6zbM+A
a+2E50Ocu8GEQv2/MIwqRSA4z1GGi+zziVzEp9WMVwOmrMWSIlutvFeC4y5S2wdC
JhjeRG1fhDv2hHg8N0ruZCwe38cbALqu47ef1zfy0Te6sirYeYIO/robauaENrza
CBHn9VN47QleLKQQTygZxMsLMQiZfIV1PqfEu3xn1rJVEtLDClm1eMOA8JukXBp0
WgBUHAZQZ3KO/aCATrZEMxg7KfrN2RSotNF2hlvAEWvRbXtNHQui0eMWTlcl+qmZ
PaU3n5GJFGh1b85s6aFhQXVxsQpu2gjvBdRZerAuJhErpRJwNdX4lBRmAn6d94bW
BCU++xrz7flY17Flo3cIBgzicjqkQQdin4drDrFwJ/4rZX8/RrbpLr9efoIeZqDy
ORE5Y0Q3j7h/Wj4IpP2Y9oxaCXLymk0+K7vDz7sDNBMpHYBDJoHmPILz79uGtwYc
/1/xAZeK7ZWzJiXokwup7SukAaG+YkWzURlOQyU2IFKjSh+kFRxUDtZ19IqylpK0
7tCneEynXkuU7EQSFlhf+lPAAizUnsu3eFIhP8Wwwd2I12E5YFm/lqM/FAV/aMGu
cZf+D+LbfAWRItg6vlvp1KrxGogZQdjVaHx3L2SuA7vsY7nGRgOEAdUqgQwW4hzB
V10fBXrWqB16TOr49ZFikEHWRkgSYWwzxFZezgKXTlhB92faK+WDK1Jp40dglrjj
NizSiDWkfBhtR7hckSg1tj9+u6MDCI8bQR9OakR9uLWd6gJpm2VFLDsH1yUIN2+3
YexrFgyajwWagCvCCiTPsKJjAP5ETknLLembuqUHi1W2zjxYpdNIFd+omlSUeaYO
u4is+YwkJ0VZ9FmE1wGZhKrz1cCc5JROMby4tw78SBgFxF1w1FhUsoa46jDWNha3
VmKQznJ0MUTNCAGWJKaX2CVrrGdlBWupXnCBaPgFDkDfM89Su+5KOFgUckAZwsbL
6Y6/v7zTGCGUN9AEGNFsflf0Xl1iykiU6IMcpIWWvUi8QR+6mummoem2YzyyGfRE
VIKwK3IL+w7hXcm7wVZi4kC5ve9O555pXVJCNMFMmUwkl/dYy0QP48FFaeM9QbeY
kTshHgWALsDbbRMU7t2W8t2/nFu0qKjSiz/Wwjsio4jJdEPrWI44Qmlh82s+Bnis
kxiyx9ccYCGCVG4560R4wOygg1wBQyJLz+I6ZmoW4hetN4hRg9U2dTGHu+G1eZAj
3I+3yfsrUMdzOF65M4AWN7cU+uEiIpFslkQLZhlgPxhptF+AGQWG66+mLhfd09x4
/XhZ/xGUIvBW0NJt00FWasBStI9W9w3v+AMT/YJN23Oh6S4IulWRjdNFFcVHrPdO
UO4FtcsN5hzeo7z5mOnPKIan2hUNvkz5fzXuhPv2gQtvuzKNakDKzIukr+2UuJMQ
FqQk5vE4Tgv7ArujG1qTsjhfvZEa3q+OTXakk7UIyLYpiv09iN9nxAnzT6ZcYGA+
LjyT1wIA6CUjRR9RI79FrAXRxDiPdteYKixE5rRzZLL+OMWuhlK72WLfHGLyYeOm
RRsczxB2vNOQXjQl4XbafJPkKOi5lNFyvfr49Gs/+9iww0UnZ122uYhCVCHV2INi
AYQzhvDAslVoAb2mA0G8fxbXG5Y6Wt3iO2DHGJ4E1ZExcGePl6HixIXTqQxBMmr/
S4FEm9W74gwWlPQSVNf5/aOj54zpde5etlUtjB+m+11W8l3J6faaOR/+cLyVyliC
QFIV6oVVSArpChPqvjdLfs1ZbAmzzs6A8LVAOBkFGL6ZPetEgZ5oc1H25RSTInax
pKOl4ouF18eWuMJq8v+a8wTWByDqaVS2grjK90FauxeAkFpIGVBlSOZuMJnk52Db
VcVSj5NVDGZ34+kEVoEItC6yT6xjKdh3qpomVwQI+kStK50aWAsoPANZ9DcpOAR+
iT5Zxf9NkLjG0o0pEPO8Ctt5KALx0S15EhqzFyCXU828TiI2qZCLVrGzGwZtuzHF
ohBOlwdTHCCrni4mFNZusik9Wwei9VD8yknZD9ZM/0AGWjNikOIYIoa1t1pFjnvA
2ZKzWZdVovOBu+WTp8XWNbAYgnONMTQBKwSvkWhnRFFPIJ8lKwTDvXBl6zHDblLu
ZJa6eGrxS4b4HR3ogDQfU7asv9p/AJnST32FmEuGsO3E3/lPfWaak0ed9KaKD8kA
VQIvEtxumb7p0qV3fE+/dHRS4aDchPRlLRr3HD/904mnJzil+sw8dOpLBdiNVfyz
EbWoj9ZzqFoYEkfFxaQUvIHKLNQLRXGS1O2WhRAxl9c7J1EXbejnQWA/dPomG/Ap
o3tS6944cxZadTDrcSnj5vhqT9d/UpUIk6q5kqhdYyT2iLTY8OtEmNIYPd0UvBHK
/SKkxK7+Y5ea8qFMVqOS9fsj9+wVpNwSOSgtTf01O/9FJZzacpV6NGDBT2+lgC7S
582/JIhhkZ/yE+7bKQjnjyoHyHw09oEbpDU5PpXnIQx1ppt5wZ+W4yr49QWXqG7P
kxyaLJ0QDW/w0E/2qNfA2vBgvNfONXPHJIXaqOyrRIKAXEBd8I7UvzYHrbtpgfJP
o1x/eBdvR6cZ1w1t8dFxqAkcMkTiuupcCD0QF+8VacQAjCLSPM9kJhXQ3EC19EgC
7Dq980rr2LXupKuyHxIjfb33Oe+PEXKd5a/2xAECrGurwGRivFB1jQrDgXg51xQB
rwPBNTRlc1ox1FWHvpPbpw2NPOeIers/Xb5YR1WdXgxKnsUOgUWM+rUgUdlZrCaW
RNRZXSbKFVxtbSR/USVRqK9igjoLuEEbtYE4uiUYw1f7mP7MiK/ai96b++G7uxc3
tKGOyiU7tNBpfpeng5TYEU9bZsXJohY8P8Bg09W1QeekzmZLGgym8B4F/6ZHaczg
9tqnlqBpRXOKCqQLu4YX3Uxzp3QAiBUDmE8nnTJxyep0PEySWGjP1XbdOPppTC7q
9Kt5RvTFHxWYJTAvbxWuAfWRpFnKOhhUYXoKP1r4LWD/vPMFvHd0o98U1GKU5v3N
+mRC695R3Kn/BK4wTmkQyopFhur19Q1hAiMJTGrF53ChNA7vm6jAX4td83C58lbi
a7VASGCA2YaHXdK7vGA19bmbQUzjjj8tJ6m1+o+mmXHWLE5YifEOjW7wH1N3nzum
G3TUeBbki6uBGq685kMY5dT4+co4dJ2OOzQMhwvBrjbmlydX8d/uW2+Jx59AHohN
fJceImGQvnXmZ+4FynieD4SGNkr6NUgByxdH8NYAsz81HnH1A5fqERvq0LzXr2xE
jfHWXddnmnJqKh3v/w4jxd+L6niINMb4QZI4fpnFu+o3INPevCeJWpfLbhIK+yS5
ri/e8xMjPDnkbiP4Hz7X0lznjnOK+KY6R3L977rVlqKOK3BX/cDg17JnX6yHhCKp
DoZIx7bDbNMQjiI1enC38S7XEROOLIFfC6RJTw4syaKrC5yPLIEgye8R6YREux09
bAW2uLV7PYykRie30C1JEXGS9SWn4biabWYX+vLddRDOcAPeMtV7EzPRN3ZkQ8vi
WrA7nPsn8hw41Az9/PZadJiIdmf1E/3A0S5rKFB5suNel58EcfE2wanGJfFjElGz
B6FoyRhYUuiDihZaZEHzkIB9TgdDifXrMRFm9OfHSMR6gxGyGeGRihongSuAh3Sm
hUKQ5jZSeBhM5V7A7xLl2nrrZeetmVU/4t5h2lfLs7XdCnCVP+dxxacUGMgbNeU7
DxzfMuDdmHfIaFUtaX5qZofqFv2bgZQNxfnEqM1Rzlv03BcvMaEw1wzmEoT63QtQ
/4leFeu32ubHNm6wLMq4b/IPjNMGnWO4Xsd5UNyI/sJeu1FvH55Bd0cTzrm2TLuX
Kd4HCM2qEs+MfEdXklEeZtU7wuKTAx6daS0y5h9+2XS4mt43xbGAIfouEGKeSAVV
+BE3cjLBFZbuDJqgo+N2h4higvD4WGjBmzlxFHvAvhm/6NUhwhbqTebQWQMnr4Bo
XNR3XKwDbzTiwG4WsziMkM+2aMaEgzBSXNGk3n7c+jhvxx/xR0FLdMIanSQ6FO8A
n1oWK87tlxCPoIyPmeWc92zF0wBz/4sVA571WgaiStE2JkZnuemTdRE9ULboc99F
PSdz4kn0OM650JTIULm7REoAXnFLSLzI8PQ6bQiiykLz54SWHg5QE+iZU5MWFlrp
1a0pugHh4UauBG1gauhYBfyBOJ2HluqS2vGvh45VFNHQ6UxLExqrx9anZHqd4j7o
pnZXn8tFPBlzGr7Mx9R49SmHn4tsMfhjjb24ZuniwVTfvEM5Mut/3QFS3nBF+C3Z
Tu/+vZIy0sHApGO6YcdAhrF8AevQqxSosspN9wko8wbi/o3p06tFd5ykXYrTALVt
1xMuhNDPjOgx36v5gR13KiCPAl9Lsk1vjDuxGGp5UWzStqF6u4tZXLFOSVaN0mHb
9u23c8lA8HFoXgskYP6C8TeL+bNe22bqraNh3rCymtXKnW+lv6WrSM2K169t/b0O
mxtokufW8rv+VT/YqRIKievrEe31ktbgMq9//+W27h1ksCN7LVnhVAoGHiHEMQGh
dsqBcJoUeuYon5r+ktIW/WsJdMhLtqePqf1a6XChhJr9qIZSHpXBG5MqlhemTs8M
WVGNPqJHasOF4hhYOUhOhsEC0SbJgXD8+8VPjLvFsCnSNzIkAj9nzHa4hsEwt543
TojGlwZLnuEWzcYZa8W432C8Gy9wHgQi9WEYs7isse/K3w6TMgSWAC7KZIzCsuYp
6mPTYSM8+c/tva/L9H9VM5dSOEhgidnTtjDarFbXvohoF7qpIZ+6+WFBuVXPalA7
vUV5eJD4woUddhVwGsOGjYqj6Jl8iQhg906o3YJcx6dDRnjkG2FU0ArzUTxg2/Z5
k6Ahf7/6PbHpAMVM+Bc1g14QCaVrE0ZwLpLh0KI0XjukccK62Uynnll3JkJy5x2g
6mhfzO+VvBuO/mtbSVqKWahanucUJZsnv24UK618z9BRX2CHH9oJ+wug3QiVN8GM
GWUCc7cj4AljenYUxYjdlZPWIupgRhnT70pyvLVTn/uB9XeUwm1lZ/HJl4jeWyn0
AtfdubuqZkO5xLcctay+pbBIy8M5nnLvpL6q3BYv2VKcNTaUFkJgHgDEY2IisHWn
o+EPSkSh3q4JQqSQ8ZFzywagdTQ4CJEkgdQFXYKjhs4lLnRoXjMNKxzVJ9mZ1gcX
rjfXxco8QfJA5hAnEsIz13KAVq2K1LZP1u2iygf7c4P0Xspv36X2s++Oecl2aq5u
dly2SkZPpT0Qp3wd0ykPmUcMvEZL7iMsLeaITZ9s9QRXyza0Quybv5XfcovE1MuM
ffQ/3/SQ0kc7CdY60Pbk/WR0AvuWh17dqt2HtqRr0hWp14Plqn136fJE8lqd1b5L
BPuk75yXcK/xmXsO5hTXiNntOrjQNO8AXJnin68qCm84Y/B4bmDbiECHgWRVj/UJ
OHeSPPcSxILdN8UWpGHa9D4V6KoTGJRnmbFLcpbbFpkaF1+gGKDQCYcE+OXHVtKr
QyRistPZkkqNnjHNu27/zxdzba0l9HTRA7kEMDv8g+u/ElIOq/7IZyk6OPemwCPf
mBOKkOf+/RRkZmfN1wMt2tlpJmWKazmEywWV0mqf8KQkkjjaeIqbqSzF2hcXX8HE
coD4onpVzycz430q64/1YyMl3GTEzbd+m1PdG7LxpBABpibfSbUE3sVC8i8F5CaA
83Umwthod6s3s3NCmixGKOuZrFJV95q7G5Vu547dYWLhLziMRRlhfAr8utYGzGjB
7yPdoP+uc0Fn7bcPeajanltdcfl6HrwMveJUDTPtreShQdmqNoUtaNRI4Az5s01H
YzvB59aJRK02xRPd7U6Y3anOpwXTmE14CYV7CskVDJRxRNO2ih7J0H8FIJQFTZFb
o0o3SK3lgUb+0nnDsk6lBEotLOfNh5bsGrVt6yqIa5xl86PpcrmYh9Kep4bShmwB
7shBZIv63MdXUEHqaA2H9Y2HlHzUmOhD4YvZuUPIsdXtxHQp+ppJ2/qA5NuDHUxq
7+L+41hnXIVkXCCs/52fY7+4ZZ0dfzI9S0gjElbe659jduWVHpljEEnDbOmPi/na
dFT9X3FabIZEUsEz7kEjDpbOy+XZe+X8z8tsXpykNiG8/vHjGU+xp5S1qgroWD6s
t6F7amo+YiKB4ipFz35MTX5oiA8W2JROZ5nmmKInoFehREh7szV+wfQRYtO4yr9w
DKkhCF9Jx+5+Cu4CePj+UdJ8Htf+lIzX9Dpg7ncg2c+ws1O5K+8HtO+OyKBGDz3O
aFrMnNyRMSU3FOvo3DUMIKqq0v2sguwHZ1Y09zouc/kfakxz3cqDhVsZpCFWhw+R
iCcqg5I4KdoB0Q8+/N+jQww81DXKcGPNiHkWwGn9NutiSzXCus0JTMJe9p+gLb4J
P4041s0NSE0sb1mZH2Q5nIiRD10wcbCki7wmldmwIUX7u5ibgTQYkac00tsprLR0
7OWbPtJdmweu9tj1PvdBhWQzk4vAHprB9S+/U3jJlEj52GcuQzVvQy0nOkvrnNFa
7/HaTWYfVJrnKisDtB33PV445LzXHhiafFfBb1qBESpzKol04/S42tzLlZDKDbnc
B6XkkZqLHKYhzFeaZ6zVrK/2777SwKs/KWvxcLxImK3eY1aig7rDYqvN0g5aMhkU
CMozgeQ9+37oZRSCObTyOs+cgE1ZT1wcbPX3nOlgI+uv3kvljx3gSG+sBH/3snlF
i1G4QW8hfTUUEgBsACkCC6rcLhHdtH0cKW5pbgNBMgHagtmZk0eEp6+8yc+xLY4H
49z5sCF6GH7mZtQJpu+ASn6Ky7p34fOm7SS3Cf1IdJhSGIhXW7nv4605zAk6OVU3
VFaFtGfNl+/nltXiH3hg+npO545rr80nc5XlJU/31mPJjKcQb5CCdHiel8tfJ2mJ
TKTLxvYeHl6BqmNyzREjDS4tiIQi0EX7wuM1tHw8oCDDuKDomuACw51zBoC8Gzm5
Z3Eo7y4p9ZCHGPyva/DZF9Mnk+IRCMW3c9SuqhWC5+FzWubh2L+1f6G/yS5hPuSh
K6BrzfaaVGHQ2qz7YnsIwCN328B2F0slkwahpIOn/Y+CUByByEfkqxOtOQqWPEvU
OC5GBJQD7uNzg5ZX/1UIEbzrCygL9tI0EJEnxVeiLl9KjDzr1v4OERK07w6Oxnjh
0zh3e55esLMW5uWBIvZWlCdrOaMy1+SreAs5qdy0MH5jWcj6Xgdj9/EB/fEyLnEt
MnxdQAJAsPHlJai6wBDg325Qdfxmmygh1QUWPRlwG/YhlBBrxi0aHrdXYWlOGsJC
rsiIgBbdZ7cePIJmjRG97fyWnUNyR17/tywwR0HzCOZZcroBIVp7UjUuQfRibPwz
ZY9cJKdjLXdAFdjdm6sg2MzSPgy3vRDyAUzv1VO3A/mNv23IFDfoB2jNSg+2BfSx
Ro7srp8tjFMF6oHpuDhQSzyW8BmK8iEfEThIDqaJrJ96HbNcTHEwKxxSOQFadC40
28fIb4E6rr/7PTjIme/VNYzXhmLFGrjGOyVHPQqrIYAHcmata7H6wBe8vahHT9s8
FFJmqoOn/vnDkN5dDm3gPOYMO30TfooMUW/tLgAp1Gcjf9NaTWPlTodMojUybkyc
XVtLM36gScPduPYbfMFbiv4zq67Dx4YdYGtg4AeFrhvlRgdOwJxO43MhtmhsZ+jQ
iM0mR4TFmMyvRKYVfRxNqsYX2OqGlvI8QVQZLPicESy9q60IPhJDQgO9y2ZxLAFK
CQKCnTMJbF82RO4CjJV9pBuCTHPDWP8MCZidGXbdlY7yoE7bZW2t3tPL1LXHMpE/
fbnaoWi6wMFsFp8vwf5peHY4Ilb6a4CD50IahiHe0fAdBh25TVmmUwpFaSzJksrt
QsJHEm92Oz941YQ8J0+3YhL0Z93YWfEi9SP1OgjhVNqq36egeSsIV4y6TFBtbVXb
Or814bm0O9Zqq7C3FXU2grL6Di3vVl754BzvPl+QyLIJ9IjSRwrpDXTWCMZhduab
gFnu1akjPE+RE4XqpzMnVr8JkSQpm5gBtw2buFXVHaL91JJJEW4BCTZVB3NvIbIq
dxzTRgrbwDqP3GtlRfAn+Zva3aM5HdYJ9A7vWNHaDyxpPHYGjSNk7iukwQU67hCg
RPaF7niDWg86kQg3Drw8ty6cgKZVVLb5tk2SbFQ2lrtTcKwvVve2XqTPMErrvY4p
0YZD5/JAw3LK3iJYJVQVyd2YRvafl9sgj5ehB1Z869pWXY/dNQSBOBwJmOh4JtIU
4xeeKKxaKYXQ0FyJNl4wSMy2GduAtW3RxTP05HBbU3Y4TjUagKK2ndDZaQlb41By
Bw6oIEAZOycpjl/mKhQt98gyvhhNqZ0LLAgHK4FpY1wcMPlCsKbHnFT2EIg9wf+z
TlBkI7H8aUFljh8SUQ+ZVNqz2NTjo8+ZDhA/KeyONnwjEJQCKEvK/ybZ6rrJmd0F
JGjXRZ/IgPi2n/9+jfRFbzxPz+7vrKe/fUQjfS1zevU9wDTTviSFZhqQ69Ho8uVW
7Nu18l0MHB9m5kstQnXgA4XLjTUFkbNoL1x3zxZGBih30GwQ+hOHNk53RNgb6lRF
BPR9jltNwO3+Fdpqet9Onb/fgfXW8wBewEpejIozoDz440cHO2+cqwd3hqRxQjI3
/68ltFrMwe524BVrtyKwTQ1ijb4pKkw6YM+hk7zwpXYddEAo3/ZQcg/k8nzjm1kI
6g8K6eLjbSObBU5EzGrSaOdAYivVDZAWC1gjwjfYMfr38sFlbJL3XwRdXm4r4OvI
g04lVlOz1cy8vpaFnFJdn/5dX5vGRWK0aTgjH6hwuKOqWWWf04iK4C7N4BrmyX68
kbnjBJjDRH1yr4cQ6yzPLIcIh1NI722xycw30nWtdZcmuDs5+kC64P53Iagl+N8+
RBDsgny1cmyK18epVRCTo2tigPRhPHY4GEe5aFcFV8lfyeaWWP7RKJN+80+ogT5x
HSCV7e2GyMtl5TrEhNCUwMUqo6cEYacLCJIn3vM+/5zSZ6yyGglUZCY11o4NKrvx
DxBSq9hwg1xSfZOdsNx746EOsR0WAY9EnNkFlgG96ttUVCL9AtxzXlfJ6mMsJ9t2
xqyKVodB+gMr9Et0iaHxUNd40ZuaoE9W23bfxA8KrdyeTWuVD1944F8mp8EE88m0
GH6a02VEiDOxHZhjpD7gOQCCcqGzQfxLRjp8PdvXyBMPu8iPcO/Zdt4fXMfL0+RH
5kN6cnj88H10FJl1DKjpjb3IQiFS6+GLVntUiYH4Zhj7y4Js6dkjAmZ51AKstkdf
g3cIsKkMeEw9ZKj82W5NSA7UIcQu47/PalblIR/ckGNfH+9SxTWhn/DA7MlGoprc
PPe0SdQSCtbmKsATSvprUob6BvN4g8DXKY78YNzV1ohZH1x33Ca0bTQBmTyyV/rw
M/px+6RY4TU+NSntAVzfTITXNCEdi6Qo9BzSIVhg6+YL9mo2CxP+tnRNHQHgqStW
X6ama222uLbjSr0KT7ArbsizE3GT7zBgtNUS7jLmdBL8WqrHaNIwwANcriXzxuw9
gv1VaCxeaU0+GdYext0uv0BMIpfZZ3KpkS+nIuA4zhg5Bj0IIKBT1SYeTIHYseM4
tOQjJZoFaIdzSJXiIMRabAM6FVLZwP5DpzZx2gDoeEZGFmv0UlfQYMFNatHafLV1
+QkkSkp2eG1MworYzF1ZsifVRJp6SfDtoucYmHJZ8gCsvZRJakApmwTJ9nnk6YW1
XOZtDq/H1ALM1cAZBsAE/5dWqx10aUnWdTWezg3Tt/IO8z4WiYd240Ae9F7/4r0K
fmd9AkYdjyZlscMw7gvxEqpnDg1E1PLQJcJKHd7ke+jX77s5hpSV/PZrQ9TCxJto
dje/C6DTPLEZFYa8qLoymQst1BDJM15hmX++zgkRC4OmzqbMnP9Vt6rBd/ZUaaHS
YAEgcK6VWtdPHCdrS9UEky9fO72IrBKLQKKK1TpAp0wiDjfYJm+BWEqRmWI0Zpoz
JAFXNB0DrOIiordTukUC2MBs4XBhwGAvr5BLFchOjRKmLBbkbUYVBLIAGVTY+ldv
GLG32xT8+k1z2R//KvoYerWVAmKZHdbhLky5uxm/k/AwnTtyrcjZ9AWbix1J8V/l
5sITFfs35L4UXu2FueTVsgy5z39xNMIOg7p9fZ2D5kmRMDc1D23TT7wrF7B4G73W
m45UoENx5X3S0tKAxl6U2zTJx/y3m9JXGfIoPGWVKuG4kK3QjqIE51JZzxbqLwJI
Vh872wHvtaCXVab3nlClEKZkxFn8wQvObPXiHBhn73YeDwhb+FdHoeLhHwRLul8t
Q2Kf8U4SPZUS0oeOppIb/DECTpPQOEnO/x9GNtPdO+lwDmGnLP8t1b+uxTgHIT2I
jffEbUe+CS4sSpK1gvaz9tsK0YJQ17L6JatlP4YP21NYshXIAl8UOcOP1PH9xkXY
E6kiVDHTLhnn4vh/9K0s9nnSXbX1DUpx6QvpZ0EJ3oTFTw7rSknYqsMPw1gWgyBj
sxRXuxEKjDN5YXCeboxV9GD9ld17g2Ffi/AQ/ZlmvUu3KcsAyZoywU6mwHd3MT8D
efqs8tSGaOwMhizmsWuvqPukObMZhOpOQV/BIUTWI8FSRvd3MNzyWLsX3OKmbq0N
4h7k+iAeh++tCEX9I6IJXDumoGPDEsIDbcgHS2dRXOviJwyvyHeNZwXiw8k/gjMX
CV2KoyqmHPzIePO7/TSGZvQ/LBfa02S8u76FHpwy1IFe+slZ5+iXUy8Y4YRUaMp7
EdYnnsB3nYp/a7WNbDRjNcv839lzkcZIeWKDt2J+/8lCJuzdOcEmLcCJuE3gxGoQ
5TadXtlXkpNa5Jlx2aNTDFGcux884fhhdhEZSuVfPSF1ghe54bY4JqMyg5D8hyLR
7kI5LEELVdHkC3vL38Lz+2NzjiTNJKYBshmPq4G2me5ea4agmFQmIIVoC46+0ptg
buKMoatXE4tZMVLHvKZffjVk87bNVDABFcAIG92Sn9gQd5fhmjdVQSPvwvvjd9sw
6FLZpnQk5zgFIpzmXfjMJpRI4oceQHz808zQOzasskFKyRFHOAq5UPo+YvqcGWsl
QufP6UFAUFjX9PM6MU3dk6mRjLDwKimapuarlsgxlO4TpnV8n6mvskqxdQ2l7WLo
A+TB0D7H9GBDjxbNs4uHc33djoxkp0KcUQx63NSmUXh+NprBYHrCibwkVD2IQGRW
lW7gLwObC6DBtnR4B6CvqOnS0dmO1yiJiIPnQz7yFhsraeiESq81Ba1R1A/3cvGf
H0Fggs8jhCRT5Cxtufob/1uDbA2FJHgHVufx3pLtas5iPiCzKWou5+bPZYaWTYy3
xDu3Ajk6vRvN7f+HslpSWuLElRoRoOGaNM2y2JkqpCnpAC2QxoKoa94c8EHEmx82
i6YZf4OnUgaBccYoEIjTvF3SIrXnBxPCFziJjhUOI0oUcbGV/ld1xa37LjnD2eGz
Dy0Ljpz08Osf53MucZzRCDirRPm//j9tx0Kx+9oAuj3yMCP7gDDnaxOY4AeXzoDn
okxjK7Nxaa/u1YJExuP8une3f5entkkEHEgEJSgjbVB6jNs4yP/eVAu0PigLR+EI
2+g0x6nNtyY1/OfrnNcBnMGReqalBPNlv0Wvlbg7cluS3/VqPa5Q4QH2wmY5yd7C
TSM2OeXss71h+u/Q9wdCwj5qiM3H6UDGQLR/5F9Or5KKMupZhtf+MLJ7O1tmnCc0
g/eMAT53H7XVctdrjwTR51KlveuCsoA7xBnGXpIr5Fa9r6tCphjwAEPTPEoWSi98
3yF8QgwqdCQeNc3ZAofeBZoGXrYgkUzXD+YXRVCvLkDhg+gysSAjesnxAfEnNRhH
bM90ktPRZW+0LZe1T8J0EljD/f5kkT3ZLznxq4fQcMyoGr25M9XCB0S1ug1Mnzbu
hoKv5wCffGu5Ry0kzzmOCgsJduh3bwp2WzEiU9FdsJQbTCAM8rZt0W4mEd9zKeqH
1jM2hhLqMXu7net8HkPIUt0w38vWI52BVeVJ4zg8mNPMzM0wTdiYx5DUwQejyiQJ
CL8gG6cVe1ko6ONqx1BBYl4MCk/S3nyz0Wp90B4JTJ0kTmnwm+hkqzHUXogkPiCm
Z0Fojs+9YsQMV+rgPH7f7RZdVst9hWJjFRUOK0guzoOBrKkpQoEteX6CtHDTzT1D
94bTgEm33f6kZlScrn07xUglnUv1Hxc6GNd5408yH6vlmAS9g7gGsVDdgjc0mCke
7oC+3GCKwii9nmvaJECQBGDH0OQjp4KSH9I+WnBfAKPegTk7GfVdocqIKvKk8nmU
kYpnQxfGRK4/bkvn3dzIa+3/qcfrFFTJdP5GBrpQKqV/a2bDRal8fKdAiYM3Y27L
v/Kb4KT4n4IV+6VJfoVSChHA6AIvJbS02CbAuMHfoN1YLMJ64anNX5vcIb2644ae
ncj6Esxy8Oh7kIH1Kxl5i3a3bP1ijM0UfTzxLf/6f1A+Q29W+5XTJ7zk+0aQbw31
vgekoC/Mwd2XspK25+nODTlG4izM2AT8NlAiRD03RaoXaRMgQTCI75t5Mfxk3dHO
7DZPwyFbPC6IiDvzPoVYzkWlBO4u40tTnSKKCWY/I7b8EQmEyiuxbIMeufXOZuT7
Mk5/JRSTi1t/2oyUHpMwQaynThpF2GrMLMnneVOpFBkCrPSjLmMt2QBklbM+FaWm
2CQYywhJjQaa7FjjIG1C2VPh2CDvH0+e1jyePJem1Rv5XZYURh1cPR9+695JbGMw
i00FOxNdJ2BczzSxQ02lPtdt52KMmO3W0P4laqRWFUVx2dSrvwpBxramMm7gBre5
SQ5sIY9wCsoy/l0MELWPVaWh8nAMAuUWI4Vs8TKpciNrwLqv5x42vP6PVinQ+7Mm
QA6Zi2ThelsrS9vxwAlje6ZmtdkO4TlOH9AAfmXBPm0rSd2zFNbQGqdLvZ2kTJHq
W6nTwpeItRp0hTtB8WyfRgmYR3IE9I0awNcwBv7GPxBk0CGuf7EptF4KHbiHQOgo
OP0SfQ8v48TIj5lxqRgTWSDU2QmV19xndlzs9CeLah0LBUEBz/M7UY6DYjo1b105
gRdxkwVrei9t8p0jDP45ICclfoxy9BegylrE5ub5rxLSc1IAdCPGpWyYveV56M4H
aiGk+URM8gDqm6pfxKrVxborrQgCDzbH4u015DgkTsd5g+5uLSaw1GeGiuQFXZmw
FIHbfC4P78qXJDe3sNz66i395kRbezeKC0D0gzmU9+PqlHc3R0pQX1LThwG0Tb7X
7FLDbRESgL1Uf7tIEJOghe7rUzPwe3RXh6wZ1DdwWt8kXaTD5pegumDn5Frn6COM
uOWITubyHLmo4ee8Z0a+1u5AozCPmKdwA1hIhwy0VL/yhswKbw0qPA9DPPXedK0p
im6SHSF3AVftsOUcv6uJtP8G4VWGN/VWOJdp8V8tLXer5tE8F/d0XsOZPS129z+t
XDSITSsNIVXQ3hWZe+SoTYlEytK/6c5rrhS0aVv9+8CKlBkYfnvVX3fWZrDpE3By
fBFXxx7Wn5g9BHbuF4ZVF1oZ9Ydfe1LPLj95o2V3DyfgkVX5PS6xjRiLs8ErC7sW
6yb0KtLUabfgaP7g/PtEPrTKZAIkCqXAsHiDTSi0m2vcFsN12oX0OxbgaCeLt/ZK
1+/5PGjZjEiJcGjy6ENHkBNyh4R0wTS2YMLJNBXNiB3o5QBCT5i1rgw2RhPkdO7s
iP1mwa4Zw671y7rtSTLNClrLs+BkWEH9McrMxM8cSPOvtLHyn+p4PG8ed5+gV2oj
4u8Uy6WRu478F8vLPg7IQf4ZbBGXqRNxkG3jmTzaddwBlTxoChUCNgM0RGTKUS69
ho9riV2OYMZVdhSMK3g0B6unNTbaLabo+Rk67+IYMgEhjYyqRgfHJzs4OTd3LnFm
M4E1sXX4fVwAr++zWNWecmQOCW/TF7IwGsgarj+50JHxs9nD7NS65qOoo7UvLA0b
al+R+nppSjj+uNUjeL7muiVen5uNNJ6Ahf1MxIeF+AGC7LDWea++78lV3oEdC0Cn
Xpkt+Mx/McrozeLEP8COGn/RoSrr//eXthfOHZsj8ehuItM3ePiF0WoGqXmnn6td
/80+R61yLD9BO3lBgPvemYRzfXTjDAab3IF8Giic7SnF/dSgO5sbF3kB9cq0Aa3X
60hZFn/zJezR7UngDoiMYCVxycEjyNnq9GnlrL9QU2cfs6IN4Q2oGCG+6wDaJSjK
Z4QTvFHthwaF2YUl+uQtBcmHqc8kbFrtE/eOQp8nl59ThWKGzg1CAhccJH8ne1wH
vMysrYXSW2LTnbo0zGnJIcmbKn7B5vraKSPpcvbrhJq0pJAjBq8EORPWD6tABbyz
3u/iMJAOjKXDD9XWdUHlSBfroArIdRmMLXRWFYEFgB8f7UllSH/vVh1gWWnd5AKX
qRRzSGXfpNDPRGMbwngTO/gJqOchCSA0aiCv9fYaM6Q5HGPQqVh2bqWc0iFTC/LO
7AWFxDFxEfm25SE/fu+Td3HD5F52qcCGXPcgAmI7WPO904h0j0q9bgQdqXlJ/c20
uDOWrTUaeGClCCz8qVC5fW4LhSYDLjwJ79wGruwMq0INcuhV0sx+0r4EPQn3Z72j
PwW6mTUI0MyrAQsnHOxb4v9HvporSGa7M+ICRqrMnA/gDPh8eIrkVKz1RCZs/EE4
VkKGPU7jCp5E/FzCRI+5n2fnu44K6Fyk4CnAV+G3pFKjkhA1X2fHHEW8XCm90E0D
w1pv0bmG0tO09Dzjj1Ni9G6BCuvOa8gPfawExZ6dWt5NLoRBxwEiduyE6oPD4ckl
+fKJphwLpMrKnYm62YLV1r4EtXtqu71lp7EAjXGZRweplGbCKAtH0M/yCO1Y9Iqx
YkYwKrAWX22zqby4pxUFq+ff2ndrquYYrlfbMNWy/WNsPU2vxA9bWniWwW6n6d+g
NAyJxYbCFDcLJGKWdns70TaMVi2rMJzSvyny5H9WQlrWO/Oi/jcknC7Q54ENJHqw
GsIbRB9+7A+hAb635qCFGSBvN3QcR9yUtVMcFyCJySoGG9Pu3QVE2x+4RoC7pk+Q
B2dV+ASyXqTYP59aTCx/ppHcYTgeLhw7SBmfUZYHMKT8w2wez5h7+PHfaQ51ER0R
LczuAWs0qiDV6rQ0HXlGgnyHSZSPx0d8N1RmhXQ9fILgokpqQwabhwTu3fwi+bQM
aGcOQP7cezsYcekwbZ7bixDoeKNFymZOvj50zQXxOYmU1DhFTuHX5znQphKzzI3z
UbgjkpRKroshV9KoxrwIBEEw6qevj86WafXfm654NQImZjVj56xlNLwQW8NFhmP6
nZycL8mm0hYwN7RPQ03kob0iceGaBeTP4swf5URpgmgnYheceuy3lZsfpaF0+eZD
AmMIwDM8D5mZAIpyeEt226vXkjzo78yyOnLYXhiQYwSlSd+Sb/9XQt74sCUSgQEC
7IYBn8OZZIrDMfvkRGfISnd9jThqU0uQv3rnsbxda/v7iCGWUp7Ll4uxHN0sY7pt
x0C2sabKR6i1bJbmdeIXJ5A/Xilz7Or6KgwN4UR0mGtOtysEuSP3x16NYFOZAjUa
vHWfYsvQUHYawjrMKYXEdjyzZ9MZ2FHLJJu1fQI9njRRL51IzG/7CKMPIhnlfOrD
4GkN2qmQ//1zY5Tf65Hdc7HNVkwIxXSX6V7rrS2OzvPojUdjuO0/eVJ42d2yfcE1
CujRasfzO0qUzHzNfiBEizfSE3FSfifa7D9+VudRvjXC3jde9qWJJjRc/R4BQOSx
D9TrjNq1jTuz9WDa0s2B9K9XcuTkSUPa6FoXDoMEiVO9xXsC6befjwmAXL1RWpKe
iZWQdTT4fWNJdUA8m9Z9AqJOVgMQw1wsMH0rVk+ijol+0g846yhFlu7kJYTv3F9M
IfvkT33e4KcPIkaY8VAL/Ndxwgiaoy36V8qElrcSSq8pb2vSn543t+cgCXKH8pNh
1OFGIwf+cRzk13P11yID8xtIpRA9jCsD4dV710S9axVgJdqntSa3bBRmfJ2QBNEw
zOdw/2zvMvMrdJuoxfVxwg9mDtobWAP1w70+Ynudyv2u3vBfQJXPjS6S9Ti+auF7
Jg3G8vMIr/21vaB0qsR3WEZiyVNppdkE7u9Z+LcCV3kev28G9JVeaNpIM6HgwZE1
9eWQQk+uD1hBqJ8H1qp+UxBSCksnQCnDsP6zRi/Igqir3DFP4ZVYo2RbEqE0a/FI
ToQiULD0qhzqJwfGiujWCurMRyR9x6XPhLoNCi00d4qnKxsrgzS0fMkjQB9qWb02
6Cb5dr/6gKfw2ocNHeMLdica57LFMxWju2YRF5whAUXXatcEW8Mn/jEpDK5KisMI
I4ujeKofUyN8vfpWkr7Yq6zYl/tMk+JK9diXqTPp9hRKfn2nLj2BkCi2ljcQwwZ6
MaXkJh9dOPRl8T+cbdUev95Ni50CnhdBaE9RxxR8n9XrOGeoFHFv0z5Mfj+q8zhU
3yQjAojuh6Mkrwecxjm6IZHy2hFiV+rGstz4iETq6G/XkXr2Gv9v2ODG4HDZ5j6f
mL4VxvmMXXJ+mo1b6mObMayffvByOL/aOePGQjaiU5lF8nmwdBBTIJsHGTYz9M4O
KbbB6ql06nhHGVbCTir2JwjM5N7WNFARabFWRlyBTKBtaLdn/zQ3hUbP/hvopPrF
RgR3pJHaxo8yZDzm/J25ZTflzGoVLjrEPE78kzsFRF0nn+6eQEtQXAw7Er7MFALz
NPTASGjaEDkFviijIUu/rkNPwx6iLjhwJS/TEeTfz/unpW4X6gY0RuOJOTfeWIGw
G03NRDXwURrcCSrE0Nt06lazzjToOVIxG6bPs+iOJAmMmh25PC4XXCtlKHT35I/9
Putr91bN50lswHPIgg2iXJb/+O1FPVPV30K0aggyS5uU0c4Pa2PfwyjMcZXY4i2b
bBQ80zavhjCqQp6eR5q5k7Qkg+44etsyK+hoSRAtW+8MQj9bYeftDf+Piw3S6yP2
phuYndgeORYUcVKU97X7FXb6HaVcDyLsb0hRJ8yLTb/YvFc9CcQ/gv8myTkS1hzo
xoYiWX3O0+BddHlPzs1oy7whhgOhyv/eGQ9zmyTsa3kTLJJNhxk08TzGlnyZ45/y
0kt45+ECMig4D0aQX6IY6XET7qP3Kn0Mg7t+uhKowkDpkyr2BckircmMZOqSDGJi
swGvdqwU+dwMsB/C2YwTHIsLnfu8yxd1ln6oQ/lrLwF8dTqsRLqdMInDPBGLf1hE
19l6aEw/rZAWYibtpQ0iFHhPChfLLd8DEl1t7RP+q5XhA4lue273e9gg2IYtryXc
9JSL88CpUz/K/Kr7E+0CCgrzi4qpeKYSJkfQkZpQxy9IXsK0vZjAs4pyRV1CZJYG
1vqTOlVuX8yZuxxo9MyoDSaLQYf54vR3+88fHi2a1pOAJrhUaqOL4HI47eXj/tzv
+NjNJn8lfAMxZ9gr3V4ySjJNSMgfyGZ4J1bplBfB7FFUUhkKq/wliHzeHopsikFS
l+DiYlVPSQ8YUjc8jYWtSBjeOxx5LN1lCePavKBkKznT4kUBUMZMeaHwhEK5oCn+
NpOgBiJfNQdj34LEimrgjA4I4z8durGFAm8jAlL5L9u/3eFjyRwnbrrUuW9z51rd
qK9XmRtCJmaif2Nk7myBHeSeYY+0Q73S5naJ9DyI8pOKjz+zJ4BfFnB/w+fNO+5A
bTQ0NIZVY4RBM2/FGUF4AoJrZqmyH5co+HrbfnprdzNEdDc6kvTvd8zXYkebdZjO
funbBVw7+JeNx0IF+D9kXRkV1oV2FYHD5v+YZGV4zVFn+1fk+qslPVtXHZup7cry
YcuCvRIeu9s3350wj2azqMazZken1bpvWAIrz5dA3Jq/tz+D+g81hhGrUlDx9bRK
F9b/gGUOI8ME3b0N4w2dW7CJisj9m3OJ3SHnWFR1bUftfUZmgO1JBQnmc8zI4EZY
MRcIbmxKnkvu3w3cKmfADntUK9D3uoxXAJctFNCgCmDdvIkt8k22X5uyF2LSzFQ1
k/sLz14vxqfXBMuWuE7hlM3SlFwAuxem3ADeuoua5vHlXI/fQJeZxInQf01TF65u
4P6HU7G72KdYkF0TFaV/o6npO3ojpYsvyEA7sNBdOov9rZtIIEUksuq1bfTzaSUW
dqCAuZpprzI2FIZY5f7PlW0fqZeIjwe7sohxD2WtFHuFeM30/pXvan/E+lvTywv0
6LRadCMuKl5UGP+WZGtG939TgHcmOFXScQgqG5BPQis9VzSZTfebv7O8mP1PQHkz
r2BDKwP/nuDQOUa4/wxqgXz4Dwa+i9PczmOCEOv/ibHIypkrJlSaWEkbwtUX8kKG
HS8owpWY6gwYngct5CDmnedURH7MqWzcWEFGmdioFiRwkk2wvteXVbDQFVdQ2ruw
kb1sEMp7CJ+65YFRbL5mcZh190KM9k1qzfaKkIrwn6/2EaUbiFkBDykVf6yFABr5
8WOfOodlzx7dtFoH0sGCN2gPjTafJe8thwLmsPYJl155LcQ3i7HUx/4adozDSW0y
dQH/D0pa1utjVGVMX3Q0knTO06yHhnRmyxsfjqxtjJcJvxWQHrDyPqddOdxP9gxN
O8JXG5fRz7oyLghEjdet1LpPIjBqy52j84tDEcC1A1jgvo+kldBROhPMx+txOPvF
zc946hDWDG9+ceJ26VA+7pJDXGE7wC8+8pEAZ3GyuQoqAbuOlzQn+DpQrO2E2xRQ
79iDk5ZydCkEfSp8goee+zAPWJ+XZMZprqmCvTfnKsc26jLrjUjYJApR4BK+d4zg
2KkWyqvfYkBTei4Hz/YlfjaIZrVv2ptp8qKZMvWNkxIQpAlPN37ZJVaHsSDELT4R
w5BaDTeO4VVofGbtU0jdrOJwbMy25NoND6AmWWK9ho8aDd0r97rt45XOxSRb3HLh
+vrQUKu5ELWGYfIbs6PCf/L8lISdilYo0AT7FOC04bfJCy1cp4IIv1t+JZa26S2r
xTcEd/3Hcv85FzvzXQeKOOweKNXvWZNGsXIdcVvbNxE6+GyQCx4Su4zqsLnZwll0
SggyOPqx5kCF594WoW76kII7K3WaJxsIWrzTw6/7IlmFNkLWpKaEfR8N+TQ89Hsk
uvwLTimvhyvCxDMHTlChzp4OyrzdN0iv6od4MZEAhdYHeznfIuy9IQ2646BxYz9u
u0mLdpYyCvldXHYC3ma9Df0X8BMk4te2cCVbbvbzuwTNwNyELrHd5yEbkXwVMnoe
Gp/+vWnJBy7/PqLvak/BwHG/jHI5UoCcTNoR7QHwwrM1DMijKHstdnExjgUaBCja
s0GdGTABRRyvea52nZ4PzYz3GNyrRY9i/hM+4uysnimWFQzNObUJ0evQOnDjyL/W
mADoDVfQupmiyRIJsQRSPe0P+9ZLh3HdcyS7UlavwCtMn/cunPeHv1xiu4LARjQ8
p4X/RzsMFNYbiA8TfV8dK7GeL5PG+FFVNyb3ZwboRSn3f1AQ7tI++zhWlZQqxTAR
tR8o6cB4izMZHvtxwb3ssmUfjKYQ+Vy7qlQ3YzuXnm27kOCk02g65+6/MOqGRgVa
2wa0HjoXGV+IPPXSvFqDFxTwnWScvM/Io9ccyab+LiH10AY3QZKQFKtfLmyDzCtE
hXedpvUxfdNgjluvWVxxTaQdrEXpKlcBaSvrQJPiH7W+TXl0ukycKfbwtXF5WKyo
g0TXBnnCt70+3dL6cL4LS0uK4rMjqRzzjMQJKD45zPlHEoDOH6CK/9w+YbHF3nMA
uuyD68DhEBxLFSbBRq/x26hvHs8FVQSssG9Jf0hZ3H/ChGGXkFwV5TCVeJR2XREH
SCGUTcPmylkWkoWH9aznRWl6I/2B5B1/4CgRgPRBZY3AW6zWrRodP7wNOzPpyUEx
SHUosY4vHPfglqJCcVjJ5s74xVVOM9J38uBt/+TqAMKnYtUYLjR4T6NhjCPV/Nw9
jrRi266P4SjOpPpO8CbmamGQeUzUhGcu6Qyk7yAfGgzHi4gz/2TpJ6l3FNSRPf+s
45NELgj9Iyjdp7xm4kj4IytEAMHUQ1pKXN9XBQxwzyR/r4gubxa2iKR/MMcNqYQ5
4TtqhM03EMsaBnfogT4igynP/BJSWARcD7PNq0bqqUmphxhdC3QOGJ0vZ82H58Dc
MZZ1Lq7Urc3z/4XniRkS+7q51XvmU8Ax7xQc2LJ/gbJZRh8U4tbIPPShVqpwNT6b
7XdhZV1Reyv8P1y0vrw9INT0sbxvgLffQOYMP6GE7PC4IUDfBNGTawRNepP0odms
KijztwsivGgMFi5VdX4AUsu6F5yAMvxOkP1aSI6m+eNIkortFiiykSURlfRznGRL
vHPB/XS+PpjhNvai5pGGRWZemjC4iDJ3voCxJwZcn0D0AN+WBWEtXeiNCsjhkddi
jYCRbLymE1F11WgQkKgsYFXpJPWn4//xUPa7b5PqvnP7EcQibHTLQXcemDqCl6b2
fLZeAflj4dV5cjBp9tHkd2+6U+SeeuDbBgcl4KzRAbkkkKdtUQq+ZnGzcFbwONvL
q9W1hJY89aMspEIt23PQ1pC561g+EXD6ZzGBOQL1Uil3tdTlqIfOJxsA2efX+pxm
VsIvgoYxRo36A8XwPZVPaCUm60vHsSlD1uJASrPHR6YS9aH2U2E2szGSw6Oers4Z
U0v2FEL8Vm0N794iRnlnOB56ItyhBALS/B9+3F0t4+AgHFwT2TQVMoMyZrQK/FxJ
SpwojhbPDhAiSECnA7J7FRv3BlTphMDYgLHnCHwl/+Mg5VY0K2zTwTAwz99p/W0D
TtQBm8CqfIUQ2erzjpxQld79iHUW+ViKt4VF7n5b0dnbYS0eH0SWLLZmloouAsrk
CBYjHanxsAVyZgX4xCVQeiB3yCDtvjRPvQpmpW9EWiDJSM5sxR4+AVoSgtmEPiJq
BoU4RrmaUMnijb2sj9Ld7ReFohwHuQFjagWEkoASHfG2c+QlEIdo3rGJetRGc1mf
9iY11Nk8+z8lC7h50h6ItEsFJZzLlTp0BQvrmxyg06+dZGMLEj8bpAddn//J661M
a7AUcehSv9TbZn8lNRRAxY32N1CnkO9uSL8j5pMt8c6aWHVyKbjlQF1fFdTWMm/Y
qp+EK7plWMB4hAxDqVJvzq06EApJf3OIPkMYzaPi6Ebsv5yDg5ur4EWq5kYxhsK1
RM2r4CB5aGlcqPgACloljRGrRxBugyWdYeoOoWXlWeVZxUrKvFcmK7VoxaXDsZnQ
FdNzZCXpGVuvh19mJc6XD1HjvC2OQ/koYEWBNwN6MbxM5Tus86VxLb77OexGmRzE
/fbSHxbIos0pLGt5RUWKblnPA6KrZM5oV0IGtpzpKpesDMW1DwMldjf0etyIdw3V
OkEnvrDL681yUsmo7oR80RwVQCQdtEm3KTNW6rbBEobCUmyPISJqDDc4P7F1GQbd
2JBdRcxwZVidtyy9gUPeVJfJg327Di0K+a21pt12f1KlKtgPv8koq2KXNOKxT2Hv
WXZ5aGLkKMVi0IFO/emcd2Wvpn9zz76wkqB6nXg/nl4DUwH469RMLuvBzIElw3Qx
XyF2rxc9UhOaHKzpk3c1DrY6Ytj64hKbxolRzWsSTlBX44cpZc9EwTG3YNSkanEG
WdX/c7Li+Pu2Yv/qfnXpqV1CtuHIsmV29nI+2kfe2xeI7JwA8sPQemOlDLhjfkjL
riA/vPm7xsAB2auNqMNpATbpBYT1uKNoZvNFY9KhhvpaTRZN3N9D52pGu5NusabY
LlbWky/UrY3zgCPkTMR5NxOAQiXCPY7D/1Ndhyfxc1C+1ZBjxT1dOA0CrGFegz8x
8KYNNxGVU//0G6fJLaM4jvbQoG/FcArSV23q4oMNXslrrtgcVnmd/tbjiL7DE06K
QyahGhhUeImQgu8xxmkBDzmlvG99HgT4ebTkZKcOyHppL/V4xLQ37MbnxOoZmwfY
KjpZzNbFGQz1tmVdEAXyQbIZpoM1oAG8BBMM51g9DGWUX1+pV1SSfHJCj5Yo2rXi
vGlROiANfTiRqIyTV3m05DnV4ExhrHoCBus3An4M4ftDqvvUIAKPJRCNe8kmP456
BqWpNrMpDbZI7lkP9i5winlek9AQOEqbold/rupS20VEcxWXyPyYYiRYYEex2em3
czIB7qL+G5QkhW7cmS3s0R4QDFC2oawmQ02YgOjzG7jsEmH2tcAOCP53TOmt26Pl
FDyueQTFbcjAKsH6Lqyu7an26LpA2Q7WbumJbeJrdyhdf7HQrRlpE1nE5A9nrjv1
aeXr1rQFKgdWviC2BFFmBI4u+EdAw/TfGWeSTZC+pe65MnrQIY/+9FJnaeyYkASM
SGZ/Nbj0eEa+0s0lUNUEzcgT4PUsyVX6nQ8OQEL6lB7FMCdzibtP+ZX2LlIUptE8
7/jP3eKeM+Z3zWIDJTogBUvLCvrQUaphrzB8+Gjpwksc9PjpRhpCx3gmHe4kvSJP
Rw+jdfWVAzQHYEHyZfTFYJ+Ec407S8tPSwX37HK1T9OzRCjlyjSnzvnY2cjg3zEs
nrmlrCjeeDmZt8QQXuSrKRXFZzFOuwlnsfg0e/u3cXB/fyq3Gnd98mMizEQFfZw0
YLhSkRs5bukHEgN46MlYXT1Z8/hhFqi2+IepjexoEeOO9yMrBZMtBYPFgnlpUoFG
wTHAIHXP0YeY+haiqPoeGd51VjTZut4s1+cMGnvybN3T/fzKoAnMJIFIFs6htqix
lhbdwA0sbL13Kvn+/qm2lSNdGXsNRCrLdDwiHIWnNEHUUWDWsUxX4n9KAFyt8ZhF
k2wp/h8Y1lKOqsIQTS+bXef6RvFLw6v6b81+p3Tl+E0NgMCO3SKZLTEsgV4jBaTg
W8m5qA+oNKk63sgdd9f7m/hpQkrK/KIbxjrXEx0AI0kAEPxZorLaybg/K/7t+PfE
r4gPgq7ZtxoIzQCBMZGJmoKGeZzKe5GmusplmMJ9wQZLtOUAQ4css88hs/kNT0F+
Bgv8vSbC485KuUk+yY5tm6AW2DuhCxBgTwhyXauy2Tf/dW9RTkyAMSPuAOiX2S3n
4Eg6qQXUiW8qFikiRmzSoZvtnDULgzlBYupSxe4u6eKea5YLyjxeU2TCLe7OQ/al
trJ7T2TZzBJ4rn9Ea/bLakvkATGZOFDFKHweMzWepB1Fsgeme9pKpxidd+0sSjLI
YvfNw32IkeqGpQyBBI6wFpWEamWO3lZT6+2eByh0B+uUPjmJsBXe+qu0UneF7I1x
Wj5nCVkgJ6dssgnM6aSkUjzGWKWF4g2QGB7OAQpO8+FDhQsHU86/sP13SX8lPEFO
OqDecQFhBr+olJRx4len/pQD/PfGrE9QnVGBreJtxLlDEUsWRC8BSjKUAEmYC7g3
zC+Z/zrr1Ip+JC6+E1N00+C4hrrz72bXx4zWfFFuccvNw7t49uxaKcuLfTlG/DQs
BUcfH1OZxE1li1YOyB5+ubKENSxTbyaCTKgOFQ6HBOVq7K3+xGPwhVF+tajxun9D
/Wx7H4Y83Zev7zUez9BeCn7RQ0wjxdoeEmoGgNbTv0yGeBDL9NkJMe94R9IDib42
bsEu6IHBj2NApgv8ZE9XJD69LbMTatkKqcVYLmPB3gES/A/60oCoxxc2/0vZ6NIc
0ceFSuq1pVqSVyKvjPxM/Ku4zOUHNgA05MtIjKGF9ftPOIV6s7MnwUuDeEMfpJ3d
gLJ4eR7TrQywtKd+0tAYdgnKWG1jlN2RdXzqSISSzktVIPHQi7J2yhFWzBC1bTxX
7mWi3y+RrghAopxtelaKf38k0o2nAJyWcxAi6e6gVPbXGe9E0O+2SvKaoAiftqPH
g9YTRrg8r1i1A6lUcAklxLnY6rWJii7D2yz3yRCtWNY7sLnEsuT3aZGhKnm9epfK
hZaW2/k2n8BVu408y4y9mO/ih9HmnRKQK8eWBTNZM/ugmm7jv3aPFmyAr+07skj9
stFGz50DoeMU/i+qXPibzHN5Zw04/JnH35qYm85sZDcfGDb4X8eTn0qInZZnDYep
2GjMz6EKH4WeAluuM4agFNhxkqBaIDR/DoeMNB/nEpdOXyIaejvxyLi23Ib/DXz0
diD4R6hCtHEX+LXrDcVA/cDu+D3weYhlqIiEwz0c5qIpua4a7o5xy9ziA9U7Urrt
utLqOcJ+9wn7Z6P9WoPr5pgKDtPVnW264Jw9SbLAI/t0N2WqzRJs3X7g/4vCCUY+
BVYWb4lXyti9TfC/h3Xe3Ut163ZkB1v/6mcGEb/OKZ692qsoDJDA3gF7zvXrM+R5
2i5M1DqDvzJigQGyQhCFNjl66QJmBxiSQMAGy50CvKSTrd4CACuHtAXJElmfAoUv
BwGyxLJt9tYRW1rt2h6qdaOgXWvrryow+n0wcVohNxMBFOs/2gkwdiWgtW0SxmCC
A5V3JrsYbx/XEaotVPejdn94j44BIlWWDZRGLH/8ZUhWqEzcFxdDY7a1chq5ENjZ
RoJRYu3N3EndT+81DoIYuNP1n4QKI35qO6Vt6u1UEwr8WLefq/3gG20vZ2KmhNYl
2X49HfJ2vldtJdxCr3gDo2RAFQxRyyYxxzs8Jh3hOU8dlSCHkbkfQ3skPv809foq
ijEZUtt0+JnCq9uWhrsyz1YSH7CqzKDcKpDu0FJpP8wTmVP5kZOAnPgOOP4S6YPM
x3UEFltREQU/CIqbHwuJWAj1pHX26Pti2mbDn+VY+1zLYIJEryXSGRCd3d4okKZW
oRAK4GUq8BH5/IHUxAHGB5fWYUVAvNnMHtnuQ1Hvy5jRubnwq5m8h3R5/qIcZFCE
5s7PlSXTULoQTZd5UxdS8YnDOsz5Hu5/DgitgdU/b3SoyrSCkJHV/8h3zXbnQ5Ix
3aAWDbz+zxfpn1cn1KwjXlY2Gm4JUyPkVGT+qo29kL07evmxPY8v1yONNyQv3sg2
aUVAXO25Fquqpl9vXa5/lrK1U4ggbVnGjixsgsdIr7kkQ40dECoH4eW3EgtREwEW
Eix20ufE5ehwOeA0pw69LIxOW+NNq9GrmPeATZJLxug20ZUOqDe63ILgbbMAFiA1
+F9Rrleets+TSKqnTpc8Eikrw9TsstfvfcajWo3A09jO+rF4ucp+f5Z93ZTNCDHs
/Q9F6trg0NP7jrz1qwDYVi12Uyr+kUc0R+yfrgb/YOGY/39AZJvLQ+HJ592UPXW5
/ab9EXZEPYiFpZtZ3VrxZh4Hha48aNPmFwL0ov489skc8F7+BnmEQPgEqtJZpLUh
UPfv/IUdmOdlNawgB211LofgDqZdGSeDCunbt568wmUv0JsJz9/CwZ5cLFP2KUZM
mdxPvShK7ayAZ47vfj9I3MmLvbQgqQxCo0Lc956CCoK9l+hZuPYEDvHD6eKyGk5O
x1BaP5/jdS9NwOnGqaUebVeFaxG11lLEXM/7F311xrQv+Gbr7RLx1xrNISqWS4s5
S8LJlf1x1MapFlnygeQhBm+VXzh5/e47HpjNdS5Nq697XlrNISHNqzsgd/3boEad
XELAF+Y9vB6SVm376qzK78Bv2SOoPUR4BZhNwnGdgDpJZwn5RvKSE5tRF9mmaOnk
49XFC9FgmB1HPAaObZI05wek7SjKV8CMv+5M8fmygPV0ZuQAi6TvYq3tihdWv4Nz
EdvmBbhEiGRML6qJNApvtTzHw3sh8tEVL7dqSBrVC85cVreyQPwXIH/es+w14cVN
kXK/BLE+N1rehMTvyjVin19WxOqj/skXliMm7AHOyNQqWZddkyVOFbjEXOjceXhl
Rz3DF1u0cHLtXwpO7bXnqmvWq4F5SgBSpRN21AIA/JAoc4u9og3bKjNQHwiFzfz2
ZYtT0G+oLiyM/VsFjBT0BZjumMP3Hm0139YK8GgTQUpGJ4IKKJIisrzik1wxINx0
rD59gGYtywj508KAu72H0TkYcqn7W4cKaHI3ZU0rtZwWGNCIiCXfDFSbURU3DfNa
kHAGmgEM9t56E38/WB5IvHtUEAGY8IEpdM8F0FQYmiFFrdyY/ozHlWxdMFoyiql+
BhJAny2KvawtudfCHWimFHJPa1X8VPAb+eJwJ86KXqqDC+WOYoSoD7jG7+/pObNs
zre+jnsZPRyQCbqPNbs0e2nUd7hhwFtk3TeRRWNPLMzHVcjH1BNycjZCb+wJ8AKs
6rvTALRnk8YMwOyFwdNaI3SrMqewSPo24Bbu8qsTMyJ57Mt2HURERdHkVPWBC1t/
6UB6Cr3IhbTZix0WAcbr75GcEKg9R7/yDKwoJTgu4UfOPHsaeQ1s6ZKhjrtNrC0o
TMLSYF/0RLrxetRGAECancojS3FOZv8vbSY5nbBVlI+JwjC6gVYDcI2wwFUo/pli
5NIdNOCVEqOIaC//ZHNNuS21uzKo4SFDUxo4u0UBR4X1JmqnseEeUacVCnetZ2xl
IMMVqjlVZNIl/orGOGC8e7RK91hYzsroAC9WK+E7zC0gnH67lUsyX9rdV+S4ptQx
U88Gg+0dWWRWDWs8X0bPnwzPkwzgem8qi50Kk5O1YljXEPUJibCPsnmXnFM8k6BK
1b9AHK11YpSNpHSwPEMDeYRTwCo0Gh0jCdOQMjSsv2Sy98Rm+r5tu5yOZTNoYzeq
awJulCdmRFyMnlbw8zNzopQexiarlZ+I8xKQgbO5cpA6wlHqI1CVAb9FK57LBAAJ
N/BLee51VFwyTh80Sz9/DiDKE3ySRA2T8q4VZ6gW7/7fqUj0DfmE66tufJRXwkxA
5qt04jc0UDhgOXIMLOUlvYMbL429zwDp2DEpHR6s8AEikTJwRadBtEuAfF3P+0FO
WerwXDHF35F29OWh1KpvOZLykGRPknp6dmMiBwyMjAMtkavIoMVuQPavxnBGqQAX
nIY+sJuQfRt7bM04swtxYUdEDmgbu70H05/5Um4E0RPEe4h4ibn6f+AILeoeihD4
GF3hgLzh3Eg12tUgv3tx8f/MGK7sBTpUavpdPQ8j8mKY4V8GbMt7zPZnhy1aazgj
DL6aYSUg0KMmfL+DD6lW1MmhG137bPiKcGTN8x2Dr2hkcNOOE7zFUZo7XmW9H4eh
fwrswSS3xEhjwgr49kka8Z2WCElXoapQZP45hi1HdKsFsfE0XjDv0nD5JQR9iZwn
xOZXWWpr7NV8kSNuYHnFU2GvOMnWIKNEg/ToP1ICFWesu1L5IL98GFqWsts9W0Vq
cTnLZ4wBbNheGNNo65FsJ4bvXAPFKTPEsUlJ/jxI0DYH46z1GxjS3I+F3A+LBuw7
wXgagsXAtFUj348hlJ4/FaDPtYV/QLWH2EfDrTGcwuMjWPPaFZKZaopm90qN5ddb
NAH21RCsY19+bcrOBNyoU61vKzBqUetW6v1EdQNW7wPdjMKkY2d0mvwBAvIRkOI1
plmvPWVFAs+Ks/in6PUd2LPc0/25ZWxAuviOCTMZSDPOakAB7Gw1PQ9ZG7m02iBl
7Fwfl+P9EEGkIdRZAHg2MHMpqzXt33E4A9JaSl6HCXx4ZyLoCx06joV6v6B1j+ik
JswaCdf2Q/AbdUF3UetLERquzwFES5+dRuk1T/j5T4fqWBHcaD4vfbpUyp7Dae6m
5HHRVt0D3Vm2MUe5avVrcMYgN+j+X6AgzI8nlqxwyYdMM8GaS1AGLb4hfVSiNytC
GAjh/P5c1u+PlCHpIcW6kenV4MLOQoovdfRFGvjPy30VhM0FF2RcCULJW/7Jx+Vz
Ji5dM3/1NQ+C6whZGt0nWtMqI9uIWsePXcaOrXwTaNgg2u69bC7ZaGK1EDlx+Mmr
EbkdFdh1lwHH/BT9cJ8zSJkD1hdCjgyDT1AednBHT+/xgM42Zq5H7LeX1tsTh6Xx
xLrsBVwyARBQayshjBUp9DWUmye7UjoYUARKaspzriDMZ7hPL8JJKrx9dW9+EFnH
EhklqHtXp+fUBmUo11WH/eW3foQGLoIya4ZUHhbta/n+quy0+AvDX15+WErrJ3c5
cOIHZUWUrvR/JTCTPXbEja8vD+67tjCNAkzFVg5sCttBh8lV+xCBfhumk22EETU5
uFGyWbzVrBxXCACuqqwCMSkMnhZhccDgVX0YajjEAN6y0LWO/eSf9jem558ei3H+
IeT1WcVAJWGrQwJxSEx2Kr+mE6cTZel8Z+w0R5yuR0zbTd4rcTkuluMdiJXs0QT6
zF0JCbkM7mWG9P8bMLxdSuy6+bXQ1VwnDKiAfru2Md25KqQ7KrQeAW14rKt7pNWn
LmFhk+/SwkDKPnTSjGn5pzdcc1LQ/fDBnm9eyd6ISupDHhsNnaPrF74LKJHQh2S7
5NAYFLtLZRa/4Qk6IK6GNu7jf3I8u18br1lU9nNh4U7n/72rtK7mBO/ScrFdh8lA
vO6xfjofTXmsLZwReo6TzwNUZ4i3ZQPABBFWOOyBsdtgUOjyuDls0YY3cVhXKOcH
uEItjryNnvImxriCkc8h/Yq9xm8RC+oun7FXqJpOpRVPmbMSsMCZYU5ZXfaLoBG/
kLxA1EW6awr0D2F9gbJUOThBdDptNjOloE7X2NAyvOIeuKKO+CM+XFOEl3HrSK73
QtgkR6ezd4xK/dJ2iXEhzQ3mGcdsW0TS/UYiTg4S2IxLNmpG+Y1ovwGyq8/6HdIn
w2sIBQ8OKMmfsU1WJab2WSemTRFAYz/KvV8u0zRkaQJtvbetjoQbKfgetkqOq53C
NRN5m39Nqm0De5Vl/LLAf5sRfiEZz1fLuC6mwhfSrg3/CDzWtXmHeGTLQYjRRBIr
egj+oyJxHk8bKsdClkryPZAcpVtkLWlmQiS6QT0JBA5DYd0IBFbCC8Qu3pSvuHvd
q0ZWHSQ7JQ/5Z/JgcV5zxago162WlrYrnlwLCF8iLuoXtq4evkEKigHJWRNqQfpB
XCZHJrMBAcQWchk9t6m+qJlNtLLEv7ZMxcjccUYbK7iBl+zIKYli85QtqT+rI/xX
hqHRC7Gjh8S48h60rG5Io0XSqP4+Jsl7DV/jYGTwK69Lbq0Si6vziaoa2eyrEJvT
YOXz+yKczfA4UB5WltHJcOczBvUwloscZ9Xqwv3Xhr+qwFzvUbauK6A+5ks7a/bP
QDNzMViHQbeK0ZpU6cjPSsN5UfPbp7NBRsV/3IXLdq4Bzqdez5a77/UUUDu5xGZl
1hGI3sG5O6xmrNoOTJ5A+Si/Z38U6KL/Gm2h1yjdNgCU86UUNZ9WbWTHVD0knaFU
cSQnw90KuFFf2JtuunQxBRtQ++bhEJOdOX8WPB4yJg2rz95QimoIM8njWnixQSz+
7VZExOTWBO8QrCP4itYb8a9nPLc7QaQbEBgTD6Cc8XN7GKRELCRPGmDzQM5h+6ik
u6FYK3Q9T9u8hrOD+7fQFpxDz+01hkUovcT57KZaVslwNiSZOjJowUNCoeO3e5UB
2DETLEWCfE7CvPgFVBXbEkLb6eueIBwFUiyLOswcsnRuZAf+ftugpqs9h79nwh3K
k7lVWPQ1LqG8qHc28p6nlTrzATF+oBV1OAj1B+y3F1EomGSwAbs2N61P21n5oMKo
JSw7g3ZsOOhDPlAfGjSYMJgB0YhMVcAy/OFA9lAzthdmVdBS8jJrQb+b0kHYVeOH
nASHiABSLotWkDFCcFcb6HKbPg9vLYuwCuYJ3oOsBrTCOaNa0vk0kQdOCZCv9j+G
FesMPI76VqHRrd844kJJQfL2ZSj98ZjwLRxUGDkNl+PURFp2f/7WNSbwzweEKKxa
H7q3xCY2Lxzrz7lgE+X2F0rjoznze1YwAKjLXDVdVque1RC5hErtmQ9Ro3nfvT+s
OBzxFHZkg1H373w+dR6la9hkXFe/7CLgI7vQ5SnGo9erASRks/pe4uG//Dvy7ovN
9V6Oo6M6p+TovOXYNEEEohE+bTjLbnEBQZBEosvqVxLSohH4jAz6CQ5jdqgMRtJp
9y9Iy0/lKxBXkhQZC7bkdJcf0AeeqsOaU0OO/UrCk8G6Ox3+XzUQqr21h9SPFbHq
rGw6Kiwjd3EHe4UMUEjOc9GQqnbzUpS2p9Dlc0TjCuCTpMNlZFlXwGlSNXEKVQtq
AKcxhMWF+xLMvuxnM36h+EqgTCMHvnkZEVdvdnpTXIZ2kC0d1ZBF4CvYcpyWrYod
h9uNuQgLokV8gQxzP4CM7gDlMCukHWbbYZyyPy0135iNCHF1kIWIGmU1CtZZI/cK
wAZDijrzCzj2ZU11hs4On8JiLNZPVQS04isg7UXN+Rw8K3w7j+vFuVFuf3u/Yo+8
xClUn8lqyEtKaMkcOYSJx/PKt6aihidN5NsuqrcW5PCyhAVlmbJUs+31PF3KfnJL
+24pIkt22Tm7NTkD6C32AY1PtbPQ0CLcV02SmWxQIkSNV+wioXHWeWIlEO/BLktS
cIAgiTLHPqdoDjATIUx0IRCf8ZvtEFo7deWilfj93WVrcwVOtVEqpT4LmCDTsm52
jDQHAgv65J2ltIipj8Az+HWHWoZ9hVGG3BVgUFsPIrPIYXCDk1H3yMQCISym3Uqe
WR/2oCVKVbcxhO+10MM3c7S3hvTZmwbiSWT8u3Cl2IaQUtJJJfVSHKtnoEJhyMM1
dYl3SGsoxAfudl/QTm8UTzFzBaGi5ayMi/C1iYj2zmCSGuWQF+fRhN1ZJMxHmm9Y
fwtE9oP3xNelPNbOZ9xBhrnMT3Nl5jhOdjQChtWd14rrWLCDAwHrOFrGa59jqtU5
uPcFLK7v+olzUEBu/ro13aHXGQNF2h/aytiIIbawnX4FOT8bkFlw2+O1rM9Jj0jm
XpHMbHvpAkRK0U5t+dkrZnoT971ihv/OZvT0effXvTian4mP4PEKWy1Dq0Z+CSJi
svVwyRPx4UmKVFQ4cxEV/CHFMQZW4Y2ilDMmz/1G7xXMHfHXRicwxqTjFyEG5wXY
o38mSVCtPxXilr70UWHoBlyaxa/JZMTpswmxtPbT/3RhLViEBZtoaRX1DRfHvdR/
hhiwxKH9kzcBxKlK25FYayp6/oriqaQ8H7zvw3xQi9rFEne/Oo1LYwqf+DENW+r2
ntUfh/xRf/+6N8Z1eOtru9uWaI/IvikvXA4Qh4v3pNGlsGVp/yFYyQY+K9EZMhe6
MqUnvU15uTcA3Dr/5RRVxo8C65cxuJhI+TsoQu7x3qLlVx6Z7laZUqqBd2C9kIyU
AR1xaIS9KrS44UcSlkB5ldRUsegVwqsTuiBPmbTApF2eVrotVEyIbAGMuTBnGe38
l436AKmp7jAkNsaHDGtz4GgndM7GJnIUmTCM7NM+u5RXkn8tQa2zxrUdZaAO1wLR
cP0ReFk9VbZTVhkDHqFn1V1GJPam1owFZF1JxE+zhjPSwI4KaqX28ohhLxWobuLB
vQ/h6Hv3FXh4PDqS8ZPwere6y8KNUeBB9OpGx+5S+snqqchqCocBxY2sQvyNsiDL
AR2Lo8+nOoDImTCFY8LrNRjzFtRmlpSuk5SSpuryGh2qIazXqfCliTwKjndWhEDN
FdZ/FaoHeAx2+uL5KXN51bSWb+Tjx9DZGxloooLhXIJ1Q2H4lEBoCq2eDlZc6PTT
LUpFqI+sPa1QidGNwXoLQSpM/O4x5/KJfdCcNLwGW9g8yMn+7CeBjf3EuPsMferr
8uMCpvb0VX77wfth19nk7rFpOX4m1slz4XiD3UWBZ1Obc268do8QgTnEdbEmnM2/
z9UTSRWv7Ylo99qTqJ/HI6dBjEUYInUFL+C9dCElaINALIl/TSVdaf29zg+0BRnn
a7oeODyqbp5nAeXecaCVPK4c2Uwt/xh8eS/lncY8HH5so8XXmJBVZRx4+jc3uWHI
fq/FILd7OLRNdmAIzPNPO+KKsPk+Hwm0HgPD5uO7iTJC+kPapLsS1ATDYjIJexSF
hyljPL6s7ZT2ycZRicXxVLd/sXy7flMz/ywzxhHvJrTso1AdCzwdICCNkSHqptP+
JQFMJDC9msUJtq4f1PfQeJG/rD3Mw121Cvii4z1to0npSa7Quoky6PNLDQZp3QKc
/NaX8J0kpBJFhn0oIIBe3V4ozn0S/nTYIgnbz45aD9szKsRBKyKhqg7C1BUbtydt
5iNRkgf6t4AVRptREL5HYXTee3pHQ2awbURG10WT4NS4eZhxLmXDocAfQPAtXNS9
juN+2QUBytFllpY/X5asgzI90G1NcBIeKgPiY4T+8iLXnepp+apB8qI9bh7MEBcg
xGqk0g60VbW9ZR/M72GRj62Wnjk9cyThu6AnP918Bz/L18qM62Lt9piH1qH7ACgX
aOuX5+skT+X/Ym1MeVIxh553e6HXppzp7zHZ4CJqIRZy4C9PxwyYtTsAl/H+YjNG
kqaA2taGussJDfkSgZoIPip1GSnmJtlMPF6jARetQAQYqP+TBpzE/9DXQjp60CVC
gHcA87EsCuvu0YrDUHkky810GoCjBG5INqHqTvQRmrgI/DlfUTgn5mZ7DFt7wg4q
1Z18i0FjKJsf5c3AdQgaUKpLghVhdkiE+M7id/Vc6ZjzqgcW8F267vMm41u6GxNT
uqH6/kPqWhyBWZVL59eLAvWN50I/flSDng7eeHY3t4UGfdnId01tAdGz2NQB7opD
oz+x1DtPCH73uqpTNjipSuqxVxCaKDUSeP1holylN05pOcXQ1eXP/k6P/lQ9YL0k
bCnPgzJmZINjfBZC/CyhuZs+GSGa42fVu4lOKAkrpF4hVJsZQy4E+bdPAKIsSrRn
BMWiv3GO8ojEgiW1hGrTOavsUdKqtooAjQIKZT+2thfBgHKpyW7s7ubv8B5ib91+
Hq0TCADweqodvgNC1LyzycrJYxgMsoVRl6Sgh6Sa8KcMJL4wGsjAYKkhvBvx6LLO
YF/+p80/oamK54I1jMm7bP+18C3rgkwjxOXI6YETa2Sby+43dduOWIfiaDeS5owD
nrZ0Wgeycso4Tdby2cuZ6twDBvSeWeYtfDmeplUijKsVnThFlrjxBvsNpWJIUCET
i9dHDreTgz/5XuA/HBOnxLW6ERc1nB0r0GCCSOAhGPeOcFaBWiRbAU9xB6r22jDY
ANOdn3HJwVvQjtS1MuzteATLKP9fHfcdJXoYvKwIzwEmhuAe1iioFRvB/D5w/3kH
EHevGO8AGODSBXDFeIf63MnW/lLPXMAGM5rnpW+2bnn9BnwqD4TTCnBkqsBFRMX+
Z1rP2KhO/xJYRFRo2pK3yXNUALrMRUacUxQfbT5YSgSKkZNqRdLA3X0TaophtS0r
J1j5KuzKM1KNLPMDSAkpEqhIvDbHUxJEXzuJNeLDcrVsYc7eu758x0e9A6TdmPg/
jNFkVfhT2M9cOak6u/zN6kGESdksfE0xLe+3sji7FrZ2hraNaFSNbzdz8IotgsZQ
QNUK4dtYR/gLYDKBIkzfRs1Y68RmE8D/PDKsYLA1XGZqGspCqULM4/t0YzfmqW3i
zkclUIgJVhVSf7K7Ja69cwHMe7YY/afYLBGbUBunIOM/erb9LN0ieLeFYxld44Gz
rouQvH46U3c/EGwDIEt5h743uTT5C2Lk6xTP50zfaemhoc6RUQDunH7+L+XJJHEA
9AT7I9nI0+F07rvzVElWOKxUidr6oR7vgtgD/twMj5B/T0Z9jMrCRTJ4eg1m/4HN
9kEIzAeVCqa/4xxINNXjEsh8UJy7cBSqN/wIP5pArVSWGsBXIPPqu5GgtDwboB/s
vfdirKfQyOsDbKl8QV+9XvrucfJm5R8vvwYSB6GPjjLhDb0Ol2Hc+naOqYjQ8R3D
i+i8Wm5gKFN8FRDQZHjF4FUlywpIWRIHA1pnDZbgPg1BdWJuz5Ll4dWSZR8v+Xvo
29YphS5ps0PKPa0VBp2BBxuTPjN67msciinkBj4yIahu10HvJ5ZgL6dpnTz66why
fDCUmZ4nTofZN9lmQfYsSLKXwun61Ha/JPItC7Yvm53mmkwNntf4X2L/BLwMSPD4
nWpJ/vIkjVYwAhbumRNQpFhkXeiXTUFitcVLTUve8n7G1Xjf1Elz6brR/5GG9ieL
iSbN32XAjkrkPnWaF/wYB9V947d1fCXSINUSEbA9nlNSdqfP0Ih1EYNDD/0/gDpR
dU1aane+5CNNLmnR+Gah29nRhEw83DESSSpcOy3WkF8ODNWU3PI7ivQVA9swhkZ4
rcDWi/r3R6CgP+Zo5k9tyYGyXe++pUBlGHPTkWYZP2wUk/MjNhTzPd59A7X+DPTZ
Xigr+tAyQBzuojVJ+5lsnoUCMk/b3TITTVFeP098gq55tzkqSmclhY6N5sVAU4dT
XiDh4XtA/Uuv1zCou5Qhy5IV2j77HHB5xPFaQg2UUz1LbagMWAPUHRYn0PbSr+si
KTsOK4tgt7WU9b7RKlBC2gwD/l6y3hbClV282ZhrZtYczGlfXqElo74YW3/tVbPE
e4HPy1otgUB2ugJBJfWr3PGtNaBFvx+ZjM9oPm3iE41l+jA7a0pW/lUR5icoU2tF
MPoGfWFJqZMJ94kG64ZjlrtMoICV6/9YdtFIrrq98VKQ8uz0iSiGGOW6bc1ngdwN
WNDQx/l2dlRHDLVEMTAI8YhK884Uijp8Gd0XxPOtTdgZa8NurzvAebr4q2cLc6GN
Wl6wsyKPyMyDXcVOKOFf0O8YppcrmqmECVaWw/MRVI6SgZWK5yI4cbhD0WKb6r13
fpFNzpfsRLaNAjtp5CzfLsHDpgjqr81ofl33HR9glfdWPcGcNaUcKwdwB6aQdQ9P
OG1mZgRAVKqTOkfLQESVFj5IrTdvfHjGKE9yu12/VtVqqmkEpLobDlQa9iCeXytW
v6MNTn6wjrXMzVe+ONBYLGcer5Y1Eoy6soCo1hCbn0WgQpXzUzGsrzy+6T4e+jjG
mTJlTyVWgw5B5I14LRpHKUNHndpS8DKoOm5+eVYT5v4+ZDtRI/07IYq2d4H7EE0Y
YdzCxU7RuwE7h9pkic9BEQ9dyEX/3e+YYiU/iwbBC/eVT0OlCOnHQDBwF5kRvBUM
6dSSXMtMvcc46yrGgQHpbzRVQDzM4Xw63vyL0MchSw9AmdhjnMmuB9qQ7iAkkvON
qHlNsdmmKxMnmXdoT29A8VwtQ1icVMTN0g/kjbB1/HsLOwAXSTQt0u1rqcVQ97MS
N1i1f7D2W3W8k0crUnlVgXS3WHCS4nGhp91Se0fPszTSaHPEs6L7rR2NqUWpg1o9
2yBo7vP49MS9CDFJ2gZR81SZuUtTqCH9funllpo+wNyXp3BbspDHYncQhEvi1mxB
v/fWzWfl7wPK5VKUmlKa+Rr10k3/QReNs8RBpAeNVU1cyeFyy6YZS3ug9W9F7KRp
fXk/GL90zxgko+AibVQpfKaIWGzPY8t8mu0nJnZDC+K3fu0/jCN38+HiBks7srMN
oOlj8AbGWy+HXDBQVJVUORcQ0bWOUgyUfjYygNN8yqmsf64yYM+6W8JHkPN9zKQA
AnG8QEaw1HLp+QKnrLvGl9om8fidqA60iijekz9cY99INSC4ALDTx0VyFG5PdQu1
6jP1iRSodpUGJHQ3QOYasgSlV8oIjHqLaPzw+Kptnt5p2fX0qIeUaqS0xdJ8MO4c
RYsvh9HY069yN8J6pFgJm4KORiFkGejDKNynSgVJBHLOTQ8jc/QX6Sq/pMzgNcjG
HVk+82aeYug4QmJ+tYKqo7yJTyJMz+noCne3cOVp6IXBKidkBDWz3h//xeaB2k43
vCgSfM2XwTqx2pd1EV9K8cNXkMfNM6RqnKW8R5E7b035/D3tC1DKmp4yWiwur400
KOcsrxaH1ZLVBoH8skgcX/Dzn1OdTpYIo7ac4jjIb5IW1QMcIlPCynU9T0NWwr5c
7TmElQRZEFsunImcyS56yGa899CZ64oQj2hLLz4jq13RY6VQBCOOIOQv4NdoT4OU
ulaJ4PwsHkh4krRZ5PV987Qya01HfX7yGPMemDW+o5EPe83HmvGjb+zi0ZbftGQy
UoePUDznq+zYY/NhPJz2vZUdjdhuj6uiTLDWdgSSNhXVoVBzekB658/LgqFAHLJ0
WXxa5n0WQjSqRzJW1hH8DnRx6Ljz5IYFjQmNZZfHYiH/o5lmhsxSi7TKia9LMTEw
cB1Sm0Sw+DxI2wMhTl/nKLMVbMwHPsdeMZYoZbZNVK5Mwek4MkQ90LBK5Ipg75r/
GpgyjewbJyBq8cMkHJTAofQlHUUVbAE10maWyHBHo0tN9vIZlqSZ4vwVpOc6SGQi
K2c8YmYCyvJwX+2qdM+2mdP+m2CFj7LvAiGaoHC4avAKVNrEgUYDIU3AhtdPAvTS
txjq4AacCuz6H/NMrDQbxSShI4ss+ngU4xK+tfTDuCMp8V9S42DPezSMunvmENyX
hPUZelquM/HMlJLCV4lUKCKcnYMHOCDwAdgNrOXteU6Whu1PoBrMuJ9scoOqF5Xi
EZ3pd7c9glybKVlUrw5vro5tBGzLCQX2Obgm0Yrh6Dggp4lIMRCws6tfov5mUw1R
QDEbpSqab8Z/hg/t8Aw+e6WoAEy++o1zMWM8EIh1O9bYGA2ta2Nz2m+venFww6A5
77MsQXAktF/NsrwjWorVjnV5u0eCTNZnnpjGp82AHhKaYSoFmGBD0RsfC/6lyACi
7wfwMIZ0LDVJrS3VKoEUwQkXi5NzC/wvUndKVPPsFMD1Me2yimHpfHkgK8M8AHeQ
lVHheESXqKDjqYrHARccfng5MJHpWdAOQ+ZYPF3mFmKL0dhJBiaNhFMBiHh1cZEk
y8CTORIEBIjBrGxTQ9Y8ARoO7ZFdt0EWYFgBg/FHBv4E4dVZH6RRjWZNgpCldWh5
f1uIOdr5tAfinEr/wGx493rYzee/LEHUSopb0mmWwUZK3lEmU76nOaS8JIyvY4ng
TLaSEsA1FWBxuuyHKVvt9R2HN+kp0njiO3ouVKGqcp+6o7mR04Q31pYb5jnw7wU6
kea72qVX+RNgX8YPKxoLWSK0G4btNUtQD/VWfbw/0Gla+aUTLDb0GoTsr7YTnqfN
SUG+fMjZ/4nLUVQTQGrAGPkZECZkSCxsJ8Mg8UadF5pd5R7DI6zG6RbDYdfEsMTH
yOz5Ilz8FtDAa/wq+naROddrDBFurhatFP8tc2e2HgTOfhZhZxQWFBqAKvMr59ah
FQBr44i9ownI0A87SRYKnoX8UuWbLx5VWB4Bw1ZOph7KCko4gp6MSsTG8Ayav1Iu
zjp9JsxmRR23QxhJLcjepJiEstsUbnNYi7iv/NA1gpVk68+vwyQ72CocoE+hPCnt
jP4IGLhqlVgWOVrnNR9kVNzs0apRHl2fU6XWhLiZwmCdDb66kaKXQ5gv/ZmADyBU
pNWRYTAtTREWOZ0kE+3RgpCTDx+G0/5ft7wiReMqfDJMoKMVTCo+vno6r5R/chEy
hl8dt5HoKXxitCqt/aq2Khuo/eTghhQfky88dmESCc2Jjx15YL75nzIztTP4KFBX
VIsYOu3PCn8KZyfNh0RTEq6ozgG3uXvU7Kdh4jFWChNO3N5fyJ/p/d4sBNYiBGRk
q7/gisvlhNhEdt+nGGPbRazlK7PkBZMByqCUeljJU3ddhUa7RMPmoAUvDhKnssUZ
vgnRWgAzY0GJeP/fKJUWhtSJLY4xVvyGydxt1sdFO51OUfU530d4NnBHqJqOsgrz
UcdACvSlViHLjiZJ722J7D6jplwiwRjYFnUbiSHMOAHiV93NdI//Ffff5dlp2mr1
fn87LPM8a5kugCpm3/PwMip52XX4Qb3CapZxiWGSSDGsoEiWTv6r0x5qaal56/5J
34xaTI78eQ/vviKHL0DyOKJgIiriPnCuy/ggXLHhYVcwNYbcriIgY/ebS3RFv44q
rgNRVmFa/4J3dPjuYYlakpWImWB/dkl3Oj2hq//lMOHcyKpBmhZJVZK93snXhkId
Cdai0nk88CmTFo+Yn50sPgQCVAAQyreZGoZLqnTLi5OH4ebY5nUYGVNyIb+78iae
XFcewAJz4WA+fF2UL7zxHfx2szEMhuvKGZi+JEISfR4JAChHsrEBxJckJR4bmkdg
kLNN+SKbg8Ufj+liJuS5TQLcU3w2z1sgE/IIRG2piMbiu8hW8omi7mORZQmpf1bY
rGsttxlzT+S9n7jPl8rfvjShJGOc2odfCYfqc4TEK3OKrfqrl/TWP9Q+DcZipaeN
c0yVbuAYShXzyT2GLnmEm7usUALalsADX2mT4PqHYZFxAsfMwpIQKDQPbeccKzD+
olhnogT11V8CiNqZIF7q4n4rRw7l6ENOenv5L8xbJbh/qiC4K44cNXMSGtHI/W28
IVfmgcIh+Wp5FY32NP9gxMx1BIEMWyfOq3Dd0TnGXHMiBTLJJb8fu3wq/v6x3DMe
WIAHDWFM/AXBbEFq1w05TOB73EaXpYjPujL7fRPWtBxzS0ixbJMrQJqJEPWutXjS
2IE3FAGJBGZ3o37yRUtIlUV+VTmXixFCfhSxqJWVOyIZvVpFEpOAcFdQPB4SW1qa
40i6IxZ/ehhDfUV3/Rb+7MjDk82mQIoqEONK8LnAU37yzPXFDJP7Wb5PHeBX5qFY
W/yEyfQHoSzTG6EYnICRwiMKAwtY5PDdyZ5/10aGjDTO+osge3gC25aBll3SJoGc
gVID8/WVfs0kvMfSh2Y0TI6HJ46z1I7UT9hysi5dbOuO0uQ9Paw1+pOMDOafAIhg
8hrWKKyFma2v3ezL8/o6CK/W9Zg/qDNdo1VbR3H5JNKG++tEfQ++brSqzQZCezUn
q4rRp8H83iaq3UW5dsyiMStexDWG7ECwiKYERpepyVs9Q1WeUWy/ljVbgIM5osH4
Tkrhan3waxE8791d8A2RaA08nLkgITmHTJmHpdBMD49wD4GaEPvsU9LAtUPqYf0T
NDlz62mWrLgN9UAVS/jSixfHmDqP7v3CnZ2LIps/90Pge9jlVEjIQnuaCmv0PPVn
t+83cY9DHqHIEkZG7CO3sIrCRQXfAwGcfRuA7Jzja7YATx3cujs9FlyClvyx296C
VcIMohL3aFgBg390i1D4WasS+oPIU6H7/KolCz0eT2W4K9yweHs3aqzLSqMo88el
47QYn2OHMsZ7oMRxMBvsWwnLbArmylWp/EQihVnLMtMHz4kc//EFCF65GrzYUFJ9
mIHcwazy4TVsZfb7zQkytPHxzsMRjWEX06rBYGcGcaLKUgUKKZsufK29O+PxjOGy
tRd4MtzOWTnkALgxQ2GC8o5rey7Hmsi9xQve0FLFO7JK2vdBo7GVG8UA1F+XM0kM
kL1wgFxfUidyJomITRPhdzYc0gXX4gb8WtjM43LAjkzdq2/24fmq34h2rXTq37fQ
NfompE3+entRpcSLWNEGxUENyH0bNy8C2tgdJWlmzLk9kiGO3uvydKfoUyvr0mET
/ILcrEjFSb7TSEiuxmWoo0xLp3BpT4kFcBFWz9NZImdb1i5FBY5M2b4CqFccddss
e3HKOvALJzMF/IKBDTniT0KKbZhXrBhcUGjz+q2vIDBxjlhrzP5BMGc4TQBH2ni0
kLGQqDiYLj/S76ULXGaXtBb3hjhkb9OwQ9lI+v8FXYaN/7MsL0LoD58nSph2+IWa
LW5fXYDp3lzfW9wQXblWlOaUXus4OI8NmuKX63VmVnS/SlISPUzUx7SJAQrsAV7O
cm/rYpV33FUmBNzSw6gcAiHJb4BC6KRg0dYV480V4v/8vquOiJCbL9dDTUpUyX9b
eqLAni1fnXjvbL0Is0BRAOXN31ibTCSEGT9TGPUwhTPsndxV3cPecxccWKfn4rNd
TXADg7T2SHZlxU66hjXxuc+r1b4A/ClXSzzyOmypnM7gXtoj7oGNx9kFgnrpl7yK
P664EJG7u1Im9Huu4Tis5zt4OLbVygRha9VQLgigXy3fw4H+idA5/kNAY4iEn5GX
1Dh/vdWdOEQ+4jBow1yA4U1gcC38v1qmByNepThzm8N8y4nv9HIagFuE8fa7dvuC
+WZrtSN8yydfdhg+9IMPsXbQ2A5mVXRKHKbBmAayv2XEFFcEhtykXiuW32WZjxAR
4LGFi6KTT9KGpUzi7HtcvAP35NiAUUpj+5IBMX+bvZdiDFpnAO+EkwYXDHBuOJaH
mSK9+9f0nE715yHpDVr1zEIb86SuNae7AIRblUNT47LIALBF+5LRO+DqX/OLqCMX
6ykMNeTR+kHUZe/KohjaW3D7R7+E9BuyEBJYVF3XVIK+DBeRQy0LBizHv4BMO6BR
Sg0xiIM2Ms8adV7ZPEqPZqNa7tES/0V0EzWcu3vzn7AiRLH4NS7Ny6R3YzxfDSOn
luW6XAvuoEA4AZhaztq4GB2z6rDRiXFj1eTjQ0E80ylghuLlG0hY1YBhnY+08YYU
9f8xW7vpbuylY1SBqPksUJfsNTKTP66weFOhjTEX7MaP+9dShb1Br9rRm+Gw/9cD
/ExzQILQ1JQPpc8wPOu21JOEjIa9G5VjYXEvvcttxaxvr8nEbhWke8+wu3dIImcJ
XCORSgkcSXDzJy8wCSDwiZ87XY8uYJm1Sn/249gms8eMXt1TnRfbhxTl/3iOIE57
7vdhDzYObSAjK5aYtYBuj6l1ntY5jI7j9yIlEEyX96Vme43fgLHtDs9/8Fo7rrv2
3K9EmVwpQVthaSB1Ls7mxnUTtB0SX0wPbBNAFDlAX9Fs2oP3KLOnF6A7HN0xqi+O
lxMhkr96tTWrdKu8JnzxOLquf8cyFIGrnuQDDYfB+a3EDkEKIRRNAlHtcxNgt7bg
pUPGxH2oox0Ki/vWYkjZUKx4TtxCN6ZQQqKBrN4eP4ybvIne8SCU89r17ColJ8MX
TAzg0fgjDn4O3KH+e9WxdQO08BQWkzl6ViILunzrxlkZu+w/7tvDQGEOu00OuyHm
zDgo5P6xs8zOo91uk9ErY2N2Sly6aKjmLvoUfoQoeYkmekR1h2K/9ezHW+8E30NO
W87EQfVLw2LtIzr8iVA2OpSEquqhIbADN0mbwMf90wVOUSuXRRUqaiPSlWUGprvs
JYOfDGDZBOXiGUIzxXZo7EnK+DzmsZNR1sASSwFSG3FCmIDf4uK54n1qI2OusTYD
DQRRgzMTSVtqV3XN9ZWSQoR/I1WuVE62J1uVk+FujL3IHb1WFFmzmE0osuHkE1Bf
0q84zsGeDrwO2iVlEu9uVfezKC7PW7JQgERv6IvjoAGNIBdEgCkWHE1xGfvZH/Em
HEaKBd7+MP+ifxiNCmCv8LNJ/6N52qLlhc8XcP1ROGZ1oXufk8e31Cygwx8+gsXW
9vlAqZYRgFTUF0AAXSJyOCOhrZnBB/gSUxoEj39qLuuGroiQ78GLRow8XB13TTgb
D6g6ydO694H7zVmpey/ZezIfjW/rcFuaui6wnHYvVuYrWs6XV4w31x5qENTdk21S
YGYME7cWT+M5Pu9ral0W36pyXrECvkUEoGHacFMk8DUpzHGtbwETpwKTUDzx+aXR
rrf8SxygjNYLWtj4BM5z2p+cfgsqThelinzLnSJ1YSUVzxWDI9t1sJmGIa1ppwIM
MRd+G0cz9YrhGU9JZD1G6TR3NCJXc0mWMp9gnLi02KiU8sBv1mBpYqTr5bcIKZCW
0+vGA5Q0JlghVpppEVTpt2CEVD7yEUBUDBGBghGgE0HKEvLyL5aJPPoEGhaZ+zCp
XK+OgPqlmODtwKNp07FCn8yqDcUr1+26E4MtXF4TU2397DDCVyiykslJXwnjOwF2
7M3yeRyLlcRzDUG2Rje9Dz5WjBDLQ94YkwmQosTVMs1q1duPV1XSw8L7HVuzSemo
IW4mh8Y84UrR/Cpcz4GbShfez97qx66/qW3SeoNQvRMh3F9RLLOd3ec+XO3qovTo
EaoNB0NO9G5XS04HfdZT4+girIdlWHisScFIN7VlDDjk/0gljyaSgvNi59OA/EJx
EUIGF4XdJRRTzejq5EBfbH4dorogotE2WLyPJbHDZGW+r6OCdsKj/e+BPR6OO5GE
g7B2K78xWSVlz/IP8hqbeLqaVRl1LtKD7cAKP2PIbFg7S/UbNNNWtkR9vEtm0q8A
VtYGZqAueuwSXlfU5PKhFPdNiMeciqKpuznE0vyqxhNVKr7jJO7fP2IAr52YU7Eg
GdtvkC+464Lgti40B4InX/PFjPf1skQfE0Kfu8grQCw/4R8yfuu3Lr378usP8GRZ
iYGv/kqVUMJH/WHaKePStSWJIF2P64PKgudi30CBlwtBRz0K2aCZGKj+8w2t3kOy
lpRdSqki/vzZ/Edy3Y/JOs2yabw62sURE4b0y/1sIau+ho7ONzktvvZHDc8teosX
roIAo+zGldJFQ/ZOvJjBdl/x25+50T7wkTGYOwohFJ2RFDo23BKAhFmDugrM+5Wf
NPa91RDmF49g7GfVe70N1qbbis7IxKZEgwAd6vXKBjABQSCzV4I8wwrMQz2KPypk
offFERQqQCYvHzAMzTTuroiknYJMpyhccib/sye1LjOfE9hrOQ4WEEkRd9FdMsDK
c3EL6PUCHNe5PBlEFxGWLSfLKnmvCGAufk1vkfXLKv/nd35KsRZ644iNZZ0/xPS1
H9weGSu9g/oGRjXconEZoO6Ax3+meDVS46pUU/ZSACHsPkQjMRR9wQ/YUolirn2Z
qmUwLW4GHCXycUQEBSufX43THCATIlb0coyL7kzzdHtTkGSQLWzFaPfGoOlOK+bR
+izYbne/0BdfO9oB+eXArB3xANfZdD4KYrwuJNyeFU0DjhjEU9nzPRLrMCrq0YNk
3mC6UHgzhQCSkjIO87YBDNCc0LMDOyxroKyxKaXhrd5guayOSPAZn4wVTJtaYYPE
2EQDCkz76iD/vUpI39vjdMrzFeJdDn31maw/IKPTayKmHBM7vjO7zetyHdGzed4V
Q6cjAskeJoF+ohppnc8GJs8rvvhYKnMkxmOnM9YbsBA+xnsop4Smvzm2l2YAE07k
vrf7rDzRfYIjD/mECV++MEri/snBSCsLUBLPbNPEAlD6Lbfs9VqxWQ238X56YBxe
J1T970/pOl5wGESUssahJie9oUpWEeRYSwNGpCZ3CSo+6ueyBmEQOVw6hmjFWBQD
jlACcOhdUc5Jn6qd9k5YnRKMUdAoU4E/1U694QRBh/yQgAmaAD6BWyBYKh9Mz5G8
OdK6mu4Ctzlnq57DgiheuaMtlMTg8Ri129zYR1kAE8cvA0wYWy+KVqcrB5uY5cmi
oy4j+lgxgND3W1EKeV01Xx/2kRmlFR5HUd/44dXFLcdpIZmqTEAhKnmv/kJvP2Pr
SoKDbazhbIYySFesuXK9VP4VFNQBsu4e53FgrfDvSwQBsDHzJOQhs4N5LRPniJT1
tndfOFJvuyhadS4DL3HG2rYOlxCA1jAFMESK6Gr+47pqw/f33BYDg9ZG2nanjSU+
9Q2hwejeFQqMoENGFICywOTaEsrIyVDFh5OCdfxXCCKaQ+iEs5v41v8+qBT43n5R
W6nHj9X9+pERDkppfUfbpvD/E+++9ZKbxpHEferzbLZrDryEjezc651DYrkA1KBi
8NO/mynu5uZXfEdEkAM4xyAiIs98cI21ImXbZOe2+wzTZ++eWLiS1PGRG8CqtZv+
8S13jRk4oXp3SSe96Z7NcMtxO3NI3a2WoNo+4zkAA+bgIfKKKRgLtPDe4l+MD6hg
T2o7nC1SStVKOlwD9Ko6QhAMiE3Wz57OC/dUI5eR1s/N8KxweSJkv91t//4ShDOy
Sm8WVvDuPaSmNQdxFaML9u1vS8pz2JDqqGb71oOZGrgBCDwWItlXZmTbS8YFWTCU
0DuLdRiTQwppXyn4TYRrEcTXs/BhMbWg/BAxzLThe1/0BxFHoTbjGX4jb4CouLFv
WxnLcjoT/d0tFi/6LKlZdAw9soFU/ucBzEsSMCRpt2Mikpe5PvP2Yrah0KDQaWGe
9ea1AFr6lgnYYxJdX6CIgB0ddw1DS26e3RSBjF8XcaJyZnPm0aNrMtzCbLuqKA19
XBaJABX8tRzyQjcxI3PIUgP6lc1I91fsESH+ZNj2LUV18biXaUcNM/Fh8LDzznB/
VM4rJx3ZxBFOw3zxaFZLrNe3Q0ziEIk0kqmgEy2h37QSkyCjj9O7jiZYzXRXmO82
HA/AYWaKCl8wGsT3AuYwkK+okusqSsztmXINPKU+u74xR1FCYYKfvF6And7d6dCE
WJK4qkS+H68bWfTUna/8tSYn6QXuSrfwZdROjs1zhsd/rPfYIFEiiiad/LVP8IIq
ueGBj2eyliG1DeCX/Qek8CBQyZOLqhyPSTpLxTKvJvyCa5hoV0Q8UcwSY205MKNc
jlxVupKZ3LlXplbmPWtLiUI9SD4QKa+1NGcU8WOCsGkGSgHbFYL+QvgT5oouM9Wv
8IftOPztngrc4jQPbuezE8TlXbmfbQRXKPtHCIC1tqdQJW4GnyoeA8QoHujBMPlk
ca2u7Gsv+0cUkufcpXqfNROZXpm9eWz+H7fRK6cPOe+bEBKqzCVbVRshI4zuDLg+
ED519AiWt6/yMpQJe9eshk8HetQKnd9SvTRN/V7p0+ysUh0zkXT9LBTqUafLzstm
LA5K5wCkWcC/ROmMNACAxDKEvrdufnwH6kZ5b+yoltz/C888w/I1rx4eycfaLVFw
zWPVhccwPcDMLOQW59aL39R4N0882y+qsqsvbgmKx3Vz13fDOD9hRneX2BHjOcS0
ycV+fD0w8uUVNjzb4gU0tTzAH2AfuB9l7FD8lVoCoYjKXXE1oQV/wIF9z/RXjye8
F2D2O7Ijc0CWhNryOKJJ+U4D2oQN9ZpFVQSXvltN02byotyzP2QdbJ61SDhuGpJ6
NbVA8Jh4l5sZQpYNI4zN2UBpUxOKa2W8/j6LjqyWsP1WyjsHLG4T54to29Trv6KU
gsNYUX9TEDVSY/k+Jc6QgHUu3neY2GRPAZOA0kI1oGyO/TGElgJAm/grEoFDnRSI
lI1QpEA7ASjKwtfECZiP9kp4izukeqKFt/Bg19MA3C50vWQKsPUvrH5qdj/o3dQI
hqibxhxs8mIgNGr8E6SgrL2ylx/4ktnwnfq3vPDQbbgJosahK6yaAzINv+suISjc
+c8qTuthxFOjFRI7R5Y+Afy8TWed1tPKz3+79sD76+53Vs3jH/FY1Bqm5tJPbU77
+Ul5x8cm/BTL0J2Bh86ToDAFB5n2stD10PKYvX763U9o84zFTCZINF89uNBDwAo1
Eh1twoQRiuEthjWibaK0biIBjYwaA5unuVYc+l7Po0jXFCZ3C0s/K3R65JNmeqmM
znTs5MMdWUG7gBG+OCyb1bXZg8z26mqdabM6hdaDWbYn+6zFeDJponkxSygT7E+B
2vC1nRhbN1BkDVhPRKMUxvSrRROX5JPDM6cMAzRHNfXQRU63nd6eFKvTZ4O3WJpu
sEyLDwKlmf4zFJJootGQPZN+cOCZu0faoRrp4d8WiLvW66f1lfihOL2hmoZ280M3
nA9Fp8QewA6GDZdo0GJKoAWxn9vyEt+lw4f61FfXTjrcL56hbnaOk528JlvmX9A5
XhpmQFffUp+IJUP1K81gSHq5B81SzanqSxyDoCMfQZdtnBYsj+5A6gXpG/1BeSB+
NV2z7GIzYLo2SrZdnztHOHjfvJPAi8VrR2XtLV8axmaKXArt89IqGAuqd4JYl1BW
2FJZaYAZGdhNjbQwfCh7Jq4mKVjJ92gcyIyXh/OyTP7UnTNQAU2SJQz7vGYa9uFP
ZtDUIbmLigCSxOBfDDtOZ1UTaxOzFa5DxRu8vV3gQCKjVC0AlQfEmzPwt5hQeek5
VFUGv3xpzxwbCe6N0DNB8cYWfJdpE7Dfu11wOqZIP8M5hKEmH8LF5pg5PtqTJ+3Z
KwSlF0U7jP2Sx6Obj7zn3V83P0KN5LhYcE2RlnTbJ8kUDEQsoi47HUmUdP40LNE9
t1SC61iC2KIZBppZO8xqol95yZiV8QHv4yaIcrwKgaRHHLLlcbg2Fcgpd/KUeU+d
zCGpRUCtud+lwDg2gnFQMjPX2UfoUkgGRqESbygrhUVCRx6BUMhoT6GczIag/GtG
XnAmJNJEnpj6tfzt+hN+a6aKFNrOenxMN324O0zgztJQoNClM/hUY65TkGMoDCkN
ieZNenReeRXm74qn3xai0jaZSx17HQ1n40UHW/dD32iL9lqYXu3stU8usdt7/JZ4
ollTodam402or17XXvZWPf3aKruIFkNLl9VBREvriB+jRyvRfJr2jUDNit/dHGvp
wucETRM4oW5EJfjQ1ltNZBLM/TiML4OE+pZ2QYk0pskB2FY38jbKLgbPHZi23Pzt
QK4/lXkWuJOxenPR3nHkn0Ea5Qx/PGjQ7C2YjiibQAO1oni9FV02mkxQg2TPAttq
Cm67Fct/mOVjJgLU95lwmTKsDOU2AiX3pWj+SiaKqFp5I4b2eQPnlb4FytNXyJGB
x8VHlw2O2pgjYs+wXKc2LLtWhvUP6I0/s0wQmNbvMErfKMDSZXrGF48dV/cd7nB0
y4wZG3tDiEXfJqWOCD2D+AJObKgc+Tm4k12uMia/nr0D2dWk22qSnw0MB3YRmkKH
EDude1Bo4uETi9jdOPcLOTSEpUxtucWGVrPZo1+hYmjBeQQurubpktTthtVDyUGq
fSgPCLzfUpSPcyRhSzbuzh/Y+RsFV1DYdZuP+9sfO6MCorm0gmeFrW4QOGX2suD6
ozUBGIb2gXC6jLdv1JJ/qg41bGrlT8ENZbgqPWPirdB421M6qFlNO6/vlDvoZ5fY
P+3Ena02gmK2brJVenaSJgsDKzB5R8wzvp3jh0ENPujlmQ6FmwqB47rCC3FUlrKC
5aV5n1fojoLs9Cg9jhZVonD+yFTdz+QJEDb5bJ71hyIJ6T8oZp51Rz9n+DvSb0t7
zY/hxrcB+mmOdJfGXeXCgRqUHe7BtMQ5scX+8+6+gZQUE52ydG6uITWMJ5vp/xyp
LYyWb1l0DxcSidiorSNkw/JOIv7x+6mtWrzu1tioOc5NRnhgWnSZZCFopP/hJpAI
gOL+vw2rMMdcmyo0h976eZ0/Bf8135VxNLOn/DEPmRWUnvY8YEBoxyj4hwJJZ/xL
0PP9tJoiCVFg15evwKtpaKSYGqpkd2ARILUPrzuamesl+zGA+ndrdKMczZMm+TiU
s8lQGsrmRfM+m0aaADmEInlvWgfdYI4lVYmw1A33QCpHmyFW5X5Kzqcx10ZzxrZ0
FV7CmNkd+e2mmTF2lAN9EKpdo1e+IATamPqWMKrZiJVKMZj6LRGLsIvdfoMARIgI
39EW8ND9+MevaQgJWYZnXIZaSKkMntDyXD99B1FZg+I6DJqmhsIMBLIopdOu2/B9
Sqc5PDzW6SHd/Vw/nKecuhQk8Ys08Zt5/g4kaXJTsEgDX3i2aDWs7Iax7bOasLG/
ycI+bV+0j8HiJvURqbWSi8YoIoNturnJQIzZbhDrOoTsDxVfdGDUhvPOJ68Ph9Zp
hDS5hpupO6PISY/O+aHVmbVotg7EScM7fKv0St0uFy5BDKxRd7VNBzxtyEauXscW
DgsNC5SXcbO9Wo5QxW0bySq8RRpw1bRPrOTpxYA1vxM2pzorM/6BKYw/SObaj1dI
ODY6Xjhp8iqb7i4xHteiTEQHqf+8v8DX3wEML0roPlXzG4fc8x59tCXmhzxvTHCU
DzuQoAELpkDlAkQ5L//KYvpozYeElCmXr3vmehBIiVkT7RbKPd2Ij5Cc5Q1vnYE+
SMM3KO3HvuTDpohlkdZEAmDmJ6guelhXUjmiNsQxO+ZE50sXV3vE0ytB4yEOWjVj
Ha96cCofkvKrUCvOEZPutn+Pwb+e52UJc6pXWCAaS93Gri5lceIUDGg1kW5fyGxR
G+mMpcSJ1Pid/EMP6NlDf4fkzhSZWF8vqPOJ7/50N3uxRxW5tXv0FQ6201Dk2rh4
oqV79ba8vkRBmMf5Txh+r2txoZxNb07c9qAUmkTHMWU5n/uupPtwNr+Ujl6gIqnG
/iT3KzTt/9/jp7oz/iiDG6xG8Msu5isvdwWXko1yyaQrNG/tEoqqZNAMDA9foLeI
EA6byEUyY9SQN/2Uaxp7CFaW1kwqzrhC5+91pbl4FLbpJPuoUZd+CDvnEk2QrNUF
67I8woL4b0CzkktN6n7wzzCLIfRi9Daup52dIEOeJ3iO+cw3bAtU/Skvz7GiHK0V
Y61XvS4ZF0xtd2MYHi0yV2mj560ATFo4ncUgS8ilVFD4QFDv42v4lpGRGMCEV8lN
nmbnLZAYMuBKWYVfpvsfFPIQKYkfgyU+89ZOqtJefpXk6x4LiWXMaZhOvFx6Au1s
99eyP+zO3xiSgN5gN6kCL5SG89/EL3eLXVG5GfUBCU02VcMOu9FmwsiTqyk/jqSk
bLZkRR+OMnreq7Nz73q6OTnZbapd6FdHQNeyggXx1qws/bzZ+EH75I9fEvBtp2XR
X+Dez9Q2iY02HHR4PMw1OJfq5k1ZyOZKf/MQmouO2g0jW9qH5pY7Z9UepHrBULv6
Pf3hXMvnaZ67Jy266MP4aeIghO5p8Jjvd2FCKx9GwiKhZX19G9HjSZFzlqqtP1dn
GJu+DskC1PI3ACeYksr1hZKN+2CIEZVV34yPOHp8LCSBPDgZGJ4qh/S+lSeuYAJN
/4PTw4sjRTt69plMaBuKuDhdXsu1tcEjIxxzJFFQSX0tvEXLFeKhwlaRuGrpG2bJ
5zlnVCbSWFHoHO4IaJITVEvyrc1DOSVOP43c7psufXx9Cj49p8RtZjjEXxYVNpjv
7RbjO6qm0KnAwFKvvAH9pUF6sGIeSRU/sb1rgrNPGR+js9rnZQ4+cwVmieEscc8Q
Zc0PPOSYclyxYPZkyEnV2bqIOdImI/EnNZBCzC+54uvPKZsfE8rRk1Toj4jBFw+i
Vuv9b5V59V+SDIp5PYEV4SFvRn3kPWglDKPTHFCito/ObZGfacMC9uNpdzid5cmj
tm6SYfNGddMtw9dUI68OHk2EgBooDC1bTm+9EGD4h08oc2r46uVy8HwLgtsKT09j
GkpeSr1X4lz0V+CVlzjjHvSihliajPiP8Bb/oaMLoa/E3TGvzkSGN1IuRyROe1l9
uug2sgG7RcD/wnBX9WpKXNNJcxDtP7VwJ+NDOwX1SYr1asUW68Jk2aV9DQz0Izk9
MXN3Jo6xYVA2gIgY70zBrwP7dWszhing9QjqED5AW8Gqd7q0aB2/ugN91HQvKVIx
Yszq73Iy00RTIei/Uq/IegKryx7AxCJ5eyVzOJVPauNE8IeH5u4/lEyxfL7+sQER
Ntel0cN+Lkl1vmu3yAqeaKatSG6vMtyQ5ByXaFDfPFLDC/A4bUVYp2Pr75GQ/QBG
OT4BOO69qIl6s9VP7K88DxX25mRJKxSx+qLO94yZHuewRZhkb6OpxFMO/GW2v/pa
gkZPjM43vrDyckfq1UZnD36rMx3txcDi128IfOSqhkG+fgs5bFP2IceXkuU6mRB3
VwuCDLmRd6GjFbKHa7Cl/CiHjIrI5xC6hO1xjmif1dqo8XhPBEEWJ7CuqlP0LexK
PmVwWFsYElji6utuiZEh1gtnpQC7CRgc0wS5c0dJTfDq2l4FUxnNGS0oUA4yom+l
5POkgDIGc3yUuOoZh6Ku2TiqAcZjZTkXtwqv2CiqZ4L6dMUWwqMWMvBthSHic+mn
xT0Ew/vc+DUvZI1CB/en8l6XDSaYSc/m4IAfbKLOO8XII8cdaLFkXdQCW3u2cy2w
JoLvruc6LbhN8euHtWUFgy+hI7uqpPqbAt8/FYMJAVIrO2/qvY+xZQ9M0P+olxoM
0g1bqn2aDFlC/XrsBDbL2IcsyOUO2bLxRUK7qkEQK+T0DE1RgfXy1LOVc1wPxes3
z67wikoa8Z5eaWl0smAbmOzIseLaZuZSphtQtqQXsxMJcskHLyne2EzBJ6LWcYrn
oFJFqhqkGHRz/0cRt/EiMbKd2iPYh4Y7A2ShHEDyCE1ROr8MSWeqrsIuNxisZV9c
6oibC271WNX2pbUsjVQfI1LMNCtNvADSqQ6t4E81chgJZCj/07zY2xvekP8jEn1Y
s3BxswFYWiepUndsyPlqrxfZ8EOLz90rOPbCo7G4h5HmRFMEuXGG2ujvNxKZBFDp
nHWWhtzRWqFOLe9fNte3ZFevn7pWfU7r4TGioEHb6sHKeVnDfMeq8xh5BzZI1B8g
ABo5NxBF0QOqpCam4lQfdi2zd1rHR3uYRpeIqwiZzO1wKsW+CloWK+XeO/ImfNGO
MDIxOFA2lB5usSXkYwsFNTbVVh9YFXADjQ/Dbvgnjmo7qweQD1dC0Jf7M44p39R/
9aBGNlyvVTg8rw1V7REUaCKXYnfufAe5OpHYRf2S8mwNF23Ww3V36zcvh2lmZ+lB
ZCXvAGDlJBMMMkuZ2KLQ30EfpkJwvCC1FRfTnoYiwewuiL+cZKCOfY/80AsgNXkh
hVvwDuesoNI4ZQvkp5PyW49ttiqne4zgzc/Fqfks9kjRVXru6Dbhz1t1uJFTKcXy
NaSN/kjlJH7+CwaL9ca7tLFysg0YW0qCCWUhNcMWETfSwtCNumb8pOHtoUzQQLnP
6t4Pl1i8wDpM483+Tf0lUhOR33bmh2VWfGheKYy1jfA13WICNHAZNMuaHualjhoI
42XhrcqO1J6KKrFkp2rnqZ1mMqOmeJsCUP9viiVpqJ2ZuaxOGvicenVEMvJdi2hD
PuAsJddioNqKNAQQWhu+teAkn3AOGUkp8lfD9qiSgYgTWNDGSKS0mfJCdPmCikhZ
5oBlW4EuOcMPS9i5jkW/NA8H62Zu2TUDSmAro6jqpnFfFlX1Uu8p1WQK0oqxdoth
sGnjU+1pqZuYoK3DRMDUcwVmlaBkTfo/pYDhPGl3mujC6OE7ekDJ7Z4rwmwrhL0n
vdk16hAJSR8DllVIK2zRlirOPSp9lywtrpxQ3GdAqdoHtMSDYcDMGHxYpwo9PAgE
nnNyA0DB2+Bb7pl5jt3TSMPwupQgiUcKC5oktr5e6EYgjJ3cqL+peyw8NrcyvvfA
hkNU+RBrpNwFp39TJ8xbzdlmya4DKBq785EE30S6hiO8je6YfQTyiHXgCWrUUT1z
eiWyI0eEnFLHPuSTQjhqSF6AoihMmyxkx1LkmiLAksQpuSz/KyNv0mqurAMDG7cn
heepEEFeLS8C8UC0f9zap/cXlWlCdEkf1YtOHkmIU99NZSx7t/kGb/eUB0da9ngW
7aULye4E9cPDLYySQXGuP6WOejL7g8Ndv7NEgnQBwV/akAFK+lYbjGwIheZ5BYs3
mZHnrntkhUq0FmnBrqJ2ThhZIFAJb+kGsPugY4Kr/e+GSrLxQxQwXOKuzZQ/aRZi
+BimyJK+iYEPZW651onQZzENiMVf7/F6TSVKuNjeGU/NIAmjz6exsUoDGlcOzLGS
d/GqWq1delk9alN5zp/1rcu6IAIuHJ+XVNtQpHbxQ7r8pSoNPNqdAEpgIoVJkhrW
IahfdcGWb5UAX900yZ/bQaS9FcOP/Okxp51XgTwiRYYjvBnHXBcWxft5SjUPlvvH
SubAtfI/lBaWxWmrv0u1rUlV2/ng/5xMRD1a25hn46Iz0g0OlW3beuJq0NEXbGKH
uFMjrWn2CRKYLmSvtTwIgXObocAp+g4xKQt4nHdoHh/dhgubMyCUqMA3fqB7O2Xh
y5NfidxymouVgQ9dhfTNj4im8kyMRuy81FAJUKMpiU4s0qMLNKVbGWWQLDFegnhh
fnGt1qnaNdIvVZ7Re8p5ZRNYNpzYVmvkt1BYWHZwLjGFI3V6vGHFNa8sgrpq2y2f
L+MwfLoern0GhfszXsvPwEBTu9zdukKzxc6bjll4feosfBTmu0RDYuAYAMTpLNYV
5/KIF3+9G2A1gHYYsTFBOeFCiZp1JYx+e6UdWqONzkv0c0jRGb1zJNwBgr3Erev4
Bxi8gK5uN2RHHXtsQ9THaFR5DOoTGYNgLARfuWp4WCkznNZauwPnP1c2qacYQ/zb
yFVWnTi27m419ykA7l8zfiDhKlyS/6ymWig4j6SwK4NtLpts57uSoUEo1u2GbaJy
5/RmS3R1ZlofU9oBWqYd3+p2FRplhyD1Xg1HdFQRuiDr2o2ysbUcgpiYJRo/olMV
Nt3uc/mnid5fYfgvq2o7tI152rAl/Z94hoMNzP81t/Bpk+CTq3i2hLbjOETfKsq7
zUjZrpWkLpjB7mmLmLHxY86tNqJrO2jzmuklA1kE/isCn9ZGxySozpnHwAajrvqi
TuOzy0nNbXqadzSBJp6rJCObZndzbWgvZj59SDq20u2org8t9F5RIwSCO7sVslbD
wm4mUWiOIgqkrkoCT+kPoil9TxrcAPRW7kP1GHg0Z7+3zyznbB4F6bpvuyXRgX0k
63CGGpOi283yXKDiCkIbg9k9rvENUgQTw21T2nVi9c4iK15dwlJnpJ4io6hSEpPh
f9PIvpxlXyfHLI+YxHmnAYymfa+Xps/oqjvRwvaVbH91A9z7g3WeTfvfo3AyzBjA
oOtrJz1s1m+RL9c8M3f11xOpe+qo5DqaMvSigCxLfRVp9V9PP4qryn0Y7fC3iYTd
pUTqHeJkbdJ5a+5RuvQGSFFRgN6p7UhCtKTRlCONT0ijA6IS6cQH8u1FHmbVrTcF
vLb7nVhfy300nXdWbA4KVq32ncKe0XmLV7HZeC112OBnAFLKE6GYuZpe7azRbwBW
0IqC3Vjn5Q8GpPp10O+qcGgfAbX840j+pr4amNrEBdozBIeGwFTh0jamB4JnPl3X
vO5UNF14yjV5f1GNEfZKBdl08v4L3UOGHudqIXT4N7opRyJoKggn8R7/SW5GrIPn
IQMjjcHx3+QyXtVI7FpBRohbwJgN7VO/h54/xPND5edba7budilSPLkUkTl5IlXa
ee7+I11fOLtQEMJptm8dX8e3vh08O4o/FqOBp8Qx/9eY8GuLdTDzvK3dD2XKbth/
atFnC/wGszQNeIL7Izw02duKguo2TeXARZV/sJYETwPGuXtc1QIRzXUm7wcpU9A6
j3+gd40HgGdPdUvKuUjs6Sq9pMwQAyjUc1NQOIGygTVMvGWkc2ZKd5JHfudBBE4U
ws+bdJ6LQ8dLoY9aWzzMjN6Mbk62G61IBqkggrBKs6XMpxPs2YsujbQQix3rpNXy
VKORXJlN6jFcGIvIyU7GhB69Kt+5VllSDzdMngAHvj4lC+Vo6oWMGIF++1SEkoTT
sEpNWwEnU84KLmKzSdh1LHGAh67iclQgqBq8zpE2selEX0XsjfBcBYoKuVotOpB7
wPWg7Bw0I9b8Iqto4HK9/jyeYdfULGfysanPObGd4bmfr51q19zyyWI5++cetMK4
1TTengyOwBVVCI4KD6uEAsrE/nSwrzvgeLNHWajXkgY1vNJfVJi6rdL/ZX5PKaxj
PSoP4JE+cNtGkSi2ZD0nec8vvKRDPAxaWXBL6QVfIjO9owLihPKXg7GAPxPYhZEH
7qAD1TfCJUfB833qCcjQAkcos4iSl9kzO0ivoN9iFaZ2QcKsGlQlpX2128L5q9h/
Nx0uB9kIw2ScEcgTJXgro7KHo7i7qp6JSLAPlKud/ruccCjLDjGbQr7woIdfGq9n
SfFr0tix0I2ephOTwZZfNiQ7fXy9CvM6C0IQwnltG8YG7TYJol2ZnaF5M9NXFlW5
0498fSyEAGipzVC03YkurZGHYE0rt3hOFIi+NffjHJ6h3Smj1mgD6D6y6pSXS4PB
K1Wd9KCvNH5D0YTeYNNV5rz6iT54OG7eanXAfryBPDJCIZZOjoixmaEoRl5Nu2fL
lgm+uFOEbcl3y281S5vY1TmmsYc47Jb9FtJeXO0dEFZ+uvTS03EKkClRNJLk5Hbz
6NnIdR3gmnXLQrQX3xYurF0QfkZd+jdfadZ+heqf5+sSyJaSdc86DhZMNOrpG4Ke
+yH/d7r/lkWo03aMWAqcKT92B7svvz0vtVq/O4QbgrmxWErwDWIBwS2dMmXGNCRG
hQN3FhLbMSc5MR2op20rpdm+wkSMa6Ules/vu9E9GMYuN1ZeVKIK5Lo6pwviu6tm
QWoxkFCSU5LSyTbpNLRomcLIQTbNtnedIFG0d/VcC64J1Xa++EMPD/eKzLznGqNZ
/ZYfVH+in4SixhpqseZCKnDfB8CEcrWVsiOjjBUn52N0Efrda4zMDTFDut/8l/Wg
Ad08UGfcxhjoPwQ2Jnz7bfFZCMZ73ejAWh2b40sc18VTs5VI4kX7qiNFTgUS9L5B
pmTYBtG8kGS0hK3UHEgpUgYNm14l5kzyl9W2xEMfxiBSC6rMG0KahZ4DGbfDdVEH
W5So1tKsbkME0aX6e9lRkgownIXOG/B2nmRJV71KEneJjZ7EQrAaiuSJHqLiZEuy
unKqr3NDFQLIVEsNt+tFGZ773MIliWCIwV75tFBNLkTSg6rxoW7nPzar9yL198WS
QolEf2Lp+JorpQaMTf0DuLsZBees/t+LRvBd860i6MDKGtWfnxqFhZi8JN2J2iEH
fW5/To3f66ZkdZuljywQtf81+FpgEidiJS+Iv6kPWV+uyXWovuo0nZjUt0ON1ne9
zik9eHe2tlRu71qZWoPcwAehtNo//Prk7VVIPR0fPU3uhkBZaRuGFu9ZjzOlgbNv
RnrBxSlwyuQCWYVfnRsWdi/Ex10r+qBgm1/s82uJOaGSzQBolJRVvkUlbraF5yHB
5TV96yvdgK+WcvICdu4+p/XYrlWK55EEJf8WxXnqn21YwmYB86vIR8IcbrySjcgI
bXxSovAjif4uFdXsN5O5UsVz70hDQXZEeNxolKm2Kv45ZdV0KWWCdWX1D6NuDyGk
yD3JD0mFTgfOPnz+DE42CD8pyUaAiCZ1NkmUA7DGW5xmQYsWoLwc5qaJyUHORkSW
Gtx8gHCkRN9iVar0ed4A6XFDBrMMFi7wyx7Mf8gkmmLRpdBSUgerKaxKsRGnjEIi
IBv4vYawM9nStcze9kaw3Adhmk358JjvhfTBOz4lufeTpbedkL+xuW4L4ZRuJU+e
VcSKgyRtYNycpNLt4LiW5ZxwY5DKNVOqPDO1RCBqGNBt2cSpJiEM3WcVrsrHjf8k
iFFbxjgkP6BAH34ryb055fOBYlQ0Jz6ETWtd7yAoAEYEQm75BjSYz0QWwK0tGOs3
xDIT/udD27IXVmUZguWpEWaSOhNXv1SjlhtWDxteGG16l5BXfG7qE3iKHxifhd3g
pX1lwY/KBnxAQ1GVXEebNJzeTfJPlDqm7X+ZrkE1AqccwLYrcrrM3RymQSPQuQLZ
ddMCwSR8yC0d8xwaMumPDOPi/SROKuNMnftOWpYckDxAnLQTgXHK2C03MV/Utb4n
gfS5TxeEqAakIsj0YCEwb8Fd5Eef3X7I0FiWCC6bZx8D4uBVbgAY3bsxmGtVvoz5
dzligFJxzZvMqbTKVV3xSHQqCalTQEl4EAFmU3CPnGMUjh0n07P3m98oRFpKiesM
gU3IO+rp27+1zya7nT9/PPgazT7Glq0FPirTb/Q3TVUmL26I2SIwzUTPoCtEuu0Y
q+C9rDbdxaM9KagjynFBtxVUSp6QKSjl4TTL928eFwkZ5G146r2dU6qB1ru4e4SN
5ZHziR4hIar1BtObxbqV/OGzQDG/MKXL4VEj7sAzKKA8kBAJyUnX3PtgiLzk1nOH
4H86U5I3nGr9ulcfpR9cBujFwHlwUS85l5vIAujzw62KYpxbUSUfyBy79ei5OkS2
tAsWCW5YvXYUVXa1UImskYj4mcjAGQoLVI0EcYVm75BFCPB2VaqPrr9KzUDADPtT
IMWiu7rSNDwTXqRwNyzkxAh8pXWXuo84hpn4I+4Y4z9PG89U02hHHDHC9Q0i51KP
8aicgxif66DNVSZ/BYP0XGURhLpKEjXN5T375b803G+iYR78zp10v3zRWEL4RvaH
6HybPEUttnZTfQ+LPSl+cTomljP8A6gcz25LkazSeFq8dX1+1a1t0UcAoxNvM6YE
aekQyy4KDn9Dm3rFQgCaiSZfQlfifRGeQrKli4zqwfz43Urh2LHEfPL2sgdE2baT
snlyS2nA1oFF3TbcP/MGjDSVfZK1XxO0xLWffT9RUSfpp+q6vJ33/Ojh7i0mux+h
IWrIYIpcTg8y3UX2vci8IdZzCp2USl92i0pKGCrKtFxkzFO8WLpImUeV5RsiTtnA
PzZ0JdcQqBoDOyW2Czc75914pc2oqm5TBOExd+h4NgSLY+azKhxXL9237DFci3b2
NTC/D4qFZ+e4je85GXTHzDCRnwL6N3XCFXT3jGXeWo11Nhlun08kSBi4jOpX7ZCW
gUaV/KevBwSyTzEGzjrgSzvJT1QNKl6C6CQuP+YBahnkIz3vfTOygZQdbDGANVN/
bqb3T02pDfM0efNlyDE8jkiwfF7IlKt8gzzVlu84fsgxIsYTPGxuogTL6H9rAGEK
mfz4d2SbXRCYq8LT2LL3/VoJ7bedQCHlf+QWDPGJtlEWgkYsWy+mEBtbT3d0vDc2
fBsyvvzgXi+GvshwLC4L16LU27O6TJtXuxFpD1CpJLpC6IweSgx90t1D0oB/27oK
dlch+4RJc08v5mzs3ZBFIPzLmzElTdPj2+KYpUKWra1DS/lgF7dTuOkti5wTcxJm
KPhEqe+rS57EO6POLlQMrVldFSI0b98arRyWxNIIhsRLk8qZcwFwmViGkWkRUrY7
lHuiaMLrvmiDjp7Wk4cla5UCm9Em5hDJ3euD0V9pvGDnksTEEVtAh7c5cOR0iYqk
eSwkys5Cq8N3yEeQx6v2Ah4cEwoeeok5O+adut2mCOrhHPswEGtqC75Ff5wK20Az
FEEmziUmZKlVj7DK2YRgqsfrr2aTFar22/Y0tMcmOvtWdZpjXLUbNCeoTcwC2wRU
VIDEmn8714zS1uaR5XgrCqqBwNGFV3aRgVeBY3ElWveB7sh8prhGdMzOm1klxnrz
Nj2B0LEDHwU3CUMXqsUO8jdufeL60KBhLsSnE84tpKZk8/jqOzNBaziF82r/kHhV
z8s7fgjXrKzbf8MwcCArdlwgXexuM7R2yDhmKDQfphZcoYifwqL3e0hn/uJXlXNF
HU7xLcS2KILUhUk01KKb+YgI7Pmo6ZrFp+6O0PBc00XoTy9wogEElkVprCIL3oUV
ob+AK5E6qHMIfY4D2aGgTUaeUQM4z1VeMIof3v9iRUvSw7jNLte2yL4gZ+j2yNj4
THpu6s4rdQ2+Dk0CJwMGwwLIvGcKfxhzk48JYG36QfVT7rLLCgzJ9FMYQnIs8pB5
7JUUgeTLDHvWhA+TXxmR/7b7RWEHp8OEJxrc15UdEQrE97lwimxuLeNQYoiZIO71
PLLMdeZTo+7PQFyfJwAQnXsimqLwNasDSGHOkYZdIj+6mU6V7T4rgsEXLTJyNA2A
ZvWhTc4U2Lr7nLdByOEfMElc0BHscZMqIOjjVaKFu36yPFvjMjNpxQrgNlqp1DVD
tjd7b5TH5F1jY9zczUdSYoVrcoxeHoX7RmDtezAnOQtMZDIY7fMfsiCJVU+hmjB6
/k1J9O2eXNHjYE75MVGB5/qNawpExyJf79ZmZ4XPZLTU+SFqnJgenKGzLK9VECw6
UpEvUabmdQEYvFeAQDagFuyWr5urTRRBczj3qHlacCEPUaf6IejvmumhEbzOQES+
hb4+GFV/sVC/UWeqNTUilBgU4WCtqPl8qXOISeABVUgP2K8gHCCJwaaPDIOuR6O5
2sghyNIVURWJ6SQVxYU0bfWohtvYdWoyrDb9GVUjcsXbzcNuiM8HG3hRigPMznD/
FtdT785EgkPyrOVqKr32iqwrgCcO584QM4GDm0T2MNTEdeRNccCL6vna7iykYQy4
VjM9C572tdsGnQZTxuNv8UvNmc3ldkvYrs8Wr8ezShfB6c5vLsd/ngzHlK1froQ9
zmwys/cTiG/vg4JefUBInwG3CTlooi8b+vB1VfalYb3Xxrt8WLxrjDNgr9XzHhRq
aRzqbUc09ZfIQcnbDfhsOwQ2jxTgHfltUdKXaU4wSI8Aneohm69IA/iHU8MKG505
Jf20U848DccG9kRId48gD2CeauSGXTWTa2UKErHnVxCCjIHcL2xIk3C1cQm206iz
au7Rhx3hoGjFpgB9sIOeCdREK5A8MCSNVWhCA45QrV5p7iqx4CHAiy1KB1ZbuJQL
0Ak4bk+U3aerZOvENjNRR+WBY+U8k0O9Nji0kexHN4G1fFv3dAW1rL9ELcLWG5pn
zwmLu+3n5Bes0r/x+GF6UDvpZa9PZF+NyUMiQ3Wo2pGEI2P70ZAiaB16DJ7anEUx
eFG14nVoHavN5ginYteT7Oj6EvIIK6ClOgri30c/tZPChgzDDZ6ZGnAgc1+SpdOo
/kN95ffkyr8JhFmLPzfRI6krmKq33Y03B2nZ5E/0mk1/b4GLs99TWd1zh20XwUOK
fK6IAC2jsKf3ELirbi15ufzvWdLEZG1aokIHs00BDklxSWPwr1eI6ErKsVQRRDvO
JkXLN1xoWyqxVjW9UhLupruw/lBngB8PE9MoPYI94Uwgm319cvjClHcrA7UEUskE
dydtGNw6yQPxQ2kHFTyMk2rN2lGCEHvBj/3g47rzlNoeU/odISpxFs6tnH+vxJqo
JMZ8aCpTiA2ATzrO+/ak1Oj+gh54Bvvm2Ph1TnbXg0jEiOFdqkSyGuInVzpROV04
WFyRVeNejNo7C2Vv/xs4YI/I1dqY+NqLQAhH1Z9KPMKTFuB3ouxQcOF+YZVrW9km
gfcV/uyeSK8Qq76nIrWRQiK69yY8o//2msNoDifi7GK5IS2AgkHH026HOzUq8QIK
vLY/lAVuri/TnZwr1A2TRA43AoRP2wZiCYXwA2TSimxV9Po/TdSyD4muoPPxMs9M
zd0l2MHh66QpOi2DvS2dgU3aIL/WjLheKbUYYD+qCBl++F0SAsrvC05JIy3Tknu1
4l2Dj4kNPPjGWjRUUtIex2Qerh5bA0ocDITxTquow8T4d/WWJ6IhvEefgohvNxlQ
Ut5l27KKCZVlh5tdFVkZ+yFvCEzqKF19q4B4q9xQR494/DtXALxRqVXSvN3NMCXq
v9x8ZFeqKyEI9ObCW7y5H/zIclEqjpj1muIjiPWb3s1wXZbOfwI3t1BhHuYj+jEv
FJstgcZZS0uMil8Ghpc5M0qQMjelD0NNp86N+iyPiFGeQpKkCuTyVgkwT6dholti
H4R8TsApu1VQAwaxtH1fG4rUBJhDUhnx02y4UcJF48pNqwL+quHSwhVaCdjuon1r
Qcx+vl4EJFpMZPBa/5MTphFWFY1rcC6f2NnbgZRfuEFkbMkm1UU4L1E+W2+Dn1VQ
cjzeAA9yyxuwKzQZdNltBNyN9/kK5R9ye3Q2DQGaUHx4tqHN8FLCUzQWztHu8g7F
mG1yITIIN7huuJw+QIHQ4RvYV9Xcsyyke2D/YwZEffGowE8WWNdu/QA4eKUSSNYH
3RF6D4OLcblUxwOGdHF6cIS1BWnt5dHgCyG+Q9nzF8XWU72n5XOlOuYHRQ/K9Dj7
dcD0q0S3TKlOA1n1RXgbMlfGmFqw1uXL3bKHe5FsogqQ7A4gX9kaXF4yrrPLwV/t
PMMoS0+EvqVlT1xIELgcc542xnFISCz5yOy3dkNkDoQwwFNj5DwYy9UVaElNNbHl
VazcIoisgtYcnYR3bGjUyvyDAWb4rLkaXAANCWUwjvSjEBepeUaek5Lnt7CBEoU8
jCjmFeDSCsFKyybKQ6yB80D5Hd5ZyiCnRjLECjoCWDSis3q71Xf3TF71jcyJizkL
o1HQkKGfe+aGj9h+pHgXG1tTXED9g6L/KkBS03KPSeXELG2jAR8cT+jlNuc76rOM
C1Dp7t7MMdNCKqlNZvH6RYtVsVnnYZ3ODyAIyARxj97DV28ylw5lbQleOnIcPFSl
6Cux80qZXXyOyQmngzaLicbA/D+ReGhnc1ttLaaB2t4cI0P7N8LzhJXpj7Zj1BTz
6GBzwbE1BuSEgOcv5DU0ZooFa1YJ90XXe0xmrBN8dZRjXsHwguxWFp+45XtzsKlH
tikpFEeaZQ4PEA1rmCQUFu6MaYAZ3IOYlOjrRQGvaUrH4aUxKGsRtJ8EkzSEAdBx
uewnbKhceNO1a7V4XBDwEshenhCydC+y/ACbATU527HAChPy1dRdE/QnhoXk3g5b
6c7soJacLcxKNU3Eo6CCjpXOmYNMzYm7j0WCXnConpp2Btz7uBfRr7LlKoHpUZSb
xaJuvuIB0w42HonDOR0YJ/AJ8rr0efc8jtnoFooPSTX+Sh0yZVigIgKc0UwdXETP
L/ujkexx5FW81ClwCp2fMEw8lFquFDoHMkpmFLeXEtICl81HAAzpdjf4rKmfuSn7
51kQ1udZtSoHQ5Cby45zBArsTy18LKfrCJHp0xZB4JvEg+oMxqC7lyY4yfQmOjql
QBEPJzJdin1ummJ43W+g9YSAxgspj4I+aKBIdvsxhWWx6ezF59aW2WM7QO3tuwhc
Eo2HPrAo4N5YzMGhVpH6pLm+S+QXoI6+mDX8DZ7GXFwplO3kjZfRNkfKU6g/TL8i
lFlghoMS2SNpPj3BbcrHnxlRkCE5dwP5FY1Zi8SneNaJhP3qMPjZxMvQAxxw7epD
gLfBS1YISyMbh8mp1uQGIrQqI7EgLJkVlQnM65GI3qAz3bxa/VfY+3vimkssL8Z6
raoWIfsZ8JetA0JqkmNYsKHxMrGwA6ULjweuGZsdTDcVGVOoyIaM9l2YPrs7WlNW
4HwAfcrP3Sg5z9LipGkjqY9uSGC+cgtoU/vNaSVa4azLtAlZpKsqumOGHWyYO+Xi
bglrSPGhn3E3ZG/pkWme49UcnLJkZjYd3cpOBqz+6KxNKQ2tVAWgoD60cGamYPYC
72VOcj5ycT8jn4HXWTfZfWnj35GTnckOsgpupM/PObpuHU0Xcyos5Qc4rk/THw+O
XPHJGDIIs2MGEBooCpB0ZrcVDfIjStw/kiwusHazvAMV/Z4R7zrq/u/1Al8+8VBV
BdmiVZvdnad8rw7Hk8+KXN0hOjwoWw4nV1Y9tjsMLkF6gC4WvR2xGlwrCFdiYomc
Z7FtwXMQjyBLXqW/xXRXiRV2WNiS2dxRpa+4k0DesJr7C5G2pwpOhO/Uys1KSvzz
pIPD6tVzMt4JC7IaL2NTtA0s1Ua3UI+tTgRpE4Ezv7X2e5N9V9AJCqHoXbG9k7Up
O3ofz9Eox1C9nooyeLp3W/PI6aZUlElS7GsOdEJ4xTs3ppvHT9xlwPrFwu3EFWIH
ZbkB0HGq67iMVj79XJjUFJ3E69InU/JVMjJl/F7aWUw7OK8mMOV19Ae7LqUAz0E0
0V8nXd0o4M7B1d1H7wBJAuyBmFggJN6CgcsX2SdlENnj/T5X5PtLcswghGm4PX6f
He8RI1odyntjt4qGOigCRj1vNvVEocYOlK3W9loxzcXslZxQ40B/zmv4TU1QCS0j
aqbFhda15nyS5zrskShrimcrIvlHaZRY22XsCT7oAFbyRzXGfgOSH0iNzKY8DWgq
hUkvIR69/sC+uCKhVhBkU7+2QaKsqk65SnM/5IO92dzzhyEtc2oypH4mL2qpVEg8
9PESjeE5VQfooFSpU5sCGyyhInacY8roZfqHVjk3CwZ7fAqF8IbYtAt8nQuVxlUl
3mTkgKUrSz5HeVfLEq0xvQqKHLVJolyD+fsvxXKHL8hO0EkN3tJd7Kyv2djIWFyr
I96+aQ4nribK6sJIz0WZpgQOx2WZX1VL89WYaJhAtttKjyrlsVX0UNmbhnMLNxp2
TMA/M4tM4/cSG66332B1Ou2FNKMvtZUjPpwMOtAMd+Jze89Z7YCyW4RFk0JSePHq
bNatfv9lGy1CwXZhqeCRhdvCB9Ii1iAr7n22YWwS2g1z6b/1ykLv9dldPXT3ggy1
PTO4912DcA5unT85mN6adt5biS3KRdN8lzNbLT5Jv6WXmrCevGEyuWMF3qNggqRj
3HqoW3qvfxSjzy9uVXWw3OdCQrhjKJfZX9jZQ0C3I5rB2wvmuT+r3dyUXX6sWBzN
2gubYMkgj7Q3N0+CH2QVEfC4OFtJyGq+Kd+9IyGfZRNtQHQd7UMBPoXszk+O3TTn
imSt2+RT3GdZYYnvX1hKf0cC0kxq48NkRnSK7LSRl+y5UZ+W6MtvXnKgCGHwfwy/
TeGaUwaQqAYg/MBQDI9lNc+JMzfE5YZ+tWn/tDRB8LhOlxBTSK6nh9DDDjZPzHlt
1peMPRWvCe5EDaSICipnaxavdBrL70+/30fcWYUi2tKZXW9mozIFeMiMeO8WXA6s
s1iatajn7N3GgQzB1i+6Y0sJiHHv75H045QyEGnP9LO3cvXV58qAVLyX09VD17Jp
5g40U+HEd2xO92B3nI6h5z5L8XGVO68ZmVRgzGCsJIkTTWkM12N7GnKg2qdjDexJ
8da/d2Hz4k1kd0NXMX7x1qm+vWAL0ZbZcsbTbkgoGAVuTL8WIwlKBdQLN2vLhjYl
IjabqjjcQZC+R3Bq3f0xHG+EnOthbw2YQy9f/Cs6xRy6/MveWk1dleXc5+HoeXSm
PqVEfYxUQnie8cdGa2cln4WDS132w3t1Wjng8MlKY7QOtckbs6bt+gas+cZ26Spf
DoQqgBVAHYVymaGCE71QB93hSDBU8ic/9V7JFdgXqhi2xuXm20Vp4TFjGTzza2tY
WbIUnzBIaxZmsdRbq80XdZL5JrqvzzgKsXm4FKymIIY3ny4CGEeYtwJM9KFP8Lob
3a1SgrmW1IpziMFMkbwT8RVarzrzURjQXR+FzniRN9Nr9Zs2y2kA50Nn2shukq4D
BWmz2u9der/9dSxQJSbIXvpnyQojuyI9+bOao8+zQqA2fxCi5QnmFiPnCUFrOk+3
+XfnA1bpQkJi9QbmV6uE8RCpCED8VVRo+SHs2Uanf72SjWUMkSzTysZsK0xg59fi
tRLSOd5Btegnl4NYKGo/OgOfLXm6SxOdZQ/P3gJjAq/ztI/OZ+d0b6eYEaYIvkZc
TpA65uyeQVNwB5fPkY41yy2mIqkkFKomWlYPYVm9Ln/VhNXvZmq1f0NqEUnWjumG
Jkjn0GJ2gUHo/hg3K0MccNvdx4CHT4WKtL5Zq4hve+EwGNqx7kPKgPrfvx2fwtEr
OIM6QO4fvZntDHOp1NVglmYacgkepqr1NXuqVaceF/BTg6DIRNHjwW371WWwbhBA
tZJ4V4JPi4fLtnPc6dIM5ffQH8OpLwteBw0fS1zgqDwGLkSft2mpVEAHhL3B+GWw
rtXFp0uLwOYceCmvaS0tKiVnzzKSyQZV3ZwI4J9782nPxxqlVG8/9SMNwLqCEDmb
CPZK8aEf33VBFP+oSHn1dGWLwPUcVoLC4HqttHDgbI2IKSHes+AAWlNl4IIroH9X
YClRtdVZa+4h09H6E5IjgLLwh/VJTHtKZL0KoAPB65A4+2sQl0A9P48aJDVC9uFp
BCSU57H8BAwnlVa8bBsIAHD2L4jl3CrCu+baQHobXmRtmXXwXds+xxcx+Fy0nrp7
LKG0XSEKERmFZ3mrwr13rUxoW5lAye+HOh6DsXQzVRKiyWLxGO+nAy9RKZqQAIG4
NaBRBxORph4yDp5I2bt9W/vftu0AWlrVY3z6x+LoXfUm45Yu1V4/yfTxVfacGfAX
GTehlhrRCF88u13CKDggdCuUJlcWvefMp4fldzQjBPg98H5chHXW1LlCZJTfuOK+
uz96bup+TgPrNzrd0J5KjnmGCIa8RFZLWzSbZXPpjc9vyCnVVOiifE40vVdmJdmq
y69je0qKlGv1d/7XeRbi2PrfJqMFUm7dZ7pngWKcxxHnR14lWauuZaizceGeg3/J
lAkMVraW0CCehbTgwRm8ma+7uPbeVha2oAhmXy4NZxtA5cgmdAJ+tC8Q5mcToK7s
Z/npu/K/PYkYe+zDKhaN91t6vF/WuJQNphGkcVt5M6eYs6mT/wzGO49PWK9u1Q26
XtrxWKdJB9sPTJMhwLi+bQzTrrxk0nHJTX2BgNkGBevxez5G3UxB7UyFlAw+JSYp
pX79eTIv9k6fEFx255aXRSZfVSgbS9jLopVqLIJg8EiM47qZs7PW60U6yY2qDVrs
92DPUKyer2pRN/LcsksdiTWpzUjihzml6yRN2VR61ynYcdun5RlvbbwSe/ILBAlm
GSY11/i3BPSv7GJHeJudKwo0XWa80tZs+EH0ya19WAyu5PDHYzb3tnQsRlXmq0pL
jmnj/qEIV7ZWiMzuDO67glYGMi0N8vrYA6W1oy/HHYF1ug+eRNMlHmzIC32nmWlF
YtKvN0NCYs9mZe6FZSI4aO+a4lEGUzRtrQO4KcSZYxhigc5r34YfKu0mRF8rUmvh
O/aZTB4RPVJobJlQAjs+ng3RxtLBl3U+fImgqHJyZvXcd71ZYOL1ky+o1mBsOnzz
WE8golSMrmXxYbNIMxexumJBa7CwHZlDEpkUMJdOsDfJLkqToccg3NFPOz+wJnHn
Ub97sZ1P4apiCjJKDnmw86h3GBUfW1hmf2yaqYeYgzWXR+FynSo9o/37WO6FpGnT
GPRXLlSA8+D5L0two4YimgmQ6DGSUiZtzHSzFvNqX1xnw9bhw4VL3jXsVg4oJ2zH
S6/+J9S1RFnL/Xf0YVCitKxrxOZsqVPPKAPaguqysZ8E0mkvNfPYw8YyGsmDuM8m
WowSh9Jw29HuxNDJATSOQsQot28G6rqX8IUeNmDy9BYEduV7O4lc6P550BVt7xd5
M0vmlQ2bKrj9no4lvgpSc2aWc+MXyWvdYGMKvF/8Qy4Y+gJ/r2zpnfSbSd6wTa+e
54iFsSbhusL3fEGUFDt+sEaQ6rM6YI7fSq9sz/7aPXg3Sdktu8p9q+Y3D9DHqOwC
YnpCvJ95id9Peq+j/4DJs+7KKvu8IicUW6GFSjooTYekZqqfWIngFj7anoo9VJ/h
0wcFfW3nNK6Oq5IV3r6VrHjazEoAlauPRqAza1AQCAY82W1FFK3AQkYxjk73QJdN
BZIx+F+iniRFYFEaX6inzYWWV+BcFMQjsFg0FNds0qavp6D5RIp/wn8b0w8vqpqW
ys8hF1TEPaScBTSNf1UyVctnHYHSStKbkPj+dkrAxllJS0a+xSV+33zgMZZPCSnI
Fsb2i50GcYpqMvH2Zftu9hd7O+SDRt4355tjY29O8pFP21e52FiVgOMl2bAG4sid
ObIjFJC6EepVs7ehrrJ4Xc5fGdrObbznSxKt/SBd4NHn2dF+GpPaurVv4GOYdldK
3PdWAlCtAdFZO09fj+kJki62raebkwX2+JSwbvr2gek+M70HrKgzFDXYBIMiNDVy
bn7y1HJirvTtDjPfo86LK8CEzEQd3N+9LGhy0MfuvGOacdnm5qQ7mOpS/wrtmMnL
6457j5HJzm0VvznrYqRoKcIxuzG8rQZ6/8Pq2b2Gzm+soUoypoZuBmtxbu/qcDWY
CYdW1WkweY5WBvTwj3dUN7NX0ur/B8/p2JE17VKMnkQV3SX0W1HeGc6GZKUJuSHr
pT3A85FWcK4u/HliXf09mmj9S2rDNpvTfPCYefTQstWqxh30jGPov1Ue4lPRDrF8
30481dGb5ke4sBah+wrQ4dd2gBXllV+UeyF4u7TIFwObBURtfpREMleQz5VQ9p8M
RIxuzsWGVF4/3haySIfaStuIDia/VB/TcrgAh//KqyKsTwuPGwSPhQbU3uAHdtb/
ySfEiMB4PHKeAsvND6JOZqsa1kFpr8J54wwZGbdB5ryNIkhV1oLPSiuX9W1b1Gca
TrFKRx4vb4I1/srsZtZc1ciCV9IOK+9hwBEC7p5Ut046I1c/CDp3qHXF+UTpDWGT
d1U3xXDWLNaFlynTmCRAdKfgkgQi5pcwG8+x4tfBV2Ba4RBd0AJI0xxsbIuSQ0Uz
zRQHTN+oaTp8ib8ybBIPCGYb5DBhny2fOF0LNPOTGWjsYnDAUFYYyJDXqIlYemib
jH5tCdgMm9pdXVZbkiVQqwnFG/MfuZj/y98u2ZJGFM5obm4OqOgpSGp4ehRL4jsz
lrIqekYGdiKswEV27PFAgyv+MYr3LFoFuQOyeTqasm/X+rS1+wpLsLQx3xM2uq6n
rK164AP6R5pWsPiR+Sh2HbXwPjkgUrf+fmzY1IsM9wTuGcc9xnp9kCwz2/ux+Mlk
4IfI86PuXMKENtg0qJOrei81YZ2xEThlg/kG30fVKvHH59VGC/rGp+ELv8Dz1RCn
Z+XYBJzJJ4nDmdodfqJzJ9xjZQDYgnxAVV5rykjJOU+hb6MtZPrIgZMZg3YPQyP7
oiYuVNyr0yAHDUylQgrVrmL8XlVJbgj3j0a6tnz/yVXU1TuunAcwjlnp/L7jY4TC
neC0K5ec72CFd7Xnl9OYLX/KHkjDiBavmvx+lNtnNE/J0442Kwpa5A9YB0zqcR3K
yaMkbg91SgT2KQyjoI0MNT53gyAPY9LCPxd9LYfCABAcWgkcQkAwOgDA4Wx7U2Rq
R3fKEjKLSMq+IVI0Ttp03Opu4rkcSIUDZu9PrO4p+roTqqnmVslJx9j8qEolitzK
kud7+Spmq1ArWZHcsW5wk8Enx0kkdA9aEdRvoAcjiUYTyNFTJZU2O9QjE+vVYZQx
W17qR33A4x5cUdhojN1MUAQNztw9mYfgaiovTlHRp4OlGN29oJ/RClpcpsW2JHe1
KB0TIpcCB+6ULBJsVHcejEiGKvmW44rKx5PuYEznDVDjEZsMpKtZ86CYBaThlVca
+bvkLBc6e+iwdmmdc37cxS0MbgsG4hPDoiXT5gFIHaOzLenkhWVSU/P/3xW7/Tkd
2AZ+FjSe17BmD0h0pPMVaDJb+2JiHoQICvSwkwz17xs2ihoDRnWYrDC+UNsgemdH
A4Fu2ZpQFwCzRR6wscMmdC//C06GycAlk3vULf65aPlLhtijfBnbtt6h4SXRWVl7
IFQLeFBQuleuty5/p4m0RUkwz2OkQqCFt6o3UpnyZ3ZEnDPFO5i1BhTb5C9cMV8K
kT2BeZTMUBu4czgJSuE26X0Aipkz3fwgzkNx7qvbneWhn+hpCYq6Ii/VB7MkIVC6
3Tdr97uOpGQ9LDYJHZfv7tS/ZXhiNdAe1xNBARwiBqwwqiJgna34MuJqLi5OhOv7
A3ozW1TFc1jQQin6l1a8mCXuqScwuYP1ZyQHcSVU8Qy0tPBJfexI6iptCPGvNgnO
suJmgFasACAUPB11vw64MjXuajaT7TA55bMEjN+glNy1k3U3ziTTFS6RxF5ysqHT
BWzeJJY5GEp06XQ8CM4E9HU2yDuTT/6NCfFrd0qKd8V2CtFrVCKjZ3Iy6cDw61zm
uT/38nq7PV44IXAzI0tZcs6UxeownwDURkp6EWyWDbe76Xw9TWcBY/7Rye+8kntY
bi7VBhic2YSXNaAy8Hqdd0uAt/akRXPPLGrJeshYxBlfTd/LbxO6UdhcAMq0Kkfp
iFFJ7s7BhmmkiULpIHs4bX/sl6ORp5vPp5nCseUoH3Ed2h2CaJQwu2aLHe6mnC3P
D9VdU0su1shlpKSH0IiVMB7xjfRc105rTOMnQjMKOXCwan05zmZ3xgnW3AuQWHP7
y6egTC9M4YRjC+n9HikWBzJ/QH0gvwhJK8a33Hm+0Y9kbIEFGxJjVDSD4h+DuEku
BQVN2NwYe14RB3olIMoSLUOEWlflavgR5+IkETEQbURd/s4OX7BXdTMHuL5ZrmjS
Lz7AhhwhdGEBGW9wGvL4xnvSoFcDmGv6rSFXyYWIDYSjwghOhfUS+8v/Z11UZfm7
beSwyR6BciO27Ni0OijfnizTBybqatzYPiL/0rqfJMikZWXLt5lsgkcR/RiPbu+n
HYHHZLeHNgFW2g9V2Vv/hnvMZc0P71/r+Y7nwmT1ZjYXAHoXPOxPZezdpAb/2GfS
A0jVanR1ZdMZvVjZ7pvnyTG3kVpmIan2hys4ld1MBiO/r6ZHRBk59qoTuUGGtRZ7
c4XZw7tuC9Fd6PGLtSBRhIq1soCvk9DvZBE56/cyheThf6RAsbP4xbQXh4lY30Wp
LRjPcY9HuVoyjbXCaelRdLERhIoMoQNXrse+3I6hQxnMQaPAdNeT4Q3bOq/26P3C
CQJ+W05D3tFh1nzlW0elgOgB8OLmLE745rp+PNgORHE78yAf2qO3DtaeBdzJPzSX
KMASvkblUmeMlNt8QTTS6MFDOQdbIpu8tD1xg6KukU/mugaBP1aiIYZgSX3BOGIc
YM5vQhgw662TLrOykhuU6sIpNabFKjjyK3Umk9n/V7Qrp83vEaSK/xmXbU1NBp4q
N7yPOB6S4TweQvON8nUcwiB2b4cZ8z0z2CuUNrB0SjJD7Bjlj42H2hvAxPYzG8Bu
SKglsNM9V2fyb7h5K8eTMWPJokhj13xkzDCylBhWXfDl8RY2aWEa4pCEaLv58gyu
ViIUbfO83K793OSKGe/YtHaS+nkqNkMF5szY5DJqBVZ9DOxbKNFobygT5LZ8RKF/
d1o/42+DdLdcqwGHVJZQ2XgaJ4reNhaa6hE07GBAHYarJ8izlBKcBdAQlppQ9OfD
OqDtUP9HSOxUQVc3CIfpTteuegEFVrSrM+PYAtflwHLEB0OYLcev4Wht1MTKLu0U
sLjixXqpL2riOPO5f38Kuq0YaucrkQboon32qRDx45bz6ronKCQDqKVIT2SWuIxv
z/A+XbSrap3MJO0671NHhJm4CY0tMi/VUKoHX+eggoT+hv+soVOQ0FAOpaMmBW55
d8ggFe/8F3lKLwjRfF58RF5w4kTZNxapeViUYjKrVx2q944dQdzSBdgdWqXwtIyE
Vm3V9cJ89Q/UYzpLJPjatBunxva/Pf10mFRCi8c+UO/eN3ZtKkCCjTTfS1OKgmAR
WiVhHkmeHm5IyJXCIiLV9l7FesvnaYuMUiUw18xgx8VkugNGxDMcvlA8bIJs3Po+
WXhtlrctninQfyHKMm4pz9XYYDtfa15fbRrPRXB/w9OQ+NbLRX+3NrqtLiDKzvy1
eHQgBs+PViADnTkuJxqQs/p35EHWnuZS79P2tfPWSnhz61BaeJRWaipIleshvQzv
f1ue5vEVHME7yLpCvjml+eFaTHpDSsZFRm9umB1wGuvqy/Lb4wKBsSJ4c/jNPlr8
PxcbTowuO0mXhBVw9SVY+ouMt1ue2mOna1MVbx3VsBgHV5JIS/RA4SPNVr7g+oFp
CVv0DPZYsjkttJXGEsBe4x3CDRnGD9bNjXbpUp6tVy5QynBzmGUkYN+zeNkgrN7f
xZjFb64CkJ4MH20jBJWQUzAkngc6gFT7LVtZoq6hitpp8TPRh4vPEK34bIXxhVOr
9P/qV4ut9lqM5ZkuMnEEZFg1ixvg/19+g+YrhPlkCGF2vaQvuYgTOZv3kGaWddLd
CUuajs/J8YnRmI1o1f/U22RPe0aIEo0Zys3oGU4vRYi7i7WVhw695/QL4eH/Qjz6
t4K/aoPsQq9Hb6mcZ5dr6qpO8ChPpASGrr5SfCE5mwBTehV+6n3UXpO6EmZT5+ZV
A6gA5gIx+Rty1pOEGVbtTL1suTHtbpcd/L5CYB84ZezZHaOod19XNGET1WHDJ+vM
kaoUjUIM9MNI4B0Vz6I1auGhPqJPlrEjP489ERF/zPLkONiE908W2Yn/QbE7Fs4X
EItD8jfU6G6V/6AnvdN1/xsWxt23jxgEd3DLFaxFoANmkAt8caBxq3PmY1hGchxi
bePBVFS1R+2m6IBXCOrMUnwWmkXLQZSTeQmRNTPp3ZOi5xL29F501ycRwXrnHb8j
bBYx3rr/VMivv4aKv6dWHC9WdqkLG11F5aG3rvuYSxwfh9XZ3Wn9mtSA8PM3bqUg
YJbSOzRN2gC7EWRc9AGeyrYMnJyu+wGfVPVS7gZKkQ1QncGLCW12beEJGkhGRmXU
PZ6iD2kXzsxzpevKarUgYWA+tvnUwNInvO2JIUFmnty8EPkaXseBzIWYP1GB/dJ/
Ywn154SpsdPCEafMul1knak3xQHSPvJs80crUY//0v+s5XUdMa1Hr1tA/n7Jpunz
Cn3dHOmmcFWX39y3riBSUY3kl+QoSzaXGuZYstBiWvsLkQpW5K3lfI5K748eQO+4
itStxqbqLPgDcNltqCl0OZTbOsDglXV/C3JnE/rhjexCFvRykudSWk3CwWnsNKr6
6qY4nIXmKJnrSfHqrzwoCq1yCwqkQNtV2Hk3bLOw9tn3yTRj6/Uv+XrdbzXNxhUS
+H5SgkYUCamqDCEtrTUqL3QOgVytZ13LiacOX2cUDPC6gORHf7yscY0dV4GK72cu
c/+HtpTUn55VltW1rHe0+kdkcxp+pGk6NGdIFivjqR5UxWNi1sjgdOYS3AWvk2gp
ValtOAR34V0pNR5mNJXAp0tA5zIcIb5jixI7CpZekUhpiHYO7SxhA1Pb1eBp6z5l
xn8bPzZIZxd3+B+2RvgArduCYo/iu8ieXxhlxv1CJmE6pDr41F0ARp6OzzgXu0P5
DkIiZEaxqp6b3MgeiqZA8hnK0qo99wlaYYTwA/8oU5RvTq0j7Ya19ekrR/m3zzhv
eInbOh5P/3uts2B/s99YPjBhbO7PVBIB3VOUqigdEffDjFX1p83Niu7CtiNgz75O
9vRu0Y7NdTabygSn17mfOd3gJa5mx9qho4ntp8hmRXrURLF8VWypCospwsL2RKIa
YdoOUqLE4r48etgMTDDE7SFOj5OxCIjIOgehspoiKuDx2s+08u3NbEEdxoHUz50K
kBNwm+UNdjlauokGEvIxSGTkagvZZjQF8sHswM0beIVcKwIZqTnuDNebWpYtlNSq
qiRVzaObq7+aiIqLQmwEzReIkjDllS3Bjf7mvM/cV+FR5HAk3JB2ZZkjLIvrCtSV
XbrGyHfPX63VqGOsGngtZ9dwoGC7BXs7CcSWQ7s/O4EQHs9RBCFHtHAw/sgV9UR+
rLCX8+yX5ZBJW/ttqHLv615AW9lNJilP1SMsSeo3QuDGejOyl9uhKuDEUTWElxl3
9zk/venJUenkwmFyS+i7+oib2kV51+rqc5nD8mAft12uHo4Jz0c22lFMTe90MWQV
hQ0WhPyBh+v8aZpS+6ZXKFwyW+l5BcKc02WP9nGnJiHZL4HZ0tSUIkWqkw8a74jv
BjmU/3C3vsUckdyiDflipwsn7leT9NYLyjcrJt6J0jABKVGONOpR68WAuQ/Iug/m
vKLb8+41c0KghHOr1ADa82o9NAwM63ObdzuC4f+EEOVmQJAyahBNykZnA2h91/I3
Y9S+9Rb+imfcW1THQfqKEK+F4rVAknZNniw6Js6XmrRLVuchoSa7IB2dridylK/I
A6o1WIAfkBY3PH2/B5GWzoTq52XaWfhJ/29R60bz21DgTBkyg1MDeU+yN6xal3DO
VY3vUtQ5jFWdSOVLi4vSjJgS0sWQtPRMPB79vTPWRjyy6iEwZnZDAoqVmrr8Aqzl
HzTjdoKD3iNSyLEwLzU0brAB3+xpidiYR2iH/9x5WC9jWMDlEpqmS+KjYev3x5Fl
SZdUbW/ESTj1omRqaz/y7pYG3hiqbwo4jsakDj4A6COFrghunde8JH7+1bxUuHoF
fAeHzwDZrutvCfY9KJsWQERfj3CW8EIywb+PEJgs+cimaVEyrYOkFz3oXRpIZUf1
CY7eFIYgDCXeivKK4B46GbePjcSRzslljtF5rYA0yVkcb2Wdoclewki6tRFBrPmU
hQ2yzeZik7OAX2epMqdRtHxwZahP3+nhSPO+CMWLbI6Kfa9gKgcMtdei9qYcbOgU
03SqWK6oysuJrHapHn2F6gWVJDpYX5gdPXKlB/HN6HjHP8JIZrq/q4GSNIp8RMVu
ChJ4mKSmTJNwr8xKonix/+6DESsw9y6Z53Ixi+ROs+xLAxKIRtEuGTIvzs2wUxLZ
uxlReKjiFdUoX8EU5gzdXMzkWp3nEzDUPUg5q5yjogiXuXJse75Tc+Lab8ZuxrzV
2J5mLpMH9aOo/XKcsF8KLF0RlK8hF20HlDTYuF1M0qVTojRDXsRSFVrEZob9U8Aa
eo5+fTdoFI453N+JRxLHgFDLFuAbGzvHsS7kTAGxcvpeW02f2BbxmzjYc+FxWK0M
rtfL50WSFK5XMn6x+frJXNdad5ClgVYthIydPRQd/LmXLWf/x5+2pqzQE6fy6clB
CIblt+sUqEzKtbzVaMxL4s+1o1eohblzz9BiJQfui5MLt3OIWMBD6DHUUadq400I
UNp5mIoSVKCdklipY0Ue9hr9PLDY64P/2246LlhZTF6x/XMEFQ7/ogeLPOsAygJv
y+LC04uHvTHGfV76khu0Q4Vnn6/C7vYMZOuMAvtQHh89ukcKAGOYJn7koTqJWdNR
xvQB4xagS7KAD/W7VbpuKGBRlw0rqbMiyqpU2SdJD1ykNoDh/6r/EB+ysoWVT36l
BOhAo/3QLN6yuN8kE/Ly/Q68krSMjxlxaJ9+jav7lbmk+i81fCMioGP0S27PQOfO
LFGruBH2ZdM+ptFQnlgnnsN5H4UrMxX7mDEYdtRjQh9iZlBxc0rDJqLhmWaeH1+/
AZSk61QfV92FaOmgY3re7+raS0GK8SBH1IcVyNEyPqjWkrONQujJh9K4SYypExTN
mUT/LngTcEu3ViiHYdcPST9mqPyDBvlUIXsHXzBKfOoh/g9H2eCg6l8Jfs0RdevD
ht9+AKOc6uR592v2hyENUopnhokJkxowucbqgADi4IAESn0J7Yu54ZbwO3NKmu4H
7cOZ4RUf5tUcrOODFyZdsq4s1uZnItW1ACSa72k4S6uPGMaoQv7VZ80znJvAKz6o
ueh4TEaLcka04/B4dnenAtxA0Onlf9fyqOwH//ZeHKzmRx7s3SqVFjZFEFgKGAXf
tkcWhjn/DAqyOinEQHi/48n6GswFlYPYOuZ7PGR10IQiFnO1bhkYfC0Xc9vVMr0A
/veJ/74DOB9nqye/KijQgLrML6AkwCCaSd0r9KL5etV0O1DCwQTCjjirAKKa5RSN
3wnr3STxT07WipKjD/wsJcsbQPJFoOXbnZRidLdGH/tMOx+ni/S72w0XhE+CLN6W
yJQuRlzIFkup3Xoidp4Co2EqgYPfj/RSlN/88YtZ/0wjx99XZsrsHuTA2DOgp/uw
qk38i4a0otaU5vOGM7qSv/ekH2ReFlbok8n5d1Ma1/xW9ht6O+fZwosx0tGE4MWp
/SmljMpnYDYyGxHpIwo8JcdHyg0gGztPzrLNgeWta9EVkG/FItMO97Pw0jYwDWn7
mbfQXzZ2UYNqG59lQrj1j3zOpUngOy2Fj3qK9ynkzI1q3ybkJi6C3eA2hvMMf+k6
aROHZMMMH+ZvWvsTneUoGaq2ghfHMw/ISx0t0e714OPVAaHN1EHy3z8sHYJHWRan
ldooyL/b8x+v0rEMdlvRHGX1wmUCB0FPn5PBoj5Zz4IEQE0XaH4ugydLWR/4a8ls
gmoe2Ui8Y+tNATgdlFe1UAt/8R9cfDfl0mavu62CY+Rrw9xjzFEzZHkaX28bGmz2
bo9KYzYpwH+Y7gccuXKVjFnu+yUmUhPDpF6otWrIcaX5Dar+ZBEh2GFM0KpVuiUT
j9kJQxyAQCE5olkv6Y4Ddy5EZah4QTtujwTmgE8Lvot9xeR1Xa7aLraWbMVGoyO3
NPwNgu46TYadQC9oIxd4ILjzpWy+g8I179nRq2SYAmHJvWDGifVCzxmB7/xlTrO0
mShCJr+maEUQ2eT07ibH+m0d6F7yUtFQatax+Qj6h49UPZXEu9CHY7L5MCf663et
9+J0TIxByhqLty0shWEcdlP5s22Bpis7cKKhlxTOUIa9lrcsq6PNWRXVko+Qg6dY
osyQwXAXmlI7KhX2mKgFMlSjSWrRDgxT75gaqBmCzNkM36SMqDaN2pCRwNEabC+o
FU3RgVMBO6cfy/tPqL3YWS0MtOM0JYKV3o5Pvzn0bZvFJWN5aaTVFPgLW4hM1G1o
LpYmd95mP9Jng8e8l6Bzz0l5mBJGsneS5qBvb7Bxn8YXv8XhO7wKn9bfb0FGWRSr
qlwIDYbhBBUoz1voez9aQXHlb+iY3BCcdMBoPlQExwaw59pdYQdOMrHl2BPVybVh
bnXvarR5OuK6ZWFztiNjSfu+8S0MfkP6QSr3IjJyQXXDk8clvpvyn8JVcmOXODoJ
26SzXtxoA20mnFdjmOdqPwGli5tHVUVMchjmYydKfuKkqHyy+vCgEJSZHqNjxn8P
1QUdbUjO8BtfNJVwKdYrSMyR9ycQi6Wp1uTrGDV8op0pmNgx8pbXnCRopqknHFv+
Zy9W+gzCz6tyRz5LxfouF9v8en4chbyTYKF7MN6E+wYNQMxrrZJzvB8nchFuOwDL
Nmii89gyheYO4KxFTXiY+Tlqhgy1teIuEsvHRVBbD9ZGICveeB10rVFSe9qlFAc3
5ja6u074WMn1iXK86rCxskb7CdtwlV3Al6/QjKVoewiXj76YaWo5+KnO2qIFtFR9
Qq+lit9MH9HN7mTIJGf5SQOYASN9wmIgQqzF1uaqZ65QOcI7nmfn0OmRcNurlDxl
766gf8rQIZUcabrLaNvtLFTqC2Uu261MaI1S+VIp60Ih0oyVcl8/AXPT0jKkz5T7
M9zbu2QZSIoDHHafPQkMNEUSeNjmYKvf3B1jk8E3TVUc4nY/c3wIYakREZtID3U4
6HrMobwyWHraV7krwLfNe4T2pv5/Bor53vGkm7x99bNkkmi9bW5Co9sGKfMM9zX/
I3v4gCjXfoF86mNAiyOgyn42VzgtGXFB57m9/SG6+l2YVRz7ga7C3CYrfVYRIRoY
pbdV5dI+A+IX95XVTWdtQVTtGBluoHHQ+4kyZ2lLW5gesCyu+zcnUiCKoKm/0WmX
k7Q1hg/7pHdQKx5MQJWBw7Vs2m6Tsm6HS+n0HPzb5RK1QUqTM1C55zhpMhiitcDb
GAFZ6ABCqKhzDaIlo7R94Q8y7lahhRL3L+E6nhxrLf4izf7OrhFBw+gJAatDOLMO
Ib+sjEh6Uj4gx+y2xEOe2Y/zqgtoaXVrcadsyG1pBE/ddyGtQ9iWBEdE+DmbeMz2
VGAomfa6A5BiIMDqpR1bMzvrJfa7oP2ONcXiqeal4vA2i8DURBb18Fo3wHtAIHhg
UFyPE9EWL7pwSl4nuU3Hnz6a7E0Q82gyony6ftSC6k3iKxmjmqe8ovw3pPbapdJ+
gxOzOh/lzKgz8WMOcuzetBFbVrLEYVOPbNH2PR/leKGsOUtxPXZciL+yLaf0ZTiK
qptmT/1Y7I5tc7AUs7lGtzVsFRDqmHPAFmCRBtNO5uUcECYG4mUtMTYBHwwLgNhX
8EG0+1CJlfA71nsZzawefTJHWKssQbQlMM2f/Fjd11b9Q66ovm+/1b4agQu+jl/D
/pHFnVTzAOcJvCZ6VoVEkji+7Ym+i2Mf96IoDZzrbbalSCcWSB2t4iiNnqtdS2NM
dTLlx7ap9UJjHxDAsT5Uk639nSOlkPRC1IbZ5s6O2qsrWWcs8JJT4qLY25ID9TkM
7a35fNOAVbol33Ha8i/0Koiwi47upx38seG6CKTW+PMC+texYnSYoY11j73VCmk/
tTIqTdCpGcIWFdowo3f7K3Y0MlbeZD4KRzn7F1gmNYkoWJRQ22PJ3K6YQFs0C1Wn
7DSxG3gn3V2L9EIcTkftfgDbK6RLFxY/GHIfNttO45xITMmkxhNuCMvwJpQiGtKt
cnadvIyaQelKMbwyAlwm5VWFCKQv1jxAGII23rQ6LRPbon9ufbflx0Sszr9bDpSs
UTOqveIAm2/uJ+lXxokBCYtKYJ2wKqVF71z/xRC4RDPsmOSJUTYiXeAs3+WbBS2h
CT+1EY8hTTO8Uz7MKUoIPiJgFVmURK1gKyJD9OeOBK9r6G06h3X00PihdlzO6FGq
521ekz+ttv/jqKzniiBi+bgFbuz34flvioK9KBftumOQdCYX3I7gRiZzLm2WPa/m
gYBCEANBHrGgeX06egEEhNILzjn7wAGKJPf5iofnJcUhBJDRmYwM2kBvIPvL4Dn4
M1uh6DVMFSUI/XcANjE2rhnF+/XARP5dXdHGnq06IlQVuFqrM1uhvZ+jJvD87TVw
ldZOywCDqm453ANlCnPgCCSrj+Y+75rd5bqekUXkwQlALJ43omWGtEnEP0Rzrku0
rTh3liPf4lRrW+zavshQUasIPfwKpI68O+mZi/KTD9ekxE6NmFGbG9U4UJGIcbfu
Vaa4okzhiVnaUbzJVErMxr6/FrVpU/9L7NTWXIsoHOVRsY+4kZX9ZBkMthpeaGVg
n1NwN0EjOAchcMCcGuSwg1To/c0UvYUio8/Ed5tzNh2kA+MBGPpHdN2gT4R8UHtw
ZgvE9NGer91XNKxuuLF1LOzs5JC5/xq7wTgFftHZj+ArDNkb58fUhXSGvRyF5R3c
OWjwQu0tT8woknWM+/dvTgccjktkUbNYpevP5gBuvrTxRryU/D3zczXhGsv4/6iB
hHCB93dbFIvm5UuIpHlkANTLzb20bsyUBRZ6bkl1fNtz2e7ks38t/5YqAnbt5yK4
w9YULvaT7H8CYBoip2/2/GN7UB9w28Z7nJ1+I76DtL/0Gf3sOchcPJfxhHKlRbtC
asYR/jwGdjrKZFPtpoYl0gWUG3TFK0qdzbYxjG9hMMicWvd6eMj0W+4bGb7q0sxP
1bd5kBpo4fK3ofzcc3+tSoPaOQyh4KPph4WLvC9IHQ/xjhTMGuv1YGZMR47u+q05
g5vo0TjSEwEWUsl6CnXcGS5sVRQwyDg3ZYlachHdO/eJ0t0QvYC+XMzgRduNLxkz
RKhc2B7rikaZOLdaa6IsMnoNfI2c46iilKUqgEREkIfx/9x1dwC3ssqdBDugzOje
l26JEqSSqiIBAYRHarMdU4PhM5tTsziv/CddFW4NFSA0fzgRFbGe/h+nZso2vdZ/
pmouOFAlv79lcmGym7LvwhV/ztlRErDalzhzZfQ1RVsV0be8t4sRtINO/BqyXiW8
8sI7Z8dG8Nze4xIuDn0RUGZbGCnveG4VhL9saKnp5MK7by+iYoeteZlK+Fmawmqh
uIVlADEgVuSc5Xk3BSDbAFV4hXVhuvR2hbeFeauc2oR/E59wI1ZEUIhyOaGYqq4L
twfjd9a/EREiUnfwWg2xQkIT6D/xxap558FSqFDzK2zaNGD+KE3Jtc+pbwFAMu7Z
XWNg6XVua6hvtZudFm4beDkKvxqHj7plXiQmhYpMXO/0T81bkjNFud5zN45MVima
2nd/jpgz7IAteiuzBHNsWaLtrZkVtTQNj04dnoTPgrqvac5LRbZY7wT4B+B2NApF
9Yhu14yLyuHiWAWy9YOH0IAQ7oq8OpZvaIyBPilu6YD1KeAbwgo+Ki1zfBu41XB/
51k8bd4wHefiyqsgsGVplMCMejN+6js418gzF+7ZEybASOb7us3O/jtEv8v9AWYv
hMry+Tiv5nW5Cssfb27BCcdtxRDkMTWYmbezDB5NqlOTaA+bHC5l4Z/wK6gqyiyz
5xTl5RIoOWMT3qPtPtUYKRtixf8Lz9jxbANtKoLDa+9rTQ5ZNlwHl3eXZBI+9jSz
hm3mGVudlVUkmBXzMbHWgXtUzueuPz2PAO1cgN6/IER/GDN7TbUO2A6VNwJ6rbOF
ph7pSjzubxJ7nkcfpyHemEYdfls3r3O3mW58YtcrjcUBS44u7+uE98BqtR5Dijq/
a5SPxgIlH050fZpggDTymFYeawMe0H8yPwQXcF3Tj3qx35sCH77/B1yxNFotiLg1
y2cGw6XsDDVGqmydbAHftNKr08h1JfYzCcyWbKZLk8jLFuKzWiNQZxqvAL1ylqqT
iLo9ATdrLBRuu8cx96frCse80RcrVjn7WGOzcx3BwChL72RZcNMEdljzAZ1FRlJo
a2PwgyRJvBpxT4c25JjfH+EQNyfcKN9jPMwUPBl1pCS5x83Z+DTNMCg0B0vUIotB
scoJ7iU8a7FBmQb3dSHyucUbQgBezRqKyHETznLHRQzKP57uIuk8Oxt93mpb/Iyu
b3/syhbRnnjl1HjPdIASyagT5VyzqB2FqEkbJwskBjoTGu3aWjat6qIt1JSsmffE
l2Q/uEuJtuc9WASRsfhkbtlrvlT2qC+z/1oeRU1BlqxwugWm8lSyg/KROpRITWrE
+es15/Rz9vbPf01kF4t2nKBWTYnoYB3+sxyzyP0Zf/lCYS4T4D+lrd9JxVwubYra
w+0nUPrdGSpUyvliwDtKAOPmqusKBNEWxYGe5V5I5+Doh15F05NE/CQu22YbW64a
vKOCkY2jX3kkMS3PlREnzgF8XHHPzJ3iL4vMtYph9QFY/XxV8LItHbaapsLH8BNM
ryjyt/40kVs46PRGJXZF7A+8aYESy7ZxmBZ3jLNDY7L33BR87rzdHFg79Qrj3N9h
mOi0sjgEopwmpOxliG04HD8G+WmnzKuxmL8FSVnnXaTN0VgoZeCMB2KYf6ZbfHSB
yUaoMVLg1uztGLkw0S9zS27eTb7Wb8fBIEx5FVl/zF43cv0MyQjiDu1eENpYMc3N
jfOJvhTTnPhTWueV0SXqmNzt6uTR0uaG0uQj1iktRslc+6OHwc2mJQcZi/mhqT6T
GeENk2moGo4lSDf/rxdcmoMG00Mvr54hkzhm/O3ird7BbgLzxHqchjmLPqSyiZNa
F5Mjxaw1kDks8AwpFfpnrJ2+xCvuI/xsPohJaEwGjPCDN5V1X+L7rFtk8XQOi+dQ
q8d8XhhPirSChANPy85tnMjqMy0nVS3OJc+lrQzZaGSrdrSQ7It+MxMBa55i7ffm
vu8JwdwTeMNoq0eIwg/514yzC41K3v7zK/9KoOUTiF8Lx3XTDBZhGdoFCtEWPkCx
m6EPCo85b9lTJMDmry8iJ+Bf/1ILWy8/5OXda6uYqDg9SZo2u6OCZtWpCVKTSVJy
/bhaYnrDPPIFlNSsc/SiiMLOCq4Fh01GYbCp8KU98DaX/bxu/ten3bmYW/IMn2SB
xaLPxBUAUFK70Bra0XcfaHNGrgInKZfJx3V4yDK/RG503TwblGgajjiUuyox7D4l
Y4OOFUJHWMdGNS2FPYIGVTQYn3WpIebi4usBDwGy4quFtFeetSfaY2LB43isAsaN
QABpr9RlmsEqpeJ+H6DbbIAk6oVeeSj43HzBBp4VDaj5XT4TOqwcGxzxcXr64igN
gDyMr/jtYmdG4b9F1mNXhqgYsM0AL2Qxa3AgrdSsMeCoNq6DFLau95gLfF/8uRTK
POA3S78igpV7QMRH5SyisFGOvufuyvpwiqKEy+rSJI2ooIkbeCYsdmPvaFU4C5XY
aF2cg9ObwtgrwAzSDS3bV4nGgT4XDzRBtS9HNNAV44Ij5XHaDTZ59N43S7+671+Q
+WI0RdI+kjoQM03IGwkUamdbe37s+uuOZJt2ecNHrmUbzLyDLILsp+KWmK9gz96n
phk+qOTfVkS123xuyrZi71TLD6uFvRYvCO2usZgxBdc5S+0ncZPjNSAzhdhttukf
9xy/7LuxoQgl8jghBqful6T/ZnK0gsK53JoOclwgmxoU7TgFwJFSOjR8tjUOOeLl
JLUI4o1x23a4/sBqia6EdlnTxQxaFPv4iY8MuY8oaCx18CKP84WmwrmUutmNXv8f
BOs/xPW91trmLPJJRz4VJgKJYtrSjGS10iAQA46o9/wq5cUMUlGOVAJO7y0bTyAw
XaCPsPNH8bFWpx41Aj3IGIr6ptoCL1MO3Omo8JrfukA5nePnJwdVSrp5icbA9M3E
ysCOnJVbijbh94ImnMoPpfr1RAvvvMrnAz4sMHUUXCc2kq1NBuda39ADoYKCDVVj
qZKT0ECIr/30boEMshYIQkbwFblkraecIp5jG6V2tttVaoEEd/2zCOVaxYKX0ht0
BjBUxjD9m/hbBtqhSiuF5BcDWEM593pJG9afHGxqs94G6wZEKIcaDeXOEd1tpQBO
Ggk8ph58T8xjOgF5XDLFhMqy9WpgQCv6KUKgk5viOYYVSTEp39PE1up53TCs0BTb
E56ZR4y/5kmgdyYd0oKeYmLUUH+4W8SUODY6p94ejefp/X4+xKGHrDXPuRNfg/Wn
tyKoxVbaPhYqFnZCwL46wGQ3jJQWFqJgeyVaf8ZivaUaX/Hw76wOTkpWZWBHfudZ
UtMld/VVF9HTsycQcMILDUhSrlBDzpsau6CX2hCh/j7Hq7YLQ1h4RGWAtzWgDXqI
hoZPafGSxZ+zrVtF+tjq3AaKRB7JN6aABkYCzh2an0u86LVlq6EYdSC4wthDhlix
/YFXQY/Z9/XSLtIiyJmrvSgXAKuUabfl9HfAF7HQzX4pmyYzigGrA2QgZR8b0k0M
trlYtW5dmNyhneAofJfy0WoBf8fxQ11HzX+Wzh8Lq2oVioYTwBSlzrjpp4kESTiw
8bGWGdMeVtmNUiHukkFM88Ry+OAAh6u8V+Y/sIW32HxAKBgBkcE1YlQur9ndI3gO
chlmDDgugQw4+Qa+SkL5nhLZGVmz9CTLEw3xC9URtc0iiMv8uRr0C+URTiP50Dr4
/AQGgqcY22+QMa4MElKqkzB3KRVwXXbzJWMRJgejU7k2it/TBzMDtDzN6zN7aUEF
4Tt3SAqnbeJddXpyUVWkxFFPT8kMBRerfdzX/GZfBk6qXDfFQYuIVlZculXeMpvc
/2rlTuYmXQK+g8JAehxkC3YwuQ5XSS6R8ulgiGDsDHMqH5bT0WHpPTvIOl9xEkKE
5aXIeqlUroWlmAxgbBqTzO59Kdnn8nIS1cHjBp9nkMcG6AInbH4jTVYk8OVrconf
kYhtf8GOccT+AqvN++AzDXgS+NOTj1jRvq5o2AHQYyjDUMtDiD5kagQ0+Cv94p5e
dDj7c/Yu9A957pOmeFA6n11OUnq4l4i/Ju7EV7BK0ESg+VmZty8RGvJuEXe46KjF
at0hXbQIKGwL+GPUaF1jlfKZAIU1ynFWBtALkQzzrffg64qPgrm5kWXETmyIaVrt
VMsfS1F5jqx7QW2aIRnxDZ2Uz/duSM6EGe+3vkeqPVeW4gv8mZT+B+NSY8qYJZUj
d0X5Dbkq0Rwe2Q8FDoCMoQDD132tdvj1FUI92iyZr1ov+TGDSIepRjPKJkJuhpZS
1ynJAj4TIXGTyBNfRS1AqHWkAWMPFOZlp0PFZrJk/8U6/+PS091NNVbWtdUfzWJX
XNwS9tsbTB7/1LHXjtqRwQpBDLT9yf/YfjWj+Kpnl5q1Z7+MILbGBpvRF71kcyyI
In7VHmHUj6StYPnAWqZwgV2lW4LFt+W50CZLOW03nSVU/qLGothwoenIXBMAZ+jD
iItT61l4PfepsD4WK5fEhDsUijXY/h+7NxjFPNvQDTSzfmpK6UTR3JvRgPlcncrP
JKWS1YkfuiLsV86nceGc3ZXopvN9+tt7yfMPaNdsxprynfZ6YvuOO7lMSDHk0URY
ZcZ0KVGgvlNPS8nmXw1ZEKkgUaBRIe/Ix8kHELiLT7CObR33j+NRVuA3ctZOVnp1
2IZekX2y8f9i2ut3/gZn3X5dXD2IqJoCEiiqN9UDssi4RWsT3FkrlQdIeH3dCLSn
YMuCVpsLh1UqyKSqQAwbGB3eUuLQPzLmU/aXXp1N0Vv9bnhrVcFBW7IfVH7l3EqI
aiwCSJxGBw65spSnGd13sJkR1YOAWRc+OR+9eSVsuHzcPu1S8dSZV2b4nFy/sK5A
UXfQCfdhryB0hD5PABMRR3K6K/lDzpg5ZIZodivc/Ulytfyrt7vmrLCkBWEoIuJn
JYC1hGRB2/IaHgdULPap5LU92fDuTduwsMRddH9HB85f/tt9ROVkGsUWiECaKoK6
VskBalOg0uucGSQAAE4kKSbUP2qhVHnwOs6UmO3qaJt/VUsUuszdq+Fzs+wJqzSo
QZkzhez/1VIBXoIQC1KaIsKeOEHiFmdiE74Ltj/QTAWwAYiRMJBS5HWKr8pNbUVd
g/FZklnSpO0ocnoW57vPMV7D+eOFEYV8jYyK3erdF24XmyzE23UUDZzjJ98ItzGK
MROIekBxXtUZZf8o4H5aEYtICQGsO7PQbvJWAcrlErARFE+gNZb7tJQ25W/bZwQp
FOBfEdJiqS3++7VsQJTP7OUq4GIulKonR+WUXhxZjKmoUJvsX3+Bs1vHTm5zH2X1
OwkaT3SdOOEduAFtCjaFovVguSSQ7r9FEuCxG3DqvsQ46ovCdVB02zTPpMpTSPAg
ftgccxhoAZbv2FGj4HGGR6TPWG0shVsNTUXTZxpUYra3VAguhRV+Vkm8oWbeUN1/
iF42y8i3b7CuIleDZp3dOtXQfuHU5g7veeoB0aI0LYT8qIpaGkzX6IAksPdolzdN
d1laRNSGKbzk4KWm/xCF94esW4TaRQSl2kEUygIqLVQEwZxWykmwVIGyUMtkzXga
1vmmk7gacWfUN0uEXpRkj/eQ+zmzigdITq5CbiVjc7/zYOT/38qfmgZ3daRud522
s8H9nAppmVmCHiUYBXznCQAc6vQFIYreqsTRiaRBHgVAmwLIT8XR7aceyhiONgPm
NqUxtYobSYVPIQBqeTczEcgjwgNFqU18Py9aKdVejXIlF+DInM0XErsUL017LIzp
pnwxcxPVWEqnYSSGWv2ZHyazBwIMsXqx2E4GiasvMnL/V0kvJpImkqPsyH8TdHcZ
pO47RuWUF2ShcetJvJsZHkSY97uiiA884aCE5PN7T2wkUMBQZzXM9xjiXWOUtQ0c
Mpu/0vWJUa5KF4tgpXxn4tohZ6aTQKig5I2gi/3XrEe0F+ZZ19CzKs1oA26aLZYW
cY9KYgxVRmuclRm0kr/cxvik2MmmZJJwRwKyZeeWgiuNaDuFOMa0awHwAIu8mhhp
qzHRNVs6PE+fZ1NDtN1E4mepuu7ylbM/BPHUjCSfaLtD0GcN0keDCukjI/AwwRV3
Lfr2HkW/32VJnMXe8e9NEki8zl1Tlvgf9uBKKfJZgU4lgZCQ1n9xIHmqPJH9GlS1
z4cKrNNlD2gOp6my+biVy46V0Y2TILcpLxEzkr1Dta1Cj1sxzhD1k9X4jz7gI9mN
05t/f4MmJxlfkQ/QA3e0m79AvJL5QmfyrqXecAoptQeYMMZDq7z7fGREVlsKFVXS
L3ey2SkeAokWuTh35xzCdP57X+cTkUevbHFylHIjsaQn90hndHs5tmSYoTRDpJoX
Pbb05f1L4CdETQ/hs1S+PwrxDKlwcPLL+Q0NhsxbNV0gmrAHLIrxSih9Qw8pHoly
yOPe9IohMdznkXZX+9x1+QPINx0TZ0w+9fKuzhjYRdjZC3nkiiFbdFPlS4LMtYxs
NCO2PyLdZg7kJDJQ2HV9OgIi+c11txpHaFEQb6vLPEpZnMl+dh8y8ZQ49IVEQNxw
riE6ZkR5nvugrbq2cmdcuqRjSgVPVcCkssT/fF8CbJmoigP7V+IfbFvhHtwBRmis
ZQVIsfl5AKxiMKCgUpIJBqZedknnk/TgHY4jHW7xQuatDgKB845pUj7K0P6EwCGG
yyjcUU8lVbMSsEMsbwvO42h+LXwEY/PF+BIUajOxkgSFKnoh5bZ7eQuKr0Hn71ll
fYR5TqWG6pgxsCazEm5PF65/0X7RGDMqqyWR2d56UVyRZCoihel6DCF9ZXOZoU+e
oUSxli26tp/hpR3kiA/DoDBIh1l3XtiN0EcwCrAqtiKzKTCOG+ABXsSl0SGJx1d5
Ee1CqnBynIZhPYQSIhYtE/c855o//PKYua8TSR6jzEfh0/TkWNYiOkVODJLGc3q5
T6tmPlcH7lzYqSj1u2O/7wzgEGcvq3b9JKyD7xNlYBWXZ28ApW0C9vo/ZyQrGoLx
E7HQlFZ6sKG7knaPMyK+Augjv5Y1VzWFHpuK/rokkSIGcB4pPvDI5FNTJxleDi5+
Gy//ORM3ytPntjhMDxVPNJgzIsv5cA569yE8Nb28J1y++sWbNu1jeQWQdlV1QxY9
/so10zqHYeNVvguW8lwNx1HmKpiID1YW5NlBGdAh2rAe/ox1G5HXqHb21QMGfVEW
9Th5z3VmhuajLJGwl/f8MYQVti5MY5pL8c+NY76Lw5bJ4K5k6WM3ZVI8Jy/HQTnc
WrNx9zUsmvzdYWllpuMuXKSGalzVBOBPpD7p+9bww4PZLCntDH6/WwZKb7rND60L
qa5rR9DvmDc8S/Y0N5jnmBtoe5ZGAc0GhMMh4IFKBw894Z8CZE1CCxdZrIQBSriV
CFsx8YIqJ5nQIGZUk/elxEy0zRLGOym6Px1D90+SbcrDGD8ezSlByd5h1ZM6T7at
D04HmJFv3CXP0abcsbYyGFD8WIBQ0J64gnlJqCKLSuy68uON2JcEZhi04lHP/o1N
wcMCrE5Nvg8drOdsh/se/OMMaL7fyFL2B2K9k/MTh/CmIylvTeTO+BqQxcyHsOrd
VhxW3zj02wFokXMg2o1UO4P+qySWXmt2Bn72aA0BPimMrcme2UJwLmMYDlWf+Xob
9vlydOtZft534t7HS3BSowGgjKRn8OIIntOE1rWt/au0q1V9Ts5IGKoJ6FK6babs
aJaPZtLXcS1YHNPpVb4XQSExucfVuY9zg/0cquorLBkk0X5i+m0glUTAqZ7Y3sl6
5zxFx1sJnuwGuO5GX0htHBVZKgOoC42VIJla3CsNxawdjVuuOpNibuB1n4oYBVZT
VvcjlUXT5W5PCdJAz3paK4BWk4qyIhHQHAfqYZ05gb2HQtu/wBzxDVrZcSku3Wce
AkSXWVJWrC7MWYBh4LunpnP0M5crEuHdcAMTkfvOgeCzGkA/l96+mB5Dz9W7GM5A
0RFYYS1b9X8R8U9rlrMmPNfr0U3XQ1zoLUlrjixpEMNQkTl2MsxYv74mjbT7gnI0
CTlIV5Kz1xpR/Muj7JBcHXpi3r120HSTIVxW4vhZl5j38uxTHztV7mZjCJq59y9P
sGLdcq5Jai6jB8XhYs1ERfQ/n0bf7ZYdjeE1CjxVJhrE0ntBhwplt1UjCZ6Mr4Is
YHzmzb0e8nKRqAI/YAjq88v86M22GMTnU7gmz4iHor9n33asE8MhRkQrckVP6lHR
FE14Wm4W1BKTZlKp6nb10Nayk1Xq0+tA7Jji0+OPqgQbkcG1Jw03tCf//HYA8E+E
xlWDfUQ/5ObsUy7k+gZ0nM5WzISK/EbfOtdds8KEDrto4IdVJk0KL8mUrGz00Na7
fNoc+gqjUju0PoSz3r84wiRlhpz3mCup0CkGvZkcuEMAMqKWaiMzJMCumhvFLF4J
kQtqbCwiFFWPGGpzv9w2ErGADVug9pFeoD6KZduPr67O1HNz091OB4GrhZN5q+/A
OWdin62Rv6r179lR9uX836YawKnk4cqp1ZET81ZLQ7SOU9RMiHqZJJT0OaEXshn2
Y+D/6drYduw0mg+H4ifgF4Ia5hqjMWJUvf6HS2tBRYEeyCWEZbsrixK4GLFiOle4
wGi/KB56cDy1UJ8bpR8/OrdBmG4gwCGOczmFlCETldI62xSKa/jRZrfttlqe5sOL
pIjHShznOLpquUuoAAP1jwSj7xRfOvChTgI0ZPm4j1nMzHy3EFQGohJTVJ0c5xl1
YKMIH2lNEBkU934+6asZpK5Mqpfbhr5WMTyDYVI3sJMB25siKht+oOIfYSsKpRdi
Dp9fltta3T+LTe1M9zcqB32uRSxf5VQK8ECVT1my4yIjtl/IFUuxWzT8bhVW3PUF
nqIZtKf54AwFh43HbVJavCDAAUAvumBin02uQ2vRcJNtGsUJcEHuywM7n8eg4rs+
WgDZf0Vr03qRn4ZLwAjEgGNyKCvV/ABIQ+uDlFXoy19/i/chdpWA6ikXRzemmZtw
ejILIulLvFqaj5sVulPOUUbkL0zfaUnh4nhxp4wkEB5PNLeyrJRbi/mkW8T3+89I
cnmStbMCgJlsLocko3d8a8S5DicbI4CPEqiodBfJaKt5+Y1bHnubT862AaXkqj+B
IoPVeCl4IgWkUoPzDxpJIs4d4zBPSaibR3M5RiCr6Ni9KsG2AyqVhtYgRcPeIeHY
4sDFanix6+KY4/CjvEnmhVmeeuCvRm9eVeBkiiByDwNrgc77oyKyjPJD1kaI/bvc
FYeF2F1h+azaoMJONo7Y7y/N75ID2xa60AOJrrEV3MEyP0FA+38C50Dvif4WPCWs
9pYcoOHwP3OHVO08W7a3kqLEKgpuXpbLHnM/H46moskoVG5emlqzO+0Ty4AjX/Vg
v4BOUStx7E9qvegMOTwahqf5kjmrQ9A8GyXrcluuu9zMHewtooySlYcqdIwKBjZP
YIJSCmd+JYLq1HVFszVBNdNDb+WG2yL7PhQaXRFn8yxrrTlvcJkZeponv0/L21Fu
Daujs3DPqp8QylfaGKGYQWmeBidUA/7YwHTbVFPBJfgaePhvxgV7slo7rKIq77rU
FbwxTkQwTYsT5T9CbjMHuSw0nx0S2EVmPzeqrntiQysKEtauG+IPDkT7xX5L0hvT
zaUzyas4vr+bFlgSJk6iA42x3r/iBJI9UJyRu7mgl5c97XaT19aa6tq2RVNQraLW
tuj6pjRbf1OTnJidWRgKY6Q2wfboP808+fKrGdNRD1f94OVEnnCCPKxd/DLumBm1
3eYbPFGSZyZj/s1KdvsUVjkncJutH+oGYEWI+gb0mAKjDi/XCQFz/aduw9bTAipi
E6PiTCQw+0l4xIRDZauA+aE8wSrnIQ74r+0p2jGUiBHN/fsJnPkw2bq1d5YX0Qkw
pyZnlMcmfq9vOuyFVpBZqxKIV5QqWdhrrMQG9DdAKq5GGCJ/9JPadM7JGsl0JgSy
WohOlqDbKwtOMhP0+ueCe83vhi9yGwXPmyjdofbhBg4I1izIYj0i4u0u4ZGO5Jmf
W9Fy1IJkBVMU0+vghW+4/oKzqdK676xCYA3rv2JtteuV7zBeGy1wVmeCiq8abObO
Lq5xfFmojuz3lmSqAiBhnag7khDGEg4rpW+1dx5wK268kc8SMOt52hFQr4wHO/TP
prQ2yt5XUyV/evTrD/E1rpBNwBhHi++Wk13B0aeeEUpAoxw/Yi1PzEPcGZTb6UAR
lDHwwiPyCsn4oOcYH6j6ChYwFoMUtqmQT7YjG23Ka+vnh8wM1J2N+GgZsraU8A/c
+cBxv22Id1BA7UN9MTDoIe5NWgLMKr0EDwUFZdWOCrkbJ13K2+JiP0TDIXbBPBAn
z9x5+7DzVKm2wKj9gFAoepP3IyBbKNJTwa97biMRNHm+hIRjCNKCYpVGiRme0MQc
Tx/6ODi214VdKlEMzdquCJ2cvJYftIZDUEE8GjsspHvVpohhWJYOWYyZD5ZuyO1b
etrF10h+hfMqubVupkxWT1JLq/K/i9eVYCnY5/9tbuNrX05hUSincmJormY+KBSi
44m0jwWL0Sm7uYJoeANvozQ/KZRjOwv5q9/0CSkZ1qiSuIDeIFbKx1Utsl/Db7xh
VI8a5LZkZWXSKEYTty4yHb/fO68WDFaIG6dV/pPMZkY1HfiNK1iUmsHKYOzN02Yp
8EJbo/CRSLv7x9Oaj6t3Q2F6ww0LkX4rHDFPaQCFA/UG31cq4SGzbZaMce8wl1Cz
1vEv9fcaHzsiUmlT5iHeSABubBj7nF/12f5+D8/VtQPO7PTia1SY/+yNgw5hGoXD
78aRR4HfvvpTIQvfbO7XiXQdkAQV2HozEFxhvISibEmUltzBTKN6BjIOuUoRUuIj
H2eOb5CMgbqFod8wPumuFKSvEGtcs7ok3lyYLg72kVeKUkVDy8jJZssIl8+H82SD
KkyrK/WXLBupd+ITrIvuWqdh81D1Y64KI3eK4NO4pv8LyRafstQrtYpb+Xg4WVuV
GhXIX5wLBDLYI/Aw5x+JaLCJaxb9zrFo/C6EAeQSD7Pk0xaUIgIy082TJl8K7ipY
ua8RvTwaX1wprHwc7NXIupO/qm+K6Ea7WBAd49K0MPAlbl5OmSngC82b+jMCpTFd
BHv5stzihU4aNpn8V60E8JdbYa9sKJ3j3Y+cHE/0Vh1tBc8QvGNQrR/dIbU87DwO
+Mr7TGAuFghmfoOStRzcoxtiyoGBMCygVg/nl7Yq7zGXCm3amFLngGZoT9RlCC2L
XyX34Jh2t7q6mZIFSl0ylP6fI9b1uKR03oD75qjOCQoISlbREB9esu2vf3oO7vRT
XLtQVb+sw2CZu4brX8ds0Y6EMOybYBIIvxdbKx8LFKRXm9UJIBudZgjt89ItWDVm
TTVTsV/gMkEbeG/IpxN5jKNn75aetWNHu0fK3LGNbBss81p0jnqgAO9mkGYUqJwn
6T4zBHTmOpA3EwoM4KpcTV1l3w5CLZjtmcfvO/oohQj0gwEooX/aHVjfavdEj1t4
jjuq5gbFGJPhxppz6UEulwMsYcY5J21jfJkjv8lv50jMZ6gaxlRiBDSIh6jhlq40
1xpNgvKfnQ4MmoCUVHLhkIejka1V2kBoVW5H+dT0dBE+hk5NBh+kcTSbUMlWHoan
fFW3AO1tyg7sPPcZZ+pFsmDClPgECQ5laVamlCETKTqyz/xfskrKhhcjlcJFfam1
kXFmCDHXWAYz4rCQfBO8mGj1rzp5bSO7TcICV2F6fdfa/dzpER9FYPD8bo+jpIxa
zaCyzJ1mrVWERiFAweExnwDJNdwNvx1NiUpNxBSHSysgTsvtFh9roQ9mo0RGT+fK
oX6+vscwMDhKkOBR44Txk1YbcvUCzARiVtFPQb5fzbYw2bKQrvxBTuGrpOSRTUB3
XKnh+Jqg/h/edsxEm1EWKqaG41d6lQSTLzW8QnljvtNs0+Td3uRjT8QQ+7khHSUL
M44N2XvG4HF6ISHSA5DmNXMr7DBJXC19jRDjbIYghl4j2ym8xLsl7incRJjErOYn
Hskxrd8AiHl7djRVGpL+pwtEvIBBwN/tSmYZwhZbVuyKb/Ogl+yEj4GSaacgdPC2
OmjSSfhoL6XcZheA7phm5+7HNrHdzQyqT11uXCLiOqu0RVVAwDJHeQq3Sa1kHvno
ehtHkHlxdjCbk4p7b7Lqm4FNYEdiigMAflf/F4iFG8o4MOp0YXwJdKdjgQXaHK8O
uPQmdTQwIATZ8VI7Iw3r1mvjYJvdOaWnPFTOt+dIg473GHIaWYY9X/rcaa/F/jeK
Duplr2UPZrh8w4OCoLScxQpy60W8Q16CvalYixes6n5+mwDbCtXuI6llmo6bAVMj
BZqV08DhgSfVNVAtv7p9hAmkRgcS5yKE79ofnn1avjWe1I6bkyb+cxXcVpxbJ4/4
Bv/OMHKXs+ebI84riUlBsuiPWON40f01CMnbutnAmUR4oJUnW4eqHKz24EXmydtb
QGuXDN1QVSlbock6JGrIiwE0zdCbXY5/l00uqI2FkvTb3+rfyXXTbQtwV/oF1DVs
3tEYr8GICwbF/RYDTVMaZOkDPz7dDhvDubNQYZT0ttCG4Spg/26grCwjnvL19CTR
hoY8ZNbJxHrqr0ySELhWXGx/g05J5St/8e517hiuVyHSxWTVhesThDUFZ9g2lxPG
JRmIXSr3/wVJa2vC7ALsMs6ur6pg1DJ1u1EVVZuoI5uJY8x/TdBqYmeMujRhfxc/
xGmxDuOzVqYOm4R8cV3WJkcxU46NjddmQ3Bya+SX8bQqd0QY6Mn28RSs+YAtVOn0
O2lmhntvxsd8smf6MN9/YZnZy+RriQE1MKFBJViMN5PTvCoUZ/M9eJbqWI5fyfR7
VMJrYBopuLiOPhtDR0mYYksTV+PL9oURR1sVSqt69XeTZlDd/1hLsGs2rmNEoM9e
VGSLbcLvfW4pKvPLXUlTN6k2HK83dvdkhJ+AxJfiAO1OEr3TpsLbOKloCdTwlgdh
TXi2Of3iYZ6h2y9ALQSxIASFtR6IMoySs3dhU3fBYXe+mMl9ZN3nwvZyXpWHC5jj
Yo+t2GKzCexDNyJFggIktghAaOSot4x6ZtqMRVnZrifmMqQScfAG/GFaCePiIF3E
Cxosb9p0RIUaxjN/3xYJea7Txy9MlqgFl4zBIz7ZiIF96LbV8lCMD11u0joabcRQ
xTYZ7pVcG6hWeF5nkrduWZiD0NCWRqDOpUWWAka9/+Xe4udSg/RoojfUCfB+6+fT
Sk6RZkWlf46Z/eClyP3NfbZ7e24kR+N0er17qaABGQFpBwQuGU9Mcg8zWH8kAfeY
qHg30SDMZFUYEdEHs2FlMoWi5hrkYQaEzWU8H/4vfKLJ4moNkB07MztdzGFH+ooY
D7lEzgrQPicBrFq8cW/f0+W9ihz248TCByzOJDD1Ds6BGSG4Z4XVlC3D4h69VIFA
wDgc/e3vewk/QauTPp4Ndviw+dcUgNHtPyXa64A29GHMaRKSQtD09dKhdoQ0XYUW
KnxCm+IguciHH58IkTSYjr49pzQ3fb5TAs/KO3flIkFXd4ZTNTWovx7Px+3EsQyZ
acwPDW1BVGl1sn3E9ryR3dvElazZVyWzbyajJS4ZJjamTHAHvdnW53M8jfdRuPuO
Aum25NaAffSMS47vpexPaZ5siXCr5UQbpqcLSErngsBfN5i0Fs4HreonGaEb11jV
SvsXiHHAd5zOBlw/9rDvLGD0VKBc6ZCEkq92hz1C2/rB9bSCyGXYutDuySiObu6A
5/Xakafdhkn15kIbzAuWajReAxrwoGGuZiCuJchCIwvMssmmP43crfsOfo2+LRYo
x54fR8VYgCgR2DoQdpus5IIS2BKQSd215dh+aZtpX40YEikcsqMZBvDC9ZrKIJKK
vcaOO4+uGTP99AB6ul/Q3odDu9xvRW0zWGglK9JaJLPBazIIfIj56IwIgUe4jri7
ziSOD+Dexm/1W423BudethnjH9Oc7/oADu2NM7Zw+stceh9OWQOJPjPLYuRHFcPt
kf+0htFP3qBFkvzF3xTkzG5Rw2rKlklF3L+UTMbq9HQPJ/IxL0Wby501tQAeGG4c
MSR8hR+8DRabBN6quxbNQ9eZ57jGz27FYsFybEBL9ooNXHHkwMlCKGte63/F5TdB
NPQnrL/AWdFm9JTjbQhErcVJlqFGmx2OcAVsVn1v5euPEwFLAszX+PlAdwqKRBmM
C1o3/D60Ci27kZYAlGRsWZmILhCAB7gnQsW8jU9O2RAAKif/HE6qUhZFZwgP0Mbs
BRU+daKpdywd7SM7JVg4FchtZ5yQuKLh+b5YUHIjIXWttIJdyj8e+NXil/NPg/YA
97ikSQ9G+rlPfUB3NIrCcq3ckFfRy+rswvWIMAgkOBYy506IroLcGE4RbzseWGwT
ux3V4Bd+MBdAe9JVyerSjv6P6XAqFgvirrUTByd3YC+ZIbZck4n3xu42mkRhfPzL
3Hq5vrzcMOk/VHrgvrmAl2dRqDA4WqGQwNzLTLPya8OeaYXixdELYS269cjQjhI7
3fe8BeyVWVOEub0//P3P5Mi1XLQPa93Sz/LppXFV57dD7MOewm47GfAI+Y9jE06q
sERDqYAyHP3OHqnLLwhhOPN7stU2Zl9MCXmfeXOKBNYSVtw9c5qd6cgw+gdaegYj
uRm328w+uOuF2U8DjClxpTblCmaHx4XJeWk5lyk5CHzw799Y/P9vpq+7mcdIqj2l
t2dEdg/p+SwXSHdBTgjtdhySF3LidajQvkiHdM2c5J4ECMTKVRZ0j1FFBgDk9d2p
8q0Lhov/1X2ZQaibp5RfOLT9mqSk1pAkFyzxC4zz5NwRdn1NzHH2cJaaB4UXp7yo
xmRJ8zVM8g2QlM9b6sUWG7XOEseWr1JG+9lLHKb6tRglieiL3x5Dzf80bNsN4aY3
BjlceGtCLF7zJGQMOYpLEdtpO1GSOkG0QRqPDLKlNKqvMuoRDPEQkh+WLmii3dRq
kKi7C7tXSkxoj5/NCXHi0wG5b5aKLNsYH858w5PAT6mNG6s/w62fFeFWdIJNyQ/h
weE8HTHLfSIWxSUKrjrRB9/Q2wufOG3M6QBqrEQiaAqeisjwN5UmuxRjqxwlhfYz
0A/vublasKHPHKq0XIJCDnaW7Fent9khKImtA/PYe/mFC7ElIiMfTpeCE3nKzq1Z
92WaVvQl/mX0ErRRZEZbKv8z7kAqy5goMQD8viRbSWAzgCO3lCSlL0ryEvSW2tss
e814zGVr5P4gcvmqbqfjGMUjq4u2KZ3+sPFJEMgP/2jYXYwtFL0fOnVfgoJq2JMC
meW2gq46CIyL/0bY5aMxpNNLDNh427K/crRIDbxB/MBKoguBSynx+dXkW01GNjDd
bLjni+zonCYRZySsi6WzqjzMtyX7JfIa6EdYV7Vw9GY5p0sY1MmXrKMTlEX7LDLh
kTagfSkO9khKdu96q2vL1i33OCwnHb8flOL/h6BZl1xVdLF5NkGueiIr7yY62CH3
jEzT/TXKZKyxkAkxj8WzsH/LZWAgYBm4fpvmAP0M1IH6MucXIyu035QONMLVvSw4
rPGy4j/YG3YhIOmrqw5ICT8uYeCBaXyPLbsuggm+ZZUQPqBtJ8JvDaR9S5UEytBV
HadjK2lZMZRwpYhJT/woElNkPnW8R+Af9HxZSVAzEmnQ2uTQCBM3N3pkiVaok4gP
EGSzY8kt1FiyWWf8ghhvfBf3KeV6tNOd5m1r/VCajp/ci05QtsbI4KiXIn4vkao5
ZuXzSuMD44Ax/rRTk4/dVA3ahot5MuXpGdavwnsv/ZkgrwiMp7vcWc7qL1BYwW7c
JUma/AzwimP5dK93Xr9YEGqSquu60mx86LCUd4RUgNvK3jE5+d4yRj0nLn1dJ3Y6
x96O4JHb2hpxRrVtMrpZG6UrtEK/NI8cZORr1lzmBNGgRs6SC1Eu/yal/n879UFg
lIPkbyCfqETPfL/Hj33w4RgV4lHQM9rQm94NCf+lUayDD0DLI80Mj1IqhclhuTXQ
ENphSStxW6BzdYEI9OVxSTgzTWrcvSiSGnrVhI5m63SnqTGQsJnYKXgG7kTs3QhY
QWNVAryvSx3ta3eHtjPWDqGx3hhQ0tAKw/Yzj26683M0oJQoXMDExENtRCOESyN8
E0oCpsIV/b4ytkw0kLgVaMv/Vf/4dtRvhNdyPwSVHdpD8mQIudQsiAjSHK8OWbtk
7r0aX/CfcxUSlRAC9CDNkAFnuCwrggDFuzEmhIIGn9/oKKnnhke/zLXFFCaXQWUV
lGhdCKdEGGSxV3pgcn4tj6t4KO+fJCbEybemvBtCSgPqqHkb+VyVDSK2gka+/bBt
iPAXvOu5QSpbJ+a0zAw8/KTlBzcOsjkxKAI50XtGb/IbVQJv/LmWvD4zK/letDef
5vChBWbk+gRz6GZctTKkhh4sR18RJ1ZCgbQip0AS6K47s2np9uoixG4ikjUS8I3t
4vg8OXlSMq9XpOsChF87a2ZfJvtGxOpfcMXcFHJogitNtkuq4HmDCawATgjMiiOz
4KlX8N4mbkGgQmS5rSJBxIAkw2v7QH17OtvIlx34rjDUgKJUpnEA9BpVfI2MP9Yv
EvXwjA7+rLywiwKLIqBtjE6FLsvHI9PxN17vnMtN7y69c13BseT3atgomWCkaJm1
BFdallJPRHCc/UaPPd0+I5gQ1rPsB+1EQckfRiXiKQi6koiaYvDE/xE8ipdHTXaF
1QbyhNOdbLAMLvwKyyLLtVwfBn4V88ny6kzvcjjb4WuInRPO4SPBoo2xUB9Wm88V
0LvilsHXrrAj74ODMqIS8lmUJTyHuyfO0LhH3beod/ugDS9bXSXUq6cRrX495Soy
JGlp2R9WO8ASiiyGIb3YWRLlKYWukl2ebBCLBbpfSZracm0TNosrOZT9WbkShSic
gKFZK3cgxGaqBv7WnTCKnnE6oqRzpCdGD3UhBT6VLx35QmXK2rpxzAc7DvB8IPB5
+r/DXl7HtCgTK2O0MJO48VELaG+gQIDlnnPz11GHsAxnvu0BqPspD2x1LBE5UAlW
8ntIp71hp33pKwJrg8YzEtTOa0wRYSGHa2PhpoQ8WAqkbDcCGb29YF0q11wIX142
X5ZnLPzcdYaq8xleOl2HsUip2RIYPV2oI7CnL9LVNUSnqyIG/zKJkPea0lRM8sxN
/pRPEPCDGI3rog2QYL6jAmpnGO5BWs4THYlFWZpbbjFcScfRJB5Eskd/vbp2dJuz
berYUf/DumuS/5VrGkLysk0nJbVSS/xP5SgFWmdZkYwhyZbvqPSPFtd6O1t2FOfV
YnjLVBD2OCPwJDSlxuw7hZYwUwg4pNy/KnHVJOqidzj9EyHJT5iB7QOvB9BMKpG8
TXjYyZ6zjV2xNGvFQNd3Rzv/iOTcXc7WY7C4ZRjqQU0V0DpBZhFv02hPpxCLLMTs
AP9gDwDDfTet1BA4AE+UskTP0XyWzPqWAbFvIlydtRpA7oRRqO3UJH9GJagDDrik
uQDsIkTrCjdzCLOfiClSMjAUd3HjdPWHQkSpJX1S3SR1pCOkqX9kpez72zChPAkE
ukOHBJWxEJAkqliUKcnr7SE6kfrdMJnRUSE/sCokZLVNtfHIMX1DOp/tkXJ0dBTA
d0g17RHGby5x94A3doyPuXBn39cKfaAkT0YUWxKTC/qD8Dmf6oUir/ywJSX+MGNp
nWqff4bhej+zdmj5KbJyL01RtM5o9lRJBu4UGqSEVRFFJmqt5jVa3PGOwvNp5Wll
ugBO+g3RGCNxlRqSSl1hoxue4wTd3sTynb9oDX72JL4oP/+IIcMHI2nmGBjXNbHg
qhLs4LiTcoypfhtsUtdkuIbLMw3RUY6jkEdgnUSt3ZfN3bcNeJKeJFCEL/xYOe3u
kwXJMaVUoONW0lm1TF99V+p+hZhM8yszytboDYdrG4R8MqqENqY+fbMvCy6gjn+7
lkS3CCfZJlU0ZMSfz/xRUrXJi5F9+jlq9FTypUwOy6k4RI5oSsElttCB8QbQrViZ
gvF+Ak7O6UZ0hI1id6BQaAfK7N49XDlwYJfh4QwcwZ36oSWSA0buvM1OEwvaShQE
9V8iAih05R9QZhQC3e5QzSOpBNnAvUwiUe5gb3HbJNNfRO3lO0H8oAbqlbCo1zcv
+ShSel6ZUJ20/VrIR+4Kg6YHXIJizY9pG0yKEdHFtxisqxo56iWH8Cj8bPJOMeZg
NzD4etuHkbalWVMZOPUjKMBospH+5okJAVSUshJkLoahcEkYBwSBdoCZMXNpyZX0
0ykKE8joXB7LnChlzwYsPYh1iBN0UyKNOF0nSOfW3aLwtOWd1umSnln/R7fyLirN
fTluLa+m1VbuOl5MmuSX3M2wNjawmhZyfK71Jov+X1z9Ez9gP3n0MwmTtX6qiuPE
CehpYWVe1aNcWjagO3ZdBhRAxHqhtWFh2JdH6p5NtGGMcWyU88XGHYKIUoEm8Cp7
gROsd4Xy77QQJappHdAzD9dmqNifsm59HAAif11q1HiHNmB+WQnSXKbXWTwb0sKm
VAEKasQV83Olh1ajF28sKt8YHjvB9tlpYkmyzKmJn/1+6nCVSA4s4i90I2ZOy1tH
CElz4dJxXVjYRFWSC8o2JGb2414JVUZLfiXxTZon0HVcdHyLUW84SyO9iATQdvX+
0KZPKUcx+bOiqBoty57cjXT/T7iz8CaOucJRLKCoQWLBIzbAJs5vxCv2duBPHHRX
wqb5fRj1mwyDSIvV/5oaeRewl0eDnEIJnnxjQuRCXEJCign9fsBy34DgdJLTC3hJ
NVmDlRlTzSogJBonIbaQ/W+7CXdINckLKiostZ7Q5pkjfPeZEnbrhqHS6XTqiDI8
JyT87WDrmnzCTTaXC+m+BFgVjqRhgSnNM3UMklcDSOPMykb613e/E27Lx1cYRmqA
IjDFH1/KiqHa7QyJHgdmaZcPXm0mIVEnlzM8/Z3lwbU5fHhoQ3nRLDGGKhHqXhOX
XxbpauLkJf9sEHX4CUiTzwW3lECcJNHx2o310G1o8EcvIAZ0k6dAQFZbVcPHyIzk
STyU2VF/CuOVMi0GdvbcCf397n7WlUc9ih7AUWXFipubMTkOGI24XWjC/BhiFIR1
jMQpt6eUXhtCRhyr7PZHDHzwsGMzYR6m8jGoZvDQC++rz3uP2NVY4Gf14zESn2+9
cT+44Rii7D/CqOJ2xFfKwGui6tDbmStMotGugHswUamcIOXExKtlrbcnPTb3XBUg
5eQe8cmc8C8OJ8HBk5nnJ8lHE3QAvcNgF9hqwdELsIZd8ppy1qYsIXlUV7TtxDiO
/B3S14wE+22cPxUKuUl/HCmnTcX1XWAlZl/qXiYPmSarNbqUuGa7ZEfLmr4Agznh
wINzfgSSUwYSNXq2FZL7hLY/8OrOdGH6XIl/9daaKslUZ34hX/co9DCWgNZiKISq
dIz+eflbH+yS+H+4DqAriy/TM5PtT7jcjL+LA5bl/02BQu09Y21EOAj21v1xdZGU
Mndxh36f43ekEntOcHyrjq77523ZDbVZtgObc1o/8pSg8AI6FO8s3Mt+Ze/kjC+1
C6XYFteDQbPbm0xVUd/t79YbUuFw7nNqIDAECXvys5OHZCXwjvj4sjEGFml5Zpgs
1VeGb0y/KnKs+pKMwNJRs7UzwfYJOgjZYn5Qi1P1iG9ystk2fY/n8vH+qumnpQxJ
NDh6J9bP2jWlVoNZRODZVyU+btC4rNXdbf/dqIoGZPsVBPs6nfNFRAvfsb9GtgwI
kzAnEfQyt0XpnbNBzVlvavJ54x3Ykamsp9UY3r9DcARMin+ZzhpasC4XBSwCtEmb
JlUqrzNa6MMug6t2gPld1KQd9Xb9dEWa4Utbyx4BbzBkeY2uancPhScPUeh1PMHc
0Jeq2EhDEW0zoEWObaixABeo9nSWBQkn0FjRoYWYxcv8IJlnHc4qzTDU3wh07vhq
bQXd3wrQBX0dqULR7xrp3u1cX+xngMCid2Dt9PUjs2uA6budHQKTYT5P4K+eSlK2
EFtI2c5/598TA4JKtjylMUkhgnHfDetx3/cP35o8xbxEoKtMwJomrHzSbskoT4rD
a57oZvRjTzUHG0PjGj9EEQUk6bV5n6tWr5ADZY2wY3ylUNLAmhfetCMiWBdDui8x
xu+nkqe0XhTHg/CwPIioeDUaGGksxWnWY5SntMhioOZyDTufSryXjV2H1ZZddXYf
zzbofgML8O3t2nuT+XPTaGpRZUujY6JJ2+KAYYXXdk0vsgCPbtxdPR5YUTJkPZNR
/jUcjM+JhA5I+ASJsALyLP0tOfHVl1BjIbJ9zB7JKQkhlP9Kl+fFmYF3iuwEjGV5
2AoTCai/BXQTdkJl2HvzO1oao82422t4obeM4oQ/uHwAATBFEH7wkuCgTXfts/ZN
68mwLC4rcESbY4Wdd1UIeJky3OSZra9kCYNYLdGYAJpZvkoFCkPpB4B5z8KB47Pu
72ZgO7mstA+4gkYQadbfM6IWW1nP4c4sSaM9IJp3b5sQCELsZHJRKzwahDJpDBYJ
NubB5lu92n7qLv13EkWVBQDY2t+ioqAKgMH9DDoXVvKPLoiNlJ3R2AmtNob2cQKN
PDFFHdl4skHDo9NyALLgFnyMbUrBEuadfQuaqS7rd70KgrKsYATlnahgy1ksEh7S
E2b+Hnl3sc42gIwG4KISDaaP0FdKC7EY+PSBMzRfY/EP8stkO2FEGQDOyl4NGoJr
ZnueGQLJDwY6zYfW9/0gt+adrFuz1hwualKVwm3QifYQ/jEV1UJoWIMrhlx5CrOY
pJuiSlK4ajqV5HR84qsQ/zbdzrlNKzCEK4407yQK0wsJNxYiAR3tjK5mBdzF/pxp
ngOJa2sQZXHAbfbbS25/ATeNkzRIICs+HiH+Tq7+srWJW+YNF/eq2Xutjl8Z9rad
h1BuD+H0OVdfy7qBeNHA4PPS+J0b8P/VP0eZ1HjSSjBu0yX8d75ECFDGOLv6TehK
a7qs7B0DodQNSibFFs13Gg==
`pragma protect end_protected
