// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ela0qPJ+4pCAKns0tjkcuFQhTEDvFdrBM2dg8FkJbKVPqCA34qFRUPWDQePRrbpQ
4gTze32Vb9Hq5C84AtLjYd4LtAN8fcxWYFa1YBLP6gtBlixWCao+65QZzWhkDZeX
o+ohyh3WVRcjrNMI0jTXHINenmN7DIL2Brv2MGvgQmI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30656)
V4haM5gYcvzJ+PkQpB6OMg7+cLXsu0Z8aiSjf9jN4eN61dj5IMy0EdVxKz5PAY3v
MKWEZeEx4h0WHBjnCg9pEIvUiZNPTsMFBYHUVqSWo+uXrCtEKcErOzW21c+dZWYw
5ccKq1A3R1rFJbzWerM4t8SKjHh3hJGFJEE56szQj2Q7nVMyFWKR1NTT13WQUKiN
CXQ2QMoGxcR/SuYBj42D7V0/CrS6uBnA4Im8Qedqp8rWOJvNYe7B5iwm6IgkWDYq
zrW9L+chi6c4GZqMPt9guDiE0uWWMZ8VWxaBHl5chQnGzZKmXNeQ5T+5ngH+l7AM
UOmtGpFyvBpUe6n6vwkSgsEk2rAND1PMh2VGWYR7LH8CVYs3Ro8VVhalOtzgoc0v
oz1zhUlwmLVBSIgmnQcRLOJrfCETqge5PgL5qT5pPdDmnam6Ky4EF3BKyWytTK15
8BBDwbSg+UCJFsLSdo7oD1dbz05+82HbdFKhxxIv6Zmn2NQfDlwCk/FNJn8Fl2R2
Ws1sgj7hgMKMUxuD2wYtX6cvwPe3Lb7Cw54n6AW28aoCuljIz7GfdyHipPbIQtTw
isDkHmzATG7Vfjfc3FIzPPLZcd7VFDgnAlj1WwnM8W7/15jf+CLiJqCw7entexjw
7XIZwz3eG6rKpbbFfuurMG8GGwy6CChYr9tdowIUHAzEqObkaroPTqJI2gYlvPPB
ZGP4IKaFKMTf89Vi4Qm7ymywcEkSypMV8S5OpONkAksSwLjQt8OYKsnxNWBy4aXy
Pe+kiPyooW3smwKoSH5IHwOB2wNu5gYnGgRDCrY+4TrjmJKx2Z3X9qFF97/OTqG/
mQ3mhxfToePXIkbVbBpsz/5+zt3YeCdRB8pDlmGXUEkFex8cNIIzhe31PKTM/3gj
oyWb738SeEJlPpK5WEoUTwpPaykGNXuv7JTijxAronatIvi/fjw9Jvz+rLQiRnZX
F6zFticjZfR9FPykptiJDVWyvPm3K6qsZQynYbE4n7KIqhyCsy+C4mp0nRj+zXVf
AcLSpemh+jYHnnlu4/6r9t1awxplZwJpkC0hcjT+SWhpKk7+5MTBS52geYc/UZCi
kCrVAcxXafXndMvBE/heq7CZNOQuawqx2SyqGl59MDg4VN7zU2X9Nz7Q8/oVN2x+
ouJjGGsogi+kEXQuRnjOHky88CAJeH4Ls9B00iHNxQGvjSJTdwxOvofYk5uxPMyD
W9jyObv+dnd4ZEU0D938JvhSkdtKX6X6HkjSCX6+CHIibL1Zvr1XfOfBLWkzej4g
e0xV7UeF865IOVo7AlAWjfVE77OiRuFoy8s+Vp6mJ+h+HjQ1Sc62ojZWhOcI/uVS
npoCPrdcZhZSSpIIepP0VYbCEdn61+wzDs0QKrwguzvj7fryZfjOKYsS6yi8mf1U
TBYJ/kvi1R0Yyij3D4QqIcTAPKurzfCD18eZvXS/8D/Q8A5jjL5SchR+XNDhXVPQ
hcM7Ls8TSA0no+tLie3GYfrgpLBY2RfkQGXL1eAjFUhW/jLKayYW1wymapFv27GB
F+MXJTszPzsKLfQOkFTons4Y0UTgY168TcA5GdKmME1hRYTUuEVAUJRGluKz5TCc
bH3OUQHOh7iS6LZiSzBA9qdNfGZaRXdWc3IaA8ZHM6bmBfpdth2kM41gDekqrNZg
Cai5fUTg7f0fS4eRgWiaSxUeg3rlE6LhJ1wN66JK8DXYieZp1LjSxegnCWEIFneZ
5wEXiKz/RYT4WX4FjcNzWWOlSfq8bZt7ayODhY7q13/yAPzEkInLzr/z/tWujNBe
UA82XT0xKUHgBUcgGLIm1Fr/mWUIosdN245Zh/pvVK9J7ZjI6cjCvmZT+6BIwOHT
xxcy+jzN3WBoszkAZr3gzs/BXIwwNUmeh1FRyyRyr7DzQ94GEzv1gpnvbWfE6BAX
s7wYmTpn5E6y/wQlPjHrJWiit+XV6Xs6RzY8SY8D7HBT85AaNiiwE0HBgiex143+
DZM6GNtXVggzCEpWCG/oitO2rI6bqjC+F772bj5MllX83EzqifUUTjkHINol6BLs
0ZRa+qBVC51UM/KMSj9rjFzjVW3Gna5oK1FOQRj3b/7/PcdF5uN6ChYbI4dP2+3+
4Dzj3lrMzr2q9WHfSplnk8Lt1pzELRfitF/Hzn9velMbNrpa5sHvLgF++sChOrK2
ug4g9ngU4XXEsdST32RbU1HQN5ivKh+PCJw28tdFGjmFZ26ULQLhuj/842NFz6zc
tvNsAJ/WcKfvIeXbMtOwz6r1N8be8SxZOx9ae/GRbkHZrt9+O1rhYezhQIAaeBou
LNzisR2QXCS/M/Ml/XTD4a94J1IarN1MuXrZ5K01pf6YWMcqv4DoIDvB56u9N3Zk
7Xfey+iWMePYA//XIQhbB+ZsPsEBCDEm0eiSCeixVqwwyouEyybvhNRjrZ/H+J9m
kN7MBexm4ZvmaACC0qOKKndq1Su5XWLa/UiiB086u56R29vM46h7/u5Yt2j26U/M
/GkrArlOpBhas53MbQlxK0JZMA0gypX5TNMQMlJ2eplM5LASJ1DIsR827GFkhLKV
eRq5uAdA6AfCIgtYnlTI+HSMcuAurUCDXwea1M/zJ9MO4i+TevGrcp9fxfX/0Lje
BKZxuDP3KATZvSPaOJZ5QcjbT4KOeOF0IdVyjZvLhaNzAE3xz05zVAVZvK4td0eR
SMzi8Gji7xbFjOHeuMK8xEXQl1rJ1oi+2Pg657oqXaemClFazxBqsxOH+CFoq2nT
4nhsEvItkU35a+yfJp2UHy1Ra8THapgH2Ha5uEOIpP1iOlHuJg0oZAL8r9LYwWrY
PFEAflEtp4oScWuLEC7HZxUiLlGOuK8CRVFx6RbDzBNWQ3i3kKsWsZAjEDDAx8PI
dzDNiPaprUjWOGlenB8/xcubhHDlTqhMuSkjBFTrZwY8QwnEomU1XYWWoMznLDXG
wTMdh62UU8AroLgnCQFOlayjanIwlVEo2mUkQ/kyFSEpaULJhtQjtANx+tb8EPFi
UlpPqJ5amyRfGX5c7I5BWQUNszXcNrYpa6J+wok7u77g8gWdGCJBiAz75aPMTWNm
bA0OhsOBfDc1LV8ydWz93act9lwDso98ApEDL5vjvtxk1VLq/MMaOF04dGc3Lnog
mFXmhpWLlovIKLaYrHJoyyKl9hDXEPKGuvC/OjigXADMFEIs4PR5lf3REFrF52LU
hxRH80XwynjhIkndI6HVeUSXVtsJVo72Zvx1i5ruWNnZJ08Ps4d9vBnW3BptNJOK
tKFHWiJyNGhGnr4K17abNAKl5MPbATzySyJK+fhJhKIFTZV7ruV3xH6oGg/195Oc
CV6+lCh9ERrc+m7A/x/Q6TClE5aITm+nPMYK84o/e/cWHWpPZbkL3WexmJcjFsaZ
4x/wVh4Gm/cJgS0JRWN9FCiq5HCnbMDVVMZ0H6oZzPul3meQ2/MuJtoD2huKoZnS
X7uTq447vfo4E2pTEsAFQC15ASPs5bjvNqTISvLFslNYvbJvzROHzF9qD84eOIkJ
pXe7GqPV1VGS+uhcn6xr2gPJYPYS8dMqycSSM498Pkq/Kv7bYJWNd7A01YuADXuk
BkqjsCSEbyBhmWffBt4MWOw5iyZu9z6XhTRegyGPL+c+maquvCE/LH61B7AwY1yZ
FzczxMxcAr+F1vy2p1WISun2MpC1DAjHRXTYRlBujaBf5+TaK0NhmdUJYfJAbVPx
q63719mjgnz0Dx/HbXt8NsrDDyO4JfXGGwckQslL82QdMBZTa/iK9BVr4CFmE/+l
P0RuV+jsX8FeL62k96fVsuw8PNB05XqrWXPF3lpXy4Km7Jb8464awBhm8uyV3zU0
PYsa6tSeWqOeQOcZYFBUmywMw/8eIfdFD2Mek4nHS1VNQwmzUI0SjtPmCtyPD/G8
gpRAFjUCKdLx2aiA5pfeEM9NoXEB8OF1soE7BKhIYAXHJA/SdLxOES5vf+UduW/y
7HcjZVkteFca+o1nWNa408vWAMOEock4mvj2Hg4SqUh+wk1BWt+axZCIS1nfXlVb
i3kX2iXNke+Zg37putI5RlrRlgvekuRsQ1Q2G5xBjgtxeROosMppySBkxHU9RPUz
LnP70xAUu6Jbw8LDZ8QO47EKDwu95v03i/U91E4XFVz8qc2bu6OLnz+gL6CfGFmZ
/2AxWhT9RimvCmrd3U+wllu6CEwN9oUAt0skQQ1WLe20AD76bxYChY1aS0+XbFO3
GEay0qFgPQd3vFpSdTdDOvgda68LQT1suJt14NqaHHvfXJ5FoMCgYzMyDc6j9T/7
GFZTx1zJCqRJcwFW3+Fsnqhfj9fZ9+rE8Z3ROFNhEm+EGZHLEgzKEJjsG0kZhgYc
xc+lrEz2okDjdqbOhKSE1bRhvvFcnL2tUh+GlYXnYO99Xxvxeq4tJ/itu9Obd4vS
1JbMElfrXpGl2jV8z3rjCxiEpjyUNO97JCQsZzVJpO/6KYcYKjPmZq9JgOBiSOBr
DwS+1wzlmrrDLtFY0ah+LtPiWDi0Fx0wwMMbKVWP5tcV6mmLohbnPe3Q5thMPCDf
flwx4c8N/+Mp+fOyyqYvliRQw5hWbidSBMtvHINR7JKt+1vle67U/mKg+L0MhyQk
ITV+oGUiXxfyVnMhDRLESf1em3VWAHYQ+EgVwQJP7+2tVPTSdbxvRHP+9/52belm
qwlb6CASLLO10S6J4H8hBKhB8LZ+Z4H3EiqXO4ysLtAHol7rP43YRIvO6kpv96Pu
VntOmmIuBXgC30mTEV8OcXUUJk91sePEuZzSqNhUpKYupfxLDDIzXeTcf1zhshdp
KuB2SWmsqsrgrcqs/v++rM18R+v/5Bm9gxluiZwqsWXpm2KKNASEh+zvHrmRt6mz
WbtscixydWWVWmyiaumTYDhn0/HNo5j4TmVYyItrVGMby5eUG9IgdKnhYD83GeO3
d1teNmy1ogtgvEsMp7D/8RUucAQ9hwj2/d1diWh0r8Owf8Jgapjg8ClQjX4v1GKa
uHBdHEnxscdczv2+c6F2S4euz4Egl7c2A8V/spOkfJx9Yct7Cw9YNXh5Eet3eyhV
gq5eV8YeNQeVJ0lhDrVu02ipP+EykYPr958tbc6eKaqgF49eb7o/r1PkQAu7C0QR
XlI0o5KSB1S0sP2ioX5fCwqumQa+q9/MNs16j9Wf3z23tCAONUW/4tCKiPZfNWJu
ZQZPbD2FGkFqPgvYx8wyack02G18wB4QQcWklvKnHUOXWx6alx3MCVnoGxET3ofe
Fv+9tVKzD1WyimseeTdg2DtEKxerUVwrZX47BYBwSCpsiDO/9YlshCHbg0qYReee
WyfvdDwDTCCmOtOSbhQ3UpGoVS4hPo0OaZLZrs/KlG81KXmbwTRGPCiYrtP6n9QU
P5XKFXnBVmWbrDmdAICbm7J4P0baRHOC4ztEO/bSah0t1Sf11zGUZdW9T3L7+z6i
4z5j3bTGhOduT3X0jTVmNPfjOoBtlTihtcFm0wwUSSSjcvzBPTlUt9toMSE4+CSK
OyqV7dL5iNAlOj/5zSDVfrApj7Qr4t1PuqR0yPb98ewfFjhNapvdGPgUjeSEN/ws
Z4rjqNaTr5ItOkbDVTXkQBP/mO0DEFSXv4ucaVHj+0SbLmQdntV3zpUgUzgG4NaW
vLN3nQUFGTS1yUwQIFww+XmqPh8PxgHADFH1yqlpJzbo7ieww803IfrA9oUAwqdg
w7VOb9tYvsIFqSIAAlqIogBNVkd9TUO3acGH39rgRgqeAUMrbrJmtj98rLqqV6/f
FPLzK/VY7HRLhXUR1IibYlxaZotGyPkUxoNYlvxEfVr3i/Mg6vaKP7TeLviZKeHA
7xAKCZzFdQkPk8tQEFINKq86e4QKPixbbE40UOUNDJOt5jH6nbCScK5bDZ7vfnm0
k9uu5+1NERW/xc9pctnkyyiZ883eroYlymbROoWEWo3WUQa3+rEataa3vz+Fe6DT
qAsLKSKrONa9IoNVVLtcGlgBxWeDN7Hdm/oTXNTwBzYxDRVf+WsgT6P+gBxo57Fr
ykNALHlz+2UIKk9xk62eGTTY6q0o7dciS3QeyjHWi3s1pD1OysxIJ8/kYH1t5ON0
WDib3fx3zMorZgphl1V+uD4fusTz9AH4LN8/57xQos3jNrDNJJ/YzfaJvfG1KQMt
jnX6k+jvLVCXv0RIYKtbW1Q01StsYdyJY5cStgDdB0tC1T+4Pp/8BA5pQAaeKAyY
0BBXcuZV+5Vnd1NRiveEHPM1REcpA7SStl8ouFTL9brEJ6j5JR7AAj8HFngkQb9B
DDF+2HSx6XtRecleoWOvqmNHZn837X35dJFV6EX6kUqoiV9wo97yGlZBWEWSoHq9
5M9xVIkjj+o5bOIcSaKEqsLwl4BWnphHS7zQJP/0pUcIrnY1N408e7+Q+bywHhVp
ztRaZ8XTn5bQq6IlllbCIuZWgLHPVMAg3MtpAGNYwpk59aSePj3mPQ6xRpuKr/ku
ObEs5IKsOmddfYM/9jPwr1SNFiiOfgpix65pQAXXYMb/F8QVTkXG9DihS6yiYmeE
xv1NwT3zDxDMRiJq5/5T3gWYAxLqNz3vdPWKy5azKTGZxHKBSLjJqXMkGbrCjGOz
aaYYxyYqaWAbw9OGIp8PBOvzCiRNRG/j9CSZqQh92R01nHel9Nwoo/89dLEQXJGy
T2RvKHepErWIgyYFU/9wrlfiJarbbGWktYmqbd2GRJ2U7ll54EnpcSqF84MTvdKh
cEx/+RgrYbtJccmnSNcUeKOZl6fczwEtodiER1uUlU6CAtrBl0TZNwaLdJfF2Rvk
eIUtmjmcoL9BNaZ7paOOpse9M9OzWOPzDI2crcg3NcqJqkDVFYUzlPYTJYL++/Hw
r2jMPnQTfDoUiMjTe52oQ1OT2t4qwER5NXLja0LD6syAIwlkE+BVfaU1ditdt2KA
Xg7moYD5gTaMCJevdWEzhrk7pfM9BWfisE1nTISz0ntlZpP9FRLCyjyxwtuFqN/y
ni5KJOWPOPygur6QNrFMg6inJVrBthExPwqZtASxLlG7ET31OQbmvLHcTGf/SrWl
hhd8sRGUpAnMVwBgrVb8CrwOFvf3zTMf1vQeJ6KuOmn5RkXA8vmDY6jLLowGfjlV
QH3A6JAknH6LSX9BEtOQSAjKkdjX1DYu8YH2YKInyDuWWy5YxaZNAyXZ7u6V+cxy
Zv4LEi10uU+RWXi40hFGpg7W2BRpxGcfH9z5QYfDnLdyjIe5tnKaqDdc1d5QmI/7
HD17tlpUe1Yt19FdrB7WHCmFsZA6slheh+ulnuCKYCeecNNduBab2L0eFEssO36U
e+CbKmGrv3ezvJtETNA6SEU2A0f8WBIC8bRDCpbI3V5fQ6r34YHv62BxfwlhZQYm
FjR5cXm4xjweVjzAvr9pZP/2e8QUe49g8AqpjmP4zIPo3eytI6p6Yefn5ME9vixm
eovmBw7BkjIKey95KydTZbGCT3DT03nG/rFzLLwI89bWEBnHuOsgU/FRV1jpEgII
exdmZE50opTUuAjyvTC6l22NZ4IKE1sQkvt0D1Gmgx5ynl1bMoQAK+mNfRotv+kC
6fhPoeTAsV4eU3r79Ww+fV8/QbuPfBK4NbNmwdj+L/TCSsXxm9PskpVQIcjljWEB
Ywhx0EyctuJf1R8KxBgi7iXIuPqMqgTCxXe50Osje+6v5Dbpt3OjBw8C3WTpeTHv
MngXWJRuHBuCEjog70ksXpRBrc8zjgnIhH9VDk70xbLmT50jJtiUXCe4nJFr4hT/
ze8lzBWScc134xDcdKb7nPIyZtA8MC2XtaFensrmh/IPNe3NjeTOzxg4v1ccqEVG
/xsJOTFmS48fBD+Tj2/6UxE05FSjq/PlRI+7rcGnxyKFWvbuPmYZsdcLxCn+5uRC
JvDeywbJ5oE7Mox8sDeOmY9dsZlV5UNKqLVv03w9YT3yu3NdNWNFoU/LzdQBBStJ
4L04hyqLZG507ESnYhPU1DzHTNh3tQkz+50CwEWgJPh68N66+NnFIiCaVw7myoeT
89XJOCfR5J3XsVDioYqENWhj65Oq3n+pWx/Z1wRNdkXAlxPZuqRGaQvsbbpJTTqB
wLA+yXR4T2vVXcRvWC36l5SC+R8kDyEsJcLZrCDEHfxmUialTY4kHmWvLkisRQBO
RTghweKEIw57CCaIIq+cPPMtQPyBeKqJzf+4PGYXxp3+/8k+q6UaBfhmJAo8zOW5
BCCgDGJjTwzd4MWkDl5PYHDOw795N6zA4GdIOd52Hx2kxNQAhwaDh5R8eK6+ike1
/oa/5DoirJi+LapnBCnndJ9Xu+WPROCLRHpRiFVx/f9rBuzK2e0YPte3rRmymRUK
NObn71PdQ3tXTrZCeyjyAhFTi69bS92FBpWAitK26C2/2D89XbVdfAByl+WnWSIE
Sxpnjvk8gHWVGg1pV9U0Hu2oJxVe3qQQYn/aXrjjW8oqIVEx69LwwWjXQu5T91m2
BRLfujSpwb2q6bDdZTOyB4N862hGn3OWn9q3p9z6buPtxup6ihRFqBvCJltnJ0hm
TDOrHfOoSZDwUraVv5T3XNm+6oiSkxGwcdgaFcsQQd2Rg3t3ZmVgwvUab/tZuKv4
ZOmNbi5KfISSEr62abUEeK8MwSfbWmybviyZk+YeoDGN38xIQjhKZudyP3jdRhW9
x/vcnLH9h9Bzsh2TslCtSfPk3I39nzYfnIV+AWnOnDf9Wnt6sdaOzFuNV0iHn9Jp
UxgBdpC85kSsXXZcv5j8m65UrGEay9iQyDQgnUf2Qgv6EA9EOJqV18zyMR1V4lyN
L+EX302lnaMxuCj6nHzmoPnPlfk41w3/vuoDaKJl7DplbctNMdBnaytmVtnDms1O
txFUw77lWUpXfOxqENOjjEAuNUQwebBiuCU1J2CNwcx4Ey4uHGVPrYyZ4fUJD40G
6WRRa9VOzCmlwX4W8iI7cc0brUNg+iD6Wvm00dqvpvW7XnDDMZzsh9fB1Skf8Gc7
6HYby5gpHD+9i4vhRGmlIAJ3HN1j+YTpYzuJuZv6gyRw63Ozvg2S/g2V3SY+N6hZ
h7FH6ODImOSqw8rF7WsY9QHN0m50h24f1nnIuXc25iI22Dh/fUZMjND7P87KGGfl
MZKR0oKH8ITRoS4n/XwEfqUwODGtZQX3SzkvGzEoqBvrir1q0x6wwVuqSCbQ9lkI
Zs9XPn7ONi70zu/vQnAiEENQ8QN4p+WHOn9xuDundB82vduuWiz3z84Vw2/36uXN
QLWmXGozI0l0lP4ttNxEbWu4q9uLOdOxV5urul/dScXkQpvP9yyuMnPdW1OcctUj
SwPCkh2Vd0RcjSv0ewUVpAaaAPCFuDXbKphjzExugTf1azugvz305fWbufFsrJrH
yYXgsxKowz7sP4Is1BIfW9FNVFkMDiDVLTlpJoEbDX4w/7XOGWvfPGjFpLf9h11H
+WrEPMw3mOrobugM86QdCTBeYyT62DrDDzw7s1RhHxv1+oh9W84ZQq2mOBsI3vWV
gkWDX+O5nCOPumBUOsoLKz1Ng8zKei5J/RFG/GWKbw8pDTw+S9hs0rE4Vezjou9+
mfe5IKch9U/lbVnkQpKyQ0J4dY3UOn1OOddxERrha43jKzym9XIiwDahBhwGHVYw
N8rXvFcLAnpZLH+gYM7lkt0KqO/e5BjCCiKF1VRqQjReodAbGR2RdB1s8srODsXR
mrvvpXTsfh3q1HHu74TMyV71IPqicmWi+Yo+N+bKkozktyrBiYiUzjP1FwfBHYDZ
CdCLsUWR0wnL+elNZwY8VEXVQro9wXUB72F878J9wEDMuWw4jkqUnrnPQ7I7TgzM
KCGABxA1FNjqBaWcEJUVBwLXcF9uIAay6b6dDJ4OzIcLD7mIfC7KQwdcPyVRSq02
3cqR5YE0lVVAZ8fZXREWAlv2hpzGP+y4ftbsE2PLxlk6rPm7oYCfZUKRNNC1dtO+
PfP2bWdh8nC5PyjqPHrxKbmyTKHjR0dS64jQt/o8OLG758vgezD/oXsCHz5OiXxU
pMpy3UHMZLvp7ofASJJxk2ZwR+OxpdEn/gcQTYO9fHEN5G4m9L2F15rNVDCO3hmT
GHy1+sPCQLDj9gGWjWB7j6lPo5/RG7hrITExjhZ0ZLH4ndX4IuYW2tlXDU92k9oH
4gQLguc8oVUX13vGkk9dHJU1BC4b8ZDFqm9NHUl9mNCLO1MjBNYpsRwwY79p/2h7
GcizDL4Wvd3FYJc5bYaTZlXQrtcTWiqwFqo7I+EWry7V8hjsqIebvOaYkuAz+3Sq
4PL7KkHyn521A6ziLtezDnRgwX3QERNOKjWwfI+I1bAbAPahSPsqDGCLF/ZuJ3tb
Ta0oJSjOqSdNW8cldfEEhjIjZStsOEguHDZAPe/Rz0mfnYAoP9RBAuqmmIILRbce
F+TskrS6KF0B7FQCSB3SWTlgoXnJHXi6pnI6Aiqw1fw7qJ3VSCXL2UCUoI5bQ4ir
2wxoJnJfpNDct+rN/gO3IilxIfSDz6T9nouy3eAXapW7Q2vV6GEhWcpZV0UPy2PL
Nh661zhBOOG4xYmkkhm0I1K+4DZAHTx9HfTJoMkPqzWh1hwko2syIDPLs65/u1fQ
ZnWmp2lo/t5B6RllY//nYfH0IA8WBalXCUghCGSjO7W89Vz2pz6rcqFZEueO9fXp
GvJ/y0jCeBrusBggqPdkX1CiWLCh8oOx6eu8SX66MWW36sO/ssKJAWDJunkIk+hs
9sFyRrGYxOfL1AfODioY5yRmjwb5yYvAqg3HSzhWVeG3RNBw7U3zNnZrNNtS9Uix
1tPwMuNQxK7/DYXlNj8xewL2YwRe2CWZeT9wpM1y0eTZO+NwYAOxzMiULorgNqhY
9ScIBcM4H+2evLlqKmFkJUIPQpd4xwargfOHlzS83c03OnACaDbkHnbkKOLQsxGC
uhMlyuIb7mojLn9Ow3soIdpblB7rIWOxqQyI2JNccpz1ryL6H5t6zsnoIeTJBl3Z
V2NVil5hZS8uH2mr8QJYkO8ortqYQ1Hpt7UISKNAamX3LDOVB5voiyPGLHKYmVJe
V73NHvPhXoCWLFaTv9XKi9z/haqOXJbB5rN6yN4fqNBri4ztBjY4qvtiP91t02VP
iIV+/zcyqtKSGlz+7TumJnYhokuxajUO0aX8CIBDvwTDiICyW+HR/zbv7c1I8ObE
y0Dm22cvQMRU+7zexYUvFjl9s+JXztO0ZO6LekClq6fapZW6qx4a9a6PlU6rKxQd
TPby2dUCyvzN2Hrv4BvPiQaVcecqx2EwQQ2MaVFimI6cinNiuVN/BlTTxfDi2gV4
cPt6VlpzDZA2wtEW/LpiGz8a9msOFfUBcY3l4y/zJfYt6ASuyNosSueUqsQ52RNx
clPIcz/5Mwbxosi5OmdMXRPBGYugtavL4ZGCo74eU1+qdjDktUUPlYXDSs8sFMjH
XT6hdbQu0E00URfPjcpKnkSmmjMYK7VjGYRQvU6gBy15V43X2rl2uHBJULSn1zEu
4ftsXFuXlIvCUKzj46joMu/KIKmHc51tvgCr4/jbSGFe5R44Vdf0zyMKBdcNjiAg
r8i+Q9NiWMmIPlPiaz9z6HeXnoNJcLb2CSFtogml40Fs2UizmS/EOEHjfi3/6NVS
6Lk/D898bIVOP2iH5W3r0xINb+UoSuU0zW8zFIWIL9jmu7JxAIoi5gd2x+fYv78Y
tQVyn7XD2abOm2yzPhP8U5ALWCWZZcuoxr/y/NgJjUHw1hhOnILvHohXqKfGkar5
sJ2TMPSyNA0Fh2ztpG5sdEv7W6R2nB4UBcpZC7y4BwBbPqN0vQJWHdVnuWmWtKn/
2ySKkn5YKIlnQWSUQNn+8YlIANVh6k4OWiUOcMJPk+7OBgGczJ/N1Nc2Ur9s8h18
pdKRRx4iRq2CaLyC5qaYffvoKeHHgeNWJ6bWCaO2TwLTc57eee4iNYHXmlCzYnFR
kJPNtTeP2sRoSP0RVs4VP19x3YyOHWb5JJEb3KNyRhrkpLcD119XM4HWRdrMHIu1
F0ovnZDdrI5ZfNwSp9wOKLt8jxt9XCx3drLWHc7Jzyf9M6nqd3vEfFRN/UowGCMJ
xcScbWRGpYWC4LwhxvCXgbCJezyDCJtId9n2IQ90+c2ngz8x8XlX5gqgeQycZzfg
m/8TnUvhMGt3I2m37yKvBM4cfk/OkKFz9agHo1j0qEAUUkCOA1kRGS4MhtaBMKCc
hZ/JXt9psWAnUq8jVXCpQIEJrLzBz9k6hHqJEyUUUKI7qk0/Afof9nbhPvETfARy
NcD8LOErJDVtn3SUSvJ+Fy1is5nj8D1KTkXMbHwPvBa1cIQx/QQItnURbAKh5c4x
41vzNcXhBXeGxhj4BeHFmgWzUsNvF2aUWuNpO3Q49PbqXgjzpiv5my1spEXGBvmJ
6CACoRrJyQncAbcRYexfyHuA4T2iyTNFz5ev0Jf4rcnUquO38dhLBZFV/cAH4/af
2g+FqjlRbL3Hx41oFnZGNYLT+bqFse7KbzdOylwnbiKz3bX6K1I/7FIzJMEBME9L
8KfW6NVWqGP32o+rpNXfLUpXbpBUs+SJo863kuruvRKPOHNofLslFl2aRhNdhAjN
Bzcy9vEO8InN8692jg/96MxrLA8ZChEd8gQbF7lx/h3XdvjABnYLFMAMkFz9UDS2
Ry+ebKProsGJsQPUeBISlewy7MokIZOdkQevdi9S8pCJjWojgrb0YuN+wKTWz8+I
bz+3zdSM4yAwAJU/b0nJV/pf6ity/c/067hEuXV3kZvTERuHk42YAcX7b4WACCdt
xozTe0FTKT92jSIFzWFfpivoGNk3wsUB/UeyDs95N6dZ9FN7Opraa+996KCls8pf
0S0QUHSkzBQd8QOWwb1rAW6JRNftN2jMm37+lQHp5edf8hIO9mgPeQirYATpGtCY
yDVO62trw+1JGqvoRcfCjxljRuopu2eIfFCInNM63cBfNcIe3UJFdqlwPs4xuL1o
/TmkfGD4MzwYF6zdHbYhA9X810/HofaozzoNGK9Ppms/X6tjoEy9zZ/AFPxATCBe
9T+opcagCuWXmV09Q8RdtH3JkgjiV3V1GreFgAraPveoH48Wo9BNGEOfeZSGH9xY
N5eJP5sCEl0jthJ76qs6JcQr8drYD6wMgDuXNv7Q7LqI63RehAGNTIb8Czpq6UiJ
XjWtYA97sbd2CX7pglOe9AzJ0Qhosj0iN6cVtGVD6M4Wm3r5iywkUWL7HTXxOsk1
aNPhN+iuIVkFdS/eXyCmibFdQNDS98cpNzgNmAyd/vlEgHtcxwgs7RWAp6j0rVhe
GbbYXuw5ALTNPfTHURCrrv1qiPK+shULKtvmNbmP4GRaVc3TAVMqWmbwcHcN54A+
0wDUhOez8ck539r9CsKjwVRzzZneAlsygNlz4iueKFt7V4gFZ2ysgIwXWgN0jbtq
ECGx1tBDaHof4IHxdcOvTEq05jgQA2UjkMfsfzPNT226XtPnrqNpYkHiXyTYV8km
TXXZ5FcmuDWg8kdz7ibgbkL4BlzWJESxHDm2D8UpReTfP/buApkYpEPdyEgvvyJO
kxIE+4mFW2kPqHfZAVLro1psEl1F/hUORL5HGSlqMToC/5W/2BsOzQqvmpYi4hjA
z9zw3L7Pvdz9sDuZLE3BOI0x9Tx489qu7fCs0VK/pUA1eVFPN7/QG2vsQ+qpbDj2
yGwsyJNe78g0KrjV9g5Q/n6SxEbuc0Xo5L9e26tfz3qGv0t1aTo5ywdZJogXti2B
OCm2hmZkZSqDRwEUFmlRBntqpDbAvfCK5kdyCjrYLI0Ydk0xOfGPiP5mfsMjFAWX
KlVBknN41dRQaneJd2CcMCNkmIKnahihoJ35r+f06J6s9vpstAta/L5u4rtC+8bB
Z11L8p5oCLVb9/sWazZ5s+F6gQ/lV/r6cRLbtjWCXhVfhDWNw5heuGPydzHtuuI/
DRgPSewADClnNXEDKFb1V3Qc11nZQZzEGnJXXB43+DaClvB2LEMqSU6d6a/rHY+w
l3+GoC7xgFDwJ3FCgJNmUB8J7rgFuf7Jv/1w7NgdTCPPnSuAaCABcM7rJrWkFLNn
OZXLofKig4z8FHp2GsaluumYqDV/JVKDyVM/VvD8ERAYkw1JbPbtHZ0/ja6sdsxJ
OtO43DNq4aUEg0ZWBEEFKIrud7IOUagXnKUPEJjZV7S/bgPbCarZHfnRv+liGJ5a
lY+njB3iDWmREIeAucl9QRGxysgFwnCSNv6cWym/rOtnAJRbd0tHqbk6iqMsw40I
hLbTHxYh1u+gLRDEM9wOKqF51VTP9QYSDWAzfkXDDAjVJf4t8pUZpQe3grJ3CQmM
uTZXYIGSB5JyQi1WDRbY9r5H9tf+UJa1t/gqusyelHhb+oh/Uhah77dOduMdKUBH
AC02faMs7qW4rw2uuLKbPbhuS3bEgx1awTEwrK2ZYtk2Mn4F8kObL5gWIdLWD2A/
eDY6w4Kaibc3YfJBw1QUCJN6Mgii9o/8+e+lDDmXN3QOLK2G6S1jzb0WRCiJrVek
02kSWEYTL/hhLnNz52EvxMsr/XpBVDCT2QKeqc2brGCpJv/I10nAg+I7FkS0Ljn1
zh8y+JTLBq9ud1wE/UlERFjSUHorjlSy/gje8+4KTBU5x7PAo1ervjHSXp7C4XHH
XzV8O6YwFiIu2oTQPyYnfL++lCFEEk+vaonZGS5twSaAaSkZlkfYU/fScOrIEPWJ
jB9rCJaNJXLfd4OGdqLp42vBPeEN7jfsMzNIMOeWvq8tnlwvlUJ4SIED9KaWUdn/
8Sxuy1s5Qulbb8Sor01Ondl8quGNJZq/H1tQ+3j4E3ND4d3fjalRAb0qJ1cAv73u
syG+6JJHJvezkKE4izjG67Fc/INVtGedz/C3nWvlh9xjwMdNun7T7YdmHPcOEVyD
m+xOrA8mPWxuQYFVu0EiNhvZ7yS+JqMfQ4801/kaywq/CbUN391PQiB0cNDM6efm
r/lfFM3zw5RTbn21XS2z6rnYMNqaJPLXgM2TsFYGsVEm6+nKumGeKiVUDtQgUziU
QKMBDC5gOV1SEwSm8DY77QhZR+Z2fcHtdYBGG8ZVO2F76bKStU6zNzY8ueJxVEsI
z0o0bkt0RA2uaWl2+Hi2ZtQFbkY5zkBafcuVTGpIsvRotj0GYE9yuNbdm2rb2dtU
FWsM+zOyuPjiflqudHPxMzVfXfBZ2BGALrZ4GaPIqt7GNHiTbij3WpkQXV9kUfrc
Xmgf3Aaix4TN9ewQkjj3gAfksahAcEmNmlZy2wTZcHzz1ZUJ/C64OuSAcQlcJ/ZC
TYyUVrKmg82v2CL0o2eaErzF4DjQfMxobs5a2hl/zPxDDzpv3S07+6m+kk5vXJ4h
Iu1hka24WGT+C8JZSr+rV5bqUL2BnecB43pDgNer0ML0LkF+yVOkIPAtO4chHSto
LQvUI9EJdtIG6Ug4JKVB5IewclKO2tWBlXpa9JegJcQkM/bmwnW67YjGczwz6aLv
u98uIpBK0ZAT0rsUZmrhysltPiBcbH58BUDi8HT3tfRKG3qo+KvJ5eHoNXjx0e7+
pKgff0ekwpnr/cqAGx8+I05wIogASvymxnrJFG0ZlNI8xaZHhPxryIdOkDjvT90g
/CS6EBMagl2xii/irwZt7oTdQwwXLp7Xg88IE4UmVsQBizLxzz3DsORR8YrVECzx
u6Ep42FLG6itc4NAIowNZ0wVlYm7d6aJE36efIXCgBBfUiY0dn6IAdhkeOHvTQJk
6ZtSoJpNnt4cPfl+oTHXmujmiaPIJDbK7KcLgu+xBxv74expih/w5SRhd99IhvTj
nik/F6kxp4N8JPHjBDSwWARQu3jIu8vbNxPBaONBEF+cSPadf7J+pJ6e323z1j7d
kKFTjFehdowylhtWrTG8a5rjHSP8AHva+Rew6BtTJhjvQEP3a7b/pzpGWBoA1mU/
LCn13WF+CBRW/xuIb0AmxWnzmTyi04EWNp7h4Tk7bEsXjG07QtQj3WLWQh78l5tJ
8Xl61b0zjKvUOBmSvk7qS7vxK2MVAPCjTJz7qhL8JZBQhKHIb8yHU/oj2bFeC6Uf
fw3Ffu5Yluxcn21rSkHsb9U8xIFgurSl/GdHEKgjfDXOy16HkYPlZ/LbRD86RejR
4IWsDtzvF2pB5F0gSQ6ZzOkRzsmB1ckT0WKdVCP/1CCAbqSRKGe4AoW/3O9opaCp
lUJVpI1YjdSAsufXiOKaAaa0Dmc/mm4AV/naPz1zeiubtQPV7kfAqeJVVZxl4bKd
WqeqIrW+h2q3FO+b1CzO3TWbSmMmQyMblM6K/OtN0jD4pRJHZDlANud3b2lNGcj1
/xiUgMXjawzQ48F+zw+6OL0ef5n+o5RyH/gNtO+IIjs4SH5oGwGmQU5snesneF0x
d1Mk7PnVNUO5bZuTLBjgYQI5GLpg+5oFMBhSB1xkOZblvulWiYhdqAiBCwwxou95
X72to3oH5/idORP3499C0Hx/2JH7O24c3UbnqRhh5Fqroz4y0spgrFVYaWwVD0/F
kiJ5tRuixYHwBEE9tPdt/2+9515LIg/i7GvA2Y72DqbWAKpW8u1jZeqkogUd9my1
bUd2DLEQaQvlLuOSr5pndJKsEgvdq6GOJ9r55GLNKl3IrdGzdHmagdLNlBkdqkjv
6SIhtdiopCt9rEqUWcRRU8zEW4+8h7L7q4M2ZQhkuwj64DK39kqfh2KU71jTg6vN
3QGIz6pBnL07eMHK8ev8z5FpmS/KAdzhsdkik3a4qeQcAvXmXaKxwEsTC2cVzc4C
u+EpIb2+TbbwDAcbq7CJnxJgIBxBzuDzuVo8WVFfFaEQJU73liJqi8THW8bZz49G
lgnyDY9+nMDY06b76SsHnSD989l7EsIZVfSb2+JE83E1ashZE3ak+Lg0R9J8KbAA
64d+Lp616a8dr6xrybYzb55qnD3Dx0HJcfbAh475F2doLic/ogi/PE2cUDYhZ0qJ
4knemtuMv11JnXVq4E3nOeWPxN7ILopEodyBjpfZ6rJIFQ55R4XRtYDRCe5XE5mD
LXUH0gfe+l/z6Ib/Pu6f9HPQ6pQIM/57rE6SV/ofzMQABQmei1mG4r+e8TtBk9lZ
ZBJ6eShCgvvrY6Ei8/jEs3L23NvcyAPGnqK/5NYX/XWY9msqEhIYX8NyRptI32v3
xguavA5/q/9FeCqztmfk7XGx/I1Z+O4jUNVy3tzrkY+BFlDrG8SaBVVALeabuex2
okXY3QeUmN/GLnE+ocPXNTZO//U0PNF1L53aw99WkOO0jYGz1F/KCzMy/KhVbNWN
7ualAsuGK/5OXTWPMqrCQ0k0e9ytLtw7m3M3+no1fP0tWJ4UucpaqY6SaxOEh/I3
iwul3eP9nfEPOAcfEeg2h4xgCPaGL7JqylbgBuuUwQVV5cOvwTslAPyFsXPl9lwl
hf/ajWRX0ov9Qctq+01VeVBtAWaoYH9/P+8L92IXUilDfrMnoHmXBUY7nEi/2lTw
jnbOWdhqb3zV+9+lr6sSxdzoaLPgl6ypdlwoMHgHk9/2QZyK/ARDc9m5b0qU5Of4
lHrgI8t+47fUIvFZgG6cwC07scBVvifyEB9phTFOEoJRb/9pGulSFN/HB0Y5NIAH
8SdpICx/8hbOzyy2M0Ap2XqG2LtJQKndF4GHNKXd74oEEOCSsz43daP935bfZdVa
HVokhXBdu8gLNCxwTcP1oY+T6eGeUV5gSfG2uoEo4YbgBibvdXDVeWnX2hlNnyxx
wXIVRw8wi52DFrsJNaUTS/f1tj6r+bJ7NnDqWDl16zmcSfurMbd8UK+KsxayAml5
AieUZMJvyYxpkt6F1jKV2c4xkMhJyOpZTzEbbYwJwKlhVJRtnx+u2bYulBmu2zNu
uU4IaYEu1tn3gdNJKqUMQ7XF6Oj9Tej/+gszg/N97Q08NbCQ4ZcXe/NG2v3XXoaK
bUuidpIGxUy1gCLbUxRh1VBS4CBU+kfboDvc1YsChvWCMa/zuwV2jwbbPTkRYke4
GyQiNlwI/VqYCisVMpL6+a+9DFeQKNaZuLJNTqfE/Mgb3iwiR3y9B26efgwzV+Hd
GUb7xxAU26N1IVbqwrV72NskDsLowVGeVkpj+UPboe8Ltcl1SrT9MBwaOTd4aQUO
ErymokgcerWvatkbWyruQQw94s+Ej8nHnsT9mH6RvWbB5Cj+jEiTqSck96k51ydC
vuZPdyxbO4JQjjsu8sJ9XbhMnfBFOXhnwZ0Tc8fas9++es/OuGqOvlnMPpynCFyq
BmC73nv/7S0HMpIfAyyYA6qoIqbQCxwvvBdq9VaRApD5Ypo2wYliMSWfsQhSOFIv
shE9As7nSOodOtU1gWOyoY406VVhGtdTW/nw8OIpoLjy1L4CQ4Udku0d3WR0nvdy
BDhcFPjLhxAxyRctirEV/bScHNVJKW/dlxGa1pxXgt4UkQhh8FVhQ9fOFs4ycgMN
j1YJBQKhZ7hHdDBUXynzYqlN5HGrrKlHaQW6X7INu4LdzjaH5WILeaY9L/ia/4xj
GfS3HbD75QAH/FYPluH9uBlsgSrvNO57HVqtpPobuTQDZ4fF/j5S513wRV2cN2Hk
HE/sOrdzbIb9qC7BKBQPV9AyQKafmvF8vkpOV9+JWmI4EvZd1SwTKHfJLUZGY3j1
OwjKrLTo7+mbkKDsjIqJ8R9mnlRTIj5BiW7REhcvRYMw8xgFDuyCzS9tj5oameBe
TaLwc6frSfwx5ryXARuQDSFRcnYn2r3pR3JPaozGCuHUo1fDlPx86e9Hg7lAFb5k
nkuNx4yXDSs9o/dC8BObOKlSR/obc4crMoCoT14VAbyrV2D0l312Rxou+Hf/mMwg
8SU+G0ZprxzdCBr1sUOhCvipSxJsC43GcqIXVa/LyJxKCH5Ndbxo0ulM1l2B55FN
Kbs/+04kSk1Z2pn/59Rlk31GYDQux4yedxvWJERQwZf/7sZq5JX0jmdvfcjXDvC0
X1h9ZmPlp81Yy/2qIXmw21nzCIaSE9iYmT9q2CB1txDv7YdY7lh94KhNQGmAos65
IlcRaRaQVzL2AAA/Rk/CIxdVu3GVgIiUQJuI5UDpGyBfjW47OteANpOjUsWtr8fL
ALbGGJlhxdN+IfrNcUx8rL64crUrV9t82CxIviinHNIARGgjMZgjJi8wkxfZ5IIt
CY3ct3vU/LpqRVqCAUkXUKe6BqFfCdbDvT8Qm7v+yBGYS+AM0MK5zJDFSNjmuSnB
biUbJlwDMtwoqlsRjlA/hw4feTagX5jF4o4iNu1gC7TMAuP5Le2w5Woqhc5GavBj
DcGV61q1D6z//MMzrFXDp/L+iag51gnGuSGjaFPVg+WnKSlytha3LPBg/4eEBpR5
WbZY+s/Ykho4BuoKGFMWqAa6vGU9uxraWUfxc0VzzswCd2nMMNx0Zmi1pmGHNite
1wMWVSkarmoINglMqFEc3pfHErzMyI/fHZXzYmesJ4de0fXt8jLsez6SppfUe8n8
vXbQtBsf2sf2OSFN0LeyTvkKVqZCjwxCO6vUCKvBox8MgtywZ+aIjfsp+xyPpYEU
ZDbib1PMkFE4HWFs1sgf8Gn4QTNKDv9/u/2SzTCHOeJdZiwFkjwLl3x/1F2O+rmo
L8owgdvAj7oWs/ZfJN79wXGfMbj8Ibj7uM16KcgcljU3OowanOqlGbELGfDOtjQg
haR+Oe4QqUXX12bQOQ/u3v/fWaplHjfxLDqc4L7i9eKv3B8oslRWyyOLOrBkMMnX
lgfY2S5ZShs7DrtVCVSaViNxiX68xPUyehrcjbxv90NUTdkSlF+1yFq+nj8YxQNH
/e+ptS4ECNADq57dVmmRKDqs00tBlsBT+AbSc9ACE9Sw+7cfOQ5oLDIKUd+VWs0A
JW6WhepF5gEKVl0j/VdPgVLXAmT91wigSvMMbbpYtfNxgt52UBT1W/3T2JM5U+Ye
WP4PP9Iag+Ov1Lb1COfLjEcvgxA6EzVVw9M+Nms5F9G7m77CsYxk869d/sPVTutB
hbTMm5LHmYkNXJkB+1aC2JBLDVxhgrbiDxlfvoDkEcNY3wjWB+eugQMSZl1f7yTM
od3MSWLoWHhPVj8gawpojjouGlMmZ4stZiTi50J8XefXT+JuEpVTr74wr9MFxH1g
8EY2aXCA44qhApIvIcQPLLhWyeTh5WSPvosFwPY5cbTaLeUdFJyewKsLk1heKfgs
ldV6hejC7OG+gv7plMSrlhI4zjqkRH4cthP4hrViEer9t9TyrezGmWt9rQRKaVu9
I3LzKUogrAvgnBRaNST30AKuOZVSQMxcgE4o+RihtbJcbQiZfK10J1faXDwVFYOH
kQjHF+kGqnrLeryX8/kDjL3HrJI+AuRTW6OCF8lcrE9JxZkV7XGNviVmyq51SZ8C
Pn5wEWQvTBU2D1PUKwK1UUh8iYm/RNMVJQ8N/bkVVCP1roZj42OHXOCW1DynnFi4
yeLLbYdILGydf/VMZXCAjPA/tHywLlRFXT65x15obZtuTmm+4QXxgG+4BLqazKmE
3e9X7zRrZtezjYaukxK+SlhFFOjnaWIHxh8lGWLOd0+kQwWbtl+QaPii2DhCePV5
aZ05E0V3oRZvsW4s46srnBqPJmWMeiXsyD3p+s/g66orgaLjCiVGglLdRB14HTIt
IRXx3FMPzW09mn5l7Khy95L7yNP13cSF03D+e5eJvOQhRFbrEEs60kkwgviUNWt5
4GS2oG0ZUpynoGCN8IdJfOyVvGsed9vE+3mpspGQ+zC0CZeClKd2HJuvNucjQhYl
Pebe6zKqM3QQajrHXeWp6FT7+3v3/rvQk7IZf+AlfXi2exAZmvc6iGpVdclxTI85
U8XbVJwo2bywdhHn3T3NLkURZ6kP9RAvPOmdSi3AVauo8Tcq+WlRCU6NPpjBct0U
yLhmBP/FgLm1orqW80yKp4s1vyTLM5ooLHhHgZ4FTdTyKPx6SvtRKAxU2y/A+kM4
b3l22KJOnD+kvWubTYVZELHnq5lPX7w4kSSdOqBkwMFankwcYRYg1hVSo4BHUVXz
+BX8MdcNdm6iNyVGaAVQ0NjgAh3sz4Bg3mfDAV7TVfBTLlB4uJ4NRmFTpyagKHh6
HcKw1oBJF6FIU2BsuGk/L3Ph5t1JjlrkgOb1l4DaqaXKghNkkjy40R9dDgvH7pNp
rnuOSR8MsPQMxOvPUe5jcnp6Xv08Cf3zgmdcXCzlRI3nKSs5BIwwqSO0L2XwZ865
M1lbebXf984nZmtkYM/fT0YMVLStIPeoFCpvCUzUPKmOWDIWwu1JyZAGrBwXNOU1
Uz7meBDyu25uVUrjcv9o38WO/MjFTs2uk6YUu8UDPAITl2EwCeTObfEzAZsx9H1D
YDDcdDXMRWwXgOcgs3fuYSEegtAxbwC77nJdrBHvcAVGEVJvHcqw9JjB3I4JcCVK
WRFsgx6Dug/hSIV2f9KUtTq0vEnwJgecS2eQBRuMdYnf8/O4B9z0R5/kvczpmKV6
49FAvs1DaDsM+PpngwvGTXhOfooWM5tSZTVpiKfSqA+lKEY3m73U9h214ojMOLOM
Ci76wPVmdCaIYnqUjD9s0wF7XDjfvV1V3zrF7sIvTrHVY24tokIjY/6q4xpGfbAW
Pgl/6f+8bV5WukQzrlTzexf8qrXgeZ2KKbVyg1OVhu3+8p+RdGCGJhHXfycZI+qE
4tf3RNCNPUJg3J3wR/pkRHjCLktDrWsCHhESS8gd4DDtcxjW1ZvYCaRwHtHfXKX7
Yz4o6/iccp9VDP+9U7DA2mbOOcMn7yruO/qcVjIIBgp7g55NaV8cG5f3ovMEMhyQ
0lsN0+27RVQ63ST1JAWHdEWc9wKifAkFoeq9+bGvb0XPEHblJB30wDDcHl+obO7Y
orP/WH9mNl+FZQ3KGjCtkmgcXYrqzAiwOu3fElZGTc8FVby6faHSI4oS1ZP5I7Fe
6n+zbNonzOjbf1vqNlCZBuJeJzni9S2ONCnd3EBRiLLbb3OYkluqctrQY9Njcjio
w8btTib5N/BwghpE7aDBOp1x4u1tEm9ZtwtOj6vXt6EeX9EHjmFOh4XcUxw0XQBF
JR8gJA63ASw7gRedYSWd7sAgXvgiogVOOn7xQ8H0BT27gEizohyCaK+olvauiiA2
F7EU+4hQPN5rnuY06h1N5Iu31n5xCjDmaoWclwyShWEaTR+zHjaiLOdh19FzQu0g
Nmt1x1/HOsCk1O63mVmlGUedT0nWTjncdlGtVxYVY8dOYQY2ZdBAQyN2rZVfrvVy
XAq3ZW0Sp03OXwlhR0gWr1f/7Upt97CjAu63eHCSTwvaUBuq2OO9+rTZ7Ih/ipq7
Dy66DYq7TiVndCnsKQQLZZzYWtohpAtnXBT38ARYc4qdj8wn7o3x5Z9Ty0G7SSS7
rV4mJDEEXw1n01/gcKOCoFlwS6dOcAhL4u8vXZXGzrWFRsu+VARTaFxceJKbVcbb
wWXQ3//Zkp6+acadOiohXPIrwI8eec27+fgliPAAVZoeTj99SlTPfDcDMzba8Zh6
bRlMIK+esIuDCgvrV7wbhgKrxwWdmot2Km1IHkZDeqV0xcubt0zRvvR6k3dPquaD
vrnzbNbYRFGcOS45FZ94XU81IQAJPOcZviOscjU8+AyEl91dSeiBe8fAPVaXac20
cHaQKuR/L/ozOZfFmDbtcyPHzGUssvxvncBRLpzaHnbvVRQrhNSGKWbBFr+PyfmA
k1qr+t1fHW9/w8U7++TX3Wk/9ECyXc6K/P/21RIR5m+DOOZDhNDEvzUmd66iUwZy
WO+gk7U3EnPJd+ANRbIfpvdqfAGnrqhJTWlIQv6iWUDpJ70Mp+9v6xywSypf6Rrg
zk7aJbyalcY/iceaO9Gy8bWkX21+EjCrenGSaifhhZ5j43CDus6GTO2r/7IeXe6V
+qlO9wZV2P20nd+A9Utn6Iet5KwlTpO+6akkwMbHz6QigwXFbTzDVrkdZtYs6uJs
DqHSpsRuCqFhWEW01xiT8WHMsj2HTX6vuwKw6KYkJatZLmxdC+9OfaJr06vxGJo4
YIT9yZvFy5SEsJ7q/vOQxcddVZhVUTGfBba5xKmafmhK43/0iJKVSJQUjwaI60DY
7/ZYARHhB/Ke3dzv6En+4tf7XyeWVw12AK8ofqUfSdimyc5Lt80H0OnCOgS7XzLP
pCxutJuexbE5fnA1pK4x2JwrWDazZILqXjl9vDQktnhTdV+ftBPGfYK+jpRp5dB9
gWWt5R42AsE606hedob0j3WOxPmmiaTRx5QoMptaLmSTF9bl5+To7JYoQK61mCtR
k3c/51TVFzhjOCMf8METzQ7nYCqvdBIuKemJTXgJMo43Rhwzr6XMCIpFdH2wFJJz
7vPCAzW6XKYLzkoqujXAzZzP/O9XUIVi5xJX3cg8uQi4rOjG5z4fNvffOB5DiRWw
H4Q/GN7t+0lXlF4BzKBCduE930rhdxoi3Jveh5HHvPlHfvPz2zdP/nIp0OMplgkB
G3+foanF1ZWtf/tySh22sNCfDXSDbGlvQqtz7jR+VABF5Bs4bqjeGOvmAuHzki6K
pkhyDncpBydlLFLz5icA8+Ox5dgQWOjQPn2p8N0yhBF0ilPCeyV49V8n2Yrk5XuP
M4VRPV7igRO06zFrbfrUPqTnRRmfTZZga1jAzTIgLrAtHhEPr7oHvYzTKyxIyI2z
bsCeG348qmyzJkBUPc+YeVAqWLMveaS6CL29HxfpnM+Q/ZhRkSBwbqK5HiTCiL5O
o8maR06MdzSNNGkxrwuaAMmOFIVZldOILTRCwANWzscICdHcfA0toN3chA1SeiQa
QfaLzQZcLAOQAI8sPIYKR/AiTjgM2UVtqvRgTu5j/drT5PDbwZ4vNLYjWANMmZwW
ulJCG0ptHaGQUKSd7XWh+5b1+jtT6PuV8W2lUPYdKns87m/tMFRPIQOkuJqRlg+3
szdu+wj/8ea37jZibsGBZORo7P8vCucupdZ2UqP15kp7k7tPKKYHa5u2R+ie0Zx9
EFhW6j1zCkdN+XRvxK0dgvWaatZW9fI2hVK/faQCPjIseznUCixLOyoUiuFGUZ58
Z93qZr+fHv5mRj0mBcBr9CUH3JQMXsTUDecwlwVSvIOsOaFG41y0KK56xOBr6BsF
5lXtUIiFIODg0INRQ+Hs4DXBNwSfZQAjvwSkWBRWtD162/DeFNolEvXUAUGgkwZj
GTpIrjk95H8gkAJTv+ALcUmGYE6iYhzcsgaOxVsk1cUYkTkXy5rzQrUfTSQ2KxOm
yUcu2P1bsNfqdBmFEZVfOfQOFAIZ8IVQMpPfuTQth9ItfCl0W0s49Ao+yPTuYqe/
HuBVLus1zzgneMQqew5zq0G6aVJ1jGVzrZPEZzsQIvC/igIQ6PfCbUn/y8Z4sUvh
xlxZHeKCnAi/uhm3mVfdBMhyv5ALcbNYxIj6c2pcqV4PrzfS55ZCc2Byw04ssMNi
uT+TROfplvkV8UNdPeQKNA3EmQutTNTi+IJFCNpLSj3Sogbkp9Jp4siJeHnDxIeN
+N96hP/ENOxrMDwh79XB/k3hbFoTMhugU64PQiNShGsHT2JaGuyadi+gnCkybgka
jzFqSwgBsD3Ooe2V0bHs2BFS2MCwD65PmwUrsO81iq8mkZVoDWbCBW8KSd1Q03dt
cUY8niWbgbxrRQJ+jY4jCLSrMo9hw7WeTgReHT5sD1g7fbs6vNUuZiZ5Gg2Ay97n
vC8utM1drpegha/3olL8GllfP5ersmU72BndlAuYFUtxHpsf86tdovK+Pwehg0D4
CKTqtdfTGb90wD0WGjWtRE9dGl3jfgZHSZvURDzhHclWGy7Qsbd99DQQ3j3iNEuw
17t/0SkcfG400/8PiyoUqb12bcRjM6u5bQNvI1VzRjAqZvVeJIVjQbkafgL+Bjot
GERA0CSFP+dbBhbgzkMJ6kcIOwCyDQ3O13vvE3yaXOW9AZ3IG/TY3u26WnWM4Jc+
APO2yHe8i4gLCorNIJ7lSN13VPbuv1AyAn/ZuGh1Tg6ibAUpJwAAGRRceazWkIZV
seL5b4VUchBNJTQxemoaK68rxzQUX3P0ocqOUt5ji7Hy/DpdcLa7LPx9YQjcTQPM
+kG/EmIoCZowTnLOUTXLEC7/TfhJaMG/xiUnIvKDpUVIznoyONasJ32m0MHFbRTj
0SDXcmijPextNGxTBvP08U24DbJMMphKy333xms5q3+8eAyDsPbrPOb7LtSktwY3
iwnIBfahaAFpL3BopkycM4/u0ts7rZdpS3gbgtii4oGDOD7DP5yfo9WlMCCvwkxl
dvjdMX1q4b2XK8E7bTo2zoN/xrgquIU8rG+OTjOrbK5iiL4jgsNEQMXVUkxS1aYA
l7fhgDzg1kfm0SCf0S1Rf1hy2Mt4Eg/1uV4y2YSjcV0Fgt4819fIrkfarfrBZQnM
BWtA8CCmdz3M+OOckBRU6uGWYmsULpiq+rIrQYjrHrJ3vCsHclhIM7tSTaIus19q
3PWS0I1M86elMDfjAheQauqps9aem/rvSVpZ/s7fjODDTMCCAX7F8ajyoEtsHQa4
WtxeSsueMUeH1j8cYtouui+wQ9hNWRt9cCeJ80Fyza69VD5OwpiLMLipeXGQ9/P7
whA0I7VP7gk1yTDmPvIlfOhmFdjyAnWMSIN4fwwJN/5T/Sy+QQnL+0MiGBcVIsUr
pIWxBVokwSDKBK02Ij4u8+7C7tx7j96ZAw1O53GIDXG/M7SM3hXW5Jo+WF87vE/3
S2+6Wg59jk4+lEDHZI46twFgSgSbDOwv6V3LVYO+GBRb975Sv9oJUo65VUfevFni
pa7TGB+d8c9djy9jLKhSPqN11oUOjQVOzMMh6VYZo94b+Twm+KZYuHzOphmrF9g8
S9WYCkEgt/Yb99y10pHxLid+CIH9DTOv/cT4+YALwpTz1mpyOwlORIoJkkQGfzQj
XIXxJfHyNo6uihMJVVHm3hZUrMdCpk91zpP6jCPQdzOIik0dqAmM6RblVXIfqJsV
6yenBgkIBRlab6dEwdR9GZaliT7Gz5OzXG4dHg9ZkBEkIYiuf9lPxd4FgGEdLfhy
oaK4z++JHndMh5FghBYh2vwHnYL942bHoDg4t757AAQOsxi9vub+XQtHZb23/0vV
gSmePlc/kli7iEUtngYhTDkPnZEN21GVXQ9SrYDgEm8EAUVoKhMRKweIMww0AHvS
AGc4mjMaYrfeypnjpJX9w1WgczO9czr6wtEtgciDkQCINp7GTpn4gm6eM5yjlZ80
ZYKpXWBygFzHu75gBDBLCnfDfN8cF8E5f/Nryntdhqm9uBj9ff/WwnFqO+Qx9WnX
x15MKhXBi9geFfflW0ABaih9VnN1dLQxLWSJApqOpE9I2xZJFxFd/TWIJ2n0QqPM
g6o+SVHkVE0thM+rUC9gW4GcYMAVeFVUKPOz/uKpZ/PYkDZH4KFqomS9ML/3+Mnt
znDHWhqHjLBoj5UpPYLZjzwPL37JKuRlHkD9EIBbnKPG3ToyA7whmXwBnHc9YDQu
7TcBW2FoXI2993h6f+0Tl9l2Ig3ZrsO/pOidk/fG8llCQueBix/v/7zCZw8ZFt2L
2+6i0296pYSsLIZjOhjhmndS2gMyP2Jmh2Ol1Mqvr4euIAiWDGosT9LLUwvyu2dr
OfjUaSAyCL97YqX7l61ogiMYWuoTWP6yvS9u+lTu7L6cF/AyGbMiTySAgDJGNoJI
q50tw3lklTLWV3Lc0uPbazBqXhiDLTWRDo98iy6hErjR1hXEwThG5sx0ECL8ddvC
3SW24FXtV+A2npWoOxFBEhO1lTipGwlrRQ2WEWHdMDo8Sgk+70EPpzKQoZzev5SR
zhJmAtMF87TfmA4EaByJoFsaoy22p/yTVyABgiIOJLwHjGsBqkq7vTmqFj9McRV7
6xs30ao2LnahuVpkEfuNtzqMHa+0IAK/JSDzCENymEriFPQlkEficKzbzrlRsxxQ
zbEEoAKPEmyA310QVYSu9WGnEhCY6rudJq3PZV3s33o0uHuVI/4SDrcYsGFGeHk8
A7kEvXjEVqXVFlCcar60fmd5SKEoHdFbsembN5YBwXdIdNjhBtTTvXWXGnF5pepA
eZ63oODUKQ/90QearpoA8r5aYbbselzH25O9tJ8UDJbb7Td7nrVQuOOQxO2AxxYK
SXNH6jozTtlWYfFQRBEcWtl3vBnSoweNQeSqaXx5ehuYKtcE+CdzU22KRhsLi9x9
w+VkqVDjVI+CaExTvsKfbtP6zfa3h6k4zPjwHpuO2E1un2xP6GjFb11h59I8eKSt
DTWOeUlveHxzrKrcIY0ZN8cqLP2bBs4JLZ6oXspXh7hyEJYYban1dDClLL2lvcnm
THJjSLwfBYvYylT2Dst5iJCoYhtfb2ZgDhZ0rzsvgp6shMFyOywYUr8RRqGa8xt/
Ajhl4t7lCxhif+nzW8Ntm8f3A5FrIHDB1Q0DN/21OvoEW0TRWRDknNbKQcrsYEDP
wi9AyiCi84Sn95hSt82iqKRmYmzmDZvCSwk7JsgEFVYU4jzC3qxjHiY3vAs/Zx22
GCj2zBWRRDYsyaIcDD+arFyCzke1J0vLU5bxBnEfYIKNi8N1nkJ3Q1knXJfdTlZg
3SPYzI+qBGRlAQsQXpqvFikFxP2CQ/P5Vi1ArkTUNXlz2sXpD2BMT9PsPOzfDava
//74wvsQEtcdlPVmAA9CADuS01ttuJ/jKe92L6NuIYo82eTpERu0vXtKB5uOc7EZ
HKNX5ZVcpLJ99lpjVm6cisNwnw/ihw9Od0xku+Y1/0/UiQz7Ey4fMS2bbgrnVCj+
e8hQdxJpPF6BFeR75FV+umUl0D0Sotw8/aQ7FFwS1izLOWTI3cH8dknBHdN6z5Ah
8VC+ykhu1A48X/UzRm2wVOmjMz+KoecjqMYxdCrFpzhHQ4bMlmAih3CMpv3vbk7D
+yobNPcERUBKB39HM04wv1gAqfW8XOy9xf/krm/FnIUd/SXmVnS2Oe6H9JlWj/od
NfM2N8QtvkEIp/BDrOjfXUksytUm0Nn5JIuQkgLD0CNEf4ywRdQo0yc7Xh6T0lZr
airfopjrjhLZKJzv8Rnfa+7+oRAcAha9V96QNAFfS601mSXR0DFQ6Fz320zR71Yu
z2BuOXxuH9wKa0dgbyfwN8IxqGyXrtnF6myzYe2I27Nr827p6mm6+wtJQWYCTmlp
7c2b9CGhn14z471cDCDLlecYg3k4qYEoJX3U3+4MqAdTcLymVzCmuytFogV5eqp+
JzR7GkKDn79+1xpge08QcylrIeFesLNOOECLeSlmNHK9mn/IYOkCBKHC1V05VUZw
R2GS4yDjjaWT8j1kbg7L/izUF9Ysfdwag0gxUUpChtJ7BuZGQ6Z8/6PM5wpf7Xm2
HacDk/ha1cvDLSXv8bMLJ8Av+8i9ZQL0qEtGw4nzEsp6ftUIWWJJYfmihQP2ZLo6
XqIgmBoJghGpVhoPMa5Tm0ZspO/OKO20utEcsuMqfAQuHDP/yE2zhCRORul14uQm
X0wY7t5qqOyoXODWgMV12QBiKAlTxbebMSBnpvVnKCsIwdtW9i/gDBFShFNcFxgZ
qDkFkCWR62w4EP6Jp7frRUYvucbttS4YaTbahMfFBUZGpgwQmfgaPAuw0FJgJcIl
4Uy7uZqoT5VzLjVGGOV8X2hAlwsgI9EWHymiPoqGqQvYMW+X4vJpb3lcm4+zSYWb
r3eiwblnuQSQjX9YLCf+isfQqmTEpUvFxS4fWi4mxp7u/YOqpaUr9Lu6yFybEPY+
PxiDWXS7V/0YwDKRtsT/v8QJ2x9YmZOY47PdpVVZvNyM1YkY728Dzc0p402kB4qr
xp24+0b3Dz8Ijd4HOzfNiVYLwU8kB/cUA/ajNv6c5g/hk/tRIZ3IxJwp7IrsDaZW
xeZz2kSVOxV+r1iTuY/NSnbbi3j+Nx77YbHCUKfiOKeOwdpaJQIp01K8WRcNRyZh
qXyTgm/VzYyuNxnSPEoxscvRW/uQoymHaM2ujR6ORrkQzgRvY4XWenAn8aDFe2co
YtcXSsPPfIDQ/NQk+/QabYaOpUtWH3RUBxfR2tnhMaF7BXv4Pzt7lSvbRRh88q03
tWauy5vH6Q1N+7L7dE5fGz7QUqY3fndfNjQ6uu1ZhTajcu1lfkm2q0/Jf9jDkA57
Kg5y2cv2w4tdB80a4zOYtQsYuYOI0J+93tjQ5sKO1RJ+gPFRe71DKcppRfRjzcQ+
ff1yd9kWp7XMt6K3j/i00BxGgCpnRKI9T7Tmb8X5M1pFsCAj9F6rAc96qNPPv2r4
+Y1wpG4Fxf6THpiYh+W1vxALn21N4UY0OFfF8id66KTCEBvMrtrfAA1JWf8+Nu9i
8QAy7pPduFUQyqdqIUHSxUWhRM+enbdErv2KkcIrf+W0E2qvMz8zx79ZNkDthpb9
UF7dz7FKJkFBGTNsYCihtYPMlaJdk10dU3By7dt41khqYj+YT0yHEF+l3AKyT5EX
lqwlXjhHki5iMLYomxIseUg8BczUJfbCU/TsHwGKQKMiqlBek82OlmdW8tA0X+Al
JQFpc0jYUtjECrwC3VM54mg563pGluxxUXt69mzZWMmS07Dla8EEmG6qCWyiYVt/
IWtDzOXgDkuoDkqGzq71Z2yLlTotlaT2DNXmjKzZk/pv+ldcxV+dtYkccsPw7jDg
YoaKhcHFWRhDonZTLR4K4zz9nqi9PvjaR1JBLDcEZiS9FzSH7YbdevJ6OFX3kWmn
s8utaao1uj8Ty4kJFNlLRFphd8g/6Pykxusr0u1xuQ66Rn2uXfXqCVtyGJScSUF6
PEBq4h2dGjoTPOq/vH1xDfxstQKGFzUUktgdQjSvo16L4migll47gCwTsMpx8zjM
RGLXWoDGGvDxIvlyfYSaUAV4dxzJNo4fSetujCo/fnoTxLfGadZ4oUeiMwqASt3+
PE/RbiN2+ICpmKYQdNVrS2AiMBphnrQQ3u+RQMlxHckmsaa+ElUURyEfJLgi6Gbm
q3tZ3Or8M0QMtkboWVzKW0vCxSzYjznpofJYTl43iiZ0yEVTTLLiAojc9eVbOMV5
TwXsK7apghgmA961SSVHxETGdoUp+EzCVveMDUuGsPeAX3u58ZATHdXeyI6BNVkm
LXxmEu3v+JkuNWQeiRhKbTnwtsRD4Azx00Gq21FQzdRr6tkle0DxmwJ0j+6SQ1Au
OErUTZEDzarGwCW9utHOWmhm16gRFYekp+triSkqbjxO4BF1Dwv77XwY5QXPT2Xc
xetJw8EJArB+0tI3ET0nEGmJZ13YVDBwjofd7Su6zOO8weH8WY62O1OzwqvAqiwL
pOjhVU+cCIROxIHL1eMUPTHNK8ejQSa4djqQ0M5u5Nz0E42WgQNCr6Sc81pY4cC6
rdDkmMu6wC55jk6UfVsdSoPEdfIHCh7B/SGmWmMExd1yYVLrvjSFTw3tQwUMwIDm
Xcge1nY79wCrH9iVOzS01O7sxWGvFdxH1JOwjsVw+cMe/+HD1BaEmQ38oQNk/bFH
XP0F1E/BNw9OOf/p4JjF5CzFIA4vnl6qNC74gDGyh7H1UPrVHxt6zGJfc3/zhWDV
IY8rVUoODn/wVBqsFtJ2YmAHI6WvTfKaZdxzustaHmWpU9qWv4w24B8GQQqPwtcs
Hgc00XIIFGs/y9ghOZYrToSyg2ArdJpjCYxxQmAolLbqy16zKGdBwMpgYsYFWdxB
PWwVicGLHQq3LQ7q5HaUzZT+tWdatakyp5cwBYjYkYAEILzMijcNWn+BdnkzXs6X
NW4Ag7dnlpJQXet2idt58u6NZr2qtPqn9KxdB5Qe2+XrpPP3oJ2SNI09fG7ZfZeJ
d3hAqdVN7DnndiIA3YsYqjKEqDChdjvPMPg8IG+oVxMLl60dj3SxLWCwdRa9Tj1z
FrDEsaoWxVbDom84dlWyWoF9Q9czlgxs8QjUiTJaM5V1RkKv4Fl1dUNJNUQ1xVWI
U+ouInUrWJkyxmnYjPaxUpyKkYuEY+33h7INAmH6B6VVxMIGUWDfh4Vxqs03Vxce
5R8pk+ARSbwscNuZx13rMK6kv7HTmOF33lxAQN/c3vXwHFgZ8AZLdMbTq0uBvBl4
x+SQOeEFiuGShvO1luMTDMBNH/G9B775le2sKSot5H1XQZrx0cvK30fo0dc/EEeN
PTjARfl1yF3UmBZCkyhM3qepHg9JMllzuwQmvsxqe1MiMWJlu/DTD341ZiaeK/tB
jVrF1BzZuH5TIqtTk/9u7GbsApbXQvFrgbJl4QLB1/ZSVqeTkzu9nJjg5/SuXeDs
rbCfVqbquv03d1WEtB1aTv4Ni+QHjFvrcTxLm0vtWJl9f/nTPhF2hLlcwpnzOHsP
YS7lHuI+zEITst9EGLhHLBnXVXpoYqVwPgCzrVvHZtJreUuJg0GMTpB0D5eBEYo6
SqOwa8NmVcKsj+S9oo6BCPvKneTiUGG5OVUEZwZ4+K6OHcgr2qsFp7V65OGjp0z3
oPT8wfP6IGOtU56PF1QDGcaqvtzblUEoDAUSZZPrLuqEN4fau3bb+BVn6twOT0Hm
/SEesHl7OxLO/aufWJggVA101BetFRuRri2+cCP60yga0VuI3uimQMRaez+PJSgZ
lxFQY39qe4JAa9vJSrePhCOFwlwyabjr4F1hgbDkWyRPsvli3a9jKH78k7abitsj
UBdFDth/qfOSlQ5umiY8TYpdbnGSjGM06dXwouXW2ZKrPWWDaMn5npS7uVg/OfUs
hQtwA9/G8sJkunpWShcqqm1AyVGgjLnIDU8C+mI0voyC8d+sD06DLvkMNdWchriQ
aGRw3qt0VLpiCt27clwJyuXBdQ3nqanYFLkVPfr2XOhIZM818qNxZMx5f224fl5D
XhJO6a88O3dmgtankpD+j5O8mwt78yuFbQIl1QGMqTTPmz3fe3RKfM6/YXx472OU
02v4dvM+w8RlfbWEYt805ZtOJMicIJo6Q7NQdICbTBVDtwilG/Dbh0A9hG04Tcp3
v5h0QGAlN5EkBPHnUPiNQgucePCtHxnV3/lF4jMncYqem13JJzxLbfQqR3DhlhA7
tQmlIAvxOqcTlSaLGxGMYRdkwRLh8kK4cvWTxnuULZiAmKEs01Y4ATtJd6tVbaHg
H+4SLw9arcWCPN+0t3KEVvdzVa8MMDMrwPZydtXENLT9+LUxKUZYP6dB3EAYr2OV
FD+7LIipF/PtoY30EnhKIyHjN0dT0L2LHkPkmAQBscd/uTMhoYBt5t4LDJ82gYak
xYjhONUke9MtUHsvt8cWQhNZJ3Pu8TAY7DAUjdxVquSEZfkGewMIpHU0cJpQgUlv
J6au+HcPzleCBU3bbOE99mp6I3BgfIkoU2qP9ujzUBqkg6WXJI9BwCJAZA5ZJDcI
Y8iWraD2jm59jKxNchrJeUAEMH3GQamizSbH5f2bqndFJojWLVpFOVgs4dyFjAKQ
n/GltOpd2MdF70hMEyvSrvyfUdYBACkpR5s4UI8v716I0WP6rz6sq+DAJ0ndCA3k
dKL95vHNH0x7NLsknHnEHfBvWPmMOFAY9g2OBYUwryFmOY6WvK3wtmyRIiDpJ2SB
a1WC449N4P30oC/6PdHTphmQlpuUbFvcS3FTTtV6TqM/4p6k1i73Wq8ZinvhRoAh
C/GQQOlrUSv6e3ovLpopdWMcLI66rbNUy6s0+GiCfl0AR77mG+QXltfl71oz1uTT
5v2SyzWN5ghI/YLqqezvwuwxUib/JBu7ULe+kdkfN2FXwyXImo4Of//yEJBM72Zi
mnGY2PL1MxFUFx2d7w6b8nPTOpa3QlJGnYY+Cz7a3KOqQQLqdz2+LEhqiOpTsOND
h0dKy9sC0H4QbKxwGDAkx3lHm1TDYL9PedLbnE+9eJ9xXD2w+Bec3JsZ5ruZCgb0
xeL41tT4Cid0dRRGl1Sm8gljQM8Sxzj5wi6ahkm4fRiiKcV2X4x1wVz7x0nwrElu
PEogcQHyHCXmjbQyoZqzESi1D0kwHM+CdHG5oWkOv9oaepMULnhX8xexv+pLoPPs
ib4qq2QU6P7tr6EztV3xxoe0OrIL5LliHVN7A2QPsZhmBlQ2ZO1D8AcdDpKIY123
m720iIbZjU6Xc06FW+ky6xY2i4aO5ugIEueh8bkdzgoCHAs9eFwGXfpoZzg4f2jt
Z6MmJ95NunlW14RUUBqlQoilk2dB8qV1KlwndlBOpf4zOuZUhooGhklca62kjS8j
jAPRaKYFQNFkaV2G1pkarSy4McZc5ug+7KXDJSsHLTgPWJkOGPgBGLRF4SdoXGIg
XUdat53kQjoYYawYcZpfuVCBV/jM8Quf6XfOpqSmIade7hetJ9M7gzZJoncKU5XQ
Aev0mxGJtiZ2QrR+LF65/eum01j9dws6rd6NIDG+16F5URETxCpA2FUQJb1f8E/d
ZDSSa47+HfoIf4N641S5XxM+vBRE6aaKSpa/3+Sf8dTK5JcnOoO9xhdaIrifU6Ti
kY98yL4HpmNjGqMNrhfRiEg740ewN9huis374pj//T/lgMXiu6MDkEvWEfi3qSVy
BVkEoSMLcEgVDN3jjO58y4+4qRy398n+bWTI1QuBxq8WXmM9STSmqustWQFkIK+k
RCzxiXwK2whAcKLK9dfDleDmJcLxp7VPmR6zEEoEwDDeK7eNbnn38Te8X2HdDf1W
p92v4StXF3mTxtbsj1qBc51gCOQEMwe/lRDdHBYYNeJq895MRcjycxmAWxaJT4lq
TWka8z+5bpXNXSMTWeC/pzCZwwpncQ/bhe2IIJlxv87rfz3rlRutsm12fAKQRoqe
TUjvXi2WTRdAhGkO/8GXMwlt4LlT9jTShX9Y4s20vVwhNtFAyEeZTAX3+YMgVCF7
M4BohDkV/4+yypWmdjOPj0oT50Rt3+qNRBZ5d5gGKNeAUvzDw/Ivbdd+B57m0kYs
jnAVKJjBgcI8lPYT0HKKyraJKnDwUpFk7K4dmFm/RKgqnyJboDMxeqO8hq2VXGlP
TSmGRE/cPzTHRpFe9iZV3DdQF5w79l959qzgspnxGY12B8PxmrZX2PW93xS9Hf6A
1XigL4X/DNzpnBRB+XgudUgX2+6QFAdpOiAm2HJNfYLvTowmE5faoIzeehcwQr4k
WZnn/1SwFo1KDdbJ0vDX5wcn9H8z3FlJiJXhTWi4HROmnPI3dE9U7rakS0r9NZjr
D2hbHACfkOYiwhwk2LTNzWg2ag7p1xYYfm12DWgrutkMSqglegmYmcBqY1RVDdHW
1vtQxGLgL2aS1ARTuDJtaNG+g4S6mvws92xwAW9oCzGUWoFw15+F+6hWfGr3+hm0
ogb9SBMh2ZUxzSwlJybLsCg7UbBxgim9CoCvEAeM8ZNVESA9fn1LZ3YMgsqg4taS
RwwxZyDqH9S6GOfhE2WMx6CCYu4R/XBe3HIkBPadmSVNrmh3/N9bar/himofWcfJ
xam7f8PMuEdqqaTUY0ehN9q9A2hOKNmIKD5Kt/pLdtKcfA8libBUcZ9udeJafFGO
qWajHkctAaBuQj5BsSskNma3PyT+vv3IIrzSZv5rBZJGZTtRgwP9FBO96orixvWq
OKyoNzS34kktPW+3J76sTjRZbdw2CSwDADCXurEc+BbddsmRirdZn8UXE/6CJGMx
ce39822pKVRdZfFGdn384IfydgflWfONfA/B+B3Qw0H8N/Gn0vKBf+uT2Lo/OVaU
ToRmIyBEv7m24AtgpkxA90aEtf/xvIc+4KhshvEYeSepa4ekWekALxmmPgegpaO5
AXZaz7UJHfKsWWByHGPGcBwZwnT+YxFjHIAB1JwrLyUp03bWiKQT5uk+VqXSS/3v
Texcqs8sp6g6kXokGKAB5Tnu004+MC3sFWha0vuIC0tZ2AqyilosFeC0RSsrMyX8
X4JiMab/B0ShJ93gpriK22Ly7CDfIskQlIoGpl5DPyTB+cfFgaf5CAV5zzJ4ZVLT
QHx/jIeREb5hUvJzUprUjwctKDJKFr4104/OQuRXu12FG/dWQzBlJCswMKaPW718
NrIF0tnPW+Iw49Bvbq8acrXJSBMA4qA/4PAKia27leKvsZ4fwEdQ/zQyRd8V6PzE
ni/pQnf1VzvVN18x/MLcvK121/ZDjtvT3bcosoJw5CRjqeyHFrKYGbQ3/wqNCJGh
K4oKA2ZZEgJs9WGDCRW0jbmmw55pQv5Y9lQtq1JPPM1p3zcQGl/pFxpu0u4/V0qy
XEZ/kaGGkXUYx8dZjpqqyqJcuuyuU04ceH47FPDS/9Lth1SjCWGhoCTPzvTCrSwT
vN8NKBUDZ4xNJQlmz4BiZ2aRYyrOUDjJh6DUm7i0ZS3xbOSfeLx6CnuLZOfIrpQO
albYxjBsWLdyx+CmEer39f0Fce1cRPeYCmjP/nBxoxTS8LSQSwlypZkCoi3jKbDr
ZgwTRsN5xH+o1Nh+xFS0/sGpO5YwGvWnFKt4/aglkdbGgsNhnl/sOgxExz/ZSOvE
dyb8h+GKILEwCvA7AWZixiNicVCtTMNwhiAAozQHg238wHBI+3s5gT+uPZHqbe7e
m8Ps8+jF0wINFXNcZ3OFiVLyUpX+FhuAHsg+8S1Mv1d+YZVVGWlG2k8w5zlVuECh
MWLFymsCPXFqp4NnOIUpPiGS5DOQli7BE+HlLD2w62e4a7bT9q7P95GADHk5R5gZ
M/AIRqipN7wKYCVCcfeTdDj9bz1ofucCxbWQ+Jzwf4Jn7SU9dUCc80kyltr2aPSX
HLd68H9IJsIeOWOT8T8DronCiDAIqNW+Cg2oYUVfD0p2Q5UA+F9dQNYkx53H4L17
VCEmmMVxsWFMC5BwAzmYyyq6DpE3n3EGOjaqyNo+mHJmtSSPYcjtN0x72hKn3b+e
yir2ofu7zoE9Xa2xuxEE4IBw0Ht/RwRO+VjmU9SWSVgcDUylxrJGwGNAYd+vmE99
7biJcQibfnKuWWJWGZlLISW/wsNz9Nb0tvfntjmqvm4FREltxpHUiGDBcaLzTawm
zfGN6MVfJ36cOBJYOL5k+f+jK9ruzwBxaXaP7OtGi0l+t51gdSGPi/OBE5LcFxCt
mF2/GNy+8udVb1AQgUNBHrDDesCb0KlTNjjrSrzriuQseC8BQRf4t/YGg/Svg0bi
y0MDxeg+3ItQNGPIF61/nYQurqmPsbcyc6Ewo+nkVSiiWvGdM7J685eHv0LqHbwl
HWMJt3GxRLX/3KJZu0b7xrjKjt2B14N4CGWr+KyFk/BBnzvsL2EsGKe7pnS1xvgV
1PHzc1aoTikn0sW5YP8pwY3o+d9r4M0gI6emX9TQ+ihWXsUEXp+mZ1t0Dxef9kOu
DQvXaJ5ejBRexa+mvdkXGqlgRNRJx0lY3xWZxbG8V4ZTRMIzx2bpB2nuow3AI2Wn
YYVu8iVAYu1JK9kMl7TJFA4UyEwT7wJt/265YV507ejbSt2frb2bsZ7msUMgEedH
ID2XhIHO11i4Yoh3DjaBnhAUYEXGNyIMBdnTZkB9q34YgNTT/0f6ztgRlebizc9l
bOEb8JhJrWpYfRi30QJKp6wr4ssI7iiOjmXlQqzxD1gY7UdjbU5AiibbXtgW9bjq
ad62/TxSoq2dqYBdxhOVO+mmvJ3+yVzaMDLQh3bg7j9lhUM19SU86d79/jlN0eJ0
kR/QzVo5XZLwOfJzHPwVrhdxbvFXNLbaD9LS85FjB0Lx6IABoOrMU1IuAJO2OqUz
/qzjKhgLVGy3461xePNtonx2WNZgqz/ruOxf+ZV2M8cEh+z4RQI9B9nn2FDPbwWx
VSn+pZw+BRCoeJQh15EsvbAxBEKYsdwBXo2t6MabAbyNXTvhH10HKSujdlFfNP3n
+PVoEQM8Ln6/UgtFd4My1SK1pY40wMvbFxO+PB7vqydebxL/VhofFoPBhilHzhFw
4t2cUAW+06lmAKzMXqZBAu1a6k1DaLLplkheIsEKA93vyPZlTGDBxWd6TQeZK2Fo
ROmFFYcVzy7KTg43aAhrg3BxAn9msVntTurMO2Xe+qxmE03dF1ftgrEugdU5m1FN
m6QsTocmKz/xdiTVSNgkQ3u3sQOy1VwEZ+LunJeS84eDkNiewuMhE3Gll+65HIcW
BVi0FTeb/FTq0HM5opoT/HKffhzaZ+LtI4tab/E8o0rkRFmiB3M4HpYhxYiA5jst
JvraEMMWHfrEDY/VQeiBe/IVWpaD7md4Jti5Hi+1of49SAnXGnZ3fjG9xX2+kheX
UqJ1+fr/J/fjIxpBdJEnv1TO9PnKD22VVtlIpk8hSihgntTdMhMPdTAP48nwEKkL
Yjq4JYOFj59KVtNAu9lyzC6fGwG1akv0XCZAX5JVRKdqFDOzHmbmN/B7TSFzSMxr
mAn7Q1+VnqdgxHJDsgpQdSLn5bHBxz5cuCU/5whZM/3ACtxqx1LV+7HpMu3DxR3r
ZItt78MkYZCfka2v8/36TtYfxWmJTl+lJIN/OfBypDwCpi66ess7Ss9/U2aRzLfl
a3hHhSG8khY++JWtmNJ8cCmcbDNnDpoYAKOiJIagnvwmVIGeqzK5GWhY6QjByPO+
oWadkgQLKgVuhaXSASJ1SR0zZBuQnCTy3nZskvTDZZ+Wy0iMZ5QBgg/XCJI+jhEH
4WNIEnj2dfy36B/wmzrw7uwuAzjbprcnvqTwyZZb2VAYNDwi3X/BkjFoN2AEpK/m
yc2L2Dhlqn6toQjtu4HKd/GUsqqFW5xpgIPptvIQHTM+17Yb3YTKnLgJ8KZwAhrQ
FZqWNgviN2VFylGmj5Ksh4A6Xj/6GKmcIVxSyJl1AB96v6Cyl/dPSGbWFNEHV43z
LOhxY8ofYwSHJ+uO2WQHDPf3Y204Mdr9/GR30D/+cPSbbRW3v+Ci5c4VgEdpI56X
TwCMTN/yNstXCUv9uL9s0m3ImMraD9oWXim+ZPtvuLGLSNeErnsXY+Q83x7scfS8
yWSPdIPLyS/yIxPc7/hKkQEcpJsk0eukIQ0q+Q4PJE05RzSlGflb6L7TYcDjsT3T
yJ45IvU4DWzmrL4WEIU0+i/PNlRxHuZlnjfRwUug6f7L1w5+vTdseL7NEPb4EcDn
dPK7Aw05B16w0RT+lz+iAzlIHuXXt/dn96gmtV2f/re4+kZfmA9koqAid8uJlDsa
g0AAzcH30KHwPQ/+fPzYMpWxWBhcZ7Ptq0zjeUzrT/B4m6kYu3kgDEB/LDmYm3EH
J8e8AE3kj0aJVCBpvmTGMSMPtQ0mo99Ovb/weZlrKuDOELLCzhPTrnGlxx/muGZj
QyWnvo0NkZt7ylR163kQHUoGnw63KBcnoGWISpolv0gzg+70sWV01WUgTEKdoAvz
rW9f/2wmN0521SlKzlT9nEJ/rvnHxG4M28BkLqESFDJfXRfGWeTSooAmU72TJuDF
3fOA622CxxjCeP0BisEoDYD77c5P9pCXG1BwAqhy2H6sIENhqVVX8LBvzK/+OEvR
KyBqcvvEONfRa0gIgKMV6gz6EukYrDk7gMttLXbtjCfduP/mbs32fIKXgj/hl38X
du8daHIEDfXMTVLpOvSuZV82kUdIav+LvJY1OBdTxzoZBLAZZz+vxWgMVJoGiieQ
jwCDjWqvyzMtcb1bmv1pvq1PsEdDLZApBS197+fPfI6I4updz04XG61GJF/Ry1IC
1GeFqqVIkIasVdMrtSrD5EeY/gSxZUq+mmqpYAqn6sgQUUvDPRPTLZ73ygQx2fJY
Sgx5cpzTT/u3ytm5rm7IXneG5JqMGAYNHPpa2yzWqH/Iq9qW9O9iRZRifB6O/xGd
SyzvNzp9bwJUkUm0ZSqiQNvKrb6sqhRGRyEMxJJjcD5UHRKY+FyL9Yu284ELlvcd
D0Ds2LMG+GD8DGC59QM6Cfa8DeryV9YjcuRbd0Li5J5xlwZ2jxnnMv8Zq9PbCpgz
u3dA7+UD8nfgGW2Jesp1ahN8hjKKk5Kf6Hhen0Z19hbKlKyPC/WvRL5SJyvzGbsK
Fpgzm89j8dyYsvSwQaMoYmHISa38mKF0hsXn9KJHF7OHu9Q+OYUqyM7MbRhZtr/f
lmB+4FZlLR/EkyLCxJLRWQ9BLx5FY2XDNOTrNxnnYInu/T+HxzLUlNIoq4uxKT8b
Vu0S5KR8OzJQulinSF/ycsF0Z9/mbVZ68Y1+SCKhBQzykVWqlIvggJ1tRT6z1QIO
yXycZAjWuXow2zxj0HJTFXqEcAWgLkH+PzzsyzX7VBPFjjC6ZLaTEHe1o9B8Z/xq
7SZvZAe8qZQDyA6VNJ7q8uYKeMzxw0s1/1lTSyu8ivrk4LvttN9EX8+uToC73EGE
xFahnMCqMD69H7W7bP0dgFlbQRNP/LM7z+rxWpQPNMGqVgoBkRk24agzfcCODaom
rq1Ddmq7ls7sC9O7yiruCTEunq1V3teLemJIqjsgfjw8X+Z/A535BbS0awOcpCZA
x8D5Rg9C4MLVUN2o1PQLyIVLf9XJbK8Q/IvZyQK6pNzuidsAga3qOKFL9pQtPwMU
g8+jkoRBBKHcX+4+v8yGORrJbUdlo21DSP+ZLW41RstAOLJbStGsDG7gC7IXhht+
RgVGhhngY4389U0O8Gkjcgl4iVx2iH8+2cBwHxVsDBrhHIYxL6r3eGhs0ts/sIgH
KNfHyUJvL2GKEAcD9rYSzKghH9dECQfGinL5b/2hnq3Dw/dkW2OOOJv8474XAeMR
PmHZW18OfAlf9BsXlKJF0Xi2fV+fTKXa3hbcqhJtTvsP3GrXWHwuSsIYLkSEzrBp
/Zu8JTTA7Ug872dTJR503hWvvin3ym6RcEguXaf47cP+kzoNPALu+UiwDwGnUzDu
FQz2ZAFZ6nPMQl43xHiLzgK6f3a8ZpXTDyvLuI40kth16YdbGQeQdQGbOpQDxC+b
d7NW8QQTEdOP+m9zsMgCUgKa/bjgT656pw9BJCrrrGTMi4BlAxiCfWPktobsVwVJ
XdlAsfG8D9DvfCTeGsFQFaQWGGi8etrT+yKS8x77iAG0xt4HnaQ5yn6K4NhAnJl6
yFtQEgbO4RoY8FMLjI1F8eV4RmeMUj8TzqYfJTjJOMoXdcdWCWqCjJQW9a68r4Yv
+rEqQ/kCQXyf2J8AevnsfOabyB1LTB0YTx9uWMPA9THxkYIB+s2b7pCG9eIHkFP5
J+bUQDPKpFBCPFJB1nGI5b6y3Is81/uQMVz3VnPRO6Qc/b/OQoJSvQAEIkCHz4x2
qWFcer+aHzLwWmJl2f1XkhJiDipzGY9A09fLMVZ2MAHUgQ2s2wPnbKqamuPqeSdb
WZATeRZ69BYpagqDI7VMTi6uVCeD8aka20Qdx8PVPgDHQg/AIUwdEr5tc90Rv+JT
YQMebO79Au7YjkfFjylTETYflSbTKSVDHN2IggmZGEpkRGyKAgStFJ97xggZuiWf
59k/++HsBNFMj+QpssTcq7cKsSqMJBCRWl92FHzpj/VGbQvTUzdQFb506B4yXdo5
SUt7R6uEZF8u/UsJ6Qctp8qzRtJvoCYbp9ke64sJzlC6hnwy67469y6w4lYaPvY2
/Pj69v1E7gKnl11MLBPOiwHUlFn5+4CmuC0kUSjA8sTQ6ugztjek0/8rkrruuu6D
dffwOsAZ6ytfay2zQK9hOcrG65WryJoHFiZTK0l6Imhodbiav66ZSbJPBLHwKAjH
TAJGcERggilzoDSniiWno6Zgj9QLii7ZUwA5jJSSXtJdHZTU6gAH13tEvPU7kTGf
CD0Q3KoixSVXDks+pMJyCMY+tNT7Zj/uj/8xpbgHmlrT4bfe9+pzujp2EiisVt0O
MXga7FUJkUzANlLrz7lB3EFW1+F9H1l2iU+v/5RZ15BLAgkwKjcRAI4wHoDJGrtb
65PKYdh74/d1daQmHr6PelrBZR8m5+dqte40RZ73P8pzrNRzdx3GxM1Zeozdbvrh
Y8Mv3j6Sq9Ahmvi87vgBJ2yz57UhNfwsSJZkXEsvd/tLRSlVIBG/8LtQoIildrLW
086lxsfLlYVIUvSvMExOQyv0NmZbxflrjlbUiV5ujzSZdKcHTxHAaluQpwC8LHo8
9BH41DBkUTuS0zyt589OV3yZgnivJq4e6G+ZEN7oG0sYB3DT0mQS5gOHpetg0z3d
M6gMjxoTnlg5WwToyremu00ikTP8QEE7PiyNwP5HjrQ=
`pragma protect end_protected
