// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RAVZvEd4VamkJeMuFpIMkt6vDAyOiXB5zq9zI3tw6Yry1mClHv0qTwb23uIZoCuD
01OOjMZS19qSoAX/2i5siMglKZx5dgWAsZFOGywSpqmSf/r7yhzZ1clTgL6nKo3X
/drnVngUPTocQ8VNtJD+A9K+e0Nu3t7Qes/ObDB8zqE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8208)
7H83Ms4cWEmDM7HbbSoEYUJdVuwD4uQEMPdfuJvCHoMH6H92Wt2v16r/cqEmfyWQ
jRXgP0zbvtIyEKOtOvvHxF6ZchHKZ+iVML0XmvyXu9XJUHVe9r4b4YA9vf+i/BCM
LRKt2ykQJY8gYvzkZfZsTrH/38EfzOnkejbGss0tkEGmDRlzdmeKK9KV24uMPUfZ
RMDGUr1DjAQf59O8pXIlCLGlKeyelyr+l1V4p4euxdElAmCuOPmg/3lXC8zT+gnf
bbWwywBmRxQOmkZvKQ6QY7x1+ZeEWn64/lo5rZWfVm31IfgXKPYbeL2nn2a+fonX
QstsZfWibJQrz9x/xtPhqHUtsoRjTmdpmEYnEsr51fLXs0Axm/EUeo9OahYTuKom
cWG5mQycR+lUbTY+W0rla3rBe5mqh68YSrMyxkWjUgR0TDlOD2tj9Lg6jeI0SxfO
z4a30oQe8uNAi5KduANAl2tODigp+kUxldx7cEZA/o7rfsMFYSU1YDhfmrLlVGkO
aRlc0zavs6fX0MTNk5d2SjAzvVklHoIHY4N/R5wvSDHcVc1L0hZX2dTNcxo0Ch6x
0P1is+EE/mhy6M/MoppQFNpvpwf4OQ501PQ1ZipeBIUaCUj/JC+5w4ntNwTNzQlS
latm2zc+Z1OImoI7U9wLRhku4l8/puHAYLI2/jQOdMRjhdcDrjfNmzuzko1y8Gsp
r3MSKhemFI+QZ87yw57hcvb/Fqz9qIQfIKwDxKM1BHHdVa9YUdKuUbGixK7hIyoL
igZX/ciYi4v+qJYgS5SSS8ghxd+mrWk+q/cSVn04xPnxIygcCBzolfBMrH+6Dzyk
vlImZU0t3tw9esGT/agx9ggyMWEc4Mx1rtU3csPQartipQMrFXmmKvT2O0hbsepx
y2eobGtN5IRlox9N+1BAFkcwRYZ4pJqjJpqcBWOd37YZ9xQsi9nYZ1V1znUp+2Du
eS92Sb2ftFr5VvCFFbjVPIkrtBIVMtK8V+cIwymD9Fd1xI8alNcHza1BCX/Cf/OE
WcsUBr0Uykw/Dl+64X66Ui6cn7fzq5Cm9hNxHIi7plggQ5OS0BUtmnrFKtwxYrlW
TopZRBCdphVf25jLpes1w0zv8y2RnyzH7Mx/ErQsG5lrjckWFzWF8r0M3Rlh6OhZ
cSqyHnQwtOKRK5/9XWS/5Ct+Sfl1VJn0jvp0MZLKw6sCsepwzOCvbXWCWpfWw1e1
gek6wlU/1u4KVsjf5fBkUBvd+aDUAje1CxvlKpqqmOWkuoW+hGh1O9YTjH7wdjBm
BMfusLajjZdcxXq4sLf1fX+obWHoWPpoSAuO8kuLaenuD2HdTRjaZVs+HXcgYlvE
EVWDPZDMKpIjr/58fCXRHp8nAmujBUinf/dhh5zXEqHjLk86d6CWZCJ0/y5lGkIO
t8Uzp3Nr/5HEIh5XuxK2ytuS96GGbhJWE20A3nrz+4kgI6pRZ5aPYRY5zzultlCx
9jcQ9h5rRmlL41W4frYQURF5QIS8oadjbKEdIQScM3NOsdwJZDUYF95UD4KcuyTp
/tBQHP4buYSMO06Cny5W6HhsNSspxSRfce3mJ2IHFG/v2oxXjSJ8g+Kp/hjbLIv1
m0hzTxTku8KvcQ68cMYPCwkzJjCTp+rN3NqDlxAiAcA83woFUbWDl/0JYwXDURj8
Q6Qrq7NYFbcSpGvUss/fUm1+GxFJnx5jOw1gZfc+gm/mq8qfGEopVm1OadvCB/My
Xu5yKxoBWebihYBmUcfk9+YEISzDTpT7rooWtZsqTx0IFCp8dIgdhKQNBf+c7J0N
mrr9el9vMLih9q1yobIOa74pyyIrFPmnYhtHx0hHY1Y1Q+P/EXDChoSD/DUnyaqY
uFs37ADUkUVjcL6f8UtSExVjft0yty3ldFRyNzlA3CAGy9+9k4VWovpIeXtIe9Gz
NZdu8Ytpsu7iEbVdbQUt0SHws7bxHY8Lo3i4UQbz5yR3zSA2YwhFlgiyBjQo/5V1
niry72cv2wN5XaKPHM5AjYnmYhWbGXesSyXGhYyVKth4QWI5Roes+PXU/nFLSM0v
O6AQPaom8u+biGPjF43bantlGU/ng+7GlyfSQot43GU0nRI9tGGEGlyWr6njNt8+
I/IBlEh5tLoTv1/7N+Spy3SmNCWUS8H1gEoOfQtwV/4Xa1iOciVveOuKlUDCsEKC
Cuz4+xRdWHsysqFlKfnk3mm7xM6+U7zktzper0KS+VHeI6H+z08F0WLLyOooX1AU
jhL5j8AFV6IoqupMq/6BBo2vQ4VXdkZ/qrYxmVLMMS7Upd/Hf2Sr+jA9Q2OOSPyz
YyjUg4b1j2La8z904XwBluNJ5lH2w3r/cgcffhzOoh2Qlp62sCI0QrO4pJ1X0tpV
kPAzGXR8GQDMIkRG7cb7aeaXYRhGaIpTBlb1A2rNGoc+vTAbGDukc3bURz5oIdYk
cEiqgXpIqbWXTrSP/N38XN7sad08prunwFlmSkWkwaG+sfC78+TzsGwg+Q00OAhJ
fxtY+eC5JAaKDolpLgZln3+q+yCqjtTgPe+PAcYe8utBtrUMYqTZ5wjn9n83JMxo
bM0Nw+vquGiWQWa0azcxnlR1LOOduMLr1eBYjWHdezNpDkdqlLtV/W9z9767hY+G
y9WSTtsZgFI5dolRQwA1vCh1DgtMnutNBhf8ta402k8iwM9kieUhTBSPFAYpcbN2
UbTiv1z2uPvR9jmIWnfDSzty/xExzRzT0/tMKAcsAZFAkeBoH3Pu+TT3XhYKnkvq
Tm1L1BnBhGTL6tgNUXnYYTecF2oM6G37cCrr1RIXaxJimvtoKMsWt6zKDiFOoUGE
QEuT12FPPuR3SCafwOUp/avTOUhtTemem+S6Pblf65WiQGXmS94wz0SsFIxIm6um
LcPJiUMSDRdwe2f8PiicA5HU67H4LHvXTUl+tw1kBYlcHpEDFV6Mjq68I2pZ3S5j
N60nJQINGMOWld/SYgcdcZFda3ZdVpyOOVFx/skUJJSSBRrujn3gGBMyobX92/7E
5FM/VAHpRoqciaGum0KEEoV8dgsBPJAovAfNH7Z7DCUrzOKkMciMI44Quta51On+
eRmwIq0QXWIk3mj4qrc1A4W1EnsdTtfkU8g9JWQLa5sZEMPSKRkyU2sV03naDGM0
iL6Z5R87grTqyjcTo5j2wDIqak0pgJiPVSKRvpSfgp5CAkbD/2JGxzdlDVXeOQEr
itFkobyEgN04TTQJ0kGfGZ4irMuHim5en7ZzzwnPtjMPKcRb7sF8eAJA74PruvQe
45UXEZXff1YrGoWm8IHP7o5eEgMj7HtyV4Ugk8lEZJ6O4YCcKPRE6sY4Eq88krD9
G7aD8sZFRcjbbbmQN+m3Cbc+qlwJ8d6LxkpYv4NluGdMCzw5Luma6IA8UtNNnP3p
2LrbpofYYndM1TOSc0VSVlE44WYlKNHjk7F1q4eTQ4IdMw401/4y8B2+Id5HiBPc
GRYAmnAY3AwdvX0YEQLfjTVuXSxEU/nk6xt8BIdkr2pFeTUuMZB99GIuIQiZjE1B
Qy2E7WhwBRcXRKWeQbQrPGqKo9fHo0Fq8HgxlMsW6kAm/hzQHK65F1T3c/dFgJc4
+QSvNPINyFE8xs6CeLkk0QeFtQR3pHxVNa0yzpKB9gUYkmtoOVzOVZMMcnN9S4WD
rxGVp/UHC9SN0BR3QuEzsQCtX/DH+s0mVPBV9uiNUp+1WWODWhoyUxz7A3Vyb8Sa
DZkWQUtzBJs4qwoe9cd32TFBlY7USk/kHg2KPB6Czbb6As8Em/YJEI/NP/3Q6i4r
O1mLKi7lvPMgOXQ7rxTjrWMKqz0Hnj6qLDNoCdkXqzXgR/t6f4VfTvZ5PF7EcXG+
L9ZXZd+eu17VSvK+dX5G67qhHCeDMxX3GcxDcfU4crkIHLL1nJQmHrSqmKxdX1Yh
yJ/K2MEc+2rwT/Bcf1/3Eq1JEHwA3mIIQAq9wquv27T0BFwMvELzeD7sU9YQMV3f
B5iRGKdRDSjiPo/f5OiXzSqoN2t/KWXetylrR21OeVPLYL657sXE595FikYK12Ar
4zaFY4bDjplBUc9ow7e6liIsHYJcUeT3HQOrk+xtbj+1orbY3p7awHOWkxABQEi1
VOB7d/cPBDkFJ84ijuUMz9x9+G8U/noae/WVS11Yvqb3Js4po7s5yE+xQLE5o6eF
hbqQVTQpVRqmFuEzAUZxpB6+OFup36gGTxYFY19uzLIYJKfsmrLUOYok1dZ7I4Rl
2cdZ4pJFuUBLa3L1z5HWeHPzoyGyD1OpZlLryP9OqxMIUOAhItDI3vEp8tZWTdrv
LKJNADMSZkMWwBtQGTHJ2KO6koYsopCTqNRQwOInigcRIl2jrJ95CnMewKmTdIPy
zB/9uEISF+70R/FULO5S6wd09hHvSKogXk+/gF+9tVPblpfyu9guub2RRPo0VP4b
c/ysm8WE81rxUvP1HlNdJnguE40mBcfaUVBNWvCTBRrfTEAbMh4piMDW7HiyGMDk
5gM/vQ6ILeAlMgIexmo1qdnEpHkl84RNZzfqBYkdIYPz4EVVSTzrtGwq87T5OOSS
k/uOv0a91maHUAVncmioEQ/1Obsu3zFDFwKDHfbjuCY7ppk1ftzT/2WV/cdUAgwG
cz+wQhK7jJuTM1NRMCfBy6PykEJk/nIMij69kxVpp7UdeUAYZnojK6EjQXjB3Oqn
YCH4yN8bEU1DL06qw3DrBISYORTAZhcqEjSNM5eAv/Qsa5bwLHVGD6X0Xw2zFDoa
f6vfDjXSEht1irTD2KTmm8ZstODb1HemxdC+y2rHRpoDwmwmW7YPglqYpziiorC0
KKceJ339gXYSc5PIGW59d2nKRqNZj5n43XgtGxe9vhyZNAbFgtAv5x+526UETwSZ
XZBa2WkaeOM471idPPgn08zk9Q1aG8lJC1BC1YNqNLnaAJjEgAvSG0QO7bvqdI3e
tdsB45IGM4JzAjt02EZqxNK4CMf0lmb17FC2Qi2LCemybIp69pcEUQrTgd1SZ4Bk
IdQT70Vx8MYJXDSAm4fob/bMsB6X+LOTqyECOmpvq3HHGOhbN9BsZQ301CK6lFXM
ICGMxN92Db6ZnTcMjJ/SQJ2L2V2iEdn0IPePIUlyyHz6w937iGCdyTc9edxfrowS
LlXD0CvfsjQNP0o/qRluAE83eP+O5ZStkJX7c+OTRT1Cxr9MMaF9hRrkkP7BA6et
2u4+PVJBNzr+aPKD7EDDoxdM0iGrrFsIBdWisOfybnUVsSBnGb9P6INuVSuwTmZ9
JnwB5UuijtnByvvcuo+N+88b5h9EiVLOVswovSVkc4TuyLWgX5vIP56wW9PEULXQ
G86gp9uH7QPuHAEX3Et0+yYH2ZyjyubSA0g0RW7bF+dSsKQr1W2D10FSCq/Bdgho
7rsmWVOkdcCr4mDCtTOb5OurCVRE1tLWsaGo5utpO5GWm6F5r8xaD7kZkoBSZDNw
2T6ztTan6MtlMNVLUL/LCL6s9Xr17dgn1Ri2kr2VmSKgWTFZ9FCY/1usVOcDq+6g
WKpXbb/Z2XP52Lug1JXqGaHkNZuytHWVV2pYsNXTjBOOeX7slIveXN2j5HvLYqON
ICebQg6kzY5tBri6eZlBmPrFfZnhVNnz7yWFKyVb3Xb29E4qTvUbXDINKCYfw5qI
cCd5pb3b8/qHM3JdZSAPVMADK83H7jTE1yGmwws9W9BhPQ92Y/GufLH3t27txlg0
uAZZY3u+fbKx/zhYWDjVzwaQsSGlw8njaBc78hfVBjGJtVnkj1MwpodOg2EuZHeR
9gtRA/ABQBdgXgpveFepE0wcNCRUCbErWuJPTkODXGhklkkEA0KW4xU4Jk2OMAdu
S3BaHsgTGJJ5JAmpEYmTdOiIB+B16sARRCDNJoCLVBY+6Lu5wjdZjo93SC6r04t1
d2dz4vOgN/2PVdAr2eDk8GN5wORqxP8ejHvNhOafPRmeytaGXKO8FLCprfhD8aZF
L/g9mdri7/s0PKTokq2rQe6Mg967OJ5Kq3f4H9uqfP2FH/Inm8JwKBVwmvIY2g/Y
rZAbytmuhWR4zDT8Eop4nAFLWCpFZJReLBNo81uofF90aKhUk4y9lVJ1oK6mFmNn
e3cQFZu0hPgVO/S001s2qOYRryXT8THB8/Tp2e28yuPccwmvUSZIdXJZGI+zpQlD
LvURxNvjJihtHhUKE0ihCWMB7hqbN2DzF9C4Xxyh8o2ulBGGRjqaHOztrbXnukAm
Al89LebWR0MBqX+WywXs2zBkxVxNxcSw8LWiD0AHihzcAzDIj50lpGe19I6CvtdK
nj2NkCV6FXWu/lrBAD8Yu54BcSAUHyBI0jQBzsf5hp5r4n41bEKNZNBFrYfnXhUy
vgcvJeDDWAQ8xAMHT1NQf4le3g93Dc3R1t3k2KCS37SCc8wf6kYJ9wGh4VrpVK2R
vDQXwhEIufa5c4t683mtEg25Ng07jh42kbR7Ws727UVraXpj/Xcy2egM4xYWGZ/A
RGQ8M/OsY1CqQeK2jMu+a2sR4E5ICvF0c5SWMrLfOrJjeSJZurBOd98IT6OGlZVA
c22Ke4jz+gE6XMisheiLdTx0/jIfEqcPfOkiw4rFLTkUPAIJ2aovNE8cPizOr1iY
GFWrLOsOEbquyZmcv/3rCG0l/1onQo4rS/9QLdSJSo66r7+vdvVOoe+QHqUZDt44
pvHObj/MPgzbdO6OMJ2PMNqt9LE027dTUk7+3CC+LXECXpSJopdP5Xj8yXjCnSJe
6YT4CB7Fk33/rrlbRa6tA9Dvpsx1MUWhRgpFdY/huxNKwYmfE+wdcF6o1xrH5PCp
fRuTHtngP/DnDrYWCD6IORJGt9iHdYXH52g5ztrvWV6PD/MZ1kMt9/6hXr0ec4VK
xZL0psPdN22Jd+QuPnB+KTHb6ivXlXRLfuzlqNKLz+5DgVm20g7so7q54RmQOnsA
yl3QXV4y4WdMsN+ygx5suaW6F9e4vOVr1HjpfI1dhg/3jYAH8DwMpJgsqRj3mI+x
fdPYJr1EumD4rJ+XBC+6D3SjsspvThPqgx0YbzuxKNNCAoy5QZczwf72illxcAbn
qApRAwE4JXHoAtSRZN1lWaGpvOSlPrmVccWuwsXmJktksiBB3xyPieMJpHu1pA4G
5NkMv/4Bhagf9Arb0/UE3pLhI8+yfa7OhBwzEEUmFIyBHTFlHTQEDP5DNR5lmIB3
f13LVVAulrthOg246piMNONHUC+/7XbdOfgZi6nNt6CofVN2jr9Abw9jWWblN7AG
5V9oAIfzQea46m9pqbAc6RTNdwGDLlx+OA7knvWLxYbXv33uwTpdh1yp68Kn+33/
pQWu6t5MIuYMrAUWRQJaclt+LkZiRmB9Z4T8Z5/U9+X18MxzKad/Rh8dobL4bV/u
ecbNVv0CkeG29Ryf+DVHvmWPLcK+VCBriMbbvCcK5r1lb/oDiOLhf7zB9hy3+aNl
lkSpnLMn7v8mKiIupAc8JmTHNRGOgMry3neMYHeKRNJmjkouVRDQW4E+ifbF0tin
khm4WR3B5mpCzAzcu4fJr879OiPmFSeWS3suD5d/q0tVxfzNy3VVOQzA/cgnMAeQ
qybFZqagYHr9VbVTqrvpzqZoXgdq1a4yQeZXgcXyeMTSVfXFYaEHnGAusYpzxhg7
Iobf7EyUiLJKRdthIhthH++QEpK0PiLKUZ/8+7OF/1tmrI9TudUuq3unlbpXeS4D
z2o0kKSNVkBG+WCOoFCUI3rp3PNwCJix6cJz/dABBToyWrNHaI2Y6z1WbUTi+cts
cAFA/hcknix5IGbsGkm5+nsFqSgiOfHjKgwTp1z6djSY92yrK2SvdgS1tx42FGm/
rdpnGWT2N+DczFUbRF/ADWQU/9tPCLhfPRoerio75GL8NdQWCKQ/a537PIVJhiKI
SfpQlYGKfvI1lfJMJO09IEh5kTKy/w3IgNICKprv4kugWZFlWz1LeFyGKgPf+/F0
NYOZFeFUtC0ooUvbMi8rIqqM6B+5EBXGZ0KtnzS9b9mzYOjK6omA33TeesUjy9bi
kPk2y9sbq9xJwvq/83TOP95aws+Eh+VOgg6MYlzsi0ykhOMTEpGJ14mWev/ce4sv
Mn3GGUeN+6B9JmZGVlVy5K+yT/gyf0hd6FfApI7KfBP18ujbi++9ThflEhVr6uar
5IJD5kvRkQRtFwh83hOQxYwXRysJ0mg6zfJOUl+4QsMPBYWrEh5YuoYCQ4R8IMjj
xCwkAFpEzUjVRady8Hn9N389XGPV+SUClWdLaGdWtXa1iZ0coSYtlsmQxeNdoMZb
qDcsxJyjWaBgCkHwk7UKCy6PqsWSvyJo0qNP6W/Abls7jiZ/DhgOhd9wiHZBM8F+
h62WaUqf+hmRGsj6H9hglIRDpVtZQEIbbc29mFBQNIQlSuPlcPWqB7k24xA3o8oU
1UnxAU7lTMMGuTMhG0xj5SLJL08NUi25ouEGutocv52AGR9/qoNqrVphxosLRNpH
QRGlzfrWH5hi6kMfp8tUZgKcZhKQn+wXdEH0RvJZhJIqhUJQKDUmprrpKsk2yK/F
ddR3obVy7JyUFtyM9C8UZWG+bPG7l2hxa3mDDVsslVbElieuGHso8LQqoykGbIb/
LezUh1t18aQH5+5v+HVioSJhIvk0QeLuZI6JDhoCIP1DuBmVRD0PJGRzgFeEnbyS
2hJClyI2BniaC556fGOUm8pOvXi8DwfOgIOiYrqEummYduC2Uf3ZhcSk8vYue7nN
FK5iLh13GeXQkdpOb6DjzJuN9Dk8neo+umtRgNiY0OFLa9XepPAGvvxp4nUJ1/pD
IC2HdysupY+yDfcornPArdhQUUGqTqXBjnzz/7HvIloVEFkwpOHm8CfHYWW7a4zd
fyWIFZb5cYEj+jznhcrtORAOJXSmFILfimqn8rESeTzZcNakTH0LGN+Zwn6Oc9rj
KZSMSgQfnuNyyQUDVL8+IaHRqQHQI5jxexjHYUGsp9CKbdKmVsL4dw2MuCk17yuC
Ja65KY61TjmYaxAqx+VO1qP33BL5eWBTEfbnaVDUW3l6QpyPL6/Qn35DJAUprKrc
jvbETOlLfrnnplKLVNg+m0wXK0imJvc35DOVX+HDvQXO/nMcW+VhI11VVhcPG+ma
5dpVnMIZ+5VnGBNXJjHuEPu64fNrxR9cdM2bk3+AK4If8QNvKk5kTwRGrTcdhHVC
gffalcI7VeqpzfoxOP2GejkDHwddfvucAXp+7ZRMkKhPCMKYFKlYo7emH0pFYfAI
NJObbQrEHHGcQoyV5yF3Or3JWQApNabEuS5z0UwAr7dIB6znC4dVc/PkMMNu/tzN
75qPOrDrL3oAMnzuAmpiuWxbR4p0b2EE4kitAKEq0tF1ADMWFUzGxThiU0ribWSK
YKbrvGLNYzBZHP00jq7HsqJQT7+Q0yQAmxjuGM6iqc45NDQ6Zh7VaMPUIqoYDb8r
ZdqPi4qvBNKkN90oQmSjvRJ0ttDIgT1qL9tW0DEXXbzXLPMfl9HhONAat1YXtD20
IKaGGqQxvJld9NlKbQIumCGnBkEPP/DxECmiBQqAu+PwfIxpBriizhk64lVgWPBq
3eNJXI+6BmSaBjrVc8F0VHkq3iLHnBeD2lzUyUKoZTQvSdezUgZitv+eKFOHo8zm
jdEuAh8leZ1wfYjdhl5j2xJs8BwWJbGXKrCkECq0mKYVUsNOfMCHHmomosekXVki
CTibrCbOuKgKYg4GYFhrvYjbwI6aJ1r/xqYnMzwp6EXXlnO8l1wrTGTW2f8mf1Vm
OdK+5/TSY11argpGewcSBs9btqsT0dshot2HEKJRGB3CBrUd9Tqpuf0XVmdsiGEj
ZHJU6Nyn3D4GE4vhltii8dP45H3xZHjm0YuLgP6sh9b3nN/BeTACEzR+/XkXgs3M
bVZEt4hqJeNVrDun3pCk6G5IYVMbrRi6zs4PBKLXFWw95atICC3R8+b1yBF3eRPL
x8m00s7vlOvOunr69ptcveeIjor3fkDIVw3iGxnut4USEh+zKr7lJdqE++ugGuB6
M+nr3CohTp5x5dkR3OiLv7QR6/ODF+XRcgECFGPjh2sWbltkeZkG6f1su20scF59
Ie0lpgyGwPdycrYA9nsMCCE5YmnQ8RQBzladw1mqXXtYTP8XlXQ8vw4OlA1OPiql
tnE1eNV3cBY3d/NdT7AF4DgiGXOaNDgRw/z7axfpEKn6aglLxJjjxihXqM4HS4QF
y3Pf7x0uPSYpfKjKSBhk36UQIMQXkadObhyEqJx0Ld4e/c6Py8Y6enlL6tsEUucO
3PIGMVUtsnuMZD5FFV/N+MWzGWmaATxkJPrAl9JG1/bvSpbG/1GI0C9ZrLkSOQSf
726F1ZUCUFedF0vhM8bvO/EZ6GR9oNZio805+cWIgsf7zth4Ul9YOr0/k2M0FFtz
mVFdCjgMArxDOoFqnV7qaF6XZMumuYxgpyOyJCSeD/+hOMY6VA71K09aM099MOPa
/mVdWGV5676fPl5nqY+5xDDfjM06SNccWTMliA7t0MDjjbFRn+gTYB6T7apR0uXi
DIKQERn2/Bpms2LoeNRuMS2yF2bEHRsw53/IjWbFkXDk3kcWM2KElpbh/T1+EQuT
EyTTnr6hq7YDASpJtuDw95jOWqLvjFd7h8wUwn204gBMfjsoO59DWH357WdIuxlL
I6CHQFQkq86kRh/fhZeX0kHYpe12PDCtWxsqAZ41d0M+nIk06pPl4dGFO46in6A0
kDamrY7+h7v1c1CJ7+5CUBtXNyclTEomBRuf2NeY001mWLh/AP/e6qUgmaIH1hD2
ASbgAFTEI223wXLylqusScTb7iSVucS4BODRivty5p5cB7tgB00EQ+uA2G9VSjVn
Toa6xGOBwFcRRiIHmu5YxR3DQd14+jLd831P62g7wxqnWPkWQhD50mf58XOr6vsI
LV9wt3BzKj2mTYciL4F6uPWF00Ee0yC8TNhO68gHYsOPR76c5aMjzDT2P+dN2A5u
`pragma protect end_protected
