// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:49 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NiAPhEfxnZQMRm1bHfQNwP0GycTP9q7Ib83IsrNgDhYHDXqfm87KY2K15dqsXLew
/y65IhFc91r4E4CatqhIZdXr6Ba8aGolxb78xx9vw/6lQhDnd7ZS6fE4gmievnE9
0D/elYc4Vaopp7QDlq0XlnxNQTdg8Gc2CsFzl8iXc94=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7120)
CvGERcWWGQV8SEnwm17bPt69kFRApVi3/16aYdNdk54EpL/ec/Q0yiVuln9RAw9J
t0wS6RM6hg2BYvzQXkvb0PMz+mDN6VvWOp4PP73tOgZSjD76mXD5wdGdDGnGC/ux
3RL2JQVOQEzPFKIGqUDWnynbNrdR+E7tLy5MIZLLJHZr2vcBAA31C7UtodvBSYED
JVrbsGX6Jh7ghR6exTP7mt3ONcCCBydZMUtNzMOcJgXN7HUJLWJaVCKXug3AjImL
gwWkEFY+UUHO+BfZeQg8r5eUIJFY/CBQshMRCFOD2m8ERINCqNJNLvNRye6AyxlP
U7g/+jGw/OQ1Dz+U1Tausv0DS3H8xQbp16Z34qtVKha7fxb+X3dcu/NiXEpOQeX+
6zfgLy+bf94OFaezNcMHEqSi9bp5UWo0TwLlKmQAHadsTcdSh9OrjIZa+4pN8N0f
Q3VPi7Uc47z67tjM77H4IHIediyIQZVU+o5Ec/AOrd+LjGLw/AVOTWRX27cj0Oi5
xCzDp79sfZt61//f7L+/PQ332bbJzg/VZW+86mi+9PqAfszMXw7cYZai395uFWLP
3jnCzH6hDrthzANaOLUeLiD2faS9Ermg2nv8ddawy3uuZX7UJdEKxfvui76Icp+o
51lZ8EMB5gsPIxXw+Sf/EhsMTg64LMVER59nwlz3GlT1S3/Z+CxDcPqkr8CmAhQo
oZcsQulaoryXMoPxobWA/6WCIgjmh19ZFDDQdX6YthIuXOqyzK2AyL+aCy9PQBgK
G9A/W7oixHANQv1FnMYPlJGyzHepK5QGt2zSCnYVtvag14IW01WoU6MsL+TSsLAW
tiTskP0ueXD1WWyjXF3/kdxY9AnHbtgnTUEmgAo8awd+3fQxTFIWkM8VZbYffTE/
nmIKlU0kWULdbha//LOtBuW1FMbgcybQN8oBnRtue7zpB0h97Xa6qL8IoLpUC/W/
eyBCQyP4zFK23qRoxoAsMXS+Bpju2OUwa8U6d6+AN6NP5ilU0CfZH+UY6gNKlxJ8
5/c2WAbh/iE+k2ILl12J+eQb6T1LxE9SWLLbQh68+SKj2+8Sn3g4yR/MAqBh4CRT
SHZGtP6hpV6Dt0BYkfSDWrVLS7/5wIWHx6vae60bz90tIZzPmfo60aPDjrszpkcJ
EhpuGT5FWGcL6IGouKRtU190EzKRA4WSFuwbU2VwWN1wuSdKuZbksrLeY/d7V+Xf
t7/HL6XJSKl6kGhrEHtBm0gdVfAqkQJUYVJ6IVyUkzgmnLFWBiZbtgJXWJsQETwG
9m4h71HmvV2uGO1/JKS2cO6nOVixw1rrlETBXQdrnlTtHgXDocdiCCiCMWKOfWus
METJBrz1LcDS5loqQrlj9uQda47HA85fNQszIshlI6kIKQS9l4kIkYiQMTmFErQq
rmzOYJh9YriI8NmTHE46JNQXYIbW/SuAj0whJcWKlwa5df1R5ZTr32qahdoZlvuf
N7EvtWRVg+lI1m2c9eI3iQqcPY8HwXQHRKst6iAknKHPBLr96TMenTR8a82Sfknx
HZ6mcK290Me23aFFrttMBbRAXBfRPP9vuGWBNTYgwfqR7+lII1l0coRaDnVQZG7C
g0KY7QlOTtY5a1GGg7IoHxix8/ghX1iLxmyyyybo2h8qRPnPULZRFIfGzIkq06rW
sTk8EHeToKzc+5vUT5up8Srtff4ib49JXmMfZZ+HyGgg+sZ1ezNQPt1Awit5FLkt
cwxvcABfJd1YJ2p9578b24s9S6l3PyR14T1uN/brBXfLXDkXNKD4vSu1bQmKu8+O
sbJEMWuEqsF8QrJiOnmagXKAyLBTvxYWirWr3TM1tUqbMzkwC18h00j4CITOV2Fh
n8Y2fkCONtFri39zrYCWLvwY68cVnOpPJSVPEsozc73K2+1SYYsXULzFjuP//5RA
ce9kV8wa4/RG4/bSUi94NoV3PqjxrpSJmaN2QHqVPO3KlgRVWQ0Y7evWX3BVEmZ2
g/FqCgXF8q05QEEB1y/1LIsEPqp9sj+amBPVCG5S05j/UdYOYwFJ7XPEPztXrSvN
6cONrEKgKIwG9eWLfgQ59vJfTb7vF7QbTl6k/YE8bbCfVbEVTaujuMAB6XucPGYT
z9GKC3aMG/f7qm9gA1WWhxnGEb804prlFPYijmPP0xRFWOCtCWqyhKNd+yaB+T3B
B9ACZXywedcXZzJ5Jmds+3tHtDZgv21hDUlu45DcN6JtHipQaFhJzNARjXVPultW
hSyaMkDzUEvgJ/6VdS/QuOurQ5kkcFJbMMZAHSRIlfOrSKNO6zibeNEvwirzc7uZ
LkV6tSAEH/WNqYnCziSaeb4mUc8IXvqZ9Ttj+MmBQ/zAW/Vhf4zV0HMXFwshFcFf
/MHNyS2joyPT+xN6ygL60fQQbvcqVztjEbVpMwvmSGuxQN+8zFTO3TheETQQIoCY
5UB6k/mmtR+DoquwZfVybxVtw8fS5v4OtcCFqnKOQZ9pjZVPdsbgHGb7AhcChq9Q
YNT6Zw5D0w8zy6Ea+NsEFiF37L3kAxIlame8PCAQWu6SGcRF9WJj6b/9twKh/Pic
tFXvaM+GCX3MU5OYGAxJ2L/rsmDay0Tiw+5/Y+pNG1rqg1IFGS83sCM6W+nFSLKm
8eowgDCU4m7ZBOVdcKL7maHXUnxCRg07/0YFMyPW4Ht0SeU1GoLA10z4Z1uy4E8l
LXnpWXFJ51eTw+mxTBI/ZsN9xCzS/cnpexXfrEmkE5m9Cuv/mafjoKCM/AVMbqsM
JSMXIJBciRehsZIFpwz6xwFsImF9XlLwQToe9IUjICAvrSMljcJKTVZ200sYMbNA
PMGVJAX4T1py3cRfabZwClJGWySeEpQn5SZp4VkTNAGnjiIXQDI+g3U2LtE3DBYf
ZnqcHTembs+/Tn69508pYJNX+fwZyVQ528iIGo0sL7idiAQtUsdIEryWmy5ZYQ8d
KwXRFTqE8bsTjvxpz6EI9G0HOEV9++sYz+AJdAYoessMrKyVaPwM+2lCUQwCOsCn
RCvmc04gzUUAaO9HKlNbLM6waXhZ8qmDGAAUhzLYFAdh9d3ssgod+aOFJzmBrNjn
tIl4tl8sFFBbXErNh/wX0E5+BWW7iVwMnlhsN3umIpj3P8kuZh0yOmef6FYhZcEA
YA/Hn1PEwIwDmP+Td94ny08ViwKKsYvYORypXVSLYTb3HTH2ZobfgBfVXKV0ufvB
8WRkcPeeUy02I++ANXQZ/O0gDiB5y/15GBBKJ9JpKa06hHP/RJZJ+mb1tpzQLYgA
NmDXYL5XmcHlQXycntZrVlwReJ2KkGxeIsRsv0Y/kGJf/GfXQjpilzDl2wMMlQM5
zLIADvBOuVeuFfoPZ1+K+3YgisrN2Vaby4HDe0i9rHwI2cRkfVS2dDCj9uBnsusV
X5+9xJUEFug3nUrXu5QJ6iEr/eI9TTm5YsWn+InczFFBbhKIa359lu4FIe6TLJN3
cpBUZt0YPnPwQQ/cIZYGo4gO2m2asP0NNd16MaBerHZcjRmqeNTuzAkiimE3IQMi
hml+zyBPXvQchJUetUXv7X9oEMSm3U9V3/TIZP0Uxhf1Ha2L7tP+XZwugWT+TE8q
NxlzqENuOnFgItUnGmo232ERvx2OEgxGkTNL+kLv47ofNFP/SsFk6UGDvASdNjVJ
nxSrEX8uSBY+43/YiCWmVbeaavir4OmR0CGgVv5XiBEvRX/vFEYQMAbB/HGXqx9L
n+tiEM8YrkhxHLOO2dI1sLisudl9Gzgvl+ydFkQy1aDTJQsQZOvC8/C/W6Z3eNmD
job/2F0WJZZVwvfAKWHALYEdA8OCplqsnAUlkn67//irmzRo0oe+txPoVf1SlHMg
pU3BhbChk2M2QfAqAThOrR1D2UFOOws5dc03GWLmMH7fw/fh4ax75mmNzgZQgcVK
zhwMmWREXmWXci29vNqZo3Hi69yvyW5jfBr6vUUcrY3RHBgzuAmVw22+yQrHGvKM
q8QidAZbN/FLpA7HiT9+6Fyrbg34l231iMtXy7zp6PIUsLfyyMNBFq+Yk4ihn/dY
GCCp/v0KA1hPpYjT1ANa6qTAPuBt+4d393CoOCWQtSgbNVSj8hwWHFGCPA8XvRBj
OhmC2UYnbVKAdSkmu1K4jZE/LFGzzQPrewuDHOYSzE/CmmiE1ZB6LYfFw8/w9zwQ
kSERQOBmVbE+oHONu/agC0imHsJiFZ1Gr5LITCMEf3JvnSyKPcGZlME7GlH+Yr7a
wcn4IUanNCe2PoTb16aFU3fO1F/R1ulTMASjBn2mhhu7eKPain8L8riJpnNb59x4
WUDsf4+N0eCVZVQRYmd65BUov2lpbpWrIvb+4g2aS4gjfL3G7UMnHOlEGo6Em2Uc
EUkDJCwNt1FkERHgIBje7s05trbqNf/tkTyD5ZL1gavXCyitRQ+2uuss/qaxGoj4
mj0zHJpiihj1XEvSg4MGAsUQGSUO9bldq2CbDpHmaCavy1VvK6YUjwL+Ya1/kPrU
MtBb8DuFSN+zISJfYnYKkYYVvEde1zYjfRQR9hJMP+bfHMfuBQKkXusqRTz1ELgA
UTwvOtmExk0i3EoaWPglUd0iozYcSorcpIPIjD1kfVNrlhDo05Ve+DwcDQ8bJPoK
U2lBTgbjp5AiuzjR9Rl67Y2WdryBhhktmCweIMZkVrgqdDohvH0Fy0wfz7LznsW3
+UXGfnl+ICsfqjJJ29NMdWKuiV3wvA6zTpokSBzmOZTxz1EmGNtJK2rb8l4SQMj9
vs9KnWk+f2najrwvGdUfs09SO4CbvHLgLwS8lP1IBwNzM36obVKSW6Y0WtQ82Crc
fndHcEFd/8N8MThv16eQ4JImbEvQj1IeVWyzjAZcTIPSgoCf7H8H2hbFNmStJ1dB
M/PFKMAQSnITUygNwbJ/Jxi5DdON+7JEtw5h85uXlwpWmDVambOBefR0x5fstEP4
n+KytMnzDnIa5UuP79xgI1ARQLjrwxU1BHsS/uh/FA/0Ltp068iJTPOCCWVX3LUS
7zqztJDsBea1jJ2XzFZG72F7MB0VoVcAELfXhVunMD0C/yTeMiBh18Va7zfLpqt8
XjWDiZLMLxiC8ZvO+wFZ3nWuljNliYIF6ydf3xtmjInPWG6a1bnF+mTHpvILEQkJ
Dj7NBvaO3Zz3gDOVcLn50pWnFPQ4KPbgCvaV2NCjTuNK8cGGjoR6qoWVuKgLnyEU
9igqzH4rQWtSNRTwZH5IarSVmhc4B0SPSl8BjY02HN0+lSPolqtBhcsN+Ljj5Vze
kGAbwyZ0J5Z0M0I+T5lYGzljhZGk1oQflVWRlRoKqhK2RIjQzDNjG07lNbhQKjSS
2CFSL9d+H2cg0t4yLjlSie/iZfeW0kjIhLa3msJnhHYs31r/pbY65pA6cuWX2rbX
vFSA1ro3aa+CGMaZ4xlH7OyKXzAxsCwVS2EY6GVtUSKAiC6pEvgeEyOeUxiZm+oE
mlPYR9UDUmmtHse2aIUs5fHbMJobVoYOIdHWXnoG/YM7R5p7uu+V1huqVLl2b5U7
8hD36/+blZnQQ2GzxKCJwGMvX05+GV2nzNvxG+50NEwnLVA+pRPRqy1+QcIKj84Z
R0G+yM5pQTrcmfrtaJSGDdDMtInasvxQuaoSAQkZKQZTZ1eLUiLbT1288Rv2PyOG
XSVnZkKK/gdtXoOSMn35sSKkawGr52YenMFsqGqX9g65/wg8NX+BVtM3bunmU0ED
Ov5G7IF7gpU+HiqYLgvNktY8xvuIS+BMyJUi3v2N9pfAoOBYN8oJRUBOcgySd+dv
qgiNQ3QiMzSJm3RHbbcPOiGAIHekJEH0bw9vkE3kN1mlHOgRkQf1OForJcaP0D7s
+tmaLgQJbGAoJJJ9Jn+huQb20n2wKD2taYDZtr2M9Dyuf6AY6QACjFEEQDWI8l9b
lDa4E+tSKw3mzcD3tyHDTjRFF3SU2SSVqO2hlX0Dfa4vxoyJXNh+NErG5OoOeQXA
oHEKjCkXpce6tMeikf39hf23gOtVm1gkoycYHLhmSWu2vr3fvYxs2x8z+bpda6Rt
Mku39UIQ+hS+Hh+sH0n25oWGu338Yor5cihSLH148hl2UroD0gt/jr7AD4Z+/43I
wSuN2RqyptX1ZDqjFgrwsQNmp1WYJSHAgzU6B7adSMwAyx6DkHu2oLkYcslPeYIY
WSxOJI9uMq3DymdfC4IHAoblSh1KC6koW9XnpNHxjvxn3/v1W55twS8vkbELa7Hk
lcKoTYBC1v+Z45bBdCajL6g5lc6E2bLFyuYPmqHP9BS6/CPFNEpzISJXkmHkINHy
rayY0jU9nHOxGqlNc7IEK3JtV4Cd4zc0Tb0L16sh5S84CddnSCusXINktXTMJWfk
9+tK7pWGlLthtQFmgv6X7u2D0vdVdDSexfqch2xBx0pP+t0SbQXXMlfqtetLJlA6
jpzpQnE1vrK0jqd/SQMXomrfffjV1sWKwPer11mugkYcq3V5ECMfqHWksmD8lHfa
zkQBRPwQSGdLYKfCENLPs4qVuPX377d5XTwNV2tGtzcuvyAHDm0ahyRUkZOX9ZEG
Pzuv8KNTh0NnNvEU/GlGu3M6My9ngqunEgf7rIuLDGPK0+Vyox+H/ENBUm17frTR
tdyQDytDPpTyj7u2EUwr6PJ98qfRv4ChTDP7lGzgdg1d5NzFCcjGZ+Vi0zOv+y6A
pUT0ykMtahU/qqbTUzx9cF6yQ5tXbhUw4pycFMNOD08O6IP1GZ8mWqfSD7mFtN+w
GKUu7wxJdRMwvmaHnwgl+cjlkyz/BFi1WcCRwQ4CbkhsrraLIZ402ksDtLYz1WxJ
nCaLpSqwd72j04fWRXQwV8b2FpWrkVNNkSrJ8jbc57+ZsFUV7D+LZnGfKzTzkeyX
0TlhzRlDYy1+35mbTrLW47Awf3pK8O6paX3J/fKb4CF+1TIkdXItwp0u5acGu0Nz
xNGuIDcbnbmaIfqaYol9Bb06OYvqWZxoOi+7OWUEU4NyqSneB0M4xD71/nnynO7F
0EH8iV4twSOwAvKTpfTpeTkkWy8/+RgAozs4ErmbchHbhGnecK0YqX08RMGtK5Sj
1j/n2+nNV6HsHZuqvtPn8dfWnAebX8fxM8uUq5uBIGD4e7hE1kpWEI0VgbHDHOnp
QgzTaq70mmOBIYIwf3wPP8j4CwyjhSjyNbrQQKKSmdii3Mqvh3nS7bB6b7lvlBWr
Q+uPeZo+YwV8IiljWvwk/RXyrZEEagNUTUgX0GTSaULL/rtKRDvlUVwqEiLUh4Fo
muMUSnAUO7toH3HMtTxyG872JNwT0NWuEo0bZqaaORTak9TEMoiwKNRzkm8Rn8wH
8uvbnG+mhh534FjH6lqt00KsGCif3tJ5ZjWhS4SRPYLIJsrq9PRvGyTfuejwAEqU
6ejGkuwwKaOamHfxH37eSG5khW6rCubYApo691pOFkZYjB1rFLcC+A8JpWvUD92k
RDX7Lka3fsbmNG8KGNTmAenkDqWGHOtszaiTz/cW6c4FFubFnJ0udWdsWKvJRswL
83xc9ApUPkHvCL+qAbDZ4K+Nt8Fdor4EyaAtNpaGm9cDLYiqHSE3LUFShaeMFyi3
qfKuoDEzHBzPeUQuUofiDPSjeUpXXUzUNUTSqAFi1wVRsPTRi8eQi22NjWHr2Nqn
kt+wETt8oKyT/blBQ+mY2ZrCeG2vZi1EhEETo4qMTh16AXbGkxHwIvNhBj44f3fM
nH0I/x/BXLt5kZnrDmTbCOH1sqhwjPlX8k6gnJ1HnBqr3FKGbj81KIicR66Ry6S/
9J9DC78mCfNmkjSjW0HvZJ9fozmPLuStvk8m2Z0RBmRY40bSxoTegQDMcuaI1q/s
olf80GJVNMo9oUXpcB1L9PhV1pLHsjZgVobvBe7n0VLjavcp//6JPLfur7DSyQfS
GmVVWmU0Ygus8K0+YoPamCsdmLkWHZ8UlAG24sZ4mPDQTWCm076933awvzSd4JXo
MHzYyqcwIN5qlrKEAmdMS5uknfi0D1DbrQnsuVOe2EXj38OBu2/G6t2cPJpvtZUq
h+L0+r/FggDzXllETJ9RS6PgI0T1/YycZRfCtsMeyj/hZGCKw8+eF0XNPW+E0Pq1
rC8uO7aDDIDXaVQO49Hy1SyuMQOMzu/9tICjX64eoE6xAYvXbbNiNkXbh5Nlinx2
ue9GLvVnRBaUiTrqTjq55ikKNCyIueUb0Jl5uMWcXK1P6bzMG0V3W0Iso1LOlLT6
TQ0VeiKQrPzqZ+vJ/memldICip0CdkYa4qVpp3tbii+1k/gwNYiS2aJ7QcABMAN5
682My/sZXPPm1QPzpr0/PUCamyt3IQtcNxM3FgIbh2InOWTr8YsIY6gAl4rCjtKe
f/zLULp6ulugYqXOUITCslu+GBTgPorWjZwIjUveSCUQA9gJuWQbQeMYauP2ZBTB
4FDoe6jtKckZLvpzX8hgx+7MiBBswFXwqkOGQoCU1qJQhb3tkupr2mnJP46ope62
Mw88COv5oSyNdkY81Z6SS+CnyfOW4VI6gTeRH4Dm/iTbDB2lPzAHhuS7sEZHeCdI
kpP4hqAHo1gRUGm80eFMhLhrGjomsxVFDuXwGsF9fYpui4nVJnrZDr/NKiB11VEH
n2DFFHzO3Eo1RruStnHhE/F2qzeJ2oVwnIna4ZvnDCH+50iMAx8F5NLF1EmujhFM
H+G5A/gliUEgkkt1qRC0DKAOpMrkG7GeHDgfdsTsPAaAAOJ4afRhZdaZ6vMAu3vm
fyar+iiGrfw6QZs5MjK07nbPFr1qjwaTa1sm6as9gPbmyX7wDtzcw7Cphs0xg4h/
L7Hdjo8jcxTg0gleRWXaQx4lp1YPzZyDUffOkGagydBtaYPYMf8kvjH09+Yb0flp
OqzNn/ZKm3H6nIfkehrhLjFN1mRhmleRL2tXB/Fsaa5fzIGqWU7ZsvOoj1swbbpE
svMh+DSdWGXVsmQqSLRlvbryIZOf2BJnYxJXVsPB13sed0mZJhWI5uyGx8s/B5KL
NvCrMmw7ECbTuMNydnDfKT1JRBtW5LahYrDuskinn0Fb7rREJWx5wY7liFQ8gZbz
j2u3axzzKGw5hklTD87ggLNY4saYHkkixTTQ0Xklkj/1DLD8KL3nsegTQkCGvimE
INWI8GYsiEbQ2EUR4XKd36plqGWU0ZnVLwltS4y4ABZN+y+v3o2+jyqwHtkDdtnA
sET+rMxmCIwB2vr7NK8hjQlKnmHhykQjAPZwKi0PqwR464F9GIbi2EeWsbnS6dWF
ueNklv6zyBHR0sbyQIzrthdtixrAE3WWPoivrEwNlFaS3x8BT190D0IpsAZFy8LB
ci86sH8DJpGO25wUu4JfjTE3uZCyIGvckAszlJyPV3gDhryv0KnNJqkNvevfwdwS
jfTRVP44FDAB3zC5ZYi2iLgaBOjVaje4FxPp3ayl6IAAbrqNqqV4rL5rMp0C2B84
fyck8E9LDcubaS9bmqAI3joEx/8YDVssoyGSLDbLpZIA5MyXobrzDy/n39bEkKsK
llgzPIm6HnEgqqXXNnw1SA==
`pragma protect end_protected
