// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:40 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N+ARLTMMwQDYjWnHh9+psvrrzQx/lrZOaV1UlGKs0EOZxgbW7Y+J4ABRxyBLjs61
Im54mCExubw7U0FbFb3u3qxY6GwJkvoVRKfdVkBw1Q2QXMLkBVzOZqrNSBTknLEI
WCcn53l0HN4fu81w9eNmWNCq1ekb/2KlV5Iweiwa2ME=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19184)
lIW9YVC8qgciqyEh5HpRI0ijh4+sw/NGiUW4h9s1zr7ULJiUHNtXuPwoUPl7j9gG
IdJhZusdgtE+XLucu71Wk8DibTn93yNxqRz4crA/f4dojYZdNdeEQxhkJH4LzGpg
1h0J+znsvJMZ2WpNBKtx9Z35eBV2dt2HdgMuGlXyFYluVsH+bTYz1PIgAJPNsRBQ
iTZxlCiSxl5zySSXnln5L+2aD5GqA+VMVAMK50H6xdoosvqbaIJzNNvu6tiBM/WD
XQcOI/+pO9DrJM57TokQ5LB8t8kYOBIo0Dt+4ACONxrZmfqftxwXcsn7cb888WCn
ougpo61omaYekI+mMnga8uN88GgOzwAEOV6M6/fGDjABJQqEewPJ4XOCU+VihmNh
Sm+xDWTAWj6G7gCu4Go68N+NIlSit54hEe3aPmuwel/OmsP5XcCZeDE9yiwfbmDA
x/N57XvaBk4e7KWMz9PLD7MjClO0o18OBPiFMcVblY9V9sgIPixPh4ejfEMDKw/m
SY/BsGQQrkR3aaVJoCk/hJfua5SyoBudhykwuloDQNh2ulZvzD6UqR864RE6G2Sq
fEROEuyQNdP8Zs3Qik0yTMxvbKvYMnR7GGl00xLIWv0R2ptz5cNXTxE7NGNEIEtH
GryLrNW58y5bTdA6nScdLuPc+Od5DcQ2cPxyfbBLumoSIwpYtow/H2ulmoFfRaHP
VLFzctKbT4xUo22N22zlxt0qpRqbcnzZNIm1LyonaQFUtkQnFUoPxlEmFh088BFI
ICnzFbemHoA8qJDRNOinaKrxarzHl/WsieCm3qRDR6of5idoPu1dXNLYeWeH4+Oz
eC+exx7eGrvnCFjOByC84WSHdLASYDGrDZcmw+yrEfBsRpvTl9o7XatkpTj0IZGL
EtvNStWzkpavtIpksPDvcIaQ+JzUjluWemGjlPQSxqssuttOEZJmD0wdGJFvaIw9
khzEgFeFrovU13fl5MZL5TvuL7i7uxmmxYZpY9W2gTTKzVfRNAvONsnHJ6W3K5YN
+4oN8ZpqTX7lr72kYdumVhvXY5FamZpWsF5qUnZAcC5t9BSletxTMpWzOOd4q7Ok
d5fXdL1PePxGIejGtL9w8vGdbXZN9k7YAqDZdn4giNViZufcfMnfcYMQUQfR4Lt2
Ahi8ErjoqFkt7XD9RHYO7eQ8V4a2mihONO5anS47egbYP9pGoZiwzYaiKSBced6j
24ZuVIaayVUIErYOGvEjYrY8AHg0sijFfEE2mjiUzJbC3AT7ECBqL7EWYOnpVm0y
GTMdUULsyu/70F1Cdk+0tS8ffmnyXUr1e0fElLXHcnKlfoP6xod5FZSHZ+dykKR+
p72AQGHOyZxs72w4TTa3UeOkN5pt3w41cZc7/xQoDVjpPPE2SQ34clg9ZBf3+1jb
0CtHhQa4iApFvX1ohTNc/sPdNSWiKd7RaFiqqVpYA814eH8fry2FApg/py43ti+x
r8mdPo2Pfam8mQ+qpsOwzw/3C+mhDXTJGJO8PEfYU+bIqj9/rkU3qXohH8vyXU40
sfq9c/JqwqAytGI/wD5wawXw0SmG0ZPWDHZtslPWuWfOrhBYZ/1LyR8lNclWirbY
c3igrIuvp0x1byl99ZPcGUJLtbHuVlVzq9wLT+hTnuhkZjMNPeNGz9gRoltMRSkz
tXQRut51m7cMtyNgt2zgafTnU1yeieuhoMINmPlvabLAGXxi6bSfncTZUzVHBdA3
652F1DUskl6hRpdo45ACPNgjQDcVMxveKeNK7PhvoS0x980I2lM5ioMajW7aXDFc
WR+noicpi+saDztqP3he4hQtgyMS7y0G57tVCrPhjNOyNwwsLFVbKRO3FScKUtu5
MPpCK400gyuN32zrp21ZmjVFIuHDJ7qVR9HQvimZLdSOiP127G+V8Wb1an9wPhuD
fhlAiF/Q+2/TD5ca1W+Th6Zvf7FdVILfpEBMI5WWAYKtCq2vPYh48f2+xmFHhuF+
RZgHXQBqtaeDwvMMuRVRTyhLHKzH3ep2mkQxhBlYfuKhozTHHCaeV+MJENivyVMH
W4S12QDrataXwpA2TKGToYTVTNa6uRGw7m8eAAKi0xB3Zp/yY/o9bLcykXBl9QpX
1nh07dZP9NhJ6lr1Uzixz3WtHuqoj51XSvKs7sg4bakvNOCELF2D9bjswAoTG0eJ
i2I5l4RuKMpXBL2HVgU9a24NbeU21CqWprkvr+uzz150K44NbZof9KSBhDckxibM
q6YHjDUz9OwXlypTX2LJoCxwPgtRko7IY2rX3qeaSxmpbR1+Lk8Z6bRWh6THini7
tCTI/BeYvJknyZH5aam+Un3mFX24gfPnVHrpUZ+KOKZvij3EQIETb/OJvdleSCkN
fH6Nxc5gJ1DeMaXJqXpggw2SSG82BXToBQKgbMCCzVRhckAgcu/zCBqt8/10vdJc
XrI4BM64Lwsnc1bOHPJf1d0960VtkY0fSqv+FlmkK/2Oplw1438HWc+I5xuY36hx
FF+LF8AR1Mdi/QvVfrQhAHiJzojYYmg5pmksGz9olvELreTU77AjvRrNTAMr3+8e
YhW8nr3I3C/MFnngyy3zyeBhwYUhYTRuNZVrIKh+pdzCB1so73KH1VJSihgMATxq
YGZmy0Ig+GfN8ITYYs/1e1GHcva9OuSXqnaNywtYJ2iWBRRlFsvnEu/ksWQSbbWg
gQedUlFhLCkePCrvWQdefRlaA9kyp9iY8FxbHSAkoyzjduNNrVXlLfbpQ2fV4273
5L1DU1CiB+DIOD/HjbHifBZMedGEYzsUbvkg0b9rKcsKnA+ZoZa3HHgjA6EYGbMz
2Wg0RgMytMWYWu1W+zyh9NSl7VcijlkcTffOq/9+vb3Ru6ytFuN69RbP9BCIF5fy
hw5uGweQvA4VNs5Z/kwKr3Mr008N27Ap3gbNJE2z+rrzNcbeUGraEoivZJFCZunO
TAcV6hVzOC3Fqz8RKG6ZcwsNLariuHrE7Y2Mj68kFfM+S7rDds8GSIcdQ6p7u/3F
3vUTLvvhD8izWDTUMN8E1nqtZh+6/fh3dvZb8bKjBVDB+Bz089xojhmOF1U1HD6Q
KtzhGdypnLA7UmDVJ5LqhpcWvEfQfLKzDG9wpO8kSg8ungyq2mZ8+gPi7oHLQgqJ
6CJVBnF4cVF2p+xk0nCbdxYsJgZ5q9HX+fr9dtAIagWat0hkPArZ7IMqoZPnbXsz
1lUNanAksPM938oaH0pudWNOhKEQpxpUalN8MPC9NYmKOPtGepyxd4yhS8Xphykm
MMJpzeu2lu5OEQXq4rvi7fQJJflSetLV34ihX0KGGxLewZgdGNAUuHZ8SZyUt6cz
x7K+CSJNF3FFobTzM2sFFI8APDIZ/5HeANRsLHy5HTM7crrjYoU5F4cb/egvX0vQ
Bz56DulxgTsKsIz5l/GSuw+xqTHhKGgMeNJ6WicomM9bwY3jwCYqNmjif+XEjxeb
ME/ttteUjxYInEbCASmILCc2EyTV22kNEA0F8WaEbrIsgIjly/ryZI6kgusw2zh8
AZiNkx4OJWifEMXVja+gvU4S13oib9LWOlkwydzSbtC8BtkpBlh/C/hlmUaHjJxC
STKfAYpWlCk/1xf36d7s6cJ4t9+SQKxe4EuVAahbGe57g83xF8sif32AUIKBtjFx
w5zwd5TyZFqhsn1nmfzGHNkOAh6zu845GP2KUnBbcNNpH4wIPjjtVek0KzJXnSwg
D8lnwfbU7R3uay5R11b6FTjm3+zopHOoxpwqx3+QAhMVgai+UCJQxMskeyhTl9pr
KfShZCbLCmQm16FP5MKcpqzab3RlLGG0mTI1ZwFFYk+jZxROXiG/QW5xAH+UunyW
ApC4eZwJFqSCmmOJ4ODDtR83nAqaEgCW3CuYOjbzk4myaLt86/OjxH1avuwwRF7z
Lt3f/dzjJNW2mML6lC1Msqj1UP+Ry926VzNTgG+pds6QUAGJBi3gyi+2n+jTUWGI
pztfyj/1qOPrT8MxwP2sW97fneUoZ0pmUUf5VNUqknXWDMep3Ta0QuvPCQI6/7GI
BiSmm5YAbOIcF3NQkPku8Sy7YLxE8/4i5iuhj06BssLtBdfFtViiGULVd5RHtSk1
+L+Hthn2XKh+WtX6B50fz/N9Hlu5V2wZumAPGU4t9X1g+vetwIp3pSzH1VmNXLVd
LKy70j3XvUnQq8Jw2SIgfbqP/rkYe8QOSt9nXlKMTlKXhIOyFkRDzkIIRnpVYthu
YB31/SQZJp42WhPTLaiS6kFLEjfBht8vp9qQK26xVBRc5QANCE0m8x4d6PQ+FkZm
ON82UfDsa/obDmyzTklMrUHVs7MFBhCpEFGs3JkntMBQId5Qzf8kvx7Zoof6RYcq
N9yqOczhbdcxiKjPP8RRIhYa51w9aKHHro/FPpQ4RKe8BWWiJFi6CtQ4Sc/CQJqe
zAynHBLTXnsSmCaWsVaAZImDBXkelc7IpdLZAplyN7U6dRxErLWyigCw0W7TId2V
euUrGP2FlI3vJotfF8utKnR8YknrOlHLxabIx1xtE+lzNotReZy5FL5e0WJOP9yi
YLYzRKr8pChaSBY3gtHsmizQ4Do/ztcbkGFUrhj/e/clXuGhsdM7aZ/+Rnz+uBAs
Fy8QDrl3Ao9/5O5wCwzwqM7CM+bqjom/8/izJstOdHDPKjZV26DA9jFgHr5UDDX7
sJBRfi+jklY/vvmwzbOW2mGjbG4/p0n5Y0YWTmYokEO1xqfZI4+lBGKGM3laZhL7
wfcdDf6BNlnttnsHiihe1zNpj97Alq3BgMykPQRFyIQUJhd6/l0aXk1lS6xpLBHi
t7ijjFoDq3GWsVpsnyswYTfKU8QtNSwIZt5rE47XLCUT4xahOccSMGtOq9VfckVj
CtzeYIKmLKiwziKurZM6TYPEtUoD5jyqyWUnMmO9J1ynTfL6Vb6+1vnkhXs28mjv
tzTmBDpaDQpVVIQ05HiPfws4djxPqKbxWHq7x2g15jVhpNKLBN1Yl9gK96wqoDaB
x1aQD7w86mWbNFjDpr6BTstcwxDrvxOF5VHoQudOm5zAByR+DYl4Q3+wnt5OVkgr
qoU283WOsVXysgeBqIgZTZdvII8OaozOd5rJQfpQu5iva2vBaDySD43Ax+E6eMAW
G5alKfrk4u7GfaV/4FxBXjAXaqI6PdzroFjTfRoJeP3DtoN6Lx6HrZgJG/OsQhXl
niQOUlXc+/QoJIpHzn77Krf+vkQ/RxEyIR0jo5BDPUNPTCDo1wQK8CPz6vndkqFU
TmxQriv7OmfZfzjU6+L05rAFhCref86yAeLoyFT5532LnOZTigzL4M5BPs7l5C0I
GJLQvdMr6dKtgW1QYtrjVSTE/rkLthF7dzjpEQ4mNDoIDSzJqnWdhweWVjIaTwCW
zkrKI/LMKKG81Ecj5FX50ykrquQoI/PNjl6DuTBXRgF0M7ZXuHWLGnQdgQNONWhC
fcgeSMNsIU8cK+UOYFqR37HpWrw7GARS3W0zxC/K8YBJ+g01k3rCsFFRDfn5Ztpo
AOJz9vjlRTaUFEDl2A1kwLcHv6y6qtJimdIX+EQZ/RRtMRrDdaOPrRzyPqsdYJIP
0lcDK2QdY5cmrLNZjmXmj1+VUAmRrifWzLxth76DYFPVkzmyVq6iooHMuzXuClfx
WlVKdSRmw+f+mM/THAP7hDOrCh+Em7hd2m/SJxZ5aXny05r3O2katvUOw4YrL+sT
4ma1KGl1eTo05eDeDazp3ZfcZTQZOuno9FTlhtG85nkHL7dbN3N69y4biMmQNDpU
c7TtC2hJkRZ5WGhDJSC2oiomiIdo+xK9ac2+ofvFpuxBJ4rZPeJgR7YUC22czH4Y
s/FWuRfJvpQHAQs/k1n5id/4gupTztipPxYcy6hcFL+cJm8kqoCA60qMMenV0+By
c78jozIjtZaF6rzJy3R76jUKfeM9C3Bdu7hrT1ril3o7qudHCtmUOFNYy6QoPlpi
53dQMMfLkupk7vLVGGI7oXwNzHdIA7m1Gp9TMzPbncbpJ12WSl3VP7cWY/Af59pR
UUhWDeErAYhZ2vvLwH2Rs/sf6JlY9dBBdFpHkOSE8ZRuL1+ZYcPUhD6fzgkvbaeG
v33BcNTeeT3/GwR7NkVRt3fxUZ3W7mOVOR58ehXCTvlcUHIinYq/8mtsPcUorqkj
+MVm+50ZzByBQVgzUGEA+kfBVbMu8whKnFRRJVya8y/u530m0hwfStn6ugjHIbv1
jx3D+6qCPCYQ7nGdy0T526RlP/i4TuEay0CZcjWqXYPEzUWWVtCVSeUQ1cL9xlbj
R8PADD2lo6lTMrOxLWOhNjeKbfYdWQdxWTnR8MH+h1ssM2jN7OQJN7L0rdXj+1+H
UVAMbzZi+KNmsOGJLX1705+gbsGrpYE7KI0ewDjVE+pYDl3vlocvsot9YJte3z8m
PTkO4jUAUo3gZsRn7G2Yv9sYcmh7dGvggtP1kIcvzKhkUhWI4yfLvt8Pz5RTIl1N
ThVNjrn767Yow688czvsj0cZXyW4sdlCtBnB/b0WHo6kJr1XM3dXWhtYFDqeCg2F
GYjPTZDd3GF1WpQIfLpwg8FNgp31DU3FKOzJ0JkCavoyHNbRToLXcwUMK1DlUeyP
zPDDEAWdYFDF11t1dfmeojXFFr/Iud5+dR15XN7oDd7raJPkAYyb3rXBPWniYaL+
kztIdEg23aj/LwEkzifT6W5i4r4xINBCEm2cjkzg5VMNWW625hQTi8StBmFONVzC
qpO8CVfdP+hEJu//t1UJQ123Ln9erVrxz2aKQYiKaCJ1ByrQ9ydza/m3/oIDCqGs
f2VmnUX74x/Rhz1SZznZVD1uuwGj8Y7p6Hj1bW/XWMs7VVIq4Nqz6cZ+32EhHy/w
wEulPBojHr5csD7l8wAd+L/M2m5WQPt8R2yR+XwNZC4Yct7dOaC7VBE8Jk4OZGKT
7joZvKQzMfSFHU8jN6566eSRVMNciBtcTnAY6oEBCvYNcBLlNyWPPmDujuj8ya/M
hk77KpfpIGx6jQygEYd0wujbUUC0Lb06PBmhKPXVAwsgPNyMGXhkxxKrmRZcddRs
fQV0RL6ikReFOYD9M77uw6shipgo0bRNU7yH5uquS5+GKxaNw4nW6Hthk/wNrtbZ
ORjoHG4TqIIqp6uOY5M2R9/11JtAT4ItNRNNBDVkHC0pc4uRZtPJe9TYmAGicDJJ
pslX1l5/mMusDgLefaSmdoVuVEfMUqM5/t7C9awsY3hg2duSiq4HArulMcayFQE+
YZGKkzp/9gf9k6+AHU5V1JRWkKGANR+1RD5b0d+GkBNoj0bAKesb4gmQvRROFLGu
NzIh6VsiljzG/VyPmfCSAU2PnCW5R6fXlMD9vFvyKsSIAikULhYrkrhlAKoA9EzO
2FgiWWGtbN2M0/6yvGEBVk4Qfxa/vME+NWXvELAiEJeHjsJzbG84AqzjrKRe8gpq
6PHZx2l1tf5JJgw1BYtF8gADFvTqiS6sF2gmxT4xlHXRk7cUUZBW59AudRCYozb0
jItWT9UQgntUdbgZis62ZOROrJyePAG5TOf5alKUIBZy1UhIQuVDnJv3ii3FWbn8
Etk+MiqP+ypz0gIHL5wBYP6VTHK9NXRjP7Z2FvGSwwmb3LjVNFJPChZ5qk5g8SvI
UQ+aNEcfe3f0zpqNkw0w46+Kj3WIbYUTzpnW/tzs9y6ZbhGHGRe2YEFz4h5AO4Ku
a5aIUHkZviRAUItSjJRLR4zWuj4V9aXNgprAHMvK2WFXyPP/9S1j8O2CMFdd5219
Tr1uOn80TJKoRN/rDqJ15HWFBWPqaqllgfFyxnKiPSYrgBw6lz70ENhS5cUbNZPE
ACpdXZwiOoLf9+evltT6X8j9oEFqUO9bTk5Pybs31keRrWziwvzep5d356QmSZov
mu5FJUF9pC8q3eaDYO1L8WZIVv7tVBg/tXlWat+Mav8NBI7d9l7TWGS/qocJsvYr
qqrOBK4C9npqj4Xw5aiYNvt6k+cOo/bAL2hJ64TbzhXzfbnfSoFSUowCaW4ZzJvU
wB33V4OkeKa7597JHKz2mh6afyW33cwQr56KCY3wn9Rz65+FVtxQ///iImCaOdl/
ilKyhgA+MNYJcy7b2H1v/GIicRINvFWRSkBVoVmFzkSym9E5f+jDnPqmMHnWeDj3
7521ZaDpSFi6ZPqtS31sLOeLLKy0ZCzdSlWZdPHVPPsMksXKB71K7AyFU7w19Dkv
zM2Hc2lSWqU9DkYG0kHCFJgwI+sa4thXtIksRKmF6gh0iJ1gOTzy2BoCS55h+6x4
i75BaOH3ZFBE3hQAkflIoy+hqXcO8XCp3ep/Q7b/oqysNYamihPHtT+a77uR8rTt
4ZYB2iBi987TgCB1BADUmHpWlLmskfMH6nvYwWHu/FZgt4eNTL+bPIf8fspLrTS9
DnDzVlRRDGlG++NgruYAdyxNKc3837r1PNDoBsSrDaDHYGoT/dAsiXTkBh9gjU3d
WzYqTHwT3ptAtzGD2QvSryP1/+twfbsntbEuQdZ+2ABtaFHfW1ZulMzz95H5h4cl
HzZriPivW5cWEKtC6OquECsRTBNQt3d+j81vWsdalwBh5jgPYnSj6M1J3EMsdsco
ZS9KF0jDU6IM1SuRr9lSaFwmcZXZ2ZctGJ2UBF+GuKroAEkU6iYsAY0um5GxpfP1
FUyxATOz+Wdol1S2WcdoJJef4BQ7YaxFZleUKszaewrAUMwnhEDnBiR5xfxp3N4o
43wkJ0K+75eYjL2FDBRyErm8yjGJ1IDe/TwmnqTLKhUCzMXfivi7+5V7A+OAggRo
1KjS2p4/qAc8I9bp/Q1sxwE2IL0ct6YqUCY7C6c+yUBvxmTR/SrSeTtKTv7qIIxP
poaK1FTi0q9e8ZRrBzGsjWEOAmxmv1YyLtRbuIJlSErJ8LWLBzGrsrom5uubwhYL
Xs4Ym9wvR/zL7mV5P9ngrpjJNnOOlOeU28Ok9b3ygO9IZG4q8RwFyEJpez6YIkpU
6pmf66c7y9qtHbXh5fuNMyOOugJaG4pWXngBBak5gsDBNGsmMzSmcyjol1854KNW
6PQ2vd0/zifQuc1duEZlVUtno5/ZMaMSjHRAl77XIuqKv6LmV4wtg31r/wOpi/cg
XoiEQvnKDf3LsswcnrdmfMiAHmD/ns+iClMH/H+6FyrD78wb4pi0rPU7GYEVh8wg
QwJxWcPePXhTvXcsRxyzui2i3tOKHrbPUkX/jY6O53Ht/4AtokheXsf9yQvONKfY
mYquSnNlk/4KuZ8vdSRPPhyQo2IsWESyzYG1XYFV3MfY0jOJzE1pUiPNKysnqAYB
Git5hxL37eeYz6n+GB49hPjRFYSiQzZ0pmAFEQMfbOU2+FJdZqbaMY76R6GShfE7
vauRWeDwWDpOk4JUD8FNJiJgjwK5SoQEHAS9jwPuzEpKkdQ8b6zHZ5vptQox5A3R
wP998Sci0JRDA6FlGcw/NNH9A3dClXNN9oc6jPcWYEzTOWz+ZY+LPLolKXyioZUz
LsN1iLbQ1hX3pBOR9qKs9Jw55+eyjMdqVdo+kdedIBvTRMx2dvxMQlNQzrqNiRJZ
aPabB/lSIwwc9jstMUZFfudtT6jH1j99K+uZE7K3pmfbW39znjKzOvtBVgwwo7XT
OonaYKHCfBay9yEs3TAr6sbvFBzO/S0xKZmm5i4bMIpCS7scK5+RVp8y96Y9/y+w
b0NKvnczC1uEOc6CvEJ7zwgEKbDNmFaQFkh6OaVA2LSnEBYHgL4D/TvUyPiXzak2
RiOxwmVR50t/wy1kjhgae1NaeCW6vWNH2Y4pXXyv9wXarrUDN0DUiI0JPk/BxBvq
JZlMYUrx3qvcrA7jBoj7LdCdLd2qAQe6fMm1j+2FflLyBexoON4I6gO7HkS0iC8H
v/ZJ7VhLMG0ceBCUyf+4QIR34qM7wohw5ISMrevcPsuibWfRkPrFCoJaJikdOgrj
AJ0WaBQMLChkBJTpy0pBls01ixrm544Ql9LbJpT3y3ro8d6PUDgQcfgtrN61Turx
tv1tEiWIQx4KNf3K0hJgmpVToazQl9z5AFIe36yw6SSBPXGb+9lwePMt1CP10iDV
foppUXW3HonrS6BtjEUEY7m7qaSb6Ki7Pl9FIa18fRjpZurP2fyl/kFH0mFlqv2W
t+UFP0gOxDfuj+hHu4Uxck3Q5in8h+in6QdndtFZLGPJCN9e8Msj07hl+Yrpathz
pAzarSdK95EvevFPPgq+uZYqLlmoQCuHAGlcmL4uvcO8jCaTjy0sbVFsVS/1VafB
ATYDHfRsGV+2qt/xghrROkPIb0uG4lccYaYXx7aXikz0x+vZs+PRdbf5BrtUyec6
nCwCBqfg6W4datekG6HIQX9LspvR+NS6Ehi/F5Kdsx2HivtOG3tvKhugiNm5OpB2
DXp+LRPPiwhCDf/Vx5qcSBbGsdV4wgfUkjZVR/RwLH6Dmp/F8m/6Q+mDAVVTI0OL
D3vtpJXdZ5IysFo6lWcPY+W4J+HSG/GkKsvRddvrldElC2tWV5FymKfaHaEdDf05
WtEU2WsNE/Dt9Aua+2csze00B5YwEhz0MeG4ypiaQJGZD9QeYGmK+IAeKIFOtA90
iUP7IlQLumQbO0r8gQqZtJ8s9mPG/z1y2W5z5GQuy6V881cBazPcQMxliSVRDDrF
dZNww0Xrzxv/D6rL7RZdaqv+ccrr+At3Kpt4cetfGhzXA+oIkRjuIh0IslU/dkdA
FwP6qGtqQq8oM80843bS2yCFbqUBFQG9C/aqNpcRL0cMN0bGAmn81o8Isp15JqdW
d+0+rI1kwD/zewqaVgn0acBJSd8BjQR3jijzTWCTCvbBtwVFFU4voH70aHLTLquz
LMWUpMiuLubwo7KwOqW803/0PiRabmGtkt0V2PuXPPZnZgxKBn1h7/acni0XWk8x
EMVGvyNgk/d+Dr3XLujv0Tzwj1x3OlICNk9Oqa96RiHpOrdK6ojPv5dHzGhCDTN3
a3mhWM8EjF3mfojs6fsof5RlAmmOEvp1I8zddRsEkR9mimJNZW/7Mw3SAsOr6FVj
BT+IIDQYaIfbIC/9soLwDr+6h+kU39fGwOUX2lk3X1kx4zHJBUdaRfw8lsKTlyWv
9NKwTZIYsN9Ont2J56o83J+m/xZtSJrTGqbgKpK6YRQzP/FKzv9PP7jdPhohnDrs
Tm3YWV3l1qgwT6xQKnsSC0m8gXW7jz4xO0dIJR2K5h1HWqw8DTegjHCNyDWNpiHM
xwD8zMKNPzpvG3AsARkKPfyyS/KzrF/8QN0SmBQHKs9P8hN/9sTS2AUThha5xzsx
V/OKrgByFrG+N5RHD7jC8I7s3fUwukzs71G1GiYC4fympJMxXCX2FQ+kNZEENrch
zwfpF7vyJ4e3+3tqrX95XaCOAiKkLxnV7as14ZNTBZh+eoWcT/bdQkzkaVd1qJTz
Yo2sQUqnArgL9sYQcTE80rohOJKYPK1pNLnES6M7bu7BOGhXckZHb1OshdwBXSMQ
VQ7TuJ2Ko+OH0o8Zv8o1M4rKTA4z9BiYJTq5sb+fTO57qzojLth74kiTBn88jyHG
0On9BaoK0ZdQhuPiVdY24736XyUI7PI8iQRlHGYdVZyouuDVsw+F8E2n78W2ToSZ
D46SRCQB+9y+x8gZ/mktxxYl3PduNwF3JSRzdBLFwyhNfyUczkP9YoGt7gMfU2c5
1w/t8Ti+nvdWyhRYBR8lHET33wLBU2b90uw5IdMrWKPkh4ITffpE2s3s/450qbEN
slOY75E0qt/Zj6p1iul055BsmRGegnc1hYACEV6U+AbzgsP4Wi7yR5qsqMiwhdyQ
I3cEF3w3IUAH8SnK+kIRv7HYEmFOAWbrUtW8cSAddyIR4nxo8E41ueg4xPwXjVi+
I2Q0zbGOZeZV6a577FIe1NeqGuEMcqLkS4VVHMyxEfyN586KSTSumKz0y3YE1Ruk
wdbHTTXoOIdemyHWuNrRQ/aEIqsdN/tCQZRK8ewgoUd74Xmh67YhndfzFjK5ascd
54GQmDxuieZ02q6yd/VpZ3W9W9NRNfZ/TJ4aoKrtLAI+/G/PNVPQPNSq+sReX2BY
e/xU4lXwLy5RcV80mA6jiaXeWp4PToLbWDalkNPaEgrUFkAdocHQNbdMjTD9G3QW
LCGwjMYDQeKTpQpe735iqeArPkIcv7DMiD5EMHA3Q5xCV3YddbVGdwdTzxQqry16
B1Y7gbgN5gGPg3DuL+/fkZT9ivwhVDTYqhRxQWejqYhKgkdTLWun1+7pGqEUqni/
PJhYbNdRl64SvwOzQW+q01emdmGB3GI4mDlwVTabQWzzrmWF1NekBYc4RQsxzowD
124gtuXQ2kUVrGrmd6xPeHCUjU1bhKk2nzj3W9MnFSLa7VJoyVGyJqtOQvNEsQ52
v4DbSXsHazlxGk3eAcj+BToOTtQvzKCs80mV0byCGkiN9acLtx2oTnKQiqghuUwI
B9gaaxk7+F+YBzeMv11WbIZM2FJkQbS6S6/FQ8P7A5TlGcEDGTe1EtqrbUdY+DqA
85CCChK3DgB9z2rQUzmJBrnEY3NbbcEdUJiVNwWLRFe64JTs5u24fD4jsTJA8Fnk
Ak5DR8sJgf+LpfvsKHn2NOutw2+s19WojB3CsAFjquOKOgyfUK7JC9GMjy0qEpLx
rs+kfBRz7nQZc6n02w/iv2HrfkWGTU4HG0v2Rg8MCUu6w1Q4cgeDDxuwidm0qMvl
TyqbOfJPJNIDzyP+xPbviPPcnkx/blAUIWhtKEJ1qn6lrWYWZeYKQw++Pc4Hy/kF
TeYMDFdmuDE/4GxmVpqEI7pZyVq+m9Nq8+UvAgkRIzgNR+wQAo7LeaLTvBL259qm
uyMTHI+R+V3aaC7kAUpScCPT/w6R0ta4/70a66+prIRz9mLZdzPy8VBxwLHm7ask
vJzXXqlO+aqBLCvrG9HqbJ6FqLJaloYTHpgTvlDhkpB2onQNprNYF4RKAv1YrwZo
c2SEvRW0U/1jCLcUVA6+Vixajw/LNxoTPv7Vfew6zQdOKDp0YmsWjXe0Eq0sf6gH
S/1tvlGfgDqUH4N+SJOjqLbgr7BFlwAcZuP3HQ2MLjDEAqYWJdhlstT6PB4StQb/
BOCxL9xLg345E0aUUrt285CF7thkAMX0l/ydWkXhP9crvagawzjq4f2f0yDbP0gQ
ZR9Lv19pb1o9IdUS4x5Z17XhFglqxGaezp1CMkdhkmWLnKuX1Habg8rvbnTSOsPW
NN62meJFnzva8lWUBJlnlxNXVp0ERw3DDOC0oZ5J0vZG+SZS4XqPXVHhf1GL3/qH
1/GCJxNBnMzei7e//5kf+cqEfcOPN3Whbb01HBBlGzycATeW/i6arrd6PtNnRfT0
LAzvFqvHhVVoUFIN5eLUzJ4oKwerTu2kA7Cfs69+TYe9eBDEoj7GLJqgDg65x5eT
h8A40J78Qqcg3RS4v+6TwLTgInIdduaEB9xm+3SHQtxA9WZpRGu7zYMG4P/gC+8G
d2fq6tWUAgfvcbstZu7wVuKJjJDaoBsohXenz8/CTXJxquIYpAvZzcKISnTXBq+Y
miPNmVB2HLjM7lwxrrCcPoi8CFoIcL46tfwiZ5gE799jvzSk3ZfazRDI74PDv6IP
8o/JpSGZciMf94R9jv4O/EZ04oWwIr0dZu6P/mec7dmVN6/O7ZWbxdQAi97Uc4RN
u19oy3WKzux/zHPY2Sqw38TSVZfauahzWLYI7eoV5MORUrEsHuCBxijFrhD31XV6
eKBE/WumnQXIdIBqEHciWITfA1VjaM6JPquTzB2p728OjjOLGP0nPifN9uBWc8Lr
oVzow6B6BHqHTHu0w0SwgG4eH+5NLVDiMNp2iHd1hdEOc/5eIKWnwgent0DNQ28Z
pIMKr6upyXaI//BRHM4A+vzlRNka3sQwJc2bWwhqASb7sXkN2Nk9Aacn/Tgwstgx
VTE+LPtxmut8SXL7Am2734geMdQoajeYL5S5mHjA7ipmG6kTL1W46zFoAAf7jWKh
isGk3mu11ZAbQcNTeB3Dtm9H83qty09nIF+BKGFaVGuxKQiZbseX4MBFbL/lg7MU
Zq/jrOaE3lDY09KDa4ELYGqn0OAPMjCxTx6qDDH/EOeONdCnJaRpWSbiP0FbIZlF
OXDKtmxJcni+nKjutFqpcTzI0I611438NfVM3szMRWd1Bd58Zhu9KaBQAUxPT1wc
EXM4VSe2vq3KcN1RGZOjHja1bB2T6yL/yTR3nVYc13HAOxHTa4SrBxqIa6BCYnw7
LxldN5CS7/GX/5hXLiSzsjjIbsXRed4wjZmHLPzPhGJ2YrSYcakGP1BXpjq+CWvU
L1GgPdUsdMPWrcDGb24wnfBLNfnw5Ly/uLdUWJjr4JahLrLR4v6h5e90uys5BFOE
bpvRcAa6huMhdzM42bYRbQXvF8Rq5wVZFJPEHAkE2DxUaEZ4Xue4hoEEfo/YQZnt
3iVcDAiNh3t2m3VJYurf2t0MfH0WYvELiSTWEiHAfgrmXFCXM1uGPs2mCedFixZw
5igWWoTuwb3QqWAcNRGRHnSGvGLNfRJ6Llag38Tjff44MWg/k2CnYbJluO9O12wI
P6xZwwsxkg0MlrP38+iiA1M5zLPVbc6nNbz5o1OBycb+8KMpDv6478xw6sAo7vD7
vKszFTibrO4JBhqwBHR24dk5MvX+WqbX4S6afDF5rJEbCt4RSkDFTwWLdtFbLAvM
JnDFbVTngIqsrQ3HtssvEtecbLMn/gAgnWpfRSAplaU0H/mPSV9fbrFZIKtwwjqx
/TfF8mwXbO+iorogFUyM3CTYZTeiK3P44eQov83gLO0sxBFo3Dkl2zUi4lsgBRJR
20oQiMm1qDKVzqNaYLuDMtDB7GvOACrzRUVMP6p98S7MurpeS0ulPVmgLTJsRpI3
UdQQBGK5vDJ6eR2EAZrIoMcbyn4quHhhz5Bs9O3Nc5YVEzxQ8uecxLWG9UX3Fr6j
QlKYkdkNJP1Yi99s+ZrjhlFbb2u9iwsQI325zxjM/dxadBOlCgwcRsoSXap8r/VJ
tgBx9FXcMH/GY8qW3L0ysI0XcCdRNd6qh4BXAhrVxTCF7zVw8MD6TCHMIDGqNIuE
fPKA8pq4C0GToCw8kzrGGXW8I93Cm5xxTCwVjjepK+UgMV/SfnKMsMTTs1qt3fNs
8ckIWOqH1HCdaUFrMvBQlHWIRQd7ucVipfATGyy71Q8gydC9z8DZK5u28wM0R9ju
KN6S/kk4Iu9zKbnWFymarxlZ6i5y6eUmW/eo5EDTm5xEn3UoPXeHyRyQkvglgtk7
kedPNZQ3R2lGicG/2slEgFOzwNYD9wGNy+jJ1zjKtCIUiY077nB4wPQ3kSg8ExnG
J6g5pFvRLjwHVLYFEEnfgpaCW1HgA7yCBQRJsu/c35Ei0RowwqJ4GdUc/b4V3+Jn
E0Niz9DzSYYaaYKbe6FNBpmchB8ALs1ZG+T1ZrVsUJfAI6aZjBVeKxxw5xyNdRMX
qiHQlUj34XGrqrcvK/R8WNVA2xErj8P+IkLO/do29Ur+K3qztgDu4hZvXTF6ulop
t7lM8u/ovoGVKrNnVkBkCK7Ju16RFDdvu6rvYj2RwqznxHOdQSgzRvdLaeNgHmF9
vQKRsZc8a0Gu07UYNf9A+xyMv6649CyyrhxImSY8ppJ3hwyroALHhMmmXc2XfzeI
3PSYeBGZFpU915GEBYN28NNemXSkMYnaYiaizxb7K7UF3vSHLQa2SaMz4nk6/21q
AKH3Ki2QcixD05Ugce7gvgcAl30/t3/I5hrJGLFIDMg384zfjT1WMTcX/YzGllrA
O9kThuc3kqjpNW6Pak7aU8kgtO0P8pvzh7E6ZszB9nk7IaqTdPChPdjL3X+/GsKQ
DRMXoAYfurQ6u0Hb1lgdL2EvNcYT0xhnA8Qvewkp1z/FjDg+fP8kzpTKfKTQ0xLj
Mr02NoDR07H5mA5o80iRUldnen3QjvoxzZmp+tkaupnEcfmjqO4LTodAZDEU3G2c
9MdBFJs59p2IAHJGn9+s309dd8b1wuZHmg/Iv2FArSI7Qs2x0JdkfsmcoCD5kxfd
TcBobI5j6VCUb6eup4ZRyQA9N5n5eu84spqkcMb2JYamXNYOjYPZB3ZjBXjhemg/
jUISGyUeq4NaTxj0gXgHtBt5oSg7UR0pwmkaGsRdO7fc93WfXUPj+4aaos+dUlUv
6UDnZqhdNJSFLXnIXC9uqULrojuwK6iEGNrgCEL2ZMZBKmAsd1j5Dl8H4OYgZACF
uFg+k3LJGqz4JV07W+H5C0MciOBuLy9yi5ReX2xBVEBbAIh5Gy25dV6dem2b+dmp
ZnDwyAQcdqISu7ziG38VVgNpNGdrMISEhoeADz+wG98noDuoA+Wlh4YjSWG1XcU4
Pj3a5lOH+mn8TFA04bamZLMXJi77rmrBBcD1IQO2onC7jubO1OK1vC2kDwq6oQR+
9boO/RrniBB60Elq5ZCrAmJ0g7burBTrJZAgxLjolSS1XDTkYNNRtTG+WMa3kqQ8
jFyC8lEemneM+MUIqET9Z+peqY/engstIzpBiM1b8ReNzFfQMXdyS2q1FD0IoUtw
VO4EBk8ztS1zjcesnwAfEisHNxyBZ4TSONiYtZGmFvYgQPV80qbwVRASdMUgu3I2
sbQHc7so025Lnwuhpe+1QF0Zo832GwN1R/FZc9guKCGCyCEm25t4NYO20c7HZ0BK
Fb4/Wh3nzZP0qbOK45y//gQPyK3SguYltlruWJoSnji3qssr8efDKC9QcjVR92bL
jaQlYdROSwQbB1vYee3SLiVk+vkRPOZQK5cfjQN1GY7c3D+9Kp+ljoIzQP+R9ShM
TLQcj6B9QJ76cAQjNh+gK//tsbmvEJdl7keYmj+KldCQylnlrf1szjo+p7HBeD8v
Rc2Twm/vPlzxYISTgKu5tAkx1RYrusgjbZ8N9AlKwUIBQnKQs38O3SJZQkQoeM08
M/r/paEN+e6QuSReBocIKOZttrPiLRDiK/s/rs9PiyYDg8DlTF8Y3GD19YdLFOax
7r/kNR9xxfwlZQXMIJhqUqDInTUa5a0DdirTYtrpmafVgtPoItr5U3uXnXx2xVhi
+nGfMLEmSRbReBtFbWJ+xlGj/qzNiUB+mAM6+hv7VNAd3Er1nVIVpSjLaqc6CoJ7
jM7+E/5QV7F5SsaQ/T02BxZLvRiN4lG8dMSGvu+JOLQX/lpo3V6XaHYzXELmbikm
pZLP4TQNQbloGm6NERA/IEIYuKvHINkIA4JQvkGU9zvdpBlqo7CLd60ltYp5E/re
vmFsxLID2lUPZwQ++SgoM62jK7tlILZiqR1JD8InSObN11mBhZ6NDBZ6d/X8VVr/
4JRBL8h9kuomjfWsd9kDzRhIa/n21aOql+VwPrJlUktwnqSZrFekXEE0H0S0qvfj
vGsEY9kOjD/sRJ6xXehJYVZwW0x4oM73x5wAIE90S/AvBMksQNNNsqnMW1gId1oh
10UfpnMPpL7GY25SJnilqjS1oMNUMt5j3ha3YS4BOVwxCas8CAcpxXlwZDcR1Z0n
ZOWCJI64qhl1fFdIuX6ImCcd2dMuN03SsO7dNPhUY/7+P9jOspUT9jE6760eeeYP
5JZ4rhAqblf9B7lL/74FyGGlmPnvNqwT0+1Xr+9JFWnFLvHNPVbQfarN/gwb/OC3
V5GaPdDUqjVs51FmvQwdiMTHlnUP4oyl7cip1ZE+z2JVGucahHDfhnv0wOhUvvjb
UPGhj8L9O2UIKlmUk+cEDO0QZ43dUQqnVBP5bY78oRo4nr6k7CvubN3chP2W8mRJ
E/ZmyPIgTHsPXyEe0MtJylOg7Jg3MK1eiUjGDxchNkXimgXMMcgoXUbVNmAlrSat
XLD6aWGSLIXOt0dWICGpTV8bOovWSEVGBO6n1ICYCYjalFdUNcNwrViWVqsecavN
FUia/UQXaxgqEKxIOekbtMK3FC+bAP4Vj7g7uhd3dTafjd5ryDm/FBjX2bvO+4sh
2iAPeB/jMTAdR7q9VRGWSjkzkhB3vOGKABIeJpPEX0LJwiGrgcLZmv0PlqTzxCTQ
cmsnI8FlAWQCZeY8Am1EjZao7FpBJWgZWXcc8KSzY/egGDTICWvDwcAKB2fVCGrJ
IxBRhk+BhZsTGUFyaBw5ieBc05YGgWMC44IH8KiKgZmHgSlps6oQNbzGiOrANfgg
2IDVTYWM3ZWV1XOMdknnfuXN9Jtdl+MGTzy2Kjwg3CMCKPRN2T1hq8fINNdowFSz
IvZE4siKTJE8acz7h948MuJTbqE4TgwVaQWWwOtcurN6tsS7d/Pm2/vgP0vwrvQk
Nr3A6HWiXKY9sRktrX009l1HZDxHKzk6BBxvCQHt3/okhCA3Z7vaH+oeHzgPwE32
3fhn5gB1V7MjHMa9abTqf6PFWewhYBVuszhHi3JjAk0Mj3s/rcnY7vqvIHSrQogh
8gGWjweOFgPTBlIH1O0M5WkJjfyGC/fRI+v97gSixIvkY8z3lYTT66tTSv5Ziw4v
pnUd5iY++HJZ/4ZKwEN1hB6uLUuHVjpgM60m7pNOOFFcD86f/Ns2ppNsPQoOqJhG
XHCQwuosZtazzp/kLR3/DD1Ffj1vIv5ueyPP9pK4Ob5tkJFILz02dC9hJdI7ZkJg
COa7Q9gfCSEiPdoO9GmaBSUj8OEQMu8OdHdiJoFG3SZGNU7UxQScHgAJPnwntIkj
pEHtcsOQJL5fzZNydKEFFvHCXAdOxSqNA6d82NmSf+OfSuDyoqwIGZA/2jlU0BRo
4XXUR5IIQqbwK/XsWVT56YseH7IaOeCGh0GJ8cTSVEjEjDlXB2EANk1XGsYMWsiu
lzr6RnSQKmy40BZyqAZK8q9Ibnxf5TVdStepmM1HyMD8mq/2emZElsEB0xsJjeKL
F6rwkn5+nikNVW4OEhsrbXTe6rzE85//paKfN7Oqsb96iFcwfJjKXQk8nFKdLnJl
1IWtw7XrboF83q4NYMQd7ngFyt/Yl3LKUFQ8gFcvBQnzdnqBZoku6Ax7nlH2Llvh
5KfKxuPeF2KK4PWd08Pawm2CsxrJ9vdK0X1slHsGLwRBR0rh+2FJEz3hRQwpSA1g
HYQdKJom+vhVZp/KW6+/sBs93LrnTeiRIdFv57P3FO4N0LV4eLSoXOf3WhoBI/y2
lAvehEe/5ZgSdWVAJAgqiY9IG90zAgcZtZ/FdDxMqW3ZEH9EBYBDWIOPWfeVUruB
Hixj7x3o7qPGPKkk/HHy3vXzvU7k13hsEyUObOhKxk64Uv5yi9TH5n0kGjoG0fzW
jb4xsCdGJ5BbW211kxI5MLvV9RDW0OAntOP1bNnKVTzLkjM9h9ztL3DoxWfkf6u4
N2hMGpc4crfMCLG4ttGRo/5F5oze5O8zlM7oZyImhqwm4TJuedMMrQg/MOthHjga
wffKEG6IXO+fBJLqjE234u1r9mhQbIPlt+lTj690UdfjYX1zogcDN8O7/cA++q38
UyDwXtwqMNpVXKZth7nFviqD102bFXIw3LH4nNjfseABF/4bQKqlJNk8VWBnQSKx
eA8bIoydoTszzISX4SF65RE9lQJuud7BfoO6pL8NwJZkNoFxmJHIYLe91rB8nMto
/bLmmOO4SHP9P4P1IB3BG7INZjwgcFHgcoJ/vKynXBQ9E7D8lF/Qy2hcujUY1IOI
KEYXQvYsbFb5r8zjLgJkyM1qdMfIftaFyaCkyB/2yDQBtDDKhLuF0pfX3lJc/ttn
mS6udoU/9TUUKRLC3Q1OCCgXVR6ATQLhVLxJ+rEgdVkHRoVC8xEKD1bQP4izY8Y+
NyMYqGJruejpPS5Sr0fNZwClyzutgsB/Q1N/rXQY0nlDla6yfki4zkZtb/TOnTCR
1wiaQQO+gKBK8anD0rVyBBRb2FC9XokB1qGjqvWR0K29WzigxmXPWHNI59UiKggj
uXollKuRKxaABw3FtpRkboGlkA0LNygNckEx+dFAnCsdfvrp9LJOLyAAOCupGQBr
PApBeS1Fr7EkLYIKZkuE+EXuEdA2tqkUxUnSjtxxxcEN5KySutVOCQkLYz+ADbqL
IXaqxV3gEBEfuI+i5YoxTEiHxtwQT4QtT57EidKC01/14mW5NYbloCH7u98FwNA6
hBxNGSmzQ0/VqCBdZACYKEFf30iZvilg9BL8HrO0+O9ECBLa+rlbBY/jZwrYRJFp
VRgnsJ0pvJYEXdTZqUuXF56nSU9n8TfNI77BMvMsVs9dPa6BV8HwHuiPWq/pbhvj
waf4XYVdoZygC/T7bhH+ugT4qsea/lUgaLcPdFXPgIeJ23LHr+v/+lALmKaSN/hH
SqrjeLHm5fqieaU5jqr2PI5c7XB8Qpjy92jvSwlXUxUT3TOyCcBWnDv90Pv72dH+
MWDfg2h5JmYbqPkcuhZgu6Bmh5L77c+wz2TmE7LmpiMoiWfUTTlbRlDmXrgRe6Or
494O+LCs6wHkwZV1F9y7Lpw2Pb/ZeopeDbt2nMob3EYoZTwl5WxMQ9J8X34+qFDt
R+HkqiO/2bvPlZBImnZpx3FFt3OGIp/ldZg8SSd9g4TKUvdcqkdXP2uhh099nid9
1C+cNvKcRsjBKgqPssFjSUql4W2dxNLH774Og5JV0dj+rodYPtXkwrz6h2ac+B9v
+jM3O7+H3WOMtaqcdP1MxwgbsI13nVLqXY1hAjG34E+cxkfVLx7OEvEcTUm8rdcf
RzCeyZjORFJxzPgWShhwvH2u4k6Ae3fSo/tWnBx6g8fY/o7tjl/rwe7L9uqB8zEm
PF4YxnK4ZBC2GuOPYFYnmeLTTEXbWRPcdSRf051JwA7N0TbWvUA7eN2JDMVEwCp3
x72iRUqwjgYdk5Bki7ZoLQ7NpQyV79SnBL/6Jba8qGwaw20uHTLE0u5SBi4xSulJ
YE4M/VLeLeUuL2DaMSUZ/8TDrkXB/foqEX7dkC+tzw2xOofSh9TRem37zYtUN7Ce
PLH1b2aM7qDkMeXzCl0gE3w+sOMxZWDHfQUBO8xttUlhjcM1ClFcU6gwvIovU6Bt
4RaPnxI4yCuhDDAeWQbv4nPvuQ38YGgAMzD7FnGzy4o26HoKNZfmQFIlf95P1DXb
fDn/MLrhUbmN2UdUZkgl+22Gp2o4dMwZ68BknkrjJpHaVoN2wWY2wvS2B43Ik3ru
dTd7TCTHJfuxJqdmaVysyaWmBC/aMAnjdQPBcxzfDQxGkvY1Y64dgQe8XY/KfzUn
FIu9GAID1PbNYS0tYD3pRHWwzKaxvhGQCJKYX9iYCPPxqFKT4C1imHtmcbZ/04W2
Mw+An4+phqPUi9O0uuGsKSq3SyoqluvDhuhn8c8woH5bvHE/6xuYhnT435YYipk1
xy8iuGuP0WeKQJxag/266dByK0V1HkZpXNlosfqg9UIEOb7GBBbMCJ6AP6gnUCFL
M/PFgXx/3sJUytbg5TpBPtWxL8N0zW02m5auWMEx+77tXI1+8k2tOnfl28n5ux5y
YMzaA4cUqIsVL/5nyUBE/CYIFx3bq6UcGtLgqzqIyPXAi7BDFmQXHi4/Vb1FAO8e
CVi3DwA0kjwM+JvVjHkyE8pQCwugchbvVOdVOnHnlR3Hm9Q5JBPA4XEGAI2TLRi9
upAvh5c1lypMbRrL2W5cIterpB+7kXOXCzw6ieNB87do8QJ5XcN/uldsKWPUyt5R
6g4QnPjx0St3GHul1qTr7hO6R7fIYya7Pd3YqAc7Y5xAsEQMjm29VRDpVRhwxs4L
rZKJWE7I8VtDdP4qSqXeTZuZXwOVWSHanv81DBMEZIUFS5oXgV9qBfMFP1JRSVeh
IyYRy3zbZxZrtN5XJG7YC4dd6XJ4k07X9v1DTVKThg/CzFkwEKd2rjW5xf0KNdRq
0y7iBYjKUZ04C8ZfTMbPxENiiTqxQq4pRas+E8qn/AwZn/BBUcP1mvKsmrwPK23l
oSaZntdUc8b38O0RWuyORjgPJMlUs7vEkpuMBP2q7arfTTxWFPn4whufWV1Z57yx
OHikzDGXNlJfMEQiai6OcUGJHygTZrenVcHpn9di1J/3ibBniObxq71+F5y/kOAT
9ELJE16sTDPUDonYIP17gtkO2mxc7uHX5cHr+HZXCOCMEUl3E3Her/x5lKkRm7Ep
9dETE4vN8G5Ycgjz9Jbztrv26rKiE7JE9w52QctIFwxAvtT4Jc2GgQy9v/MElXni
gsc4s9+5HPUKcfMZUsAFpq+Aec4p6II1zcSoEdZl19EbpQoT4B7yIF1CRc74LrvZ
K11fZvg4AhWoasmlkifKV8BxHMOtmbhI/P5cOWB3Byfx2GSWAg8hsISJgR6F2ZG2
+si3QFLR8Jlddu5wXA982JeJfbRrf2LVfWkdj5G16BkvBvsXdSnzOuTLADAquHzd
9+XoN+7BULW/w9zC9rv7p6hXdH7+2ijv1gnwxIAjztE/cMRNhGBHJbT58pkgwRWG
aQ/9N1TGlBNemfGhzD2M2fjUodMCCTBhhgS4xvb1s4kQVGE1CYZqV1xQWhdgNevT
kR1jnEaCXLMuYX1N3i5XiawlM5IyzefQjHfzwjcU4ZmmNESW/vaFJUHfFriXpAJx
EP6Mz8HbKbYD2D0yN/IiBAF5oapnvOTya7porKK3rMMCSz/GvB8EZ1G8KIOGVZlz
zchwvRnWUfiEvJuPbtjNaOP+YGIOFAOJskIDDABHUGraJArd02cPJB0HTxChyBTS
MTABZ23OXyNmqOlO95kaJ4ZLTWNwvdgjOyuVxHCs1ZBCqU2Rw+dFnlX518FfeGVI
OMtxaX/aDtXsAGw0neoK8sWT+0YJN24e4XjwKbnZYY8CPU1HOF9rC4SiD6vDD7Sl
CwcWPhW5/HLa6IxHqlLjrnwWukqfafA3LwQs5rzn+w7hdQrOeeEL/4CRmX3wWEgM
IU7cxWwpCa6yv3oE1NzTeqg90SENt+K7+qrRhneowgSmST37n4UFhj0EKCHR6xl9
DMBTkXVNsV8H44C0//bzeUFwGzdvCj5nK269Uy1BpHkGd0tUoRAEemXNs4GP5LlA
QEdhBVEXVheLshHOXIko25TieEEVhnZIGltxXzx3cr/KTSY9/w88PMLBFa0GnVgL
UgXACoXFlak7MBT6/TypU9BXwNcAwFNpZcCliPeTFN2jVfAnbpmBlOmmVUf4CHlN
WTwW7H26/Y7SgXqI/C+SP9+FksBuBwzN9QaBKoFwrXtwxZf37U4Hxq4GFMBi/MKr
99bkmozlziLcy0Ld6DMeci/T7u4WBGjwq7WZJg9onpWNf3jNJOqatFQFl/xiHRge
Qkxpp76GxF/yYdJwlftgv0+SKGNG3T9lXDpQo6+w3yzzLWQ0LPULRQOS06+NFY2g
OOnh8jnBYs9TkiVzJVc369KTSKlJh/RJgW9hKRHldA8npLwRWluvUojPt91g9PPu
amtFWIqSCrwUoI/y3TRyXKERXhJ7oBl5Us6XoY6Mf+fpqmwyFXfViSVK6pNg9FND
n1ItAfWhE+Uu18tcEY1eJ4qoxLaoEj2A7RskOj7j1H4zuFb0AD2XW7wiXxMQ3Y7R
4x6MpLA1vs5q00SB3WhvxTumDfl+p3IE7TDs7iMwIoBIr8uQ7rEJLwZh/oWVyZMJ
h+SrsK5JZdH/fKCf8fX6Dw4It17at16Tepp0nBV7NQwtCweCbgZ31gH1uCepuBgq
eSDFMGM9tykTihM/INf8GVIcxI+1y+HLuh1LYRDojGTvgvutifonwzkdF/wnzZaB
vpAYlv1qt1OyAsjIuvyGXqx4dDSfM4YWhCIj7W04VfiSsL5J5F5Z6cqcc9pqQNQW
06zUjPsHUZN8IiWqhQYU6+V61yEo9TA+pGbW0970iYNPTyXtxzlyfbUqAyjx7RIl
KHCzv2Cq0TvxQqZYvxRPx9u/1O3+ZvyiBzgwY+NqfK6hdi6L5mm9h57YFZp+6MV2
moUqSI+i0eUCJRM8FBTqueoIag+2sxeTEm3KDI679t1nFaL/K1j5t3s2+iaikXHO
8bjl5YlRuFOqt0w2O0HiFDv3Lx5LRfhpiQLaqdPZkrDOst9cjYKU438pq1zTOkZd
PnzUVjsW9OeQJYimrXZ6UFTHJAjCjRJ36NcPhZqXsKNV9JoYvZLnySo65s+XiUfi
E43bomWEw+4s+4Xymedz0fvdwZ7oM9TMb456ieBZipVBn70ZJgoleW5xJD4MAFll
hxolIMxFcY0Ne11FpBmzGx0WJyXCjld7fCWMmqa6dmgl8jq3V0JulIzDeUX0DZHP
eZ2munnTKI7/P3ljN7Ng0gO0INHW0nbPrAFzYLtwAjHG0E/T+Ewpc5k4WbgTZ4yj
IowIFYd6Fj7pa27m0Mo6nfv3TrCN6F3Yq4+B3m9awVKxDdfLmpeOYtx+zI7/xIn0
WgmQslufQRyeh0MWD5JASB8cDXH386HCaxOBbLDfTQLWfjOdsSpzDwxit09Pknou
hjrYXSsIY3Kyu06XBXzHd88V+Rc5j9i5sqLli1s+AKOXjutoulm2E91BBZ3zQ8zF
n0hEVvnerxl6bh8ZFH3HIVMcHvhbaBkDN936NsfpMx9kNWUXEtUW91sUbuzw3Ukb
Rv/ZlgrVgKjMZZFcmuL+olNqUyp7kDOFhracjxmnnv7Vv36GFkY4p4QRSRB9w3OS
X+9LE9XkQ5w2sW3e3GCfe5iUeV+/SW6eBxmbf291x96TwlsEu46Fh9WfviFTIl87
Q0iAN6TuGze9Lk7S06Fr7btvmq7D5NnzxR5Uevnptyooe/eqwzBL6J/AWgvGYx6m
CsaUICArpt59KBA3Bx2rC+QhokQczzUVt0nWhVQlPpcbcbwQ/wQRO8mC/jxtyn+u
EYHPLesGd0zIUJ/nIylqN0qC5QWvXWtaNOy5pu6wAVAgO6QfjZzSeVB0f41z7E74
6erPOUTajNBe7cAR6KaVXWnjrhZVk37drC283t7FAOaWUPLyR935kUVNP7uk5Oru
sZ50YV3AIdO7XyAuk9ARuJJ3lQ+sMKDT6zjIg3bUEEQbvD7tximG2jYaaM6D/nwi
nkVWMvrjizHY4ZvUgcU06H73fp6a2zg6cJJnPTrtHrnMhpiFjCmgNutkXwwfq8QN
j0bcqB3nKplKPrBkK6bZQnhbhTzF37s+cfr5ykedyaEiIhUmdgqqwe6mMojkTJte
CrqiCecpyJQ4Yb27XN+0vxo++P0efJiLv3mymObaJE4ayCPJ/q7i9HpfXLWn30OX
zwmRSiggwDzjZI08+p3iBivymK09bpyI6oOR7nXh+1bQZOeDEU4ikcGvyjjkbvNY
qoQlkOsm/37XDD40j+F6+5PZYW17RUmjyEL+5GlgrsDvmIq8BkgSQcuTeuAq9tG0
koe7+KQyVWCiyeaOf8w5BpApY5b9SXBkuLSHx6YyslBBX3qzW1XYyk2qVcLkEHkp
3ldLB9Llr4S+MzTGVO89W9xl6puOnbpEjQYiW2laK9nI3SrYDPUJ72aDvdgwUaAI
3VoYsmrVW7SYOggDohrT+hFME6Rfdg4+uHlrN3WQaHelrTZtFUTz+YOOr5BB9Xw1
DwtaPSjbHTMZIpn1K4Fk9fBHrDfFdoy22wcQnp4RaMiK3ddlUebYCw0kKdrX8lD4
taNev0oUmPRR/cLUvfhOKiazediXB7TULEZRzwluwfyPr0VuJqClKTi0AJozUtOC
mIRDM5ayQjIVYx2gEqk/24DUM3/18Qx+Iy0DvBe2m2A=
`pragma protect end_protected
