// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:47 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GuICwm7KAA1yX6o1rFHj31HyTK09z91kahXkFIyzLHgmZz1W16Y14N7vOpBFUr2I
1qI+8DTnsCQGpfMsKDgBH6dJOzXn83/6j2z65cfXIIBgXmmRvIdWH3qr+GUUSBL2
emrjH2X2SL1ojoM5Vy0cuV48lZ09vMktfhkUBEQ19V0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
+I4QbUVbKVdLvKAEwR4Oft94nHxr37pcXch6rp2hRcwGdlSSdhpAYg340+rzy94W
+n3jW9ihuMLd98ej5dKVKMnJjhbHdkBrlPaVHsNr1hdz1eX7hOq6woFFXgSl2omF
Wge4YeRZuIhEI8b4MszNLo4DFsweB6nVXuEviOAxBsglAl+wZDEtSo3Y7FA+tWDP
Gd0OElPl6UM2jNbxLTHIv43BP0EIwQSdAX8A0zbsauRVdEKFdqsvg+xcEWTZt8Ju
/CWgP6CiIBfo6NC1V+nEM4j7n+Yv5SKp1cVF2HAbzQunCkEyOtSJrb+rDkVoI4Ot
7YlxJ2Fu7OelBpFRM2hTOwkwWULCllEGmKY2BhOlw9cvnWczPzBh3NSLR9+IJ9Hs
AJs4AdulIvwsZJgu4+OGBi99v7AZu0id4bFaNJmhhGcmrNEZubMEw6l4C5uXQT0i
L2MVjIf68WVUtU1wKtQ3CjczQFVNl6EvWW9TcaGij+mDQhLThf1qNzFsetHhT6sV
kRinfqOzioMQZGs38gST4Nx7fi3pfltB3I2jUl3RGQ9XUG/VazvaAJyVHhPLHcq+
TMngrKnh6hOERn0wx63xyARs85hxUPIsFsBm5OcGTWcFptssp5BoVHszeJXVB8TZ
3N2XmjI2wUpL+Mf17yGZsk1oFcrmKhFXySFOI9aWG55RaLK4VDqWL19q7gig9CfM
/+8jB7c+v/JTg0A7ZZhT1B09zULiGY8GZ813ibwimtBRDUeCx7KJPf47waVhjWcm
964Rb3EJiv0YWt4p1gUglo8WnLKn+VqY54yRfNt4KkMjbohnH4sqPUegfVJelUWk
Sd0l/JX+GEKQW2SB5SPwtnaVjmm0Vbm5hh3C1wIiRpFjWcJ/5d4qrqaDf6XWnqRN
UgOd3zKzjbd7QIoeyuoZaOCqrRO+WWCCn0zSgKtokYBp+lLpuFMIKuYLvsAV2Ube
44aiRvby0p6fnGIkOToG44L2WfQgT9ueix1rdvQvwlgr3pzc3+sZZpYhRwc4ydxJ
/KzHrccrtUxDPoX/W852ZIa/XjDZ823wk/d9ni41XoxMY8OHAQ4Ng+7LoFcIMEuA
YN1OZQbegTkJNiYGzKHbKyllJXy1x77FCkyL1FBK6L1tQNNSr4NgaGw6rWwnkTG9
f7QXteszyUJgT9JTAg7TfT3OzEvqGA60y+sqP2dbAYITOgvUGGel8djALxAswGDh
D0c1rNvx+BJwxg7kmYG9ahRYc3CLdZ9Qk0bq+HbxzTJkDbdR1+zabkzDXsmBhbRP
h3Vy78So8oYL5inFx7X/R5PqLNBVWnTAvGUuANcL4hU8kOclrX+x9wmKHSkXEYKG
X71e20wzOQjzYxT1x/+CZH2dA7sAnjSfPy2PQepRyalEZ04N6mQgpFu8fVTdgg6r
4DLYSpkxY88VxLhv1LAwimTMgICtRqg0JaOJl+QEORIy+uPuFpLU3VXoZmOmQ3+e
VzAMP19AhNaVzF9/5MR1Q4/XEnbZcMUHOkQCEzs7t80v33/jCyJjNyQVP420cXBz
38FC9cRJDMbsOQ9gmL1qsY0WepX63Hf6x7x7AeFobyXN5OIbXkrfTPrLT3JBT7TG
rj0PoFndB3dIoC0F5Pairsppfu+7JLZz+tUI92o6LkQCQcHpXMwJMoceFRROGHKJ
vFN3K39eHDKOMKRw2fKmgPO7cHR88jEmd6m16jJP+XC66C5TwlJb+LNoEH1tWZ5+
jMNPjWYMHAe3LmGegXlrK5MvdebJxs9T1NX1CSaJCNBFp1gCyvDU2XXIQOyEmepx
qliarN9AzbnC2H61QXfNHeLAo3AUU6tpzikWs4S8igmmmpXrUPEUdj3SfwJvZEFv
X7JPo52pkG/mL3giEXxxagVM1EVtoEapXqCYHGZvpNY5SYNRgdx3mzt2NigVEchv
Udiizgju/jJgk03tQUQgeS/eDSJMy+BLkdL57oAz2mrNa5dC99z4zVxi3xfyGvq2
19gj6rpsGIxjHETbGX6vGW6FUmClbi1YyGbrbd/MDjYUGv8XYTIzSpaoSEwKfU9+
sTX3tGmHrfDpExrcXY1UzuG0p+uJoIcuFv3GQxhC9meA/FKCCXREeAc3Uo3orK1x
9lXpS32wAJ6f5fjH6zaa3dP7KHikDIZ9E8waPZznIWVoKX+lv0GhahSFA79h/lcX
kZeHHgsY2Z0X0wgmrBwAb08SxHK9TyuFv9MF3QAMi2FNQAxSs8vfhOpR0XeIStOr
JqMS2nHHtByBpftodRPdSyCyq7/SAFPwq2Z6Quoiyhkobo/yyj1VLiW2PsOkC/HK
mW7I1Q8dMbgYWDldorlo5yXacfSvBPgKFWEHbM3HeqHx5ow4hJFxrNZk25cQuDHO
TGnpOAMm9iIW2QlRVpEmJ0PVfi4jJKgR7IbrMte/fY6oIg3MJH+O5N7W4KBxh1z+
A8dSglDK580M7RqiJBf9wWrj8b5zBugOCMdqERCIiam3BTdeHedi0Zi9i5Fw8NAE
Wguahk5Uo1o/LkzNYS6HQiT7M8W/a1lwAzMDNLZZR6GFlfJOjLC2GFYjk0HC2HeS
D2OvZ6YqIzTVgH5fX83ozO4nVlzECpdrPeg7pYknkrGLJmokX3SLv0VDQi+hI9Hz
0KvpnqvGxWjU7PgL4kLf3y+Z+8MBSHFOrt/4QEk5FvHR+zQ6BvcDNjsAqdzTlWGM
jvHHSUkb29ZkXVMw10H/ZG9HQX5NGaq9ACLGJusBA7NShE4eiyYARLKHt4mb38qx
TMtZd18qBpNhY1I9wFulC2hXuQAU3RlyizNK/gBUZ9Sf3i/t5Opaz967wt7AkR/K
XyZ/Vogun1WRGWdR9CnL+vMonBs/R9Q6Um/P4j6/wTYiRLCeGZIOb8sA8Mx6K4Qw
nyxcQJfb8lohGbqFVrBEzZkCUOQUhYaHgONW2Rl8SBkZaCGHrqss3Gm7eb9C1xTa
BJSAG/SE1TurR7gKAmsjRRcD+THMXKDUO6xN9Tx32y6T8CGDRpAKQlQMJ0eWjKyQ
utEJgig07muHIn4IV2jnc2srApUWkYLuO1yxmd5iSKJFkc8NIy2IKjNZTBIUzObe
SzWhDPe5kXK/2oTgvo5gd00d2MvgOpyw6Q3MxXnA8NXXVV3swN7hn1tBCw3w522f
xT9LpoHatI2sGJVA1cp6Wv9m38jgt2/4f6/HMT3AKsMtfTt3GPHIbQx8n2/OcH+J
CfLnF71mf2kAlZB0Em+QTQzkLI4Wo2Wg+JTzRBHZ+5Ut1yvXp0SDXI0ck4TO9+0t
+uolPwVGLwHqzsGyRh6N5gB+qOgK7FeB/ngv33aHk7A0LbTtqAKOg/iAdoLSB/xs
MG1ZiIhwGYdKyktNUbhPzu2Bsn6wWs0YDS3yj/4ABXK4E3FqBO2rHI9uo2eO4Jr4
a4NuKAoeVQP1PcWMXzIMqRgb5kVTGxFbPfuvxIQVhGlBVptKp2viOLkmJtJrVF1L
mjEqkwYoULGDBh0lJuHL7GS1uH9LPoxbPLXFdOlfHlG40icztA2yfYYY2QpP2565
u57SdhKg3uYNrLMTqRkM8xlSuvGPdQ5Gm46BYft/YHntIJvuar6vcLNetUAsEm99
S7bs+Jw+1EBcMQSFDvUXJFgCbmKaOBdRp3K9yyYl04+vjb549HwUjrGmwt6xKsbR
wyeycU1MYc47vAfDD23teWQZFD+fdgEivf7uOOGJpx1no0yVhjO6BTnPfNhQ5lYq
7QBZU1UrVDMip6OFy4SyIh+L5D1edTBLEp0j/o/Np4jeP3Smgktri6WVsPVzbUk9
Ix5nI9RCVDW1GFPWcxmtZ2yN+2p2NIQhpt9XZ6Y2NaCPG2XQpRxSj6ok3qj5j1YI
c8ZQ09jedjSDuf0+jh9AQJwRdIAPjqejTFMbomulwCFTSrC54NERhExRMxSsU4YW
/1qeZzYJkibyjGVhraMMV5GR/Ohs6ciO/118U6DuKkp2npxJIvD1rLR4+OZO22uX
7pjlq8o86VDbsAIn0ElakgpikgYeX/5KyL+vhN2ZmSuGCuDPuTsN0MbnrJcaoGgT
eqGePNqhbSqA8KA/i/3BYYiHsAvTuMsuUZEEQHIVZxOWsjZkbSwHRXnhv8ImVw1z
agt/wcJFWg9B//UsYLEqgHQ9iZ52q8h5x18PFQliejmhmU3Ap9MlgUPLiLjr6rbN
iqnnZ6d1D6CDA1rIjsVVdSqF2nPQISOPg+R/q8S29owVElK+94DTpJpiX8efWx2v
dG7lCoM0QLFhFrfmn0yrz+Eb3GlWr38YzZiKnzUGYmpVCpsEQw5+6Iydd6BzQCXl
UQZ1IRgtTAQdVDBsDZAORfnxXbHwtuwkxrw6YrpjvyaVMRmb8hhlNlD4Es66n9Ne
YVtif2YkCRlj2YCoZVxp+G+DTSWy9eOiXJ5aSyKpY1ho0w0CK0wHtoao67Vj3hPP
FUHi2BfKPY2VUDGNjmsTAkedZ7mH+8cFQ4CoESSHCtsab07TN3k/dCQ2N0vsD/EI
j/wA2eUtgf7qI+2yKny/r+YHRQBy1wxXFdV3Dlu/Aefc9mnDn7bS75REYryVEif5
bHd/evNUnh3QcHlZPfXYHdga8DAG29SOrZK7mSepuaRWF+9TmjlvPrkMpoLYrevo
ZAnWEA2naCUForkhMlPZzN/7xew0CCqeuG6GoTettJCEnW6hYorIbjSgmsL+n/q4
1ToFBo4mIrCbpARdve3+G54Kvzez6WHdiiLgMF4JvnFCyN2DHZ1uL3FwmB8mDl6a
Xb1BEiJTAivvQeZiJFiPeura3GAWwsmkhgYPy+FJ9MqPeDGqdBoRSrMHG+qLKily
5fw/cQKhpxgrwe9hRr2znQR3GkWqOZLukaLT2F4pszOfeIHU0pmVDWJj5z0RDFRG
ev466g5KELC6Rmbw+4VROdpNJfJGlO+apeiIhDkmvSBbcCCd+r/eR8cmnGfgDJQQ
0F+rh/nla2hwujksulrIJbGcn2sp81CkLHdTcSCoago2e3fMhtJDW7PzusrMgyjR
93i0lIzdM7JTJtiYhYRoGhzZBOqP5a3pWxRS1ea6a/WXQBIkDe/CVZyoa7B52uOr
pvTQZzySqvQlrCRcTowjoyTsXO1pcrjpkNtTERr1F/4wh7s3Eo0NMC7y1yfl/WOy
YEMM6V2Xly0DbzJNwxj1iMysL1Cex2S3V9NNjxlIRJYUEPUycOrFeaO1L33o4jS5
SJyw53IZ+xcn3C4xb3cbWpjDGO/K1jlSqT9MRWTC19ocHKw8aud/RsrQT6IRzoUd
DoeedBoBO+RbwPiRRbt/aMYtoDXuOkHjC7bIH6V7lKHoNtWRAhNYWmpbECa36VX3
x3Rdz4SN9/jcFJBgejGpegy/ePAziqMFpNbU2grBKBbHOVA323X6gnMc/W+8/VE3
+IktoNglLUc8V0vfEB+t1wPrtcaJMyQv8XNt3RSWCYVuyxR2BJ7ALXswxAxCPTOP
0dOmUIdBnr1qxdPVzT563SGRwh0PqhgY6ivAK3BeLEuy9Mhoh9t9sspbVapSeYNJ
zYzq2aHJO3mf5Q/zY/z38IkAPKeszJRHYm07uBR9mc6lQsbSzTRkTCIv8tRoLlcV
YWY2STMWGOHYcogRnilwOgubg/8+ka4TaecqV9Q1BLq7If2wWpHasdpDFXMIp60G
9J7p8+WKmPew2UNhEVdo7MweHCW8XEGUFGcfXuf9qtEMVvHsF19+cTCUgODkWJBx
Tdubu9BzcFJ+O8sct4i84OlufUXbbr7YBHfIKO/IGQaOhObnI3QmXAL4UQfPnhKK
SjQs8xCJkbKLYV6T3fzYSQay7LhQsK+R3qe+3lxd5XcIbBTw+l7sdlgh9+BjbOka
Np14LZSo0G/uAVITWlOo1MInTGWEDR3vnDqTymSeDqdEm+ZwStbNEv4g9yhkizz3
yeEIBIeSgwnGVUu47U6Q+lcB8/QfX6xBys8o/iYntOhqbB54C8AcRXOuGs0qBM2k
srXLx5S0sBGj/qbq45Tsjg2LVFuBqhZsJAwrn/1KnaDnHrScxJar7UgsJKKe+/xz
M8gRkAhfkUHrClGEIATfjvObp5v9GUejniWuU3FXpcnsoqJfQsu/5NJEwj0xYTqP
9I090IinqkKF72YSKvHR4z/2Gmv8rG3ncyb5GLhPyffLJI6DCV9RuhDBy1VCQ8C3
FRfWCBJ97BEJwCURh7mTRVUrzk8h1Ryf7Iv+xJDBNmOZWBU1jZPqLSJNQ0RkHNT3
m+PYc7tLyRVtYWnFn7H+c4qw7T2XgBYUDFoJFlnGMzRxrtgk17duV+XHOZt3+8dD
8tUA9ufCRIzkh4pKR7Iem8JE26x1tmMGQ9Zo2pHBUshNF6wT9Kdsvh2wh9cmmPJr
PK4dtKTtwPlHhE9I58tNRk2F/awvmZ+h6iHFlKb6JMZmV/lH/WaasQYEXck8fYj2
/svQZXsHQ5SSOJRKqVhMnLFHkcjv09bU0kOPYkSntfyDLtmoXqUuozd3sgvV0N3k
Z7piMxvvYekQd+cSGeMKKhiSvyYmDzo+X5Jgm6rvE/0nBcBsPAx40JC+1+3mOBEx
eL3mAcO049DJSO/cgsNyLR3HZKemWfgWvccaF3wPCF9EZHGGXzjErnlms6l2MuVw
ZzhKt4JXaBtQo9IctOuhUtQ7N7lZwHgO1pDTF8hvJLMZtL7EJohnvvnPZdYRlqXj
MxvtzYfD/2kwen2gP+Ub5CX4pmQntwn6Iwd2KUHtyPOqTQFh2dGQyiwYhFq2Fdzr
Vno+QhZXeUqWhzvbwh0J/iOXzBYat+oYB4Bg2YmL6q/jXi+eKzN3fQJergiiBcgn
Pbwmx9Cpy04L2uG5R5ov8fLAEYfoJy9BJp4UlncvusXObqf2pVw+BzWw5MxLKyiA
T4fOVIbGEnEc5vHq9NEix0spfu+G2IMhXRjhkIEcJI4PespDfjoPAyfrJbLoer98
0F4o4pY4pZqpMcfvzYURHuvwjkYb+vOeMRaR8n5LwnyUNxlUebN5JB6rmk7UCLyg
GlmTiTnvRLDT0mOIZQVPBkaosqGHK6CzwuFZeFqTy2X9iw4G80Yfi1Bgpadjgw9c
6kJ8z8oToc3EsOPlTzU/q+JApJTkrP/6dtXaMo91yFcJwKeLl2kZ3rSjiziRvo2r
NbecIx2eFL3Vafdzsp2bcX6GHg0ldNcKi4N/Cq5l+k+nsLKkEO3FcsqcX3mFitFf
HaWa8ZEJ+gQX5VbH4bE2aidu5LM3YYL2RQFe1dkDMyYpgHE1Hj8qEkdfEAFLqc8a
j/hv5VvCTQThFOH/9ql2UhvQY3W3EoI86IKct23Zmc6izvM4aS8gkcMkez85oid9
yLgO0pUBRr/cs1lo0wf/pauFSHEcxP8V+9clTU2uDs8PjAGBIRchaKCT+wGvmEcc
SEPrhcppnOTmmWg5OAxh4fBttEi9UhqY1PveDcb81+2+3w105TPNuSq4fne1JFin
hsyDwVoAj6VKub5FoOJ8SQMH3wt7/OXev8AEJTLIxJlDjB4oLu1OHFCfm+9uNX8g
p87HrL0misJKviBoCSjX3i8XX+UAtyUVvfRcXnvOAXwxts9HL4Aqi0rMdU46R/ln
C9UmvD3mgJzwiE4S4spULvob+oasfyAwaDQGYpOMOoKTQt5UvNgc4NK2rkq+vTMW
j1EP/z5suErY23pkozIsDOW70yWx8V1SQI5Rt2ZK4pdlGcnf9OY5K3+TH7tscfLW
CRzB/jdL6HMfSPNs4xnnRyHLKXPF8GvDVp9qxNwYs3A=
`pragma protect end_protected
