// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VD8AoXJU1ZTA3fXWf3455DHga10UtWl38Rqt0pIO8WWUsKZj5UZkvFZ0N6DZH5va
F459/MhgQiZRkaLoCOO111JP0UTjVafGCg3/Xfb7nyeEbG9HuJagZ0vDjOMa5wo/
hqVBUSVXCpQhHkDbhnEOfJnaUPXGBEYCRmvOkq7vg1E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7104)
IFaubx7bfHE6+SpOB3nzJtgs4g3cipW84NTkT7psTYrdR8AAy5sD/2Ce2SgyHwP4
Sb5HemSd8/6uPTujAUfw1PI9sL1rXor8T95aLRiB1Mpx9JLnzodRS2RQgsNdzQI3
jFYvxEOnzn4IAZIyvjIaBn6WLwnKzOG+h/lDUke4qVucZaJEEJYjSpdQE5p9W+t9
SQVVpXYd4fsSv0WfZRLE/HRUSYXeemjRnRnsCELqhvskZw8UYKJ8o2z8GniIyqP+
KhOEqR1CmdcQsvEpMj1J6QYlW9buFv9I+mt2Umc/SNoGaCigRHHke3eNuiVBgM1d
BZODUtj67v0u8EnQxv1dtqlfL2n6i3IcCMatAEcGQgVvwrtq9snfpbxNlw72ZNIP
i1roJpTj951cx6wjigM1eizF8o0C6/BEF7twfdAFrlWA7Lgas/2FRkJb14cooU3B
hCL1ubzG74t77qlk+awZFFwgohkueyH2X5vUV8jHN0yenBELyHT/+wiDBBFRU9qM
WrEAFixl0tp4VfUVkyLXUMUxltJjwpUu7ADE4QL/DTICtSTfCiIXkoHAUYfxvr4/
jOBN7CoYoucybEbHQvDYpcpmo5a4VTcL0vbuKU11eZ5PiZUaMP4IpIpk8UX6c6Dc
FxcyDx6KsFiyfvDa7VDLQ9stO0OeRrKMQcfpQYpMnbLXIDMZRGcUin11JphKSLYA
wOxRVsqx86jUtBk6q0SBpspXg6Lgpu6cqsWBhpwnjt3GDXsLDOPggpA9TKYhAWEL
6StRyOLQnFasCuO3MgYCCzFJwyuFCnYhU3N2mWfFrBACG2mAgh5T9xMW6cD/Qx2H
YkquZb9eTvF0Xi7c6yahd1U3w+ceTsMUcWxlzlJ+xxG+Kalxq21ND8y37XCSEKXK
rT7QgChcbJV1sMJ8vJyJdlmYsEIiARWmpXM+1WwiI6pkmJP+YAeJxBBMHb6K6wHX
IChc14kf7zoTehozxMo0gzWPObTZwwjwcUkPwJ6uj6FGx4JGfPJzvAka0CCsODgE
IHHjLQoVBA6eCmKypqO2cAmx9zNHy2JqcaHbTEwlLwa0+Y455mVVg2oo+5NSldX6
T+KbXHaeMOaH2Apg8tcmrGfHmLwDj3VqIeotrNqK0HnN7UT2JWZESrSR+l3lwbMk
fjMu0GEGKg4vu+2n4rpz4n2B01aw3pfwYUbj7MSmZ+lz1P+m1zWYOpnFxzblb2jh
WxGm1etznjZwoyS4cjnzITWMdMnL8zw+8wuOiYcvtY8LIxEsyjpaSeeTbj46EuHE
06IZfK8UaUspzpQWCiPWnkxBbmcukxMZ687sg7LaCfEmeJOdzSUM3rWDbV3o7wR8
a36VzR3wIjSuvqxNopBfV8i1nglHqtFtITXRlK170m4lTmyfeihGfCfRwqecf+sI
cgcmj4ji8nfkQ4cF174SED3srtgYgMo1PBq4GOgmVKuTRDvHxiYlie3/cpyhJ6Vw
xFXnAUxSRgGsJx9u9S1BBoFJAh+lY/LDFTn6ldMVh5TIt7sUkFao4sQIlH+8jHs/
JSYn8Io6qSqqQNQTFf05zcNW+l3NpK9QCXSrfn3QvtbYDu/5zW9+KnXUxYbdN/Yc
W4JmyvoQVL94uEk09Mj0qs2ytOoNRtkNSVGPvcgdmH0OyWloi8rWQlX5TTBAhYj7
jh9aAm06g0dAC4H6V4wWv6PErD3YZInhZDq4/0r2i/MTIVwq9lYaZqW76W1+VhQW
y9ZFs3yRh4rGlgEb2yscIJokVF7PsI112vy4EfQV8y/YybP5Sv0GUFeqmJBO5PwY
V9ExLG1YecNJE9vAtf6/o7FoV7EuV31gRFvnHpZmXT6SG4JvHZwDibC1LWoXyxix
lGJ/QnRPZBTfL1sG5q5MfFuBvB0ZYKNfd9jQzm33WLnACfbxlgsVkLJ/5El0jlz/
io/LmFJK+5Si+auWpsswnrPrXHalSEHDEIfVhQ517kvK2DB09DDWDlL9RE0/dUjK
m65XqpcTneWKjzwWmV5WCUiaMw7iYcQsPAr0IjMnYSOlbsaVgrnU5IrHsYc+AiNe
BKWvW8fszplYK7qHMw/clLwMKnmyRrjMW0JR25U3QeO1oJSAb1qXNo7O6zFtSlOm
7ATV8SfkV38pW/d7zmr4xuoxhjkTM8NE45W6QaBkffpnmligGjE0KoaXIprmuwkI
8JpCH3eSCGSlRqs3XWdRg6GQeSBqkEHPeGpKs0YIVGk4j2OF61TXNr2rf9AExMyN
PAI6c0EWxpJyf65duIjHre4T9noRfaLlBUhnQoNLz8VQZfLsoDGj2dICgsNFPlFa
vFiElYZ6N3eRnLScRa7gwdZ8rIUXcRJIr6EjZWIx9Lw/oQW/LcKu9fm2p8zyFmfw
iNTQ3MlVjnGIRRWfHpnGA9TAo/5wZgie1CQhVtRovKkDOVo/Qvf4m7K/iZlZlY1J
8KxY6wf36lQAbrWGILTfrc7hXeZwBNLYSq1WdmCy4mWD2sKE5K1/cMkVTmZ+7jB4
aCbjflXxA1ds/KntSobzRzugd9RIYmP+lb590J4widdZGfbwuOSeKb1pvfDzmf9z
tU+TXcbpzkBRK4Gp+o8HP+Vatfoewk+2tyms4GHsbFQ7vTrBEiG+UKvR00gu/zba
Ibf6WlXHxcR3O50MtdTBKjyuSLrf+nuD5y3dAclnqt493weyf04UaCpVQiZeJfTd
0hmz0nsYU9d6a3JrLfA7GOrUZruXYtXDMoiqPQCOywedCaYnZJQHoUAW1+DULxPg
1jfGYQSPSKHTyUjGbpcMBYA84+opNgZYvubH/nEYMl81S+LmMyfdd7fMNBChIWTQ
maCB5vbDToiPqmONkydTdnA70UTrZJkQcNGT7HMZkLAB31aMUSHzDVPjg1xV+FO/
AJtC7Gd7VXXPFuM1FOAUZbkC4+T75KsWXnhMyDCvOXv37SnXli2kYTIh/2afLAv7
D3NZI1hmwM9YuKE8LdSTuCWsOwfNgCW653gkmxuCrxXAhTDU1RN8ZrJv+ZFPa8wH
TFP4iRmTbgtDtNUQfbGVXHIA1LJTiPKlbQ1oFpvOEafk9HMUs88TTLIna/aZd2xb
vVZjk8SdE4ISSy3MoYbox/pA3qblQ7wkNJMUye3m2T+V/+JKMbSCEiYxNRUbT0+9
zlvQOx7q6rO9Sw5ogBeqzyleYrep9jDdrM8MmqbZl0Iq/zZF1PUiYYCMGXDQOHVL
l2NEN8qgIoCukSwqbGKa7FWFRWPY1wfqQj2RQghLN/XewGSPkYiI6HhmxFmyIFnx
3t73WtT4uwcVpkCqpYzsTXJqD1gfWF2R9Avt2bpW0cutVvgRvvS30dlzNtNOtHnp
v2GY43/3EYH+b+iO2KtwT4ImxRD+XDV1YYQbVgP+Sh9ZstP1IF7HEpbwf7u5rP0I
3mGL68KYlsY9D4n+GFhrYbD1shHPohwRj66CKq4WajLs5SHijhEtUpubO5xmtDkR
1fn4N0tfQoUAHIWn5WvcqqA4885eIncXS+ewCnh0G16LkK2Flv73XVB/j2YeiWVG
5oglglmtjtAky7e5Mqhrs6KuXMsC5aFfskufaiIg6FmyB5OHR5/H9z4nLWGiDMre
jkTTABsitO8N10vr0xprg2yJXJyMe9rc5/Gu1N3dKcwjj4Uu8mlacHPPhZqn4eUv
ZNNDT+3ZD0NpkQoBeUVWS7wBi/Buz2T5TvjS/JlqYExKKo8uFBs0w/4kserNT9J7
ZMQrU6+GH5qL7ERSRs5QC7YERPA3lpzUHpoMlZER3Z7bLU4t/vIVK02Nko4jC9NE
dOUQ49qsIi3V9sgRMAh5cwrer+T2plaPvb2cpNqVWe9tqEQVVFwvupkPD4GGP2og
csLKzITcfC/carTjOy2KSPczcfz0D98hTq3nema44DC81HcnofL0FcPX2V/+AFjI
6Usr4aaBjpr5XokQdiJzL3yxKLMEX4PcTTnQZNMzU9NEiB8rpy972zHsyuT/9WOD
Hq6zMrf+bVkHDddGfSS6XS8PdszE0VcieFX1ZslLxzHmYH51Oifd3I6mHFzufMR7
Gr5RHZqJeM7X3oTll/Gb6YNaOWbg6IeMLuroplvfXmP6jhN8HLAkPcPxwhBlFbly
FZiTG8wOtxr2ZbYFrP4tu570PU5ZbxtkKsBNewnM5b6fmlsHdO1QchnxaYFQkOuk
TdM7L0Uirc74DVmG2MrQwcIFcUDkO8CwQ/+EZuEaphNxjuDcrM+B1Figfck8vIQ6
dtcJ6MyzVD7D1jyyCFbE3ai8BDRFyGPgpFjv42SZe0lOuDubJ26hr5/V4RuVqmnR
BuQXCRuMMjJN7Hf3/0lPdciRr+BWrSZUM1eLgIvlJuzwKj+/KoxYP/8yyr7IB/Ec
SGXTTEtwZ2cgFDXRcoyY4KSJh0mxa3byHAkYpEZ/WHWmcHl38xeNsk7QFGuYp1Zd
9WpHBaAB/Q/W6MwFbvw1xmUmDC+kFmx2rp8jK6cEmmIKKi9XMay1qB1RWq2wHFa+
25y07rrrUm9d4E6zKqCFzFfqZ7dNYWinAdTy5BDd0EjeMQorBM3K4LUGDkeSpgjv
s6G2enJuFXPcfm9RwpMRoXJui30PAHXOzA+o0KiZ5703a3x7g5y1o0ObeN+3fEs6
EVzI89lsitnwFmkGfOYW7fPH2C4nrNsovE7C8r5pBYX0tspW3gy0Qf/EFTGOBw9K
DnJ75dAl0LLQnkNSKJJac2OFK0awrsPwwqpRJ3QFWT+ZWAC3fyEmIUJPp92cfXwh
Zt2vBFKJ75D7EQRN3naiCPvubbFI+IzMRIC3ZuVYlA4hiWmXolFruxkKC73xrwNp
1ywegpVwCvopP7cjOjkPa38RGqDkfiex22XEYTFqa9AnuC5hJs6yqip1ipUvbhsJ
47TP3pnzFKwK1S5V6SNUIunfDLn/+FX5czKXRBSDGiy+7o1LA3PacEc2BApAqndF
8oJhFBgMluBZ5YxfNf4NvZOYs0roCHqHVtzw1ibeQ17Zv5CqLd75W17skF2IP0Zz
KIqEWIVy10yVUiPMD/QvRFY3TgqGSC84srId8DF1L6/B79j09G6S4yx2TYaWIQNo
ZuvRbAqUndP9BltOqfVgaCbrwoQUdxxIIshjnkBrgP95/4nERcK+27cmTIoWGFAR
1a28v2C3DddlxYstH8pT+NIoV96lMRA6sGgq/1g89l/k1X4y1AXJPuD6snRP8Zla
64eHZOGSjEo+u2CbDthCMP2H1d1N4OWA62J9lFsqInP9PEU6XyUVPRwWhHxXPWq5
ou5Wtc4nLxVyUUeW1jh8hA2OmtLUtPuaVUi26HEJDw+9V+FhRqUuLgV+7NCvscmk
JMvc6Rs2AtNGP0nO0NZlSXJv19rdP40hffdeHzdmJ2taFcR0/e+eXf5alXgxpNsr
zXpMUhzyaoHLuh5lynhQn7n0mjqrxz56RFxKHN290d4uScLJjtXA0CD8X5bTwV2Q
moYq92HkIQz/mWdWoGmqWKs+nODkwQxIVDRyNyGukNJND9TYpwfI5DUM920BUupT
D+VObmKV5w4HWCY8cLSckSMZa9co2SZ4nSlD7Xyxy31Gcpem5gkYztuyv2ePMPIM
wAT3CylFc2OREQyq5qDYWkSku2NfU7Mo0bNIhXARdefYSehDOf1G5XQMKumGvIU/
6+8h2vaVqeAvbA9xW3QmRJwRfQTzz+8QnsNu/aC0CptY0lCKxTe0OJ7VK+QtiDi8
Hqpg19jT/d7sEhUvdmu20MWpVhxGbwrqCQkJ94KN0REm/n1m33kIQi3lm3u9/3zT
/2SY6RfZ4tbpS0YHVXgh2twlcoKkQIrAMp7uwvriLa9iKhW+67BiGHxUW+rMgmew
xPeXfECuTUL3l7FEVn3cASe4204nw693nk2SXQW/Em7lJSV+VgWlIVuB/IXCXpWp
x8zCSWD1MP6xlK9l67YNR38736dksYEfwfIfAEDigOJtFxhdrp9Oj+s6o8ku/efl
yLZqcq5E7N7ZVhWC7AnpU+cwN3036L/jZKf3xFzpcl8oRp6yDKEBEoVYh3zSzduK
YDPP4Rgin2tVQbtxIbw/pppIUNh+3YvjDhPTM3rVxYNDILKosnDRhynEIKhtdxCR
JcwWvnKLwxyli/6V8iQeIVsKoQcStqamJdHbAht23Vxp1x/AjnDgA7FapjO4W0Gx
An6J12Y+nHltXkn2GR1gIlU/9Xx6UPylgeKMM5xWW8oGcrky6dgdtVtQpOco5BYq
Kx1xZTB/GBO1fkN/5hrfLrqiOOWIZRA6r32J7frCwQxuo05vR6DiAp1PRDzVU2hK
aXmvoVyXPY7l+kUtTCFrJoCWciNhsUfSMmS3JadFP++Yxz8BejYog5Cer++IwzKy
puu2C6TeRcOfGF9+ZmYJRI4QKD9nAwZes9EogT9D63lPwSVk0aRB0z4QA1LVDm3n
p6hdObzYD3BULOeaaSr9tDzvCnZHoNRyz/jqfgCdD5GIrdjcd/6H51D3MlQvypfP
jTZd5TTebIKmSbtmmLxj9WVl8KvKTEDyiK4MFfKysR2uiQaTaFSMztLjQCQoF6h7
cYyIx0qevPmT0TYgRRJ5Q5EhU/mB/asV5gmEuiQDsD5xOCjGFEo6irn5+dlk8dO9
rqln+TnsjthHWlyUioXt6UfYNCm40uO2J7269o0paBgerO5U0O4zkI2dopj9/vHN
lcEK4wh4TQvXRL5kQWIE/q6hJS5TfTpdxLiD4ttXhK/ho6hc78fynTsWzKQ9rgC0
X4tbYSbRhcI9eTxf2GQ0thidA1HLxmfMQQ4oevOk5InAzxM57a3S1A1iK4jPNSNq
h+s8afyWFHhTRRSsZCFBZGMmel5YqohF9FXAZTaQUStTXLWrrBFboSly0KXUWRZe
HuJGV5pUkVEiZvYrOAw5s7k8v34OXt3UckyJm1jgce+Dqhq5xyOnTAR+1IUXakjc
HfhQerNw9k16RdImCCw4t3AEw4qN5GwgPT39IR4kn7A9Ny5kEfFBSX6InLUBTRa4
1BxB4giQQu01bqC5wEUg8SNaFUTAXnE5GvYrUQ9V7eidNxbuCsJd0L0B3MTUx07d
JvIMd0Jpel1+aQp6IjEoLXw4RDd4Qsnc4U6WPV1mq1TnSIxYWi1NBzQRnCSXYEQ5
H9KzZ878P8RzvaYyzCVWtaYV0DVoCGpHmeEByZ5E5ym/mMXSUZj6Foj6VCGHH53B
ybBpIBH7TW6TPzNY0a3NRYCVTESb16tQzpQE+u+ulz3trA2CModdtMnu/HQQCcXr
1VLiz+gUMnkt1iET1dlgZqeVC/HMqOAG+lueLVw7EVDL6Zjb7og9wq1M5lTcXsTc
ARjgv+f+NyWe69G0GwtC8xqlS7Td6jB3wTXlob2V2Yb06QPuaZYM2AXxhQQOrYcV
84VP2FI+fSQr7hF+h5TB+BjhOhPmTgUbJFJaAC64cv5JXl8Ry7EKL77UIG5SkRmf
YoSK0ol2EEMf+d53eUpf/Rej7LJW+Du2bO9z+EodudIPJX6U0GXSM4CQacqLjzoh
vZDynp/A66c0GJoIrv/Uo8yR7eRXxUOwGFgbe9MQ04Axj+Y1I+4PxWO2cSpPl6gd
manjiLGYuXgrjEQ3ompY7/sPT0AOR5B6LhHJaIP8F02nnXYKqbARgh1mg3mq5Gyr
jGea+uzxY5/x6iddHY3XNewmkRk8hUPHtfS3Cao6RpmAjs1PP4NkpumRz+4EFT4V
7Vgp7w4RWa4X3JoGhKfI38krEgOnUvC5e2LykhFjtzGbWZUGtYSvY74ZBpWcNcfk
y/XArnys2zd7AWdntclZmnE0HqjwIk5zENzcJrdcR5B0tiDvrNYz0It5CHt9c2ig
SOftihX8F9p0P6sXNfirQSi56x59wTgscagYqWzc17v+4MjTdrCq3A4OErqRcFHz
dl5aTV+q0hR99zT09j6W+vTTFnLEarc+sBu661bJ3I68ypble+XHbJEj3X3J2TbO
aU9w9q/xs+ZxH4nbUb0+tZeGfI5lder65F/eVit9+TKdO3goo62JQPZ8ZckNCv+9
0QkTGmWGHnT0NvFYbwsGbM6SaxVSKcz2o2PigmbDH70k28jTFFUQB4MNunAe571A
y1BsbzfhMxJMFzCb0kx3fS1fTHde0squDCQXjsA2IZb60zt9YyymLrjjwr9+WXii
/6iG5nnU7qTKc5M9qWfBO2mFeByaGEQ+xV4RhYX3p0p13xRNQcHKMZ2d2daokzyS
8I4hI6d4uYlrlxbjb6v2lCJo8NXkTZoq5puX4/ZDMF00tyeeK1S2kshNRa7JU6H6
4/dU6drXJSEXjuV+bgjQQWfc89xzerWm306XUNZ7HCUt9S9c8x7uypC9FyJPfmzZ
iysqx9n7ps5V2qZySP0K1RKwPZ4nWZMrVYw3pk5ix6o+0Q41FAKVNswisx7gDnJe
Rx3sM/Y6XfbsPQlrIYFU80j0g6hTMsOu799WBAoHc3oFWjZHDogzJnWSttVmwgr3
IkfuGReC8cJ7otW1DkCTQqn5jfvsZ/QeLjS8nCtKWJDT+xFVYewHIJPlndRtG8wo
dkyVeXDKdtwvLhKOxzkR6b0XHeknlgHyoMpUJf7X34O6ZxOBdpMpUxii1y+3SD0y
SDF4PB8gqRqOriCW+Vbp4tw0bxvVc/JoQdfcsD2zFkeNhcMpV7aGRzw1hT5ZzjJl
entbdyhro0r6GO+TkZARAJAB5HgPKz8YgnRIzStnMQQ6MWzzBes0x3Qe4ekSxrB8
oAlig9Jpty5iA84vniN3XidB3AXhd17rVOAxvUd969oUdY9dg9WDgJOVWLQ37oG6
C36jh5vhMieCAnQocmsVf4KfNrrbFl3So/2bNG8euYRtd8IR5i99s0biL8hDjpMc
p8QP/atyixLp5hnqA7l7RljAdnCmdvvW2+GQQnWgwEuGOCwFzDD1eZ0RVX5AvPBT
uLeAbvIcoQZY55zK02EPLYTJOva6d3D/zseqQEk2581bic/+FVhola8mcVjbra6b
5lQwrdKVJykgCWXuk+POeqnAL4rgFTQ72hDaRn8AFmdEV7dYbSs/LFR470avrHWt
IuT5FY0r3teEGGexdfv6KrGEnYB4EJQJ0H9un6KLw2GpW1cWjbin2j37je5R/Hh3
BYI/vUrjAR3vjdDRmCfeYxYDy5b6vZRltymEohulWXqYCKIvLcBELvSjBEEwNuhU
89HRGQDv0CEu/vsIDhDJUowEDF0n+BGn4w2Ijf7Y7HjgR2RMwmnR8WotG1FtDnnA
TwvaNQOpNUHUDTeX0irKf5lvtDC6z4SpfbAnDxjCPuhILcV1Abpf7PTQUsZ/s5XQ
x/ji3Yv8QxzTkDTd5I0AWdjIfMXcIvEfu6VX6QJcQvw0lqacozYc0GSVXfBJ4O/7
/jWP1Z0XiEWs/newpon+jc1cDrxQyB2KEJUyHUVLmrfm1M42dgCQL95fWc2WFqwr
UaoTvHuJCxnTPWp8Qf3leueRBECN5XJOjIr1JDe4hZFFl0mIXmSImB5zNKhY9p4Y
`pragma protect end_protected
