// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.1
// ALTERA_TIMESTAMP:Thu Dec  4 07:39:48 PST 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aa93ieytm0dqaor5k1/RdkEGw42n48CNeMgydEUKBSJbnIufQlkUe+t9Nr985Kz1
IvvC7JmfPBl5tzeEti1ebl37ha8sF2p0sBtUUoYz9Hm1qrXhs6C14TbUgWwPw/OY
RdPZ/P+Mq/8GvnYvdfw5vBBSpM8j1FXnQxvSicaN+7s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31136)
Awj/ouOzF1MFWxQf7IbnN4Rgs6qxr+kdSXUcoDUNKkX3S3cr51oPlNCxMWvdR9nP
iYC75vtuxOKnrDOcAcrBDWkMuRJ915mW1GZcTuCTKHk1UHlSgeT/NYHGjL+T7Nii
MmCMo1Rzz7SEtcTAlQrQWYjQ8zDMJPc2AUbMUqOYI3Kq1eAALukWUqmW1qirIPsZ
GcGBuCgJl3mbmo3v46h5J01yc3l4Bx5fMb3w0u3Dy3+g6zlo3Y2ob/3l6lG96pj6
AVNuNMJl9r+9cNfB6VPmzQ/WGpqKNEPpM0sf/9sUbhO/DfgLnqsDZ0st8bn7hPC9
QMaARj0FCLIrW7lrnaYdP+xy8qu6tRxHmdJdpUuypQoZKnYNyJMKE2QLx1HTzevl
p57qNQ70JFSUSfZC3qcy1EOGRS9Q8scsppsJGf/F0LLpQ7zRBkyvJ1nlytHV4q4X
6N6IFe62ltSNprXN4T7+sU/hozkVWb1JYMR9lPsk6BY4odZfA6DAFrJSeN8hcmNL
lunnSvh8szcmrhajY1MzCZdL5g8Sj+uUwbHQXSO2CB2WicKVg5OUMiyR4pAwDUsW
to3i8laoIoyOp0Ji/3igTJJxMnp4z8FT6LdK/H67Mz37boLYNgu8HBqyP0/Uc9l+
WPw/0Wp3Evcw0NFgMSZQyKhUZKoez9QtlEvhuZ/2UcKkUvPlXWbLtpN3sV023xie
dvQHyAkBmvNPaztt2zqUjAC+fZGEww++nKxfp/FKu6JTfP8LFtUpRieo5oZKPp6O
VR55jqeW+50mUQiKO3+62MUOljj7EBVWcdLc4AEfdGs4I+cJWOBa940ixeeQQc9F
qenh5o4oB2dL1p8BM+G7lUH4ikvJ4VMXFIreJVdYx+2p14PDu5S87dEEuDlvpLCt
2G8sXS3zbqX2xp7Ce2Fp5fLSFnn5p02OQSaxp9oPARV7Mnb0ApiajFGYH5kGQUFl
mT8+oh5Kd5UMUQVf+3eVM3unDL704fzCGEsQC44j2LqIIhM/yJz4+FdvzbUf+0Yh
718Spvufz/ctjmk8zbq5bLSMnjJpQ7AF5c8KGnAMhGcZuiZjQ1RsvsAldVKJ+EeI
H+nO0yPy0NFODGVu24bdwTklr376IIoCh7tsEYbLHFqQYlu+Hhpv4J9RiLdwobZE
5CEtN1IyeO666IiVeUM7z57pbGnN4OFsdpm/FiCZBMLkEq0RMg+DDGXFGtzw+bnF
O/ze+SRax86mnrZMKMi6ADDxVq/+x5vfkbBGzLxysTVP/E6NAqWoP5qb8fg5LGjR
UzqoO/UrmLrZ5M6+1R/H9nBEGEQPkmMxyY/btQ/2aGOx/e8pY95o8f6P80TO6RBy
0IQYY3jD1rCABEu/o5WhENo+9e2yZcsrZ8Fkoc1Lc2oPbZFzdCMeRClZp3ij9GQ6
1MEIHoDyoGpz9p0EfhViEpnVtINaApTA6Ec1aaw/wor78ppxiJXjVweG5yH2h9Rq
O8dmRvzAirxtOaxsOoAVV+EFh4n2vtZEyfq+3MBx4aYmnHYu69+jgkh+Oi5FUbxv
FiCLfM3Z3V+nNi7rtaKzkLw8Fo5Dq0yLlVRSRYQwV98otAQhzoG0su08scuZ8RnI
e2js4EXrTBFtLobqdXpC2gCWLKBT/hKfTsJZPmoO0VF+3bMavLocZj+hM3L81DOB
HsCe8RW+3ynKs3cQ7GY3hGlpn8Gk2k6Py4iEOeWOOJksoX68GyZWf/qu9f5VwAkN
Yhixh0wTzQDxJ3+9opG0gzGpgZx1mN7oMk4ROmikA4zxmbt9N7Ie5WEPm+ypDD31
lCtSrpvsN7vD1QB4GxuuXAXjUcLl/UggZaSIFs1zI1DqLQlhYNovnd9ddi08oP0S
6YX9kRnZ6BzDifJRal2GzC3k7brGU1on749tMMehJMBEG8Yht2f7+8t+aJyGW278
Hm6gMaWB9cqp63OVk+5OdRqj8utGB3sxM1MD6dToLTEIEmd/S8fBT21oBCLZoNFw
cv+rXBgijZxqboLJTU9r/4SherwTh0WTIxksF6menTc0yKSFPfH+Dstx6D3M2Vy1
AE9p1OdveSGH1Hk3C4y71pk9LRwhQrXbxMkieybY/iIRkUZJsR/7l1jnpedOUPQW
y9EyFiakF0hD5M5usZoKtTixHudTtcYI5HriSu8eKRsFvRKkpwgA1rwE/JObRGpO
hQhSX2L+s1h4usCwKphbRoAQU9/6QNK2+lf/2MVsPyPu2I5AnLkG7jfR/eMlKkF+
/V1+SPzmb+ZrgUpDTIQI7YiW3p+J7g5ifzMWGMAfoqHNDEiaL00iERdNzCPObl9E
rvxhz9Q246tPq+d/qVBDFggIavKxduqFw96ow+AJO16uv9BEL6GMk3LrBbOzHNBM
rRc1IcRgEQTdyIllxR1/C7HpX0l2AWzD8AObedj08j7NLWXa7beoCZLIUC1ntf9l
6CWKAMEaz9ed7RO11a8l4V24s2X7XDVpwM+87ZJ4z0/77nphk3GSeWchipRDgOZ2
rBjlh0z2hTe6//Ok4oSZyHHKXHD4eekwGwbCWq5WPWYWRKDgsPlio/CQEWI4+gxw
vtTzvFTpgGfViWzBbNvb1j8vZTCcIwdWJUQTMA6oK18A/3rnQgiTvAh9TbIDKqbM
iMXJ2Z54HyBCP8b15yFfLNYhd83GcqJvQqiu11OO36W7ni3W1a9Gt37pS03PM4mE
s4nD+e9AjWFjiKXHIazZ+rwm7e437xdhDQ05d1wg5clS7PDpbxwP+8aFCrqJ05//
yRu5w2kfHKgJl2CQbxqXO5/OutKyJuJPNVMJwzItStq7KPih3d2LOvHLQoyT6Gnn
9H96gDGtdgFMb3oWlnHjZvtMgsFZwCR8xO+MDSQdm12mJGATUSKdX4OVzK3U+WiP
wls72Ra1btRv+vEBldpdnbKFdMGiPumisp1+G8RAl0TgwQwTJO4dIHrFrPeuq8R5
iHViDPjYh/Kc8MpjrzLPsfjgWPFy5A882ivczXylY4q4+xvtgr47aXS891ohdCXQ
LR6FIIPqh8oT7GTRa48ciKACRwBKbgS/Ewcb4KMHUXjNnQ1mQDRP9u/7PfoNnBaH
MPSXees/ARklnp2amz2DOSDhn13/88gxSKFATW6ET7JVovaJZtY1Z6F5iEn3yp80
SFb3KpICH3jdbtrGDS7NOBG31tDomZ5IRNvDCtwibCs3rnbiTC5p/WJ0A0223zu3
YxJn1Rilo0OR8yBAlkqf1x5gxUEonA7C6E4LaCkP7nS/ClOhAk1jFj4pbXWrycDh
+ablhNQ92xwKlUBGnjeqgrYb0ZbJcOXOJCXdrYFT/6HWBcuwkeGee0AWMhMNddzJ
ri1lg8KkX5TO/YxEa5HMVIflGIiyrx9lz44G8KCeOMTC15NoFIRh7Hlk/HIR4DYJ
15sCx1Fp88KnQDpPwoProFYx/Up4Z0VlIj7Nf5QAmM9D1nEMQAqeGmunbVEGwK3t
AJUY61zjoro6AJAAkojVziaOOHVGp1iON683FR5A/WQxv8aSsjr/KZ1TDsjuYKO5
Eci9+HEmnqOw6JtyUDI2dqZHa10+E6fXIms4dD7yxTIoN+sExn2ZHydqBa+e3UAw
PUyTsoD0B6HF5brblIKSwnPzJP36c3i/bxF1vAEo5CX5Ok1qYXWPcEZx4Qm/83Pk
isqVBUpL9KVKghtreuRIyhgrQv5xQRtJ45Gn5JmYpBO8VKw9E3q8HoU9pC+C39A0
UneGrpDkiwcTE+oAmziIShyiIX2GtJRmjOjfJbOm8etlTViNprt9ZCG7PbHEWagq
+K8W1MORGoJbFTkDFuDtU9E07jFm7uyw/Z+xomjGUJT7GxiiOjJ7c6JlnsIgP623
OXndmLKrZM+E3iQ4qTnagsOtpqfyMZBvbLu+L1en1Oj74GWaun+f6E2wspr3gkcV
V9UaRqOBTpOIopOFIVfOTHkyyJ32GJ+z1LrQfm+HaGLDf95/bjgoXCaCUdjObt0+
vI1y4NS09BWjFCYyh/5mUzed1XezrYsBOxWpJxQm1/+cvgTIkPnszwNEtLkeOtO2
/LoNIhEEiKgCcMMxbHDhxZQ4LPdSyCrVvA1DCpDS/v98x3LxEfjz2CODJfSClOm3
gTPEpzjP6MjhjPrtUHo6fxhbvHlXJWVXBnQsSNymEAo3WpA5Lz6VPiLzkZUQ/Fn7
OxdybqzrArmpkHCUrkKTXFG3qbQhPeRtganoLEtx7k1iqaVfhLFyjkrdaJ2e/NWy
JaUECiEGrvAxvrAwnXz5/QuPSwMg95TidPnU5qFJdcst/t/GpbE7dHzSyBtrPf4x
rhxuGWWvMwsds7zYAOd9ZQor10005IF44zgejhiTuWZKCWkv51GiNlT8nT6Okwod
xRoDVDmjIwZERkYISbeCWqsIDP+Wjm9F1fhg5a+iYoFZOSnab4Lhz59ivyqDs5yK
IGCmMu4DWGMttpNNKr+239RY/GN31XVtoq23rR4rNfMTVZ//sk41acMpzgT5r9/3
7JrDoyQ7aZ8jaxS8ak3GqiOBpQQptpkv3YoFFArevh9hJN62/EBvMEf7JL/K9fXS
ySulG7CQlNMXyYCackWKjk7pCjgZ9/thShZE0duMd4F89bETYK10JoK7+Yf5fm6R
U3m4fbobHQeWiPO8Re7C73AwgdjKRd2kD9av20DpPFtRn+/jgUGZxrdlo/wKxrPV
JnaoROIPqmAlgdDPkigX9x0eVocyrSUursYn5euUX5FuwfOt1Y6+i4PhoP8cYSOo
qSyAxBS+HPPTL/cPSqdUgyxCvyVOElfmika3TAOm3TyMavq3WDWpcWVZZvdGwL3m
oSaKzD3LhgKi4/brdryLgmsq1fhGUXGQEY0pVPyO+/cOI/CzfI6wvRDotXTznOcP
g4RTEVoBhgSb9oagePM68xmmKNEUHj5SlfJZwPA2ECddpYWc3E/F6FV9+PNXwQd+
fwCv5X6vxYmVW2By9Uhj8sET87g4HFNGr9+27Gbn+/pDxyBILbh6Gog9PoKDGkYp
X9ed5+sUd+qY7wlT+TJnKIh9w80jdYmjdTYCUpLYcfRZUBUu/g+bV5R8HNHlyhIA
neHrXh+q6fuNbdI2oG48JvSePsMY3rRtsCpRD/pHK0V9TdwAVyOgto/z+a22Y4bc
1gX9W2pKh7keXzljsICszu3Hp3fBrV9w22lK55igjdcS28kslrKIoSptlXkrTnNh
1Vnoe4eiCqkgR0pxEewiM3WJxoXUpTN1K5C6bvW6jUSRJVVBQZiba2G3/sFoD1gc
Q0B3ZhuPM8VOtxjDBuDCE9Z5AQqWLwAjoMQVLppiajEgVcCon8eQMHLSZvwk0hyq
5KGhBuHmkaEamkEp8lpdMJUX+beBxX/+vovn3JptikWQx9GVMo9i7L9cYUvKSadJ
D/Jg7FpodIones8e8RAnmzJDeempT0tBIL5NElnX+SygOlqoD2N/B+05vokj2paL
UVzKniTq+aQ95ggivSUhZiidgECpzo71MPRy/7/Fa56FYGe4aQ6CcQCNHl5ZMl9I
JNLIn1YxywBrq0X5JTqfeWgewlGTPzuxFSE5UATvXNwvpk8quI5dtHqJ60kWs6r0
MJcoR87kwDboF9NK+bZQVembMuu1xAd83zGUwl/hIGseolwOYXCV2UjBC95lnsF6
+0LWX+BQr3/tsLixlxRDEegj2v0fSE5C/3tFCCy17F3aipV9TBL8/XjbU4s7cIQ8
QD4OmzdzGPl3+uTJp76VZ7iHQxJQG375VLjoBZAD42nFHulhLf8lwpxWR5zvZeva
oJgAXflqStbXIosJMVUNg78Idn3xCWQCJBIJ3mAon0TMuwD+1xusxM32uH+qmf9h
oy7taaESgxq/aqQraAQSRG77xZNWw22i/pMJkDNeA8j/wNmoB1DexzzuOhpTO0uX
wgJgdpGWz4RtYrYmvpWFNA1AzVXRVmdo5iGUCR9IfsTIzvg8sXZNfjCPpM1xPWQD
oavtUsCi7v0a7YjHVky5c81M9OdhpVCq58lY1foCpF+opyaF2QkHY+DjqvYoOQyq
k+oScxM455rNDSC89uybDXXdHf/D3YHXDbJGvcG2fxIndi2+3VY9gxnfWtjwzBki
0ROPEy3S07pkAwk72/sDoSl629ctEH9rGlMzO7Fh8PskeL/D78nb4ngGh3Jn8Uy/
IoDdMR+EBLGbQAnELgmpU9weZN5peOTbJeRK0DK7WxC4J5c8144XdOTTmajBa9ui
1mBBg5O3vq+6YUz3srlHjiXiZC/nLYhF/ASq/bSFaZC4shwTQdgF5D6rE6Ol4QQt
lqHPTOLICm2N02fpAyEqs+cDYU5mDCCI/m0pEAHoby3qgazSTGp/qXgy6hW8ZekC
TFsEyEylg0ZtCZ5ov8yogcs8bzqgv1rM2ukLTk+bpW1JiRCSx0AIYwscIF+bVQbM
+F8a+5P2Iq5Mj5e7Y+BC3MYjmrOHtFtVJT4oBEw4JI2ldPoGY3Vd/8dtIWR4d1lu
Knsl347tdAQ/PQGZDc8uJtft1K8CAOYPb1fY5izGK6Fdy3Y/ZZbfILqaml8jAExf
mYedUNQsNQ1xHYpL7Zlg9vzZhu765KiZMzJqwzOaLSgl2euQKHamAEEipzFg4eap
+1hH35Bgyi85eZuaty2oXNcKyDfhM/ioAN+0AMCfidurX6UUIUXkWwedP/Gpcslw
X9mao5IVClmw/hFynLI8GM7Aiaj1X0JPKZa2ZRMuBopzk7R7BIQRCrNrbyD7qmec
gNaDxGQXLgzvX6ApM/8Lpn860cgthSdc+Oxsl7DL1TTo7UF790PdlZX7TpzGa8PW
7KJjkyo0p9VUJqKNWGLVFKTz53gHnSShpPB3uxFnH0U7GeIyo+VpohkqkOv6kzxn
eU/hH63uMek203oOayMx4l1oph46u5umuenyMhVJNdvRuFfMtAOn4GWvt3UsgO9J
RESm2eG2SV8gTOx1QTjPKYJy8BU8XVnq2Lg3ocogOl2nyDRM7GZ7cotSzKtu+YQX
cLiwRUhbVCTCxsr/RMUsihU9hbbUMsnXZGHhRwPDHJMR/irtq+mo0CRIxIOdZE12
HzAj4SI9z9Ejiv+TUJperlVmYucyiJPsm2GXAcTIiFdj752eLHkZux3n1N15G3UD
lbO7k6BV8m9V0qgMRibAdYCdzB4+ZdHnreIkeW89HhGI8QtjRXtNbvrIwpr+/TlW
vCarsnjp4YDAiOh5LvC7wBDgBSEgw07FlA+0h14kEYeoJWqcWZDwRXy56aqXjRMn
lnFN4yN6z5vV7oYHbm1CKTAkvrF73uK/UbHc9i9UCI3/V8yq3zOFQjA+w6BeDeE1
XpxvZPTo6jcZQUYpszu5CBpGX+H9BxVWGcU9vQRoUxi6O2tUjMymcrB07vEVlZcb
NoP2jFXK2nbnDBGjAgfs+0S7LhL72BDyik1tLIlTviZhZsQeWGt0Cro3+khDyIYq
hSUChw416N73tXA6aLUmOr/HlRP+L3GFQgf/p9U2tMVAa7c3eqvYrk/Brq+yW63G
u4dXcn+LF1mth3Qufxv0gZOGFkZO2vLMxvpvQRP1hzP5my4tpYnGfrWhadMx/aIa
ywOd5f1yk297bNTdldF2+dkxb46yQnA//8wydJBG9Bs9m6UQvcgG3PtEUayOyJNJ
NxDzS2+X/iNqAVuCxakw0X/2p8bjkGdt2wuWy3d4IrRYBY+FNMUMvHj6P5NTDHbp
N55AyArkRD6ZY53pYJfuSDW6dXN3Rz+iKLqEwrT6piBH3fxNKznf6QSYX+75n4nT
P1JwT/5Tt/03lZrRqpo9Lxi568JrSsc8r7xMyN24ykeRM8XJCDMwUBHejbK4A9+D
LgsXYnoC5E8obKrKPfo79SB9YGTguIjE+V9YLomoQU/7wp8s36jqs5CuM3MTBNHq
JmNNdXKKIiOfvGqwf/8ut49i1MQkCLWuDN+WhKWidnawE9e27wuTX46HuMX4dEkL
d0QOnzZ4MULhUbuD140buhyJswoTI3pmvpXFZsOLQZhfeP3Lvq8wmgmk1sMrW09L
6D+01Zp6MpIGPAQg6t5JCXjVbaKIqD3+2t6eeTqc5vPkcDyCcWO7ChvAG9FB8Bbq
TX4D52X8NxTLmfdIHLxmcprkjxvExZcVbWTz0P0JxHyN/2+pZH7Yva36AMh2F29U
VjD3oqajrCOnYLznwqD2dT4gJwt/QDjSV/3iHvkVOb3vSNhxY9QZhZUQbxemkiWA
MRb9ADqL1Yzcmdgfbr/JyNH88w5bCAURlbLUGg5SiCp1gk1c1qWjc4aK9H7kZtxc
8fI2gFcclPRzYr1WDsbzSVQYqDKa9N1TlUlNiu0SRXF6BSkUj0BqXf5d5EYO6tOM
vQJlPu6zNhpiYCX3kngRp8XcgynBlREVxABfkGSgnxCPmOMX/Y+zy7XdJfeBrDTU
trsZmYt3vT2YzLi5pvyxcbIXOxMSbdjYCSKNDw1LJOmZFBs8TpUob736hIdrdNeB
q/nhLAZx8CuhMdcX7dzq/wBo01HRYs9RCTy6ZlxBYBFM6+rhHeoWh93ZzNDrAS/0
39NdgGmnr2iNF8VTT8XYsmG+k/DLNyD5xenRYAI+4LX1mVN88OwgR5PnNos4VAf5
iNfZoetZGYEpxYChke7+zghm0UrimPye1/f7Cg2a59heom05htmUPYUhqharQp91
SRz0B8VjTSaxKdRyksBazVWjvN0LlnJKHFr5gC/Xb0ZZFQmkBzR9fGh778Z+U1oY
GWYq2jmQtFuKVox+oTHkHZkOmY1pz2iTSOI38YBTMF9AoOin+hOlryPnuWaEkyeT
X9SaQlp2VZ3AN2bke/j40HiWiVBcmD7/nmsOk6iRxpyylaHxVg2l1pNC4dfU8UOh
iIpgzRFUdP37RgLdhAepSYRB9CN2B7JnplQfHb1GH2glTLKYaAQAkSu2Lvt2Bl9V
zDT8M5rVB9WJ7gFdqJrEPN8MyhNsxUqTz4M3sXCtwOk/RcQUkG2yP7kv0Did2X53
v3ZRKx4FbtBTd+GeormLS+ZodDKH4E1EKGH7gI0wVDMv7qAhJM9dUQbPmtoTjL+W
o7IdWW7H2djTAqHEwvU2dkjZ9uz3ujxVuYARZcgcXLMagBMVhxs5tCY7mf+18K+4
S/mG3Vj5td6A1Y4Q6QsqIfEaEKUM4fOjDw291gApF6rarxDQTJe8fQwPIgdB8bUh
/EKm6RVLHkegxL3BPlK7fWkP1mSE4otHqk8cnBwm76N9DL6iunv5SGAJyVGdPGs5
jZ+Z2rgG+bLJdJWk6Gts0OK3AGyJ+H1cgCasUV90rensfVU3EAswjYAVX9oYiw2o
dhrVGGkd6qVCrC4dCLDFDUvXLR0tOlU8eQmb4sjfoPowI7FTLIg9oQI2/dJ9pYPD
HhdWGzUm/fxqVKJKfec2F4OGgxdX4RGg2xwrCZcRjiE7dHeQHm11R/K6OyO8IvZA
iXZIZOuhOAuLVDOoIWvxdlMPV3YSfmgqZmuNPm1XAliFavsIZp6MNDVS8auZyX4T
pNG1jMk6po9Hd4SfeMzRoTeO3jDGd3uAKKHTnvcHGT3mdB8EwZAdpmK+UKLegSsw
EyKxFEr99Y1np8zWFnz0tOM0YSGQHdpMgkRHG+/yXtzucOuOi3fkzqRghLpnE10G
KSqZvuI8PHSEAb/5g1SaTczpHoCt3A03TwwFB5oW/+4l0ul9r/BDbX2gAUNW5Fb2
d18pYuofqvOP8nOrKH9P0YRQ+wdBi/saMiKTctxmihXgl0EBGsx3YbVogs1iixFn
2W282XiMUTtljg9kHEfof4AkgE7XsXcQBxeEroV1o62aYR2hqpmP9/HyePxAd/lf
RBgVGeKPuxQRGYoDingmR8S8SLT9Uun46kg2/xDYcnhr7y1n0PpsfpJZHNEGJeYO
n4bNkdt2OQfSUesv55T4Vv/6gd7m3D4R/KLqvMWgcOaODADEcFcM0Lo5MG4NXXYZ
JGosuEHgdVyKobNfucCXKSz0pmqWjXMQNNpOaRjogAHDdD64DZrnZDyiHHj3K2Ta
l0NQvZOzz8PIohKaijtvoNxFifCMPSNeErWFXzHp/rgpCd8bE/AxTyXlvKmmwnQa
nzXWNDi7ptWh0I/+5oznL0CnRduPXQZAjfY98XNdM+G6nnDJ1NYbs2yQCdkYU5wO
62/XnRLM3+gNnDPRmodcW6BlY3KE/0ISFB+gR086AZskr4fOkxDV7w7l5XOsNI0a
iOWMds7vNDTZxxsC9w2NihBd6VnuiIYtktoTe531n3uDFd/XYryo7iqt1id3mXCJ
Gdo+btuhD7hzYvEmtkhw5+tugNU622mFd1m5oIoWPukNK5D2BJdTIVxS5SLDCJrZ
iHc85IyLehoyo0BjiQAbqWU7Ge1Z/MjQsP8bHw7SJhV2IyRBrUdYQAaSIHdsq36a
mR872J5GOK1KeIxCoUb+Y9Cuv0XeUqHnGZ3+2Nsqo3h1gs0nW7y0qAhhGUyLrUCu
0+QDQFKcZZSz7imXO1aBbNWYwlm3oKHzRQ0ypx5MZnVVpc82x3ZvamUFls5O3zlU
q2QRmoncU6Vu4plisCmD62KtHPUXng6lNm65SoTXIx7jNdruYPFvM82BM7vCIpSS
niaMrl8cD+VdA9McVr9jqdfQhyygTfXucdF4gJ8bSO9vC53/mXIX9c1P1p9RfEK+
72e/6SKsJe5aghnDjyO/tRxzOniwR4gepnvl9TV+E0bLRXBldMVyb1hqkcaSarRv
97cgA0ri9hNb1TSCzWJs3tjcfN0fR+VBDk7xg9tMAzM2z1pIdHXBD3eRVT9hNBLg
I1lAZ3fEmPMprQAYtY7o28zS1iGi42KMrZxYSU7b+NtA6ZkRnHC3iBbNYVGAKjFP
QUJ1CWBRMSwzL5krOHcwSQt5aR4zfhxq0xETRsBNTuu7CFzOSF6smwF3/wgOdf8l
ZZVEG7mB2RgrNjxbKdbg9zIYQ5wbhCwzSX2wB6VqYPGZKn51RGdzdDb79qLUmj/d
XMDJhRfVuFJrlU0ap5RiQeXeJRNPQRzOw2zUom9phlBbs1qT+9hsv6+7UTwg3ZVH
YKgbdIYFlYQZVzLv3D01JWLwbhMwaiaqykphNms6bNStBGoWu5RobAngccvIVHW6
tx0u9LevMYUb3jUFnArZ4Wwmkbswt+nKOLkdIrhtUTYznVzhrag1iZhMm0LrDzyC
0uGJh3c15S/BqAyRlr18EngI5DcmCxArsjgd5pwMIBYhZeE1vhYz3tkZ2J4Tiyc1
CVOC8QPAUjrvmrY3+B4Z7qRsjbJOftcHKuVsAq51jh9hewibdZvD8kQ2Fm1bRdpM
uShxKWi9c43PFA11+LySRNWIOdN6DhuSBddnpT0zpr6m2H3JC4XLaEZe+T0t1YIe
GfzKCF+zaHIp/k5t3LnYsfFNaLazkcNyOXxLAVbbK22C20tRfv8K3OwIdVJeyY/d
mPD2u5eI72np/SGQFkCtP/wdcWoa1AWDfvhIFSrhqPI6idNQHHTbsZc63VRUG9OK
tA4D90q67rpFuz8GOjI+9clOemN6YdlzuFE0KmIxjBsY/kZLiDMRVrePrjMcLvSS
bxfpIs0Qz/gf9RF780CAUaHMYgS0/wLNduHChY77zP6SxTTOMv+cIiQEU7Iq8vYb
5IgezTwA1bJKHLjwiObs7pi0b+EVlt7VsrgFVTEZlZt4qYWejsjrJUWpbA9YP5IC
Hr+z27jy7XuUkQmAY7LjeWgeoE5FeQDx0qJPKgoypAdz56qQGhyPvaGo9bTrhxkt
NZ7Uk1XY30ipKT66NubcO5uhdct5r0c6PfPqAqiYc049WiLgjFES+RjaJZ1bKe5+
YENs6PcByDU9d20J66fEJclkPhHApEAFpAK8yPQHewoJd0A/KVulu+mE0I/JiNKM
SXRO24uVffozWp5FQHm7Tvjn7gX8GI5Q7rMxRB+vTQPxBrTFlUfype69OqftPMQu
GB3UQym5NmCXfYgQ3hJgxSDF3BAlBi9ira7L5/srrpi2TXenQUKsOMrqsLmsPnpF
QyZhFUT2XEv/6aSw4kHvS2wAcSxZcSbqRi5qH+Z0Snl2wepqMpq+01moUv2WGKF3
bw64ogHOg2h6/O3kLIS+reO4lYiq/E4jvDUE20v+tqB+nou7kb2CefJXpKgsY8Jj
OtR7b7OZ18a5M86kRM4uaiEGWEeunQaKGzxsQJe4hQfHkTuGWB4Y2Efi3Vib0YgD
D0Eb/9WpR7ZPWR4p4k7sp9qtgDPO0B0y9xlCKwk0ui2ra/o9lPf5NfHxcilsH2rj
11RaQMXKU0uhaclWQ77zr8WX/Zj+4e0XmW9xRMQKOTG7iRIHF8vsrDSdf96fkqju
UlUU9SrTL4gSEgI2R9mlqRAkIm3MQTfNK1i/fzs7H8y8ou4QBBukV9DCq0/9OSko
hSYwNkC/XqlmtIfVQZFStuWAy2AfSLTI3Sh5He/BQPG/iPOqnpyI5zDgLf9VmR4C
j/4Q3qjC1bVhuuYnw1Q02p7F+9Zv5l8hw5VP63+4qnUkWamnMkaPXjaB6Bsmq45z
/mKKmjWhluPt2IxjEddChya89gc2msOeSzotp/0dN8lew0QPKnHfd0d2NDyOVT1r
wZhii4C//09jisTci+9gEq5o8buryrePf8meAOHE6LrP8ryOOwIGimUiBsmjDXG/
DmqA3YcwGbJO6R1OqTy3Vgk71d+4TIB5aK80Y0RlQ/GQSTVXG01K6E71nSCgC3dO
CwyzbVZhy+0T2gBmSBXZlU2HL/tZflz4fuTKEwzaYw1C55ry9tkhmn9v/motGuXr
W8cGO/p7NPo8jtxAbZ+t4TXZZ62QsuioYV7y7zb7d2eiC+y5rMWQff4uvaKbMhVR
GcAG0g1hnjbroJRSf/m4h6FDhyABIGj1VBqdPEKhl1J1236k8YdWWKTl3KpU7qza
gQJV9nAWzz2Ml/kndaqTeHnk5N2F7O8D6ZK7epqzyc/VsY9pKX1aIOrRdUwEQcP1
mbt9fmYdCukTl/rU+4qRuVuRdel00bkNsenzzIv8FteBUXT5CdtBKnxIpZPyLQfH
+cw5oybPDsYkOl88tMBEmoiNwKIks9IBhLNfgtTJE03t6KXUUEoleXIPtP5BfdwM
ShLBGzqyTXxgviJjpvjwelLS6D5LEhcVcN0qSFzxE+wxkAa1ELQLfDZv0ZRZo9MS
nalUlOZ1vuoAAL8xsLR1nlUyHZxTK2n0x7lYZeDkR/JNvwsMv983k8VduTXvbfWL
8Fm2IuS062MMMAZ9+uHrGVUIoqFegIACFyH/XYF1K6kvEQpdHd4lIDfdxIIOtr65
MfFWf6PFWpnRJSVuj2YnilIZNk3AO4T3he70jxCyDkL9ZlaZtDKm0ES8UZEPDvdF
ZvYGQ17E0vIIPfGc1rSuoF6XsorBPPJUBBwYgMyFIyx8jR6AXCuKqa4+FYFP8j4W
V/3i8lktlP2XSJY+2xYLauIidfKI2PofVDAtF9vrFtWMep+J+y4fjPlbOikdtt8j
tqIpNzLpcFscUP1bj5Wv31UFB3SIw0atZKF7FXC0B8iznjjMOZtdQJ79x9NMAaib
ygHTsTnJjoiAm/3sBhovnypkH8/4sGfYONKJbKw4HXduzCpB4Jh5yyytIHAxcT/l
hvdhL9ZQGVY27UKgw50TVg7GoPkASnqZ7+GFc7YOboWIe8x9GxW0sjvkY2HhIMwn
6fQWWdgXPt3vF7tCqAKIl1L2b2vEaaIi+4ldViGz8qRZhrPSA1ky8+Yk5tD0P3FN
/sg7ExqlHVeHmpmleE4qpHQftDxPKqDJ8hM3kib2seZ1fBroGQ3/fC5NLu39Dnhu
hPsSkQRyJ9TisQaOkERApXT1LgCYQ3xTF/aTSTZbPL4uSW1kMXXcIYhllGdpb5ae
Sy6P/FMYI6Om2D9gP7rB8lHq2rm1xiAKbABA6cqz0tzastmu5Me1S8QfHMH1n+zy
H+4lGDgV+uH/KKcBCtuidJjUNwo8tCE387t9HS/26uPxRrDk8pMzPR5oZlBZtKFJ
dv/pU0y6Zw9h9vMN9EfoEk+mroRnZS2rQrm40b3rc5WKZULLWiuipSpMOtdnsf3F
j2JGQKiOoVIWcggVoDc3fM7JzHco7q7xG9YqK1avX/fhCITwpCsO5lag7ffYlJTD
oNVJJoYdogYwLNwcSXPU75bAgQWKSvYjE1+8+9YOh3zpl6PRC7dfODCe8jjhVcY7
7VAJDYoNoOwLseMF3d6xLNdQXbMt1SJ6EmR4wTLBhxeJmvWc8yA+Ocf8z//BfwkX
2dFyy7VCXWWC+tvALm6QAqXT9De5O8S2VDrC6BJEdQR+cE0ZQ0dcl/sQXWBwUEbr
LhWe3tMdGULEU/6ske9uEAzEx2D8GOqkzV1Y7Dps5uij1jIicM8OANT4oybizGPg
RQR/qta1ibhLEAxth3oHj1zT2W6OK75XzLmWu5OaoFwyJ5ceJ+IG7GErUIyI90TZ
7tuOcMK/fpQjhfQ0DJ1Yi5ateTfoZFyb5s/iKjr5Db5KYunJe5cFp8WlVbZrso8t
iBr0uxisGmtBL1VL12wEdFhRWC+LHLDC9hgBsjS3EgjuWLMvdvePyyJYg8pUTI66
XIaoYrHACyy7fTvKSku1QFdBThj06fvvON4GskKJlqRpJVvBreAtSzLCKrRPpMau
nouMgQxQBLCL43EBdZ1oCARa4jgBA30xHNVkzzojhpb8OwE3R5AjsuKAqtpUQbqh
iaJJRIhfaa61fErKINuWZyMqgiFHknfD7CZk0S1VKJjzW42m0uMTMXuSg2/UfmyM
xJDzpk5Pr5KRL8sknuLcc0Pllz+N2j3ksDL/66QKnBSkf6AB9/6/Wh6A4ma0zyIO
tcCtSSEBGuItBPMCmvJPBnzHNtw56H5Pr7ukbQPuyYBfw+B497p9Ip7OYfni2On/
m3TNG0NCBV6dxb2U5AuLUEgCfBhXsRc5tmuu+Ca5uJu4xFcmNlY3KvlnKEu6x/pU
URaU2fXIm/jP/T72ubVqyW92/dCo6/ZF3Wd3d7D9C7K0FjuA8HR8ihRpQ0Ccj9fg
fp/UpTwFeHp8BCzzp+pv6p/grvO4HZB78zzSAF9zywn2OP5xMzdOTIQhdDFZXiGn
xCRKtUH5dOZSI+besTiV6baqLxgjoJ4n9vCo6QQ3+NVCjJucUqRSPyMsPdyQEtnW
mcb0MfG7wkmj6sOvIlydzPIxPHQpHYel2mOTqdySvi4K9wuEo8iWau60/ab8dFsv
DgNH5HRP1xodn4i8I+tRWFSJdeE/gaOCSMsOysefeS8gELXMnkObpWX3dVJWf95z
dzCesHlpApYrbbq8ZfLsM7JAJqYMM9BrvLjdNtddT1nlmynOYABPLj40PyOXifIF
9u2Pal/V21aFlxRty6g4Fr5M0EZ96Y4Z31/TZPXdY1giPhWk6FgRm09m7qJz7mlP
xZyvASBEczo4gphQCG/UhEdrYsA/7nfH3NZqrWhCcEOd34tRF20vTmS6IL87i/05
jwX0qpf9+ewOwwlUQFc4uvvmqf4h5ZWUK+ebu9KSD2cIYmlbMPsMrY0hk4gdrD9s
uQqOgx8FL/uqmLpQgVFXdVx5SD7UaQJ5J8Xw3xKTKTc4vmfUhq4QPC/rLX7kAYxh
2xxTZ7Bco2X+ogkoMSdREy4Y7rZ+MdgpelGn2ek1A3NBSKpafApBcUvUi5eXmDgx
me5yzBNN6YTCmRswqhds8z7BRVbpNConXCcE2Q36v2AR8/tvzGHfv4afPC2KrjCK
2hdadF4aSS62UFw1x+iUNcUOD0nvNzStZJJX1w5mMxGZmSUDBPA7VZtiSmyAVB63
geTf5+ORO7F6Si880FLGCfWUo7GmagePnwRo9GXEfVn8pB3ssQdObs1+oyONYbMY
now7eIj/5i641LuqbP+YpFYzFfU/XLpKWUFgdtVSXRszjgspKUSQ9qGHeHUxARC+
RZreGrtZntdtuoMiornR99DGAaRG/TZiWNfFk9Up+zAeMpfA3jUqgIYE1HRErWRe
tg0sWZY1QurVf3fRxZFWHvr2HjiNNhKeIragl8ruGWfR5SJ2inA1lkrNLLFqHUmC
YdEcklRJnzg0XVweAZCapRhpkWmrAkbaFa3Y3jplW4gpUngqRQsqe0tXrnmnMgnU
y9qZD/pISUTmadFpNCewa6eFX3IksvqZYam4cb1HaWyTkMW0FkGD4ool56oRZrPt
EH21mveph/flnrMr/S0DU98JfDh7VeIqVp6SCSuCT0U8Dk7csl0fwoxdrZe2ksPp
DyQZjSFauTDMuIn1AKnk+FYQidy9a6uqABNLVXaZZTvT7PQWaedXrJPSvWjMfs22
gDExBBpA43WIMH0yQF4WhlKhASTPj7SkeQIkZeHDI89lNKRjj6r0kvcekZefd6m/
TtPM6tfbhoZtsyt1Ex+GWjONd0mmVMLxv9jH10JLRidTBDwLhMB8PBS7zVSTpaIr
UbnJ8gvMmB5X+LipsZEGl/Tr8wem12LBeQeXtVRfhDIrUq96a9JEwMaXRXP/Tr7b
OiN/wt+vInifCiiJd7sqSn9Yt03x8cPCTnwRydk+8RaFRscRBS4jC9IBts+BLFcl
rXPEdfFYMgm6ggIASE5+BUyavXbBm4f5SCJ+JKXyV1fdyQHMmDS+Zy0MnSkrkSNC
RwgruVJf9uYSzJRFXO+rishRIySVpexjr3Ofo3WRqju4fdQocWlV380XM5eYwS9W
4ePQkRvLCeAXk4Thc9A1iA7RsrSAMWZ25MPYhQ+zCtU1un55Gd0A4HZx494febhG
iaNugD4P9r8WvsaTEVQreuNiWe8SVJj/1xGKODE13kmu6zRNftielD7dzyS7tqeY
Fv58pjinOrzVfJCvmr4F03TWrSiedxJmLnKnB8EPrseIkKaMBrbr42FpK90a6auN
1+ad7x7mEhIOtYfE+iapV7SqtsxSjUyuLmmvci0rpN6ZMrU/gJ1BRsdc0bCuaGcK
Vbe2otK25KX9upuSXQp03n6QNmHqiZejIfw3ygT2ACcCutPyZpDsRCrrotFqHhzG
DB6FffV2gXFJl/vNmy56rMhuLMSNR5J/+uXtWk5aZ/2nFALQXck20PqRry9XhQ5K
8KycULZynuHsQUkDiGTeSn41ywWq39/twGvMU5sHjnCneB9Mjr067k/htifexQ2U
H385X0BXIOTCDVYq5JhXJxb5Of+muFPA5o+oDy+kY5iXUyCrGzaaxZbvlxvnLD/b
DIxgXY8p+aDVtkEPHmZRnSy7XNosJ34LW/BncTZ3C04siUQLIT6HfuD+/E/TacS5
jfxMyNxM39x0vVPPoglEYmDCpWcb1Set4rzDAjwhkDNb6Nuna3vQKi+d8x5oFhP0
+rcRdZe0wtkfBSfKxV+VPO2tyqdrkDfmmxlnCyh/RjVncDfOenNRZ9YIinVsEA/k
kFoRsKQYb4JAsHrSZgXoIYdQaQZGU9tBaxmBI5IicSDX/0Q7VqbWOgkmMdKmYdQB
ijNu445ovcjqbMm1Z9uFIeuVhLVqdWC+OjcnfvJ8xcHfWiuIzJuAtC4RekJn5fEd
UpdNli70OtlJa1MYVpdDNBR99jebmdLvArNKaiqGi6xpnmiEfFbDOSDXY+YKLMDm
rYHSy993jKTS0jzsFR6m8Dtp47tkIWHp55V2khCLHTMdzLiLzDXFK7M0dhsH3BWI
t5dvLHPciJ415zSUuohWr8l059/jbyu1bX6l2DguN9HNNZaJVEvnoIKzUxEm8gFH
dv0/DItYCzCtnkvR/Pdyc2OEjM5C9Gm5A1Y6aLOEXIMXFcbsaofQgAv2bGLoyFS0
YUXc3COKjLQ98clqwSC1x1TLuchgcWHen9xO3/sndSLrcsJSqOPyYVPIk5s+EZqm
f/YgceVNR0DFFIAVDv8zBJsF26zAgTDPQURaX5vWz+n3wHxPNlcwqB+0SfKJCpdK
c65ALGglJ9vx/iEcvoIIBAgbofVw9dmUKs8wYVT3m+uzM+9irUUKAgLrJcSD2ASV
kAnfE9vIKLBAmlLGQhPjK0GNig1psddXaIHM9Tc0ATD1eIWHmbheMG1WQ+OEHN1A
XAfTMNEfblmDK0e56qaRV0bKRMy4HhUk8oUCXMJbQD6DBzDznYl3mF1Kw6Arn/RJ
yzkOD8OAW/byWzHNsICGaLKBurdm/QgegF2EQMVcI0nHxoKT9A8cqzS0oWzisC9B
uFvGjGOv9/AdkZpBMggkqLUZ3mXo6pkatCcdAtxym0H870gOVnXUgehFAwlgig4b
A4WFVxpySr3XAN9jNWzY7u/dxdMn5GdPNOtMuDFECv81LysvxX1XU+Mi0dgvDc3x
J9c5rh7XhAG3HSuea9xXX0ewAP4mfHQZARN6YwbxfI1mouIHjFLkHFqy1BTsDe3L
PwvWUHK1Kig1KghqA8oXYYQV1aJLAuLNJCH6saDf4cXVk8mAZgskwIsGnQLdfAIA
nyudW0TuiJGu3muWASx1CCGoavFo9YuMc+gakRXPJKzcKLtskGJFE9X2psU4qYpu
wCdROmrUrM35xwHSSRcqqFd7LGOJHe56FKq6Q9WCANr11zQfLoq/01714ZOuhW5I
cDsfUBDDqECmvdKI9+2TqoAt/fdDSVFsgGdI9mT8LQqF0TvKlFFOkjGVJEkH1m5m
Xp/csBKeED+fpENlgqFDOl8+OMKB/4+JFUyYZvmadKCnYIdm9E3qBSuTop440xcx
b7bXKoJAxGB/SHA4HmZ2SG0Zt1LUIASSR4M2XIaFRM9DR2WlVzA0Shf8HSwTFLtq
O8E3Vo1l1qYCHLriuRHVJHZ7WsCK6avKRrEmbJvkwHXtLErrRnSpt5AO3q01C9RL
NFjtj96psVdQttp3YQG17B7fsNyuQFIVY37gFcqgnATojgbjmQt2Q1WKobffo4lL
J9+JKVxQYQITA83UTUh889aSIZVmBKfpjc76FrogGFDfvgHKehi4xCD2k0sQhh3O
Kz9s1rpUv6LXEE56vCA0L5++MDokGnbhVfjQxW3dpcU4h175iSXwnH+1R+Eb9p+u
JhV4b/R+tj9lHltvhNuprM5jEkKFvFwpra8argBBsqqqYsOPGyGR3+iUtTx7H0uz
ootDNAuacNMNfScgYCDpgxl2m//KHR5urrHBnkWSohWvh1QCwNJ6LAzSW1KerPDv
ygd7F9/gqbNlXM909QWvsnvXvMmRcJRVuSSUveTXsWe07WCtGVGGIYud0ggq4n80
U+5yytQkzBWDMQKcs2xpI3hQ97i9IYxPXGgl8Do6vDasVl2e8zu44U0f8mq23URi
d8OLJYy7yN0Q+dt7vrO/dkyNqe7Q2DDzfl+HNIcAIfmn3vj8FzrjrW+yM882Z+lh
BBrN6y3e5LMDTAw7bDel56k+yGykYGdWC2/+hG2iw6l/c9sfUlcRF3eVLdsRN1gf
fXbke6DVa7NFI3sCCKNsx2nosmdG9aLBOccmLsGZETOWpeSoNwSp4T8g848U8x/y
g3b8R0V08lvI0rB8cMle3lRr0SYf6Yblisr7SdQUhpfyreAIGLUlouA4Cty0TBRU
yBS/FLVUn9ObL2NKlAh+JVXyZi6v2a05dYGB60HPr+1LIhfAu+K1JIXSuFw2ZzZA
1pqBh+LMBrFhPqGgquwFQaXn0V0hPRtG/bHMfcJ0CiYuPDujUntOKd8mOt5kLXuv
e/9AZLP/CgarVl7VzFK5nqg02OSwK63/RTKYnp1OsFyAdlKJTnlZnxPQydJlWmPJ
+hKtH8Yt7Cdyp75GomCCMKlhr74B+m/b2hdvJ5pf4+xWtusCS+ovQH5S620ZHSJu
uiFftXMFrWoI2UrUqQ0D5cpAqU92EVlq+Ae9PnRJ5gGj4wWMGEs8XVWP0iuUL1UF
dNJcFBKf/bhbUfoqLjJh8YOU2rpL0ndbSupuIRJif6orJbaTRNEW93nB+IiruaJM
8WP5ELvc2VKlrSVSHvjYmM/mQx46k8qodfeCOteY8ca1MmI218LePtS7PSQCavye
h/qBFBHNrS9Hfg1mgGRpOSXHXhEdtRUpW1dG8Td2S5jxU3snIONUuFmiKK0bvpOf
zVoS52WKdi18zcPB7JGnh+PZ59kFMylaV39NZLSaTWaQaCUzv9+gWZd0DUkicQgk
DfMr0Blfww2+8OUvrBqW7mRksIwbd/RizERjSn/8pdW3qZBEZOHdcbWlI9Be/O9Y
IPg3Augspu9yUoNlFgaznGOJNX1E4aW5ji8mJHbsub8V3Ndx4inG4kHqYiAdTjid
qnpd8h9Gsp6jlOlDDYOY6VfWN7u46vgbgvXLmUcNh7Mh8HTYkQ2BCX6CZ2TyFKCK
iBaUy+GqB3UKW6COsN0mhXzvF0SuiSoEJuJThI9yzqePXIUoa+X0GUofMNf22Qdv
4gImBe4bqWSHJ2iXZQxyr/HFgnIj0XeJD5HYJ3iydmAbU4Rhp2NoWrcGoHfE6GEE
OwLQNfdUni8FUXwnEKAukikPtWFB/Q3yyAuBAGVa3Z3JNf5C0pWSzCfHSpqimgoR
j6iNHt6YIzySst+qzPkcyujELLmSRzSFAScn+bgg4l3s1NutYky+8TA48DpjSISA
2oSL+oh+z6F60POz6dixhLHYrj7tMI/dsvN7tXRPVbft0fiGjfyobFR8OxOIBNsR
YdsC2whwh+J/tmEV/czR81oaBVhP9ohf5OwTjatmwMFqfPOvMZK2F9pni+h2REmH
PhaSxnBcMEUvo6IBAg1NRQzi6QZj1cxuxO+KhWwvdyKiWO+q9+D3Pnw28EdAbPBX
KRiztrMntxQNcEK9c8UDE+8YtMTdpcPKfok6EhQPCjnQoOO9/UqrgLLeibuV5bi2
dmPmOBJmZbYJdBmuC6lJfb3YSDe7OSogtyAgRXcFk7n1W1ntvPRFn8Bc/XQEurqE
cHV3kBhQkMY6wLFAGM6jRfDb/d444hYNsNlekydrj290/huW10E5iR8TsIdKmiRq
lcIZ+2pla649oioKMJBcXIltnRZhKhArapKPhPkYZYG/SdrsH5svXuP9RYFSNIFo
b4gytF8DrJypLCvPcMI1uT1PEbgtLglFwNW/U5LL9h/CoaWsvoctF2v/kOo0zFKp
mJeuFOpGTy9TMZx59hjKLoH5kjQpughLeWvrc5lvw1I0d0RWi1kxHa8O6i6YiPo/
NbQowuBJK0kqHCCvjOA0Pn/DpXNKUWgSwcLyP58LGI1ilDyPYaEZZtS1MOxFyOxr
x9Zm5xDoSvpf0m+Ik0RuSQ0wfiyxgrABLG0BiuHEKjk6NyB7aOQ/P68uO17+imbI
ikzBtTj8X687veykofCKEKDa9/zdsyWN+dNls8RSb6aFJns/ABUfxlocGlZLbxjk
I2m/0mMe0Ceda4yWoCSHH4b9zqNImjiCLRxwb1BT+ytoPQ1jp6vCMM0hoAc6nMnj
kmNKyJW0Mrd/5/t4P3Q9sv4K+lsA+TxukvEZbwgzq6qwc2xIkC5IXrQ4kxR0LeWi
481EeBQP3mZthvKbyIX10OUqKCVlTJaaeA9eKwB71gtYtvoQTHo6hUrkLDV8HpD3
vbAxIKyuoLPESRQsUcyafNIjeu91oLOFl3mwtD4D8ZqRMcEoaNeY43z7/phzyTIM
049FwCPFq7iiUS9UwhpaZQBegPgjlzuCzVc1nn7/NHOiuKfOxJygcnBZ0WZ6BsNK
Tk22c8+NxM07uHtho/wnii/4mI+Df9rPadpC72MuCY65j4JG4+wLdYUdRnR27yjS
DWYEmFSz8QWbJuaMWmPIQ/rtlGWMQ5Up9OWTC6VukH4tDFl/1AlIaCr54dgVjeco
8mQMTeffdXFJWqwN3H+K2wPPTo5M3vlBp5zI7TJLve//5gLLvvSaCpN2b6vGsf0e
lZ+NrJwYXD1UgDcTGaZtxNdJUU0dtnyDdKLRgNSdqUJE4WJFha/jSmggEsIbcY38
fCC+4tw2RuvAxhYa+LuCOeOyU+Gmzh1U0c99aqYWSy+HltP159m1tdU6yITpqekb
OWV2kQXUDQnF8nnuHid96RVSQmzMxP5ighMB6H1iSIcYDBPMhLu2wzZPD8FEMBXH
Gaa4/I/w8iPtXMmNM70Y33Mb4zPAhZ3gBnVDKd+DF1N60HWZozxGqQDJllYjJ3u9
m7jIGhdslu20edwHN/XKkV/f9ySoXW8bCPL9CYZUWSxoT5VsMWLuI2eRYbiQTB6f
YSE/WQNod/CBO6mu+TMlbmdKHExkhCcHlUjfomxpB4SdrnQ00zRUXFN6Jw/CmxxB
bwEqGal/46GObRkPz1M7Gx4TuYFQ3smLx+ra8hwPd5fMgKAiDS82JPY6huLRsqz2
CyLzJE2uT8qj9fpYko+QBZgTJqkclmfF1v2D9D5V8GraTHecBy10euiq6sBerd9u
9K/QcQO4gH5YKoAAIAQvHHoXbdHmRe3qMnKDKahI0/zJV31s5HDCJuqUu4uENfxv
xm+4IljmVqkLWZ4T0rauNWdW/86Amh9+oz6TW8lK6R4Y/LloP9+6R5nZjn39GuYB
2J9VAzM30r9QgN3F0dt/B5ErHMoZsohi99xgavSE+ne1um0T296w6F8yBv+1xkHG
z8H7IduGMPjhkfKYqqyKo2j3FvCVuost4cf8spa2Wbq/WylbYfLCzejMdyYBeJ2I
VYwwq2UQGwco4xfVgNgVVcIDSXQzUpGBJM9YUqAToaSnbySyBPZwwf392Kvs5W4J
POkJQLNUyh/4/DD0EWlnm17nE2P8A2PqL56r1JqwRxAGm7uAe6HwzeYVGZ+xSGBx
2lJAwMMvPUZUfCUKrzMHH0qeNCX4zhvfxQBkbSCEYwwJXGwHBXRkWsC4cJ4QwalQ
ebtErVLv9/U5Okg9Qo47Lds8B4oEcCz5VOYxcXoFanBIgLqCmUAq9J1qG3zMx+Vv
r09Sp2yvEoqYOCwg+MxHM+u7fZn6BUHiVDBMV+unqapoeum3Pf0svlCHKUIRB1gA
sQB0HTYw/oWHelcvst1T+CpuRPEacG1SVyiyqRnIwv8BOlsacRd1jVBYPsjP8rVu
Ks/hdiocpGovrHQLA1GgnOSdOZh8CW+86RstFZqk7j1lt91mPBQ6cVk0//aU6zsm
OhZ6FXS1hCSVyBMhmmOIQTyuN7apAUtggSVOVX68jKXSXt1BdFf32hR9Pr5Yr60M
G9HDggfh2Rg4GA78H9B1eh63q71mO/51rQlPW+uFP1Kn2UqGLpE91sNAa2RpyJuF
myXDvwVYms47fLpjMhQVr1K8/rf3wJhskPovaPpsX8v9LZyFNAqw4xWn1TFhykwG
u4rz/60S1B9tbsW9k8ZUpRCramKn7Ux9EALzfxVqvUVJ6MAmV+00QLIfmF+vCoj5
Al9Bth+r/B8nzZzOibfoBX8oKS+elI8k5xHaEHsaMJX0EwkrINbNYZJsulLMc4m/
Q5kEljgUUjWrEN75E2LOMhWNYXlofhT2xySkleETFdnZ3T5et7PJxoNpT6A8cGXA
bq9b5EwcWMaIDRClcxLAtWiFnnJlEjGmTaLf8skqgzhQi/XjIUC/bmYpHPFzdXfp
mKPPrZ/tcsEItBsTg/uJhcu39p4vG/mRdtOO/e/E8L4QonAPw707Oe19iNuKJuID
B8vDJq+YmFL8Pfwqde1Its3i6T880pHGizCrusl+6sV43zN+DNaRo4YMEm2lsKOb
7/TC8faUvt2Z1eaHrA6AFqzgJjPs27E2YBJ7nwef7jTING4L5ns8yIdO27xpmBpL
OvG2pL5M4DuU2Pv1FYwlzHKKLM3NcxrYkUJi7do/NMoqSEXORVoLB8QRE3iZJlaO
U/FEJnPX1ecAHutkuubmSs0mBirJCTSL8UKD42p1HfVQyzgYroCAatY1KakIlmvR
0KqdgiNxlmjgm65hgDl/bA5ZYvMAwsst6Frtj8QpXPEQtNItShmZpE/kOXEYNhwo
FhquahqKeOrY9dCtT8hXIyiVXFeEwTkR7+FrENvrywVGmRwd4N24QUp9BfN/c/oU
PTfHfC7h5FpFIV3vuFrr8kPj0M+ppiPqgE7yIowEopYzw7HGCevt1LDjfT65in2G
19BYmCoFIe+YpR7reZfZ3dASQjelwlC367o/za5k9SN5iZpcPZe/vOOrPITCGioI
rVMMZFfnkgWBbTM6rj1BirrhZod4V4fTGwHOrgf/5/nldVVMCsnHkf9CCQwZKEyH
A/qXj7b/AHz70NcU5qyUOCHQ6G8M1OdUs/oOc9kS4BgQmfD4/KwciDxgbUa6cycv
GZXIZQZ+qlUEN0dS6g3T3nDjWEheCXUZWE6Sk8ZORFdUalOVG9czBb5rkUi3jKcP
IF7psk0uK29k5L9onYiWVGYzoiRRJjAp3Ph1LqF5XUF8BtsI9oTPGp2wyLPQ5UhI
gPlSm0wj80CbakZMGF0dPoDrjawRpUNxfTAQ4h4BNwfXuqeA7zzF4fC6r+xYyL+J
iI8pw5PFnSZtM/XVZkCRRV3A7aOqGO8KohnO7Wi6O1uKwSpfhcyu8yGRQ+W+NpSs
flCoCKOGYUJtac4SDMADd/sdhjnjit74w1I+BT8k3yXHijsZj5Cz1V26SlpovCEg
RfXI+kWMIDLocRIE14xLEk+598da4Ih5LXtlvZZIbmikTKDhNqEBLaT0Hv8RnllE
pgxL5X9uYxDewOYZh+0kKqoC/EqqBgVriYsmtMgNNjNdWWi+zZFrW6mGhy3pqU1r
ZU0sIm9Onuef15ljXLrCCb24mIspOQPq3AD+/6xm5xl12PEs3kcucr/wnPjcL1kg
0p7V4w8tKXOTjxF7Jz6INY4N8oBi/fF7uSn5G9THRUQIleF12PPGFP/UwhntB46U
pJKDl6oRolNKxWnjYY9ZFjx/XA6eRA5fN/sQtFOUPwiwrI8UZ1KoxyP36Cb1bL2S
5v+3aV5u2lqIiI56PuEYTRn1agZLvVeqqZ+/ldl0ZqZGWUm1HGsIlIsPCVZRZ63o
kVi1CaBqHJPaAytVL3udl5u3ZL57tD7F3NNWyfezYiDEzJ2x6OFExYcDsTTKpPor
UySuzvIAHn/iDdF9+lI/C/0WdlzCHeM86r66yUDYMjcS7/ZMm3EBod9UU6QBv/iw
59EP4BqAvGlluhHVifOV1uqaMC3naig+XWh/Vl+b1WbP+SjSuL9JNN3S6mJLSygH
1A9NRLxVsem1Yy64928YkQwu7RmkEWx+naHWWnpWEkiihY2Nz+fEElxM15toIskT
erLXT5+uElEyjPqWzdbFcir7SHyxgFSlBezrkCbjyJqND/r9HWggBqDMAsFKx+ZW
QKx4g4RYijjfgsMsOAnaXKeksmEnH3isQrwiCjsK7NCv+TSrB5SGrqBhwC7Eqx5l
K1TAM7a/spBPNYGIuZLXfjP0RgJMrG66gBv0kcXBWB0t0/MfMT+1sCFF9KWIfhGM
INjA+neZm1QzkYsAx/0RNv4wz6yljkfVkvAZf/TQvkEp0F4HQPqN7oF3DQTEG8rS
ljYVjkOUH1cazxGHcITm4wL41I1YhmIFvxtz/7cs7wAdGwpQH3lEVj/+zJGcpkla
wGCC+4FogzrZ2VCZDgctYzuy+B6yhc8XcwJXOMF+O1gdh5XFN9QkCTe/r0CYBqkG
JC7yz/PJagr8m/9vBvyJGmC9ox+7RGauMA3mPUJGkHJ+5Y7kw4OR5EdFTYn6d/nC
asGClmLgOKPd3dre9x+wcmkV2b2wMiw2eq7blSpCmEKUHboL4JMJ5keD1PfYv/mC
tSKSjLW/+94DENQfduXynf+IKAnK7/h++fvsX9hg7QiIEd9zbPy2hwrzbbUZN9bm
3iVmqhE2HY7ey3kxLFBaEccSrMXxSDbypE4kgW40sdMa+YIR7sMgsWjoz22Oi09j
HpUnBNs6JeLKhEBQeEcJ+NLZTP4utFoab8KSnxtIKvygfSuAWW0cCbmKDJ5Hy2PY
+0DDCsE4gM1fcQ5fYU3atobYjEOV48AzJ5vWkrhRRVa4Oi3uruaDA9KEZFJfJ0DM
wLZBRXOa4XsvJrrLVR1qBJ4aHiemZbiF57f0f+12V93CaCXsEL5qwWNxoekjqWn7
ratjM+gUEnSHcEXoouGiVGPYEqyEZXGg8e4rCvCj1MuC7IRkdhy6JxEfalnzrU1U
g7928Hsorq08p+LBe42nmVoUkADAbtqvZnAG9H3mMqrgp3a4ZXmztCyQjr5pm3V0
b4Hhao0IxRnFMXE0jh7CcBiP60VYix4dgQ7GTchuPIGePGMxxJoAY3GELCRhtQJS
xUxZgdHBKXRJ2hTjtykamDLEaivBxCHyr/3Zx9n7PwMlGA6QjXER7WwJ1kkHEsHU
yHPpINcIzqfcuxokSzHJgx5eZPiFZBRGCKuUniDAZwXdwjTSwJuaB+/g6pJKHuof
VtvNv0SFIWlqaLSTxjBmEOVEKSODlroy+vjsbF8iLEsunBlia0VQiquUnCq9XY2V
x+m2KvzuV21X53eODD3kB+EUXIVhUtTDsjwOKIQi9CECaWNqa9+ZOxHrIz49DplG
hZ2SaETH7PPiJ12HjNseztjnwPa4jaNKSHoKtoLXvSMfTzQhok1BEA/qOkFYtO/U
7xC8U3m1d5xBR+VUULSndfm/Vk/vH/+ZlSpHemCKFJ88KDlFM5xEBUm0s9mWNh8/
yDWD0xuKK0h9lfGStj74Q6K3hIg3Ogs5SS6X+BlXygBaVC/lOKKKOBANDNhUEm4L
o/JrSKBydXrotxLPQHNoGZjqAMfjwxmhGuDfRG9NzYapgiGxLfFMqEQn2nDufNr3
Ltco9s3tHv0SrnLSlRATYsZ6FRw5XXNZcypoeTf5mt6X9DxaeZ7KiPzKf1JXnRhH
oALuJgdjD5kUH2C+k3pSrYiL7HKeqVgOpU7xcH9cn8SlCQkipNusiA+heAKGrCZz
H8cgOJvoD8yT65lKB5jfiukrv202hIIVVd5eVSxWGEAAsBA6k9PXCH4U8CQWOTIV
W1mRxVgHCucmT0JyhaAzbks7ER/rd/92n/+pDD8Ps0zzWIooNYdWKEJ32JG6LDih
4fDP/73oUGpREcRn1vyya4HU6qAs5IL8xXrJdOQ/YfUDmZOB/EEEjkwbeDGSuu0w
UFZG2n2DzrS6yWceV5ABh6LGQyaPYCbDwo8jXBYwvT+tX1F/GhYZpP+9K4A1nQdX
eEcdpw6j2m5Zj/c9V6U5VTj55Nlij73fHZyiczoCLfFlZJOOM3RtplK+aADueBkZ
AYCTIp4agC7dy7IX0CoCIlFnaat38gjShNh3FXS7iikTVOTDGN3sh0z6krswV1wp
ncntrVVpFcyOq0vdGEX0BpMj6GTitRkjxtzh8b7Wy03Kuyylx1S5zTYpG53FusW6
uh68ofJlfaOffqy5Fed9xC8CgeZA5lCG0xUOx3hccL7lo6Tn5RGV55Np83S+4qoX
Ftp6YFXu/gH/A7wTJVnE8aYReYlc61fdbujs0rJFdwm6TF4npEW9CrY9SpOIn6zx
bTVX6RVCLb3pIAAg7SzVF77Rtxj2aYXCMb2XR5dO2p1bdr/fyQB5roG4Wa/C24O/
tRNCsJjWEtXQVmi+tc10Nj/hL8hzG/B45jkSc5gJRSA8kG3Omg3TzzthQ11eHMMF
kYDre9dGUW96wwj9s6mU56Yftfaqu3JIitF/sWW045MG44FRa4sPKmBGpCiK62CT
RBsheglRTojWF+UM5qgzwFOp48B3AxF+MXtihCA6oAlz5whSs4DD6G0A/tJuAYVp
u44lbDsbfwF5htdAl7XZS9WcAybyVj0shipljMqpVhk5BSIcAG7OG56yA9g3wbu/
DQmtND82J8Cuv9dMzuKLNCVwkqElBBsrTAUYib/XdtRrTBJLp9EwOP0FvF13Yt7R
/Nh/JQZrnHgAI5ciUwfEcQnLUddtAoIeV+qta9MjQmo7FIZp3JvyOCAciFNVrv5M
mazC9wDX6rbHgVGrt2tlge140owvZRokT3Es8zRd/hVqJ6NPTu0PuZWJigtjdnGI
MYDI/SpzXbjqGvghRFWpu26wbpTBaSIA/d9FMZd5SpwP3HLk637c5V04EV/oeyMK
v3Wy6ynuV3gYAJ4lBPcK2svc+1TwZlBoLS5Y/Hpjg7IXLeVdOwilcPUnue7oR1NV
OJPSAuwzMiDBq736UP80Nb6L37HgLwEi843BukKhz/LUjlWwgjES/m/Yh6SCw7Ej
Bn2eG/fgvOKlKQTmEVYSFZR2my3baU3Ghn29MJyTXiKcktm0K5B2nWvbE63IGc4+
c3Jy+fa2vF8LFrV3RsrqhXxnHzrAfdELhMuAfAZsH9SSZzM8XyXpwH4K/jrVF5A9
R/vWs5tEwB6clUQMO1jk0/dKRZzpfYKPuvOFWFVaFR3igukomaaSM+fzbUp8c1HN
W3wad7DE3oP4hhnB8zKl42umLLci7E7gEEKTe45/MAF4Cx+Q1bUoEC0+93b6oBp+
mA0dQF6SJ+GglDezqw62U7RyisWWRIhGlYA0jnO5HJpAsjPR73WIZWUhPUBRqOSO
olXDwr74msFdbF3P+2BjMnreah/Fuf4wxjFs16ZvpWrzb5EjXzur1Q0wK6ctPtcN
rZIPq5AsOT5IXftUqNRjYSdaJgBeG2R3iy6jZFXn4JQaMyQswQPKz0yztB920bng
4/NXnw2Fmu1MyJaMvUHxl8IgPuHacVzgEASgOlGs2A0U1BCO9bEYQXF/1lPPE6tz
r3L7+TsbMamFCyTJSiosWLW6T0LNsUDju0WjMCfxd5YEfNe2alI2wUCOR5/VyvoW
w3GrTCbJoafFXoroSyQmQklJT5jWcklcTeUs0N2uzCuXPdcC+BsuJtN/9Nklp09W
f3SV6uHSw7WpB2+CHk98f7radm0XjUTYuEPAGnb7MmBmkBgY1Udn8Ssv99dkE+L0
gGhRXZxSkBCxGlVn1Hfuy+AxnH+ZtuWtj8L1seRQA0e92V1RtUQEhixM5Jn8i6Je
vk1RZDk0BUswRpRVmuYVUhhAtZR4vSW3c/PADnyIUpn4wDfa6G+om0DhZDnyIJrk
ndg5CCizyDLRhSrwX3SIJ7JJDRCKiNEeB3F9fNvi6r1r/abnYPP/soygp1UZOWJ9
kGDX/EhGomrdkB4IpBoLu5bRHdlvxQUNTHmSeKF7zb9ThBJL99ZW8C89Pz9KR/b6
NUt8LP0kofeYy18n31PzJutndPzqZf4nvVDRyBgESUBL4QLk/IG/SAXJfC9tZrVW
iGQ/GZC8vHjH+hT/6B3bRJnH6XV/2+AJpjgNZybaYEAjhNkLOGm26X5+7N6k21/m
bdbhC+qtpI/lhIVgli2yN3HkEw9QUAJILKe0y7/yDTbCoICZdA8STB0pWAex0Gh2
qPGfX3JTCGmr8pjHVrKi/fBLha54vs2srDk3eeaZzK7KqvrfwtHRexPZ7uhLSr9D
c2DjDWvdOROmzIhPK2fO3bjJYBVS7GWOtGwayIxlqbgQXOUlsm99ifGVO9rKhQeg
2FPCUTTqfO68698is3y4vyfc5OrbxEo4ocFuX8oCD2cWPdvAhHAycZ7Dz5DuxUGa
YdhdscUYKVpecrs/A7uhQ8jdVMUiE4QrT0IdENbftM3eHQFKciVUGjPsaLl+V9Au
RgAFm+T1PynEIY+n4e7jlT9IzqGZP/OJLDRuI0qf/o1SimPhr2R6t366VV7ey6pB
pkPFOeKdXzZc2ORoKNAdgMuYTJFWPfkYK/ysPlff5a+6Km37yxrpOwhxZ7OzFQRK
dXHktuf+yY4QX29QGVP0Da6X1H4/TN7EHDSyUb3ZexxA2LOrNgCugfC6u7D2wYM2
UI9Rsd8ZGauvLlw2x31vSdSLSUVWp/d/n3sYV7+ssLMRh2rJf/JKO178Tgdfii6Q
UuY2hJSCWvqmOGigdCZfzDSSRCW1h9k2k6Vn6IR8vpMT/sBW6UwtKM9bGA4gv2ay
hAiBbXaPPjmClFb6SvcD/QTQkaGqame5CIRmCXQy1tXFplGGQmKAhdnyS4xveR3Z
VjKcWtprpT1YXahEW+u5VwHToAr9uf0NP54Ju9xHRmT5BWYGNmhYCfCMeEJcVi+C
T8olddK6unOTEwwaDI8kFX5aaLdRW68iRWz4fR2BSI0118QjgG+9gBAuQ9hxZM/D
S0yxeTRl2jeyy7DejUeSBJXa63qZnH2xcyLoruK6j3K5uVJMPBHrVRR1QFPr+5ow
dG5dbxpjo+oXzi6BnUZrHltxKtioF1fNN9r00nfkIbt1SexNT7iYmOyV+F0L6Q4L
0yhzrqxy5cJ+Vi9Eyxtm9BQlV3d+irUDtHcDqcpLm7DQY5iiUvc4zSIvJlILxKiV
tRKCNHeFLfgWsLNcGPMMfQRP9r0WfyVN6IVSIpF4qvehKlv/NvkqqTbgcihi2MYi
DR9XucTnkdliEUbEr2tmw2uA8yrwRAciKifb/XOmy+RrWUemk1mHvBlynFeWDuoq
TnWpoqGmLi+/mmv+UrE7MFGVWEgFihRynCXN4wl/BofCKpRq3C6xf8LAbBdBOFR2
eYzaMOobM8AD1WUO+2r+EgtRtABtXhXBCQr6RHkvX3B2l713zjRcp/XvcwwCE3Jg
m9xeFYjHkxOtmLezl0jl3M5ybCF+E4vWeBmbg4h1MGgksPdMyFx3utUnc7DtrPsN
dv3uxR02PJT5JSTDqocyODtWRYzLFeFPdh7+S/D/AWE74KFbF0kmlJdkFH2R5JJs
eDPhJS4gfj62v7taesPdqWmmVMTJLdR+VnLGa6tPHPZdJTjZE64H7dIX0w5WgRxx
VV1yruVh1TfZiN5KAyW0xflnj3Pg1KGrgrg6KEgpkTZUHBtO5wUGFXc/GBJg5LEe
36Z3LGA2oLZnv58t9ZQvgfOxg9wIRG1APLlVisn+9MqfPCF8czNVevaWAe76/DxG
2wr+iRKexqBRbLXkdaYz6q2zXFmmbGU5G2Hcdbzw10FoRGm7E//+CFCP1SOZF3aq
n8jT8RGbG2P0KIlSvH+n3TG6aKJfZ7Yt+3/DDlAgDWa9Hp9Qk0hW6PIt1btDbD4K
bX/Hm8j4dU38glxVBHk4kKsivY1M5IwH2ICQVIViH/qsUJ8qjZp17Iv+qOsj9OhA
Q5YYVVDKsm8SAvrV+sipjt4/AzlEJerqnD2HAyzmuTbnT6kiIqxwTj7Ps8pjBfAh
ZhOY1rX+XcerAg+MC5P3xCnTqSahwTwFDcOEWAhwSvsvigWPolisK1adgpvgtNdd
0LLiBz370BhQAVuDyglOG0KZGrRdzrP6oef6OWZKlXzELNxPZHR5Vzmbq0NFroU5
iiU3Zm0f4KaZqmsFRcDgqD2/UTEuLbJXEHs+gzBZKE1O/KjYjMsYE+pGjSYMvlz6
maY/39jaB98JqAZS6EnEX/VSeVB8SCslf9vuQsjXSr7Bk3ieyHi/aGpHUfJQVR11
TSu35h/KLoDypyLOtfQvWsSbeoud4hIrPDDl2CO+dcpgeZfzprmh0PqS8vB/kaZ3
L0NK+lxPynDdOCGMoe0DD4wu35POWFqH0yD6m0iRG97o1iigkjghcw/DfkDWMJWh
Ok+JnRYHzIE5oHwqOebEdJZHNtvHibiGcGALXJMMyQUUi6kTDDsBC1GGYQpZhfvv
kvG7oxt/RyJ6BW0xfvXbyQETLF6qMTN/ePpmGeT3lSQ9acMDyR3cRi/fApwtfs1a
NgUM3bLyviqVq1+PHP1/lH/jesqFUPN/+ymbRCsyWiCYeQLG3svEo/fQr7nvMTDa
lwBj3U9bIqpZE+HhXsZtvZniO9BRk+1N7SP6bxl4mehXLzKg9BtgpNRu42sd2CEi
dvEZUoYuGPmy8YtVEe71TefyzKFpC3FN6X1RQ9eUgctP+lwVD7+N/xN6TS1xXFnz
28RPB7zi/6S/NF6vmOU7VyCTTQEuUhwUyYL3lpfiNqEF6xmC/LhFJghmSvGt/Whl
3uLGeiFlXzP2tK0Q5jV4u/CzB8KRGbWheD4ImyJv3NLNugcZVJHsUrnPVlh4cKWF
OX118Mv1qThiRs0ZnM2n1u92oNNFkk10LBKIhgmD8t08TSZL9ZAajuRLTHo2Q7xr
gZCV+3Z7TWIlS9+dGScMLCtMceoFSBDkb2AjDSUsLFp1F1gopfhlSlTvwOoEIvFQ
UKUSWkPq8JxqbQimO/k7BoNqhBv/dmdOnWG5cTh0AgLEiR8derPTm0Auu/VCLLun
jPLRQWQvIyIkVErNZzV5m7Gmaai3Oz93UNT0+FdNYdtZJxSjj/3x7cLRSo23iRjH
gSZp9KumJROKhU4o3L3GRTZMYX4mMgbLNDtM/coQW0gXldYoppBHbApTFAgNznOC
OFcvtxHEBwcUilZOvGRMgM55LvtfsK9fUwh/Rzf2Tg+1CwgYJOqZ1iQKGQnYLsLa
bLUBBVlZcKflhwbrW5dNTyx/FWxcweP/AouW1Yawa/6H+TX9VR6czv6cJCzUvJWJ
I+7aPP+TlN7JYZjL2DqBLvJLMxcqlF82L8Iry5QYo6i4nFoouwkQ1XUyptwDIp/U
s4xWkmmjTM4q2OAF3zWniGUf93Vh7qnJG7Y8vjNuFGwjlzgV9NyTFxKmNp9Bo4JH
vsa1qQ3sRNDIeg2Q5e2yS/qgQy+IjT2eO65JLmP54Rg1fcaF/Mg3PSrWVMcYxA+z
uWRFPey/5Typ+SXHV0nPGLNs7kPD/lvR93MD6UZNreNi1e5XkbPiAaqLpBYYkjci
XcK20cyUV6rLnRFvB1s+fDn255GuyDwq2ovdZ3+UE2enWYgJ1gjyFYlqronTsssN
1YxFwThlcFm1gGTw4ThFwkawyscHBLVV5IRp9NAtv3JZLEjggTFSo+4Rs1aWBaBE
dj8vwkYSIrLZDg22RsTa1LshOkXexX1W+EQxM3MFE7ftjS7TGCUbfKE4BjucO2Le
aQ1F7+bs/O78B/P6OIhO4tB4hjl6QHEA0i7w8/IRBUK4ExezpPh5W8YxFGbQjhO5
5ZMpRvsQTDLdqz1dweBEiKuKXeP6ij1LTrxEQVVjTOzoWvkY6zk8wOsXQSu7aoxb
GTxHYRshbcG79+aFEkfdtHKEh2HqlXK6nXafnsi8YuXtaGET7wc+pXOaPPwPC4fK
Jv5e4Dt+UDqrxlIlvtJgVevEOT1g1w5lGrINv/dJPHC/mNzFKmr5Ph4HmAkWdTTd
hKJlN2lLoG5SHaoZq+znSlKEXH5s2hFJotelf/zImFRuiRovODD/BCssXcgI68XO
jURXZ2P/IBJyDcPLImVTjYJqsF7JOHPl5fWne0MfsoeTv3px/l/w4SeP7mVVT1Zc
pIb65MB37qmp9GsLzVermsMoq1mtJNY/pMWW/osWmFJNV5Th2Mznm4zLr8Dennpo
1sWYBGo+nLRgYuNjK75dlc/13svi0L4eytmoRAhhHU0K2HEwc2ycpRUSRNO154BR
bG4bi9+rH3qOSZKEL9t4LXhiJec1A2RARDbqo9qbyVurZC4lSc+HLJpmz1hIANA8
2oY2Jce4z0b+Z3I605YnvJzcL0bQ04m4qw6r+Y34Hx12dW4eWHB444Jqmojg2GrO
2fPHlTcruracct47ilcl3MszS8YRmALNpf0Y3XstufdZmbhpGPJgcio2yVimKmUY
g9yri+q5pHHkMA0j1xVJiYEQUALxba7l7GienoJ/MMOwh/OtDE7Zm7AveaoNo15w
UI8iEa6+n1D3t38+qwoAYitnGJ8XscEpXLeo1THhG1s3IGNbAUSBnHpNGi50F9rf
YaaT199Xn5BR/x9irBH6JfOz+X5hep351x+uyJahcH+xlBO0JLd9EDp8EqLz8D+d
8M4+p/t3iS3qSurldzYx3WxXLHYxCQOHCfCgTp6BOK7btv0ikDPiX4ADYTtQ0rtZ
6eauWY+h79bgMTlifH3MExyNhbTka+c+9w+p1fKTCjn9jw3hXYeDWfiHAG+KmQuv
RtbWZrxTycCRYLd42HhGTm90frrjQSB2MjhvjjiPUSraPLa31k+d0irNewZUt9Lk
2ZTI9jPmyd5Q1NhLatBnWTB66VfRPgyQ954UG6t3Nwv8i/nbtyVaGbR6pzXhMhjO
O/ewBxn5oMaoERSPPefSJctQVkvNSVXby3/7zQObrHlVciX9L9g+WM8jptKFZzjP
l4j0ZZGPCHTR/8q969Tq2hTt1/EReu2I0AhSCNvtk5CZfv8CW2PGviv39wtXUoFd
F4sdtypMhOXOuawuH0j6pyBzYwoEbzRZGQxKpRJUCF51YqTAFgJRlVL/ECzEii4a
G8Xf+AawXmZz9QeQtq7/ujuTR4sqLM9ZVQOK0RgMWKSpUcYkPoU8zxlLmrkG/Vp1
9j6LDuFG7KiF2GmQtQen1iekZbp5vRPwh07O2JD0qhdFD9AAlGWt/Qg6GEKpqD9s
nwPxaDb6+YmucLbbsr9z/3QqjAJsAPlgURhroEz77GJIh5mJAL89//1egLPzTKlb
YlJvzMUTuGZ6ThfPv2YW4HpPM7PuGPNWqn1XlcVlQeIki3LxPWi2w7KvDqBKMTzv
KyYFHv/i0K048I/ke0C8kOLY2zRzYZ95YazTiawQ24v5V7HZwcCwFFfIWv9IMljF
odNcviv+3yA155LtT1v0sJAYI96KhaYikdY3AqYJcPu9pbf0rz10BXHkvJwpTKg9
xNMdI89LBCT9NnkEg/0kly/iYkw4H3poFAvlL6HBulgfj7pRTzomtnVSLAPagA3K
kjvvC37VA6wVFi6rpTBUMAX6IxFYvkhZEtMh/Hcug4zFMP1A8gNtS8ycbZWdJGvb
4eLhVEOahCV81nsG1mYEoxB3sskhy0plnTjmqzvOvhr+uJA/4wlqVIW62zR4Ckgp
wE0KT6empvl1g6j5hCubtRCReKbG0F2m6vaZckNHy5+c9Atw4DM0XBFeScJHvlOi
3fWRX9K7Vtyrm6rXZt+oxQreAgr3kswKvmlOyyCp1vhtejmd6BJddZri3+K0dH5a
Br/v+6vrkwNDrGunLY8N0y9RHHx29SOjoi1c1ObtUrL0G8RXLi3cfNznmP6rXf4M
mGna38OjcyqLgH7wjGwHWvzoySr5SYDOTHy+36DvEfNYwklS18GHx/UnJUdjEW0M
KzTfc5/k+iv45VYLJwaasnbkV/aW8j48vl+4MuhcHx9TR9/YpNQRxisYlZMBl54M
wblTGs/D9uNZfgWsnol107gnSSA08L3YTydfTG3/QvAcVglKGsiL7kANy/R5zXpq
3eVgsGyH6qJCpIxluu0YsfL8pRgF64M8XoHPcAsKoeXzRpULBpd2QdSaPZXTVHeo
1PswS844UnMS6+3LDpjuxjmdYzRGSkoNuo0/EnLh14aOKVMWJOsX3lkQlFhMZunx
+4/domvZGc5umt7UnjCXs4jzTCxmg48BFTl6UCZM/TRz/Nn+tW+EtVJ+Ks50lDHZ
8CpMlNonE1V3xEJR/SouhyhC/t5ye8r9aKf3XMLoyHzt52mM0JdxhVo/THlhHA94
9Gzwp/RX9yv7O/ljEr3FQPds23Nr/MbX53Ybz4DfnIaHhcfxHOqDp45o5i/ZjhhA
HR+lBoTto+EMJHuHujX1KegNFUBLCQYy0ItWgSaC3sG/33adbOcYdBtwFZWL2v8b
59kdt8mstVJFueu7uLhIXJI4E2eY0cRyryszaTRMaFaR+1vJmsyQ7wquMTjE+2Oa
DfhuOqUGrkLcrGanj9Ih5spX3NAp3Ioo+wWqDtD74bfaE1OnI229l/XwrmcUBGzB
8dpNaWKLqVBYOZeb63iCl/24fdRehpcq+j8wnUf2rxicBZdsbKC/kaAr++mTZr/I
MXTdGKQ61nk+GRHyN7oX8mjcZV6OHPeVlXqGHDykZvzoIPxyoPXX92AdQgDn1mGn
brivHWDpgrm8SbPwcVigNpMPwe+RMvSjuhruoOU73G2FMtpfu3jP1J46hqgoXtp7
0P71YtlsZ+FJNFjR4MxWkSg+I7Cq50Cyia1j4eoErEbbDw9YvGfgWZB9Zl0qRzzt
bfYCGNCaWslesjGRVoIUs40GNnrrZpmmXPYgJ/HcpZmQqS2V+APuS/INV9E5Mz67
TajXjfAE0KrQuZg67PHbBdopgPlCSClspyAev7cf6knhR46rEDWibBnn9zKgosSN
5jnmCnrE64tSOtEt1w85jgLsU3HGF3QW/emUdv2FPNge7nNK59HiTVcMol6VdPwT
EVNo/7xXZpZuCkAWrD/mkzHpA568BivBfJQwvwwSQ4raacprjy9OZsLxLMkZG9a5
K64nNPvesChFtDe9GxYq/m52fCdM2W934tcU1P+in7T/14JkKpEcoD4opQ5EzVSy
u8iHPcK4nY5jSh80AijHJp4QvQ4q+QvTTN9yS16wqD/T6eHFQz2IbAdBvvK7Kr2r
mnAAQGcA3XqZdciuz80WYgFAgoWrQM+NbR//vkKqiMGVthVEfD3fM2AGuHSvrzCq
V9voC0gPVAjt06nVYEFxAvOkro5ILHFe1Fyi3YOY4wtTvLcnPu5We3jvcyVG7pNd
FmClNvp7myQoXCL0GtQRdrmVdCziS8MrExXiR/tZRaNRdJYSUZd1NMlqhoYKiteP
tD/8z2Zjx9pO7TDDvIX8Vvav/vvZzxFYciUeuzPjb0VjdQV6La1FN4tti24oMpQH
y2E1LA52J84gskTx0fq/wLZMsfUVq8Vu7Xu3BGUmI3COAkczgsWnXfgdez/nMM3f
nkoBWrRuyGubDp1X7jh0KRruwyGNlQXF4zvrn4VNcIiX1fFVd3yNIf3mICOKJKwO
8ItRvaE2hO1VmxnJsGRZvd5Hd7qnovYR4VtZehbkGKFozXejSZy/MLWvc8NRjVJu
K8cuFfUT1jijBlreSJu3zdj5Pu8oSjlHD+bzalNIsh4QqOVmNFH+LMPmnInNboWz
ZUu/OrOooGpljO4VG9cLTSvsxxThz6fzmmo61jOcJCZrGqveu+inxoS93luSVXVn
VilUVV02z/J14X46/FghozRDpP97vYlqaZsDjViDYRgGijX62jFMWliDasSN5dno
FRa89tdr5BM7SuPim+J3BJxBDnyvvOwAfvZpZu9rzi1BQ+F8cXJi/VYVWMkVcTCd
Di9U1dAhuEf3L4GhQQGqzRwY7d3AGgGey8vSZWfXbNVAGYB0U+Cuo/JZZNj3HAB9
M17BsWBs+V76HNwzysa7cutXC8KqeapTvXfo2fo8e4Qvcwme8NYn+RJhWRvhKGfv
OUPWEtrZPP/NYvjYY4+sz1r4AhALMSh2TnC6C4+JSwcH/iZJ62+AnMM1z1fOLBFL
lPatB5ybD6DEQIq5MrnxNDcnNEJioQe/8DTatclTZNVz0ibf3Eov7b4tiru5Aqqy
Jwq/uJWZ6BMAQkewaY6zamTUVmfyN0NBPUcAkoydlygP8imKoRO1OSFaMY8qcyZC
wpFZ7Cp4Z63csFC55g9Ol66kRRzHhhGwMZp7JfUd3Krk76IiQYyl/Rla1QYGk+jm
F5FwOyZJfipSxkRDGIl4uS8ELlrbXQYAqKYqsmrhxXuz1BDBh7GW0cbj4nGtEjxm
Zn1UiMOjLMeuil5nFFD/MxCIpqsOpDgg7z/1IJroieG8DRVH0h9JNLfDWCHnQE6K
dZJoasKDXONHe7yBpBhcnJ3i0FmwMxgGQahO32EJDU/aRrg9qdW5JzQHdG5ZlhUJ
wqAzjlCZk44mPwXyTOVxz9FsA+fYzBS2qNxGaDO0eROZ6x3HBAENz9bXC1CoIMfT
BsCMz0tG5tVJU/q+EjZ21Es5VOxYMhzhKEeJUeGIfb/WjVIAWZuf6twRcmMSdEwl
dfcdKRG31nBgMlLN0uOAFFKf5KZyqxTx9uwuuqYPJXuNfQ4v1RSRGXnU4NQPxOOr
wHVk82SqmrbfkS66ai2lOmATuwplOP88Et9riN/FqK8k7Fs+K3GLnLW7z80WrFbc
AFu2lxtpL95ggMXi+5KfS/wWZMqe62+5nBfeyc6qulmebmcR4DynUrhr4cViqIxg
BmW5Hg5fnw/FezBRO7oxxKh/x/+MBta7XQD11Vb11XWGFxhvA0JYylFGFN7rSHGX
0vd//N1uKZbVR4SoJ7QDw/ASPzB3FES5HyVBVNJ0vYK3Yjsw+89ied4Lz7gVx078
7juNzqhr5AZfpH9BPupVowj+w8s4UAIPyqOrPzXTy82qd49jIsMxGrBLTotftGzO
fTRJeuzZ3ELjfMOhUIEZ+GjYeZn5+WmNqnSJ1ub9fxgsmsXde8jfa7vKgKU9hM7q
qjzsyJGOVQ9I04OMvK6n08l/RdZnIoLh6DqUY+tgxu5oYIEBGTjnz8FvhBS7zaPb
CG2eVGD52cY5ry093ACamQRhT7BzQSWg5Deb/wmudABcJ1GAC9f97JydqT8Sf70E
qSQpXKkfCGYf+Vt1nc+o4qhpObX2zeEKUuFAjRqjt9h0JX0J0B37+RnAsKqyfGrh
L4fQIr0G5IEJmjY4DEHUk6Eevl7GlowzbzTKsxT2b06yTPKSUSaoqmH6dhJJp6Q7
1WA+1gycbB51RKgBSBBj6VthBNRo7NLi59wyHZAYhpbinSOWXVhXJT+QsMvobgny
FaCDPJJz3/kx5zjFJGLjZZucxgQ+jrdaFQnAVvg19ZcW+DtZICx2KDkH3muMJ5+x
GAj1Yf1xrnmNthYY2hpp71Eq0F377n7PzPmKId1FbnpT+UtkY84PXtVIW3qulsPb
g8b7N9ofcFiQ+8Bt6MAMW9RcPFrpcSPvO06UIhXSno7j+BPuIQaVgCIooTgPHNel
JytMQ3qhmu46zxsOvA2wDNJYb9+UmQgNuyrwR5xTgT0KTuD1Tb45XVnZOw2HAkLv
PZiUiExxBGdGKeMKiX1hq1Hm9TnzA5POk4DcLLmPNAw2hru9TU4w4SL/YQGNdAeK
gtPexstdIUMNuqSTBHtQy02jkxLvfmCjWT9uWQi2o1nxAvOn6kMT26ePeEl3MJm6
toO2Vf755xfZjxaT04jhxN6V86pg4XGIxOHjaBZVNk1mVoM1NVe+b98uOqFOABnY
KmOuiw9jJlvPcmLd5iZBJu2v93JgCbNiTbR7TA6qNGU8/yeLeMp3ZenE4nVHQpfm
kijsOONz8/GV53O5Y87vneu3H7JYMETaoP0E5nBHlTwtFsPvOVjzpkLrAhek5YaB
EtWzCvasB18lYu3xww1PcnHuaXXf3+liOIzs7udtS5CBUhmOGojatkZcqXbuCWHT
J/EYItoFHjSSwLCu2uw+QT8qVzWB+3kT1A2K85nlFEPFDqV7+5CR0RpHOlMpnjxe
EHlpD62Iitoj3TBzvDpK5IiOA40j/yfgjuF5GNR5v9ikvblCuF/body2kNmkcOFb
TTco66Y3lHMUUw/UgAnXcCaJxkWwkGJeF/7SmBNOfDnhVs4cvG5gYUibGrUwfqZZ
vl1NtpsYjg9ivre33NU6jfGuvPz0+UAhXPbdLrIdpK3Nxn5bA8Og5W1eWiCBxg7r
Ih0jGYULEuwjgMa0PivGObKS3+0tssPt7o+0z19xeBUPSEgLxTP93s3mM91sKGtD
LWqAMO2ehB3k/b9jtRxE/8gVA+KpvkVfYFilQ694xX5chSP4UW6cGfVv1+li56In
H4O8aN35BvH6re82UX/9GNyfZxE6Onxmfm+R0qEQHgNnGhBXSkgM0onbutTpstK3
x0Qe4XdhfD4fCB8mXhoTS1hVm7JROypr1UZhFX9SqD+HErh4SyEyl9Rf9wKQVqVv
YFJmHEQBryqg2UpQd0rLH/X3T/Me+jrQCL0FBRDL7xrkhYw8sNBsTXpQ7m3rGU+o
aJexOutYuAraygYPsJwcURhEfUohAyaJjmzeq3jvYN0SL59bakpz8l3OjBR/I8Gx
Xx4JiVMhPSilLv8kynpkxmbo6BbbvDj0BE8L4pQVuN80/vHvtnUWArgNVKJpQrXW
+lgenFRMeR2qV/Wb4HI7wbAtg5VGCIrPnfo+xQXhbknvCWWm5CWNVHQvTMqdVo3M
7ImVFKasxzvIAafEIBcau8BcyyyEnCwjlEsXNNPYHM58CR4cvfVQny3zPMn3J4w6
AFBgYFSnnoRY/p9EAOWx3mq3hKBWXzf/DaJ9JutaZUrxhglspWo+vA+87//cOIhO
nRTaAcNxW8Jv8Pavw0tXCTPajzsoc4+VvDWOkh3DlqtowV1KZE1oycfeKbvQnYz1
SxistMbFdJcpoM+CVAXnWrIwDDIZAA1UPpOJR9aGefYGprQf7TzP9+XDZ2hK/pQp
1cQ5oPReeaN4wME+SBr4YkeN+dEWorc936yLcGAhvKn93wBuhd8+4Qy+N1/NkJ9w
RAHw0amC0fp824/UCPWhYfxCNoGCqI9nQEcAWypXYQtxpDtuMNkBXMLVmAmvwXU8
nw6WwEF8oPntSyK284DSErcupaRRc9efVfrAJRQDuiJl+c4GYQlOSN5Y2oIdM0aW
J2ONA1gQLIEwRIBTiwtqqsiuyuC4X2F3G4pg6xUQT3VdPv9pg2EZ/BuZTxCS8Sld
9kLzUxGTu0XLVB9Xa5lgsKf0uccFdj9OEJo/sANMr1Ac5NsyNnQ/2KTxEhdFre6C
56mjpwfTHM99XbF+yyHn4VVoJDQD8vw6jKjleYVbIOCoQBNQ+HoGO5no+FKPAhrR
ooYblya2EYJAWYRtuCeTuVTyNZpFfVURQ3gBLkT+bNMQXvG917VjjwE384XSNccY
UHq6ZzO6cU1rk2NJrUpMOHz56cJpOzbip2dvVPiwGl3PujiiAwWgsrkXn/0dHPBZ
OMJ0AdSrvuD2RGrzy4DPrz4Zdb3eUVRKDyGtrexxb4T8tPZMjGbft1TkBYrRT/vE
GyBp6L9gvXE9NaO95CmVnUdOblu0bLKQbZ1uguapHtzX2bclYD4xVuDJTqhhoDkX
c34HI/bYxk3011Bq+fOD4ye9zo6k95f91t26yfucpKyTTj/oTSJez13KOyqcUzKx
1NP4RR/dA9t+5E+rii+Qr6KdINElrT1uU+TmAPxs0vypneNN119jr6V8pGx4vOTh
QLyX5vNq6hzxKEzimkNZ4siGR2/utbXICCj9zTjb1jExXPRbIMPG4DqgdnecYgW6
NFqE7n3sUl+ragLqis/CYZRrd41fbvbuV54pKmXIgxDC3hrHkU7MNefdqfnZeq12
baMri7OSlBAsO/14s1nTH+S6IhtXS/6r2WFbWShg48dRWxla8tIX3gRBiwt7cXvg
73VXo7d1Z0WwZhDV0tOg54o5kOmKQMMf2ap3WtcyOQg8S3EuG7L7oGMQX0nVDjKL
TGyWKRylvkQbnNiclq8TrEFHexADawB3QNDzD4pf2AucXJ6LJ5t0sgbI0tu17zN1
q8eJK/+5YbpG5XpbwxikztP381uWyTa5m2cw/ciMpcv6thZr00BfGK56ikovKF/N
UZ74dO30yQIkU0Zg1xYZTXJvfqX16i1etuTzK9PlZJpLvuCQ/il5xKxNMj7dTXYy
+lmITHsl+VW28Mw+Bu5uqBuuL/n5aP4Q7H1Oi3kkBcX/0YY4ZqcHnvtT5Ffiu3HN
j2eBXLGmnxi/svgZ5svc1WkOMRh9ii/55ZjoT9w1bmcPBxc+5oo/wNEps2KeaxLm
mLWcmuJH8XVI+9BdlHgki0xm3LHozcye+Z7j79l4AeYLRSlcmfsYmeK0plgQRbVd
pSjzBu+E7kuS3DmOJoDL4JHVUxVoHUNwM/5DaNzK6/EwOrCfbOud+5VpH7eS0rKm
4si4Qst7tCypeoa8uI/X//IAPTPCk9ZDP+VQMLmNyHM=
`pragma protect end_protected
